

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761;

  OAI21_X1 U11028 ( .B1(n17021), .B2(n17026), .A(n17015), .ZN(n20009) );
  INV_X1 U11029 ( .A(n20649), .ZN(n14836) );
  NAND2_X1 U11030 ( .A1(n19131), .A2(n14203), .ZN(n18408) );
  INV_X1 U11031 ( .A(n21758), .ZN(n20282) );
  NOR3_X1 U11032 ( .A1(n17225), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17061) );
  AOI21_X1 U11033 ( .B1(n11784), .B2(n11783), .A(n10159), .ZN(n11785) );
  INV_X1 U11034 ( .A(n11221), .ZN(n12928) );
  AND2_X1 U11035 ( .A1(n14022), .A2(n10984), .ZN(n11082) );
  AND2_X1 U11036 ( .A1(n14022), .A2(n10982), .ZN(n11057) );
  CLKBUF_X1 U11037 ( .A(n18116), .Z(n9588) );
  INV_X1 U11038 ( .A(n18095), .ZN(n18210) );
  INV_X1 U11039 ( .A(n9602), .ZN(n18209) );
  INV_X2 U11040 ( .A(n12689), .ZN(n19868) );
  AND3_X1 U11041 ( .A1(n11562), .A2(n20829), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11891) );
  AND2_X1 U11042 ( .A1(n10423), .A2(n10422), .ZN(n14409) );
  INV_X1 U11043 ( .A(n18095), .ZN(n18220) );
  CLKBUF_X2 U11044 ( .A(n18224), .Z(n9603) );
  NAND2_X1 U11045 ( .A1(n20824), .A2(n21581), .ZN(n11950) );
  CLKBUF_X2 U11046 ( .A(n12578), .Z(n12496) );
  AND2_X2 U11047 ( .A1(n9820), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13594) );
  AND2_X1 U11048 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11453) );
  CLKBUF_X1 U11049 ( .A(n20845), .Z(n9584) );
  NOR2_X1 U11050 ( .A1(n20797), .A2(n20796), .ZN(n20845) );
  CLKBUF_X1 U11051 ( .A(n21440), .Z(n9585) );
  NOR2_X1 U11052 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21440) );
  CLKBUF_X2 U11053 ( .A(n11724), .Z(n12602) );
  CLKBUF_X2 U11054 ( .A(n11719), .Z(n12603) );
  NOR2_X1 U11055 ( .A1(n11827), .A2(n11717), .ZN(n11824) );
  BUF_X1 U11056 ( .A(n10950), .Z(n11221) );
  AND3_X2 U11057 ( .A1(n10799), .A2(n10798), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16196) );
  INV_X1 U11058 ( .A(n9601), .ZN(n18123) );
  NAND2_X1 U11059 ( .A1(n13654), .A2(n10597), .ZN(n18095) );
  INV_X1 U11060 ( .A(n9761), .ZN(n13915) );
  NAND2_X1 U11061 ( .A1(n10570), .A2(n11458), .ZN(n11554) );
  INV_X2 U11062 ( .A(n12056), .ZN(n12072) );
  AND2_X2 U11063 ( .A1(n10078), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11158) );
  XNOR2_X1 U11064 ( .A(n10191), .B(n16973), .ZN(n16671) );
  INV_X1 U11065 ( .A(n17919), .ZN(n9597) );
  INV_X1 U11066 ( .A(n18116), .ZN(n9604) );
  INV_X1 U11069 ( .A(n16235), .ZN(n20549) );
  INV_X1 U11070 ( .A(n13027), .ZN(n12733) );
  NAND2_X1 U11072 ( .A1(n14158), .A2(n17215), .ZN(n18663) );
  AND2_X1 U11073 ( .A1(n10610), .A2(n13652), .ZN(n13897) );
  BUF_X1 U11074 ( .A(n15046), .Z(n15098) );
  INV_X1 U11075 ( .A(n19898), .ZN(n19911) );
  INV_X1 U11076 ( .A(n19978), .ZN(n20008) );
  INV_X1 U11077 ( .A(n20040), .ZN(n20018) );
  AND2_X1 U11078 ( .A1(n20209), .A2(n20269), .ZN(n21754) );
  NOR4_X2 U11079 ( .A1(n19631), .A2(n19628), .A3(n19626), .A4(n17563), .ZN(
        n17531) );
  AND2_X1 U11080 ( .A1(n18637), .A2(n17066), .ZN(n18566) );
  INV_X1 U11081 ( .A(n18732), .ZN(n18714) );
  INV_X2 U11082 ( .A(n13880), .ZN(n14144) );
  NAND2_X2 U11083 ( .A1(n10871), .A2(n10870), .ZN(n17030) );
  INV_X2 U11084 ( .A(n13869), .ZN(n18125) );
  AND3_X2 U11085 ( .A1(n10799), .A2(n10798), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9586) );
  NAND3_X2 U11086 ( .A1(n9634), .A2(n11009), .A3(n9708), .ZN(n9934) );
  NAND3_X2 U11087 ( .A1(n10282), .A2(n11704), .A3(n11703), .ZN(n9836) );
  XNOR2_X1 U11088 ( .A(n11655), .B(n11654), .ZN(n20894) );
  NOR2_X2 U11089 ( .A1(n11324), .A2(n11100), .ZN(n9900) );
  XNOR2_X2 U11090 ( .A(n14501), .B(n14500), .ZN(n14557) );
  AND2_X4 U11091 ( .A1(n14112), .A2(n14351), .ZN(n10846) );
  AND2_X2 U11092 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14112) );
  BUF_X4 U11093 ( .A(n10809), .Z(n16026) );
  AOI21_X2 U11094 ( .B1(n15274), .B2(n15273), .A(n11779), .ZN(n11780) );
  NAND2_X1 U11095 ( .A1(n10596), .A2(n19524), .ZN(n18116) );
  AND2_X1 U11096 ( .A1(n16195), .A2(n14341), .ZN(n9589) );
  AND2_X1 U11097 ( .A1(n16195), .A2(n14341), .ZN(n16048) );
  INV_X1 U11098 ( .A(n10620), .ZN(n9590) );
  INV_X2 U11099 ( .A(n10620), .ZN(n9591) );
  AND2_X1 U11100 ( .A1(n10595), .A2(n19524), .ZN(n13906) );
  NAND2_X2 U11101 ( .A1(n10108), .A2(n10948), .ZN(n11150) );
  NOR3_X2 U11102 ( .A1(n12642), .A2(n12641), .A3(n12644), .ZN(n10792) );
  NAND2_X2 U11103 ( .A1(n15069), .A2(n10196), .ZN(n11852) );
  INV_X1 U11104 ( .A(n18095), .ZN(n9592) );
  AND2_X4 U11105 ( .A1(n10527), .A2(n13594), .ZN(n12578) );
  NOR2_X2 U11106 ( .A1(n14189), .A2(n14190), .ZN(n15541) );
  AOI21_X2 U11107 ( .B1(n11158), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10925), .ZN(n10927) );
  AND2_X4 U11108 ( .A1(n14105), .A2(n14334), .ZN(n10876) );
  INV_X1 U11109 ( .A(n16141), .ZN(n9593) );
  INV_X1 U11111 ( .A(n9593), .ZN(n9595) );
  NAND3_X2 U11112 ( .A1(n9816), .A2(n9815), .A3(n10031), .ZN(n10191) );
  NAND2_X1 U11113 ( .A1(n15179), .A2(n10287), .ZN(n15162) );
  OAI21_X1 U11114 ( .B1(n16772), .B2(n13121), .A(n16800), .ZN(n16759) );
  INV_X1 U11115 ( .A(n9961), .ZN(n9596) );
  OR2_X1 U11116 ( .A1(n16954), .A2(n12890), .ZN(n16937) );
  NAND2_X1 U11117 ( .A1(n14038), .A2(n14021), .ZN(n20169) );
  NAND2_X1 U11118 ( .A1(n20776), .A2(n11710), .ZN(n9856) );
  NAND2_X1 U11119 ( .A1(n14250), .A2(n14249), .ZN(n20593) );
  OR2_X2 U11120 ( .A1(n18664), .A2(n17251), .ZN(n18645) );
  INV_X1 U11121 ( .A(n18745), .ZN(n18812) );
  AND2_X1 U11122 ( .A1(n17573), .A2(n10756), .ZN(n17551) );
  OR2_X1 U11123 ( .A1(n17451), .A2(n19102), .ZN(n18745) );
  NAND2_X1 U11124 ( .A1(n17451), .A2(n14476), .ZN(n18807) );
  NAND2_X1 U11125 ( .A1(n19520), .A2(n19675), .ZN(n17451) );
  AND2_X1 U11126 ( .A1(n17616), .A2(n10548), .ZN(n17573) );
  NAND2_X1 U11127 ( .A1(n9916), .A2(n16848), .ZN(n16850) );
  NOR2_X1 U11128 ( .A1(n14199), .A2(n10359), .ZN(n18389) );
  AND3_X1 U11129 ( .A1(n10114), .A2(n17055), .A3(n10113), .ZN(n9623) );
  INV_X2 U11130 ( .A(n18971), .ZN(n18994) );
  NOR2_X4 U11131 ( .A1(n11297), .A2(n11296), .ZN(n11295) );
  NAND2_X1 U11132 ( .A1(n10253), .A2(n9682), .ZN(n12654) );
  NAND3_X1 U11133 ( .A1(n10199), .A2(n10919), .A3(n9996), .ZN(n10931) );
  NAND2_X1 U11134 ( .A1(n9926), .A2(n10910), .ZN(n10256) );
  NAND2_X1 U11135 ( .A1(n17260), .A2(n19131), .ZN(n10727) );
  AND3_X1 U11136 ( .A1(n12868), .A2(n10922), .A3(n9926), .ZN(n10199) );
  CLKBUF_X2 U11137 ( .A(n10916), .Z(n16235) );
  CLKBUF_X1 U11138 ( .A(n11947), .Z(n12050) );
  AND2_X1 U11139 ( .A1(n12127), .A2(n11554), .ZN(n13187) );
  NAND2_X2 U11140 ( .A1(n20834), .A2(n11940), .ZN(n12065) );
  OR2_X1 U11141 ( .A1(n10675), .A2(n10674), .ZN(n19122) );
  BUF_X2 U11142 ( .A(n11595), .Z(n20829) );
  INV_X2 U11143 ( .A(n10182), .ZN(n10916) );
  NAND2_X2 U11144 ( .A1(n10331), .A2(n10330), .ZN(n11246) );
  NAND2_X2 U11145 ( .A1(n11498), .A2(n10569), .ZN(n20824) );
  CLKBUF_X2 U11146 ( .A(n12605), .Z(n12395) );
  INV_X1 U11147 ( .A(n9608), .ZN(n9610) );
  INV_X4 U11148 ( .A(n17878), .ZN(n18205) );
  CLKBUF_X3 U11149 ( .A(n9600), .Z(n12449) );
  AND2_X1 U11150 ( .A1(n10527), .A2(n11453), .ZN(n11467) );
  CLKBUF_X2 U11151 ( .A(n9605), .Z(n9606) );
  CLKBUF_X2 U11152 ( .A(n12456), .Z(n9607) );
  NAND2_X1 U11153 ( .A1(n10596), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18224) );
  INV_X2 U11154 ( .A(n17751), .ZN(n17878) );
  AND3_X1 U11155 ( .A1(n9882), .A2(n10607), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10596) );
  INV_X2 U11156 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19524) );
  INV_X2 U11157 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11569) );
  AND2_X1 U11158 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14105) );
  INV_X4 U11159 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14341) );
  AND2_X1 U11160 ( .A1(n10128), .A2(n10126), .ZN(n15080) );
  NAND2_X1 U11161 ( .A1(n16470), .A2(n13147), .ZN(n13154) );
  OAI21_X1 U11162 ( .B1(n16846), .B2(n16861), .A(n16526), .ZN(n16528) );
  AND2_X1 U11163 ( .A1(n9963), .A2(n9962), .ZN(n15118) );
  NAND2_X1 U11164 ( .A1(n9789), .A2(n16914), .ZN(n9784) );
  NAND2_X1 U11165 ( .A1(n15162), .A2(n15154), .ZN(n15164) );
  OAI21_X2 U11166 ( .B1(n15046), .B2(n9763), .A(n15220), .ZN(n15069) );
  NAND2_X1 U11167 ( .A1(n16568), .A2(n9775), .ZN(n16846) );
  AOI21_X1 U11168 ( .B1(n16740), .B2(n16984), .A(n9907), .ZN(n16741) );
  AND2_X1 U11169 ( .A1(n10020), .A2(n10015), .ZN(n14491) );
  OAI21_X1 U11170 ( .B1(n9964), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n9965), .ZN(n9963) );
  INV_X1 U11171 ( .A(n11849), .ZN(n15058) );
  NOR2_X1 U11172 ( .A1(n16567), .A2(n16875), .ZN(n16556) );
  AND2_X1 U11173 ( .A1(n10480), .A2(n16570), .ZN(n16560) );
  OAI21_X1 U11174 ( .B1(n16461), .B2(n16460), .A(n16459), .ZN(n16464) );
  AND2_X1 U11175 ( .A1(n10163), .A2(n9854), .ZN(n15179) );
  OR2_X1 U11176 ( .A1(n15187), .A2(n9712), .ZN(n10163) );
  OAI21_X1 U11177 ( .B1(n16229), .B2(n16166), .A(n16222), .ZN(n16216) );
  NAND2_X1 U11178 ( .A1(n9980), .A2(n10257), .ZN(n16511) );
  NAND2_X1 U11179 ( .A1(n9825), .A2(n11848), .ZN(n11849) );
  AND2_X1 U11180 ( .A1(n14602), .A2(n10538), .ZN(n14576) );
  NAND2_X1 U11181 ( .A1(n10032), .A2(n10036), .ZN(n16572) );
  NAND2_X1 U11182 ( .A1(n10076), .A2(n9678), .ZN(n14603) );
  NOR2_X1 U11183 ( .A1(n16227), .A2(n16226), .ZN(n16229) );
  OR2_X1 U11184 ( .A1(n17060), .A2(n10384), .ZN(n10383) );
  NAND2_X1 U11185 ( .A1(n10175), .A2(n10174), .ZN(n15229) );
  NAND2_X1 U11186 ( .A1(n9704), .A2(n10109), .ZN(n9907) );
  OR2_X1 U11187 ( .A1(n16146), .A2(n16145), .ZN(n16147) );
  NAND2_X1 U11188 ( .A1(n10368), .A2(n10366), .ZN(n13051) );
  NAND2_X1 U11189 ( .A1(n11823), .A2(n15256), .ZN(n15249) );
  NAND2_X1 U11190 ( .A1(n14441), .A2(n17240), .ZN(n17225) );
  NAND2_X1 U11191 ( .A1(n9948), .A2(n10047), .ZN(n15149) );
  AND2_X1 U11192 ( .A1(n18525), .A2(n14439), .ZN(n17114) );
  NAND2_X1 U11193 ( .A1(n10156), .A2(n10157), .ZN(n15258) );
  OR2_X1 U11194 ( .A1(n15377), .A2(n11844), .ZN(n15358) );
  NAND2_X1 U11195 ( .A1(n9780), .A2(n11144), .ZN(n10141) );
  NAND2_X1 U11196 ( .A1(n9920), .A2(n16800), .ZN(n13120) );
  XNOR2_X1 U11197 ( .A(n11144), .B(n11143), .ZN(n16654) );
  NAND2_X1 U11198 ( .A1(n20270), .A2(n20269), .ZN(n20347) );
  NAND2_X1 U11199 ( .A1(n20270), .A2(n20526), .ZN(n21758) );
  NAND2_X1 U11200 ( .A1(n10395), .A2(n10394), .ZN(n16263) );
  OR2_X1 U11201 ( .A1(n16847), .A2(n12897), .ZN(n9920) );
  NOR2_X1 U11202 ( .A1(n15151), .A2(n10178), .ZN(n10177) );
  OR2_X1 U11203 ( .A1(n11114), .A2(n16703), .ZN(n9927) );
  OR2_X2 U11204 ( .A1(n14503), .A2(n14235), .ZN(n20603) );
  INV_X1 U11205 ( .A(n10048), .ZN(n10047) );
  AND2_X1 U11206 ( .A1(n15165), .A2(n11837), .ZN(n15154) );
  NOR2_X1 U11207 ( .A1(n11323), .A2(n12723), .ZN(n10095) );
  XNOR2_X1 U11208 ( .A(n9856), .B(n20764), .ZN(n15283) );
  NAND2_X1 U11209 ( .A1(n11778), .A2(n11777), .ZN(n15272) );
  NAND2_X1 U11210 ( .A1(n9856), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11742) );
  NAND3_X1 U11211 ( .A1(n9934), .A2(n9741), .A3(n9932), .ZN(n11322) );
  NAND2_X1 U11212 ( .A1(n18697), .A2(n17065), .ZN(n18927) );
  NAND2_X1 U11213 ( .A1(n15155), .A2(n11836), .ZN(n15165) );
  NAND2_X1 U11214 ( .A1(n14095), .A2(n9740), .ZN(n16270) );
  NAND2_X1 U11215 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15185) );
  NAND2_X1 U11216 ( .A1(n14094), .A2(n14093), .ZN(n14095) );
  AND2_X1 U11217 ( .A1(n11807), .A2(n11806), .ZN(n15264) );
  AND3_X1 U11218 ( .A1(n10973), .A2(n10988), .A3(n10989), .ZN(n9861) );
  INV_X2 U11219 ( .A(n15239), .ZN(n15220) );
  AND2_X1 U11220 ( .A1(n15239), .A2(n11829), .ZN(n15247) );
  OR2_X1 U11221 ( .A1(n14181), .A2(n10023), .ZN(n9883) );
  AND2_X1 U11222 ( .A1(n11063), .A2(n11056), .ZN(n9992) );
  AND4_X1 U11223 ( .A1(n9987), .A2(n9990), .A3(n11062), .A4(n9986), .ZN(n9988)
         );
  AND4_X1 U11224 ( .A1(n11061), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9989)
         );
  OAI211_X1 U11225 ( .C1(n10229), .C2(n10225), .A(n10224), .B(n10222), .ZN(
        n14094) );
  AND2_X1 U11226 ( .A1(n18807), .A2(n9899), .ZN(n18817) );
  AND2_X1 U11227 ( .A1(n9799), .A2(n9798), .ZN(n11056) );
  OAI21_X1 U11228 ( .B1(n17130), .B2(n9756), .A(n18663), .ZN(n18642) );
  XNOR2_X1 U11229 ( .A(n11735), .B(n11743), .ZN(n12132) );
  AND2_X1 U11230 ( .A1(n10964), .A2(n9812), .ZN(n10973) );
  AND2_X2 U11231 ( .A1(n20594), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20611) );
  XNOR2_X1 U11232 ( .A(n11709), .B(n20780), .ZN(n10153) );
  NAND3_X1 U11233 ( .A1(n11743), .A2(n9832), .A3(n10281), .ZN(n11814) );
  AND2_X1 U11234 ( .A1(n14010), .A2(n10980), .ZN(n20349) );
  AND2_X1 U11235 ( .A1(n10281), .A2(n9836), .ZN(n11734) );
  AND2_X1 U11236 ( .A1(n14010), .A2(n10984), .ZN(n20261) );
  AND2_X1 U11237 ( .A1(n14022), .A2(n10985), .ZN(n11059) );
  NAND2_X1 U11238 ( .A1(n18739), .A2(n14164), .ZN(n14165) );
  NOR2_X1 U11239 ( .A1(n10022), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10021) );
  INV_X2 U11240 ( .A(n13800), .ZN(n20728) );
  NAND2_X1 U11241 ( .A1(n13823), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13824) );
  CLKBUF_X1 U11242 ( .A(n13577), .Z(n21118) );
  NAND2_X1 U11243 ( .A1(n9888), .A2(n14475), .ZN(n19520) );
  NAND2_X1 U11244 ( .A1(n10961), .A2(n15946), .ZN(n10963) );
  OR2_X1 U11245 ( .A1(n10205), .A2(n10204), .ZN(n9888) );
  NAND3_X1 U11246 ( .A1(n10060), .A2(n10059), .A3(n10056), .ZN(n13577) );
  XNOR2_X1 U11247 ( .A(n14163), .B(n14161), .ZN(n18740) );
  OAI211_X1 U11248 ( .C1(n10392), .C2(n9707), .A(n10168), .B(n10166), .ZN(
        n13823) );
  NAND2_X1 U11249 ( .A1(n12114), .A2(n11666), .ZN(n11733) );
  OR2_X1 U11250 ( .A1(n17806), .A2(n10764), .ZN(n17634) );
  NAND2_X1 U11251 ( .A1(n10392), .A2(n10391), .ZN(n12114) );
  NAND2_X1 U11252 ( .A1(n11364), .A2(n11419), .ZN(n11359) );
  NAND2_X1 U11253 ( .A1(n19695), .A2(n9889), .ZN(n10763) );
  NAND2_X1 U11254 ( .A1(n18943), .A2(n18994), .ZN(n19034) );
  OAI21_X1 U11255 ( .B1(n14124), .B2(n10375), .A(n9703), .ZN(n10026) );
  NAND2_X1 U11256 ( .A1(n11685), .A2(n11684), .ZN(n13679) );
  XNOR2_X1 U11257 ( .A(n12939), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13072) );
  NAND2_X1 U11258 ( .A1(n11675), .A2(n11674), .ZN(n11682) );
  NAND2_X1 U11259 ( .A1(n13242), .A2(n13241), .ZN(n13244) );
  NAND2_X1 U11260 ( .A1(n12120), .A2(n12121), .ZN(n11593) );
  AND2_X1 U11261 ( .A1(n10144), .A2(n10948), .ZN(n10953) );
  INV_X1 U11262 ( .A(n19081), .ZN(n18943) );
  NAND2_X1 U11263 ( .A1(n11715), .A2(n11714), .ZN(n20967) );
  OR2_X1 U11264 ( .A1(n11711), .A2(n11673), .ZN(n11675) );
  OR2_X1 U11265 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  OR2_X1 U11266 ( .A1(n11711), .A2(n14056), .ZN(n11715) );
  NAND2_X1 U11267 ( .A1(n13608), .A2(n10363), .ZN(n17278) );
  NOR2_X1 U11268 ( .A1(n9687), .A2(n10165), .ZN(n10168) );
  OAI21_X1 U11269 ( .B1(n18772), .B2(n18773), .A(n18774), .ZN(n9884) );
  NAND2_X1 U11270 ( .A1(n10942), .A2(n10941), .ZN(n10955) );
  AND2_X1 U11271 ( .A1(n10377), .A2(n18767), .ZN(n10376) );
  AND2_X1 U11272 ( .A1(n10365), .A2(n10364), .ZN(n13608) );
  AND2_X2 U11273 ( .A1(n11326), .A2(n9718), .ZN(n11331) );
  OR2_X1 U11274 ( .A1(n18783), .A2(n18782), .ZN(n9943) );
  AOI21_X1 U11275 ( .B1(n19111), .B2(n10724), .A(n13623), .ZN(n13603) );
  AND2_X1 U11276 ( .A1(n11574), .A2(n12062), .ZN(n11576) );
  CLKBUF_X1 U11277 ( .A(n12654), .Z(n13329) );
  NAND2_X1 U11278 ( .A1(n10221), .A2(n10220), .ZN(n9968) );
  OR2_X1 U11279 ( .A1(n13972), .A2(n18401), .ZN(n14143) );
  AND2_X1 U11280 ( .A1(n11933), .A2(n11565), .ZN(n13582) );
  NAND2_X1 U11281 ( .A1(n12660), .A2(n9803), .ZN(n10950) );
  NAND2_X2 U11282 ( .A1(n9993), .A2(n10923), .ZN(n11229) );
  NAND3_X1 U11283 ( .A1(n11560), .A2(n11559), .A3(n11558), .ZN(n11580) );
  AND2_X1 U11284 ( .A1(n10215), .A2(n10214), .ZN(n10728) );
  CLKBUF_X1 U11285 ( .A(n12868), .Z(n13524) );
  NAND2_X1 U11286 ( .A1(n9822), .A2(n13578), .ZN(n12062) );
  NAND2_X1 U11287 ( .A1(n13620), .A2(n19122), .ZN(n14199) );
  CLKBUF_X1 U11288 ( .A(n11588), .Z(n15567) );
  NAND2_X1 U11289 ( .A1(n11241), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12967) );
  NAND2_X1 U11290 ( .A1(n12655), .A2(n19860), .ZN(n9926) );
  AND2_X1 U11291 ( .A1(n14204), .A2(n14198), .ZN(n13958) );
  AND2_X2 U11292 ( .A1(n13529), .A2(n12688), .ZN(n13027) );
  CLKBUF_X1 U11293 ( .A(n10906), .Z(n14363) );
  NAND2_X1 U11294 ( .A1(n20834), .A2(n10054), .ZN(n11588) );
  AND2_X1 U11295 ( .A1(n14214), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17173) );
  AND2_X1 U11296 ( .A1(n10916), .A2(n17030), .ZN(n20557) );
  NAND3_X1 U11297 ( .A1(n9998), .A2(n12685), .A3(n12699), .ZN(n9969) );
  AND2_X1 U11298 ( .A1(n9996), .A2(n9800), .ZN(n10923) );
  NAND2_X4 U11299 ( .A1(n11717), .A2(n11716), .ZN(n11921) );
  AND2_X1 U11300 ( .A1(n13181), .A2(n12127), .ZN(n11550) );
  NAND2_X1 U11301 ( .A1(n11878), .A2(n11562), .ZN(n13772) );
  OR2_X1 U11302 ( .A1(n13904), .A2(n13903), .ZN(n14214) );
  OR2_X2 U11303 ( .A1(n20829), .A2(n21501), .ZN(n11717) );
  OR2_X1 U11304 ( .A1(n13921), .A2(n13920), .ZN(n13959) );
  NAND2_X1 U11305 ( .A1(n13421), .A2(n10182), .ZN(n16141) );
  NOR2_X2 U11306 ( .A1(n20839), .A2(n21503), .ZN(n12105) );
  INV_X2 U11307 ( .A(n11950), .ZN(n12056) );
  OR3_X1 U11308 ( .A1(n12208), .A2(n21702), .A3(n12207), .ZN(n12240) );
  OR2_X1 U11309 ( .A1(n10662), .A2(n10661), .ZN(n19117) );
  AND2_X1 U11310 ( .A1(n20550), .A2(n10916), .ZN(n10130) );
  OR2_X1 U11311 ( .A1(n10687), .A2(n10688), .ZN(n19127) );
  OR2_X2 U11312 ( .A1(n10648), .A2(n10647), .ZN(n19131) );
  INV_X1 U11313 ( .A(n12069), .ZN(n20819) );
  BUF_X2 U11314 ( .A(n11554), .Z(n20834) );
  OR2_X1 U11315 ( .A1(n11623), .A2(n11622), .ZN(n11648) );
  NAND2_X2 U11316 ( .A1(n17030), .A2(n10182), .ZN(n13038) );
  INV_X2 U11317 ( .A(n11246), .ZN(n12689) );
  OR2_X2 U11318 ( .A1(n13887), .A2(n13886), .ZN(n14198) );
  CLKBUF_X1 U11319 ( .A(n12068), .Z(n20839) );
  NAND2_X1 U11320 ( .A1(n20824), .A2(n12069), .ZN(n11930) );
  OR2_X1 U11321 ( .A1(n11025), .A2(n11024), .ZN(n11291) );
  AND4_X1 U11322 ( .A1(n13867), .A2(n13866), .A3(n13865), .A4(n13864), .ZN(
        n13875) );
  NAND2_X1 U11323 ( .A1(n10824), .A2(n10823), .ZN(n12656) );
  NAND2_X2 U11324 ( .A1(n9905), .A2(n9904), .ZN(n19860) );
  NAND2_X1 U11325 ( .A1(n9668), .A2(n9627), .ZN(n12068) );
  AND2_X2 U11326 ( .A1(n11507), .A2(n10568), .ZN(n12069) );
  NAND2_X1 U11327 ( .A1(n11487), .A2(n9677), .ZN(n11595) );
  NAND2_X2 U11328 ( .A1(n9860), .A2(n9859), .ZN(n10182) );
  AND4_X1 U11329 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11524) );
  AND4_X1 U11330 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11498) );
  AND4_X1 U11331 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11546) );
  AND4_X1 U11332 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11487) );
  AND4_X1 U11333 ( .A1(n11450), .A2(n11449), .A3(n11448), .A4(n11447), .ZN(
        n10570) );
  AND4_X1 U11334 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11507) );
  OR2_X1 U11335 ( .A1(n11477), .A2(n11476), .ZN(n11555) );
  CLKBUF_X1 U11336 ( .A(n11601), .Z(n12595) );
  AND4_X1 U11337 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11544) );
  AND4_X1 U11338 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11545) );
  CLKBUF_X2 U11339 ( .A(n18224), .Z(n9602) );
  BUF_X4 U11340 ( .A(n13897), .Z(n9601) );
  BUF_X2 U11341 ( .A(n11718), .Z(n11612) );
  INV_X1 U11342 ( .A(n9608), .ZN(n9611) );
  INV_X2 U11343 ( .A(n17919), .ZN(n14134) );
  INV_X1 U11344 ( .A(n9608), .ZN(n9612) );
  INV_X1 U11345 ( .A(n9608), .ZN(n9609) );
  INV_X2 U11346 ( .A(n9761), .ZN(n18233) );
  INV_X2 U11347 ( .A(n18116), .ZN(n18219) );
  AND2_X2 U11348 ( .A1(n14110), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16041) );
  AND2_X2 U11349 ( .A1(n10846), .A2(n14341), .ZN(n11026) );
  BUF_X2 U11350 ( .A(n12409), .Z(n12597) );
  NAND2_X1 U11351 ( .A1(n13654), .A2(n10598), .ZN(n13880) );
  INV_X2 U11352 ( .A(n17440), .ZN(n17442) );
  NAND2_X2 U11353 ( .A1(n17265), .A2(n9882), .ZN(n18227) );
  INV_X1 U11354 ( .A(n13868), .ZN(n9608) );
  BUF_X2 U11355 ( .A(n10804), .Z(n10881) );
  CLKBUF_X2 U11356 ( .A(n10809), .Z(n16086) );
  BUF_X2 U11357 ( .A(n10804), .Z(n16197) );
  AND2_X2 U11358 ( .A1(n10809), .A2(n14341), .ZN(n10995) );
  AND2_X2 U11359 ( .A1(n9586), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10996) );
  BUF_X2 U11360 ( .A(n10876), .Z(n16090) );
  CLKBUF_X3 U11361 ( .A(n10889), .Z(n16195) );
  AND2_X2 U11362 ( .A1(n14110), .A2(n14351), .ZN(n16042) );
  NOR2_X1 U11363 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10607), .ZN(
        n10610) );
  AND2_X1 U11364 ( .A1(n10093), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10809) );
  NOR2_X1 U11365 ( .A1(n10612), .A2(n19524), .ZN(n17265) );
  AND2_X1 U11366 ( .A1(n10594), .A2(n10607), .ZN(n13654) );
  AND2_X1 U11367 ( .A1(n10607), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10608) );
  BUF_X4 U11368 ( .A(n9605), .Z(n9598) );
  AND2_X2 U11369 ( .A1(n11569), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11451) );
  AND3_X1 U11370 ( .A1(n10594), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10595) );
  AND2_X1 U11371 ( .A1(n9833), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10527) );
  AND2_X1 U11372 ( .A1(n10093), .A2(n14334), .ZN(n10804) );
  BUF_X4 U11373 ( .A(n12456), .Z(n9599) );
  INV_X2 U11374 ( .A(n11596), .ZN(n9600) );
  AND2_X2 U11375 ( .A1(n14112), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14106) );
  INV_X2 U11376 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11673) );
  INV_X1 U11377 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14348) );
  INV_X1 U11378 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14351) );
  NOR2_X2 U11379 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10093) );
  AND2_X2 U11380 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U11381 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10612) );
  AND2_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10609) );
  NOR2_X2 U11383 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13609) );
  NOR2_X1 U11384 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10611) );
  AND2_X2 U11385 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U11386 ( .A1(n9900), .A2(n10095), .ZN(n11144) );
  NAND4_X1 U11387 ( .A1(n11578), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n11673), .A4(n9820), .ZN(n11596) );
  NAND2_X2 U11388 ( .A1(n10380), .A2(n18663), .ZN(n18556) );
  NOR2_X2 U11389 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17773), .ZN(n17754) );
  AND2_X4 U11390 ( .A1(n11451), .A2(n11452), .ZN(n11718) );
  AND2_X4 U11391 ( .A1(n10611), .A2(n13652), .ZN(n13898) );
  NOR2_X2 U11392 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17680), .ZN(n17679) );
  AND2_X2 U11393 ( .A1(n11452), .A2(n14060), .ZN(n9605) );
  AND2_X2 U11394 ( .A1(n11452), .A2(n14060), .ZN(n12456) );
  INV_X4 U11395 ( .A(n17266), .ZN(n18043) );
  AND2_X1 U11396 ( .A1(n13609), .A2(n10611), .ZN(n13868) );
  NAND2_X2 U11397 ( .A1(n14503), .A2(n14236), .ZN(n20649) );
  NOR2_X2 U11398 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17617), .ZN(n17601) );
  NAND2_X1 U11399 ( .A1(n10608), .A2(n13652), .ZN(n17919) );
  NOR2_X2 U11400 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17556), .ZN(n17545) );
  NOR2_X2 U11401 ( .A1(n17496), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n17484) );
  NOR2_X2 U11402 ( .A1(n17718), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17704) );
  CLKBUF_X1 U11403 ( .A(n20844), .Z(n9613) );
  NOR2_X1 U11404 ( .A1(n20798), .A2(n20797), .ZN(n20844) );
  AOI21_X1 U11405 ( .B1(n14557), .B2(n20737), .A(n14504), .ZN(n14505) );
  INV_X1 U11406 ( .A(n11246), .ZN(n12685) );
  OR3_X1 U11407 ( .A1(n11144), .A2(n11143), .A3(n21729), .ZN(n11146) );
  NAND2_X1 U11408 ( .A1(n10323), .A2(n10901), .ZN(n10221) );
  OAI211_X1 U11409 ( .C1(n11229), .C2(n15939), .A(n9802), .B(n10924), .ZN(
        n10925) );
  OR2_X1 U11410 ( .A1(n10950), .A2(n20429), .ZN(n9802) );
  INV_X1 U11411 ( .A(n9999), .ZN(n9998) );
  AND4_X1 U11412 ( .A1(n11129), .A2(n11128), .A3(n11127), .A4(n11126), .ZN(
        n11140) );
  AND4_X1 U11413 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11141) );
  AND4_X1 U11414 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11138) );
  INV_X1 U11415 ( .A(n10947), .ZN(n10148) );
  NAND2_X1 U11416 ( .A1(n11158), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10143) );
  OAI21_X1 U11417 ( .B1(n9959), .B2(n9954), .A(n9953), .ZN(n9957) );
  NAND2_X1 U11418 ( .A1(n15165), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U11419 ( .A1(n9961), .A2(n15140), .ZN(n9953) );
  NOR2_X1 U11420 ( .A1(n9958), .A2(n9956), .ZN(n9955) );
  AND2_X1 U11421 ( .A1(n9836), .A2(n10067), .ZN(n9832) );
  AND2_X1 U11422 ( .A1(n10390), .A2(n11799), .ZN(n10067) );
  INV_X1 U11423 ( .A(n11800), .ZN(n11799) );
  NAND2_X1 U11424 ( .A1(n11562), .A2(n21581), .ZN(n12015) );
  AND2_X1 U11425 ( .A1(n20834), .A2(n21581), .ZN(n11928) );
  NAND2_X1 U11426 ( .A1(n11431), .A2(n11430), .ZN(n13036) );
  NAND2_X1 U11427 ( .A1(n10334), .A2(n14341), .ZN(n10330) );
  NAND2_X1 U11428 ( .A1(n10335), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10331) );
  NAND2_X1 U11429 ( .A1(n10092), .A2(n10091), .ZN(n11412) );
  INV_X1 U11430 ( .A(n9818), .ZN(n10091) );
  OR2_X1 U11431 ( .A1(n15641), .A2(n11266), .ZN(n11422) );
  NAND2_X1 U11432 ( .A1(n9795), .A2(n9697), .ZN(n9788) );
  NAND2_X1 U11433 ( .A1(n16675), .A2(n11119), .ZN(n9795) );
  NAND2_X1 U11434 ( .A1(n10196), .A2(n9690), .ZN(n9853) );
  OR2_X2 U11435 ( .A1(n15078), .A2(n15059), .ZN(n10196) );
  AND2_X1 U11436 ( .A1(n9732), .A2(n15615), .ZN(n9970) );
  INV_X1 U11437 ( .A(n13123), .ZN(n9903) );
  NOR2_X2 U11438 ( .A1(n16511), .A2(n16769), .ZN(n16483) );
  NAND2_X1 U11439 ( .A1(n12911), .A2(n12910), .ZN(n16505) );
  INV_X1 U11440 ( .A(n16626), .ZN(n16609) );
  INV_X1 U11441 ( .A(n17342), .ZN(n9917) );
  NAND2_X1 U11442 ( .A1(n10115), .A2(n12671), .ZN(n10114) );
  AND2_X1 U11443 ( .A1(n14370), .A2(n9709), .ZN(n10115) );
  OAI21_X1 U11444 ( .B1(n15946), .B2(n13735), .A(n13453), .ZN(n13455) );
  NAND2_X1 U11445 ( .A1(n11055), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n9983) );
  NAND2_X1 U11446 ( .A1(n11743), .A2(n11770), .ZN(n10040) );
  OR2_X1 U11447 ( .A1(n11731), .A2(n11730), .ZN(n11772) );
  OR2_X1 U11448 ( .A1(n11562), .A2(n21501), .ZN(n11716) );
  XNOR2_X1 U11449 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10783) );
  AND2_X1 U11450 ( .A1(n16090), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11125) );
  OR2_X1 U11451 ( .A1(n11097), .A2(n11096), .ZN(n11253) );
  INV_X1 U11452 ( .A(n10141), .ZN(n11120) );
  AND2_X1 U11453 ( .A1(n11038), .A2(n9935), .ZN(n9933) );
  NAND2_X1 U11454 ( .A1(n9941), .A2(n9940), .ZN(n10142) );
  NAND2_X1 U11455 ( .A1(n10146), .A2(n10799), .ZN(n9940) );
  NAND2_X1 U11456 ( .A1(n12872), .A2(n10913), .ZN(n10545) );
  INV_X1 U11457 ( .A(n21581), .ZN(n11878) );
  INV_X2 U11458 ( .A(n14228), .ZN(n12619) );
  XNOR2_X1 U11459 ( .A(n11771), .B(n11770), .ZN(n12149) );
  NAND2_X1 U11460 ( .A1(n10284), .A2(n9834), .ZN(n11771) );
  NOR2_X1 U11461 ( .A1(n11733), .A2(n10285), .ZN(n10284) );
  INV_X1 U11462 ( .A(n9835), .ZN(n9834) );
  INV_X1 U11463 ( .A(n12587), .ZN(n14228) );
  NAND2_X1 U11464 ( .A1(n9630), .A2(n9854), .ZN(n9961) );
  INV_X1 U11465 ( .A(n9959), .ZN(n9952) );
  AND2_X1 U11466 ( .A1(n9736), .A2(n12002), .ZN(n10427) );
  NAND2_X1 U11467 ( .A1(n12162), .A2(n11928), .ZN(n10045) );
  NAND2_X1 U11468 ( .A1(n13824), .A2(n11653), .ZN(n11709) );
  NAND2_X1 U11469 ( .A1(n10171), .A2(n11627), .ZN(n11652) );
  NAND2_X1 U11470 ( .A1(n10392), .A2(n10172), .ZN(n10171) );
  INV_X1 U11471 ( .A(n11594), .ZN(n10124) );
  AND2_X1 U11472 ( .A1(n11331), .A2(n16299), .ZN(n11373) );
  NAND2_X1 U11473 ( .A1(n9909), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9859) );
  NAND2_X1 U11474 ( .A1(n9908), .A2(n14341), .ZN(n9860) );
  CLKBUF_X3 U11475 ( .A(n11125), .Z(n16043) );
  INV_X1 U11476 ( .A(n16270), .ZN(n10395) );
  AND2_X1 U11477 ( .A1(n9681), .A2(n14025), .ZN(n10413) );
  NOR2_X1 U11478 ( .A1(n15632), .A2(n10121), .ZN(n10120) );
  INV_X1 U11479 ( .A(n13145), .ZN(n10121) );
  NAND2_X1 U11480 ( .A1(n16873), .A2(n9655), .ZN(n10111) );
  OR2_X1 U11481 ( .A1(n15778), .A2(n11143), .ZN(n11394) );
  INV_X1 U11482 ( .A(n19751), .ZN(n10031) );
  OAI21_X1 U11483 ( .B1(n11322), .B2(n11323), .A(n9699), .ZN(n9815) );
  INV_X1 U11484 ( .A(n9997), .ZN(n9993) );
  INV_X1 U11485 ( .A(n11143), .ZN(n16690) );
  AND3_X1 U11486 ( .A1(n10940), .A2(n10939), .A3(n10938), .ZN(n10942) );
  NAND2_X1 U11487 ( .A1(n10562), .A2(n10965), .ZN(n10967) );
  OAI21_X2 U11488 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n12867) );
  NOR2_X1 U11489 ( .A1(n14143), .A2(n18397), .ZN(n14158) );
  NAND2_X1 U11490 ( .A1(n18733), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14445) );
  NOR2_X1 U11491 ( .A1(n14171), .A2(n14172), .ZN(n14174) );
  OAI21_X1 U11492 ( .B1(n10750), .B2(n10749), .A(n10753), .ZN(n13836) );
  INV_X1 U11493 ( .A(n13618), .ZN(n10749) );
  OAI21_X1 U11494 ( .B1(n13629), .B2(n13650), .A(n9895), .ZN(n10731) );
  INV_X1 U11495 ( .A(n9896), .ZN(n9895) );
  OAI21_X1 U11496 ( .B1(n10212), .B2(n13650), .A(n10212), .ZN(n9896) );
  NAND2_X1 U11497 ( .A1(n13458), .A2(n13645), .ZN(n10431) );
  INV_X1 U11498 ( .A(n12015), .ZN(n13645) );
  INV_X1 U11499 ( .A(n20568), .ZN(n13463) );
  NAND2_X1 U11500 ( .A1(n12371), .A2(n12370), .ZN(n12389) );
  AND2_X1 U11501 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12370) );
  INV_X1 U11502 ( .A(n12369), .ZN(n12371) );
  NOR2_X1 U11504 ( .A1(n11853), .A2(n13212), .ZN(n10195) );
  NOR2_X2 U11505 ( .A1(n14510), .A2(n13209), .ZN(n14527) );
  NAND2_X1 U11506 ( .A1(n9830), .A2(n9693), .ZN(n15059) );
  AND2_X1 U11507 ( .A1(n9828), .A2(n9826), .ZN(n9830) );
  NAND2_X1 U11508 ( .A1(n9827), .A2(n15067), .ZN(n9826) );
  NOR2_X1 U11509 ( .A1(n11825), .A2(n13725), .ZN(n11826) );
  NAND2_X1 U11510 ( .A1(n15570), .A2(n21501), .ZN(n12622) );
  XNOR2_X1 U11511 ( .A(n13036), .B(n11432), .ZN(n13109) );
  INV_X1 U11512 ( .A(n15955), .ZN(n19746) );
  NOR2_X1 U11513 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13006) );
  INV_X1 U11514 ( .A(n11157), .ZN(n12930) );
  INV_X1 U11515 ( .A(n15600), .ZN(n15585) );
  NAND2_X1 U11516 ( .A1(n15594), .A2(n11429), .ZN(n16430) );
  INV_X1 U11517 ( .A(n10467), .ZN(n10466) );
  OAI21_X1 U11518 ( .B1(n10469), .B2(n9641), .A(n11412), .ZN(n10468) );
  OAI21_X1 U11519 ( .B1(n10470), .B2(n11426), .A(n9624), .ZN(n10467) );
  AND2_X1 U11520 ( .A1(n9809), .A2(n9624), .ZN(n16441) );
  NAND2_X1 U11521 ( .A1(n16439), .A2(n16438), .ZN(n9809) );
  AND2_X1 U11522 ( .A1(n11412), .A2(n10474), .ZN(n16439) );
  NAND2_X1 U11523 ( .A1(n10325), .A2(n9774), .ZN(n10328) );
  NOR2_X1 U11524 ( .A1(n13147), .A2(n13121), .ZN(n10326) );
  NAND2_X1 U11525 ( .A1(n16483), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16470) );
  AOI21_X1 U11526 ( .B1(n10485), .B2(n10483), .A(n10482), .ZN(n10481) );
  OAI21_X1 U11527 ( .B1(n13051), .B2(n10035), .A(n10033), .ZN(n10477) );
  INV_X1 U11528 ( .A(n12909), .ZN(n10482) );
  AND2_X1 U11529 ( .A1(n10490), .A2(n12906), .ZN(n10489) );
  NAND2_X1 U11530 ( .A1(n16572), .A2(n16569), .ZN(n10480) );
  INV_X1 U11531 ( .A(n16567), .ZN(n16557) );
  NAND4_X1 U11532 ( .A1(n16667), .A2(n10460), .A3(n11146), .A4(n9788), .ZN(
        n9796) );
  AND2_X1 U11533 ( .A1(n9919), .A2(n9918), .ZN(n17342) );
  NAND2_X1 U11534 ( .A1(n13235), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9918) );
  AND2_X1 U11535 ( .A1(n9623), .A2(n14372), .ZN(n16844) );
  NAND2_X1 U11536 ( .A1(n13745), .A2(n13744), .ZN(n14008) );
  NAND2_X1 U11537 ( .A1(n12652), .A2(n12651), .ZN(n14370) );
  NAND2_X1 U11538 ( .A1(n12650), .A2(n12649), .ZN(n12651) );
  INV_X1 U11539 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20552) );
  NOR2_X1 U11540 ( .A1(n13613), .A2(n10731), .ZN(n19517) );
  INV_X1 U11541 ( .A(n17278), .ZN(n13613) );
  NOR2_X1 U11542 ( .A1(n18054), .A2(n18075), .ZN(n10319) );
  AND2_X1 U11543 ( .A1(n10314), .A2(n10313), .ZN(n17259) );
  NAND2_X1 U11544 ( .A1(n10316), .A2(n10315), .ZN(n10314) );
  NAND2_X1 U11545 ( .A1(n14193), .A2(n19513), .ZN(n10313) );
  NOR2_X1 U11546 ( .A1(n19131), .A2(n19117), .ZN(n10315) );
  INV_X1 U11547 ( .A(n19034), .ZN(n9886) );
  NAND2_X1 U11548 ( .A1(n9894), .A2(n9679), .ZN(n9890) );
  AND2_X1 U11549 ( .A1(n14363), .A2(n20557), .ZN(n20536) );
  OAI21_X1 U11550 ( .B1(n15590), .B2(n15591), .A(n13095), .ZN(n16731) );
  AND2_X1 U11551 ( .A1(n16700), .A2(n13675), .ZN(n16697) );
  NAND2_X1 U11552 ( .A1(n16700), .A2(n20516), .ZN(n16682) );
  NAND2_X1 U11553 ( .A1(n16746), .A2(n16744), .ZN(n16737) );
  NAND2_X1 U11554 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  NAND2_X1 U11555 ( .A1(n10006), .A2(n9867), .ZN(n10004) );
  NAND2_X1 U11556 ( .A1(n10008), .A2(n10010), .ZN(n10005) );
  NAND2_X1 U11557 ( .A1(n16849), .A2(n10198), .ZN(n10010) );
  NOR2_X1 U11558 ( .A1(n17337), .A2(n17338), .ZN(n16974) );
  NOR2_X1 U11559 ( .A1(n10043), .A2(n11786), .ZN(n10042) );
  INV_X1 U11560 ( .A(n11770), .ZN(n10043) );
  AOI21_X1 U11561 ( .B1(n11866), .B2(n11865), .A(n11858), .ZN(n11864) );
  OAI22_X1 U11562 ( .A1(n16235), .A2(n10447), .B1(n13038), .B2(n12641), .ZN(
        n10446) );
  NAND2_X1 U11563 ( .A1(n13492), .A2(n12641), .ZN(n10447) );
  NAND2_X1 U11564 ( .A1(n20550), .A2(n10180), .ZN(n12638) );
  INV_X1 U11565 ( .A(n11732), .ZN(n10286) );
  NAND2_X1 U11566 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11998) );
  OR2_X1 U11567 ( .A1(n11765), .A2(n11764), .ZN(n11802) );
  NOR2_X1 U11568 ( .A1(n10062), .A2(n10058), .ZN(n10057) );
  INV_X1 U11569 ( .A(n11671), .ZN(n10058) );
  NAND2_X1 U11570 ( .A1(n11588), .A2(n20824), .ZN(n11560) );
  NAND2_X1 U11571 ( .A1(n12065), .A2(n20819), .ZN(n11558) );
  NOR2_X1 U11572 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21623), .ZN(
        n11863) );
  XNOR2_X1 U11573 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10780) );
  AOI21_X1 U11574 ( .B1(n10784), .B2(n10783), .A(n10782), .ZN(n10786) );
  NAND4_X1 U11575 ( .A1(n12867), .A2(n12656), .A3(n19860), .A4(n19879), .ZN(
        n10902) );
  INV_X1 U11576 ( .A(n11283), .ZN(n10338) );
  NOR2_X1 U11577 ( .A1(n13038), .A2(n20559), .ZN(n10220) );
  NOR2_X1 U11578 ( .A1(n9595), .A2(n14017), .ZN(n14019) );
  INV_X1 U11579 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14017) );
  AND2_X1 U11580 ( .A1(n10474), .A2(n11420), .ZN(n10472) );
  NAND2_X1 U11581 ( .A1(n9946), .A2(n11410), .ZN(n10260) );
  NOR2_X1 U11582 ( .A1(n16141), .A2(n20550), .ZN(n9803) );
  NOR2_X1 U11583 ( .A1(n19879), .A2(n20559), .ZN(n9901) );
  NAND2_X2 U11584 ( .A1(n9991), .A2(n11076), .ZN(n11323) );
  NAND4_X1 U11585 ( .A1(n9989), .A2(n11064), .A3(n9988), .A4(n9992), .ZN(n9991) );
  NAND2_X1 U11586 ( .A1(n11099), .A2(n9786), .ZN(n11101) );
  NAND2_X1 U11587 ( .A1(n9932), .A2(n9935), .ZN(n9786) );
  OR2_X1 U11588 ( .A1(n9968), .A2(n14334), .ZN(n9939) );
  INV_X1 U11589 ( .A(n10944), .ZN(n10146) );
  NAND2_X1 U11590 ( .A1(n10219), .A2(n10218), .ZN(n10938) );
  AOI21_X1 U11591 ( .B1(n12682), .B2(n17030), .A(n20559), .ZN(n10218) );
  OAI21_X1 U11592 ( .B1(n12864), .B2(n12865), .A(n9667), .ZN(n10219) );
  INV_X1 U11593 ( .A(n19860), .ZN(n10912) );
  OR2_X1 U11594 ( .A1(n11036), .A2(n11035), .ZN(n12701) );
  NAND2_X1 U11595 ( .A1(n10899), .A2(n10900), .ZN(n12875) );
  AND2_X1 U11596 ( .A1(n10909), .A2(n12656), .ZN(n10217) );
  NOR2_X1 U11597 ( .A1(n18227), .A2(n10628), .ZN(n9893) );
  NOR2_X1 U11598 ( .A1(n19127), .A2(n19117), .ZN(n10215) );
  NOR2_X1 U11599 ( .A1(n11554), .A2(n11595), .ZN(n13181) );
  NOR2_X1 U11600 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12587) );
  NAND2_X1 U11601 ( .A1(n14506), .A2(n10542), .ZN(n10541) );
  INV_X1 U11602 ( .A(n14589), .ZN(n10542) );
  NAND2_X1 U11603 ( .A1(n12315), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12590) );
  NOR2_X1 U11604 ( .A1(n10532), .A2(n14732), .ZN(n10072) );
  NAND2_X1 U11605 ( .A1(n10534), .A2(n10533), .ZN(n10532) );
  INV_X1 U11606 ( .A(n14678), .ZN(n10533) );
  NAND2_X1 U11607 ( .A1(n14701), .A2(n10537), .ZN(n10536) );
  INV_X1 U11608 ( .A(n14723), .ZN(n10537) );
  AND2_X1 U11609 ( .A1(n12213), .A2(n10530), .ZN(n10529) );
  INV_X1 U11610 ( .A(n14841), .ZN(n10530) );
  INV_X1 U11611 ( .A(n12068), .ZN(n12127) );
  NAND2_X1 U11612 ( .A1(n12047), .A2(n9850), .ZN(n9849) );
  INV_X1 U11613 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U11614 ( .A1(n14649), .A2(n10435), .ZN(n10434) );
  INV_X1 U11615 ( .A(n14660), .ZN(n10435) );
  INV_X1 U11616 ( .A(n9843), .ZN(n9842) );
  OAI21_X1 U11617 ( .B1(n14530), .B2(P1_EBX_REG_22__SCAN_IN), .A(n12072), .ZN(
        n9843) );
  NAND2_X1 U11618 ( .A1(n10388), .A2(n9855), .ZN(n11846) );
  AND3_X1 U11619 ( .A1(n9854), .A2(n9630), .A3(n9771), .ZN(n9855) );
  AND2_X1 U11620 ( .A1(n11845), .A2(n11844), .ZN(n10389) );
  NAND2_X1 U11621 ( .A1(n12047), .A2(n9847), .ZN(n9846) );
  INV_X1 U11622 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n9847) );
  INV_X1 U11623 ( .A(n9841), .ZN(n9840) );
  OAI21_X1 U11624 ( .B1(n14530), .B2(P1_EBX_REG_18__SCAN_IN), .A(n12072), .ZN(
        n9841) );
  INV_X1 U11625 ( .A(n9839), .ZN(n9838) );
  OAI21_X1 U11626 ( .B1(n14530), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12072), .ZN(
        n9839) );
  INV_X1 U11627 ( .A(n14751), .ZN(n10430) );
  INV_X1 U11628 ( .A(n14762), .ZN(n12009) );
  NOR2_X1 U11629 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  INV_X1 U11630 ( .A(n11834), .ZN(n10064) );
  NAND2_X1 U11631 ( .A1(n15202), .A2(n15200), .ZN(n10065) );
  INV_X1 U11632 ( .A(n14830), .ZN(n10428) );
  INV_X1 U11633 ( .A(n14846), .ZN(n11990) );
  INV_X1 U11634 ( .A(n14843), .ZN(n11991) );
  NAND2_X1 U11635 ( .A1(n15249), .A2(n11831), .ZN(n10179) );
  INV_X1 U11636 ( .A(n15257), .ZN(n9951) );
  OAI21_X1 U11637 ( .B1(n15256), .B2(n10049), .A(n11833), .ZN(n10048) );
  NOR2_X1 U11638 ( .A1(n10170), .A2(n10173), .ZN(n10167) );
  INV_X1 U11639 ( .A(n11627), .ZN(n10169) );
  NOR2_X1 U11640 ( .A1(n11717), .A2(n11818), .ZN(n11656) );
  OR2_X1 U11641 ( .A1(n11607), .A2(n11606), .ZN(n11657) );
  AOI21_X1 U11642 ( .B1(n11655), .B2(n11654), .A(n11824), .ZN(n11661) );
  NOR2_X1 U11643 ( .A1(n13182), .A2(n20834), .ZN(n13578) );
  INV_X1 U11644 ( .A(n11580), .ZN(n10055) );
  INV_X1 U11645 ( .A(n20856), .ZN(n20932) );
  AND2_X1 U11646 ( .A1(n11712), .A2(n21489), .ZN(n21120) );
  INV_X1 U11647 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21195) );
  NOR2_X1 U11648 ( .A1(n11424), .A2(n11423), .ZN(n11431) );
  NAND2_X1 U11649 ( .A1(n11417), .A2(n11419), .ZN(n11414) );
  AND2_X1 U11650 ( .A1(n11268), .A2(n21691), .ZN(n10498) );
  NOR2_X1 U11651 ( .A1(n10353), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10352) );
  INV_X1 U11652 ( .A(n10354), .ZN(n10353) );
  NAND2_X1 U11653 ( .A1(n10338), .A2(n11302), .ZN(n10342) );
  NOR2_X1 U11654 ( .A1(n15583), .A2(n10524), .ZN(n10523) );
  INV_X1 U11655 ( .A(n15601), .ZN(n10524) );
  NAND2_X1 U11656 ( .A1(n10077), .A2(n10953), .ZN(n10108) );
  CLKBUF_X1 U11657 ( .A(n16026), .Z(n16160) );
  CLKBUF_X1 U11658 ( .A(n16197), .Z(n16189) );
  OAI211_X1 U11659 ( .C1(n16247), .C2(n10238), .A(n10237), .B(n10234), .ZN(
        n16146) );
  NAND2_X1 U11660 ( .A1(n9731), .A2(n10247), .ZN(n10237) );
  AOI21_X1 U11661 ( .B1(n10243), .B2(n10242), .A(n9731), .ZN(n10238) );
  INV_X1 U11662 ( .A(n16275), .ZN(n10250) );
  INV_X1 U11663 ( .A(n13063), .ZN(n10414) );
  INV_X1 U11664 ( .A(n13759), .ZN(n12807) );
  NOR2_X1 U11665 ( .A1(n12766), .A2(n10417), .ZN(n10416) );
  INV_X1 U11666 ( .A(n13550), .ZN(n10417) );
  OR2_X1 U11667 ( .A1(n13553), .A2(n13556), .ZN(n12766) );
  INV_X1 U11668 ( .A(n9969), .ZN(n12871) );
  AND2_X1 U11669 ( .A1(n12685), .A2(n19879), .ZN(n13529) );
  INV_X1 U11670 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12996) );
  NOR2_X1 U11671 ( .A1(n12967), .A2(n10406), .ZN(n12973) );
  OR2_X1 U11672 ( .A1(n10407), .A2(n16532), .ZN(n10406) );
  NAND2_X1 U11673 ( .A1(n11175), .A2(n10517), .ZN(n10516) );
  INV_X1 U11674 ( .A(n15832), .ZN(n10517) );
  NAND3_X1 U11675 ( .A1(n10564), .A2(n10552), .A3(n10890), .ZN(n11105) );
  AND4_X1 U11676 ( .A1(n10885), .A2(n10884), .A3(n10883), .A4(n10882), .ZN(
        n10564) );
  INV_X1 U11677 ( .A(n13143), .ZN(n9971) );
  INV_X1 U11678 ( .A(n15706), .ZN(n10116) );
  NAND2_X1 U11679 ( .A1(n9819), .A2(n11387), .ZN(n10465) );
  NOR2_X1 U11680 ( .A1(n9665), .A2(n9975), .ZN(n9974) );
  INV_X1 U11681 ( .A(n14396), .ZN(n9975) );
  INV_X1 U11682 ( .A(n15724), .ZN(n10508) );
  AND2_X1 U11683 ( .A1(n10487), .A2(n10486), .ZN(n10485) );
  INV_X1 U11684 ( .A(n16539), .ZN(n10487) );
  INV_X1 U11685 ( .A(n15758), .ZN(n11201) );
  INV_X1 U11686 ( .A(n15770), .ZN(n10512) );
  NAND2_X1 U11687 ( .A1(n10443), .A2(n12895), .ZN(n10442) );
  INV_X1 U11688 ( .A(n10444), .ZN(n10443) );
  NAND2_X1 U11689 ( .A1(n13054), .A2(n12902), .ZN(n10036) );
  AND2_X1 U11690 ( .A1(n10369), .A2(n10367), .ZN(n10366) );
  AND2_X1 U11691 ( .A1(n9616), .A2(n16598), .ZN(n10367) );
  NAND2_X1 U11692 ( .A1(n16630), .A2(n16973), .ZN(n10265) );
  NAND2_X1 U11693 ( .A1(n9942), .A2(n11098), .ZN(n11324) );
  NAND2_X1 U11694 ( .A1(n9927), .A2(n11111), .ZN(n9781) );
  OR2_X1 U11695 ( .A1(n11317), .A2(n17338), .ZN(n11119) );
  XNOR2_X1 U11696 ( .A(n11322), .B(n11323), .ZN(n11317) );
  OAI21_X1 U11697 ( .B1(n11323), .B2(n10559), .A(n11286), .ZN(n11287) );
  NAND2_X1 U11698 ( .A1(n11323), .A2(n11285), .ZN(n11286) );
  OR2_X1 U11699 ( .A1(n11323), .A2(n11285), .ZN(n10080) );
  NAND2_X1 U11700 ( .A1(n11323), .A2(n10559), .ZN(n10079) );
  NAND2_X1 U11701 ( .A1(n10951), .A2(n10132), .ZN(n11151) );
  NOR2_X1 U11702 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  NOR2_X1 U11703 ( .A1(n11229), .A2(n11251), .ZN(n10133) );
  OAI21_X1 U11704 ( .B1(n12733), .B2(n20429), .A(n12698), .ZN(n12706) );
  NOR2_X1 U11705 ( .A1(n9595), .A2(n21601), .ZN(n13743) );
  NOR2_X1 U11706 ( .A1(n9595), .A2(n13740), .ZN(n13741) );
  CLKBUF_X1 U11707 ( .A(n14106), .Z(n16201) );
  NAND2_X1 U11708 ( .A1(n10440), .A2(n10439), .ZN(n12652) );
  NAND2_X1 U11709 ( .A1(n20559), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10439) );
  NAND2_X1 U11710 ( .A1(n9910), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U11711 ( .A1(n9911), .A2(n12646), .ZN(n9910) );
  NOR2_X1 U11712 ( .A1(n20169), .A2(n20494), .ZN(n20230) );
  AOI22_X1 U11713 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10834) );
  AND2_X1 U11714 ( .A1(n12659), .A2(n9711), .ZN(n13332) );
  AND2_X1 U11715 ( .A1(n19524), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10598) );
  AND2_X1 U11716 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U11717 ( .A1(n18700), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10588) );
  NAND2_X1 U11718 ( .A1(n10025), .A2(n10024), .ZN(n14163) );
  NAND2_X1 U11719 ( .A1(n18797), .A2(n13957), .ZN(n13964) );
  AND2_X1 U11720 ( .A1(n10744), .A2(n10743), .ZN(n13618) );
  NOR2_X1 U11721 ( .A1(n13317), .A2(n13179), .ZN(n13310) );
  INV_X1 U11722 ( .A(n13772), .ZN(n21584) );
  NAND2_X1 U11723 ( .A1(n11952), .A2(n11951), .ZN(n10432) );
  AND2_X1 U11724 ( .A1(n21503), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14497) );
  INV_X1 U11725 ( .A(n14618), .ZN(n10076) );
  INV_X1 U11726 ( .A(n14619), .ZN(n10075) );
  AND2_X1 U11727 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12329) );
  AND2_X1 U11728 ( .A1(n10074), .A2(n14876), .ZN(n10073) );
  NOR2_X1 U11729 ( .A1(n12187), .A2(n14100), .ZN(n10074) );
  AND2_X1 U11730 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12153), .ZN(
        n12163) );
  INV_X1 U11731 ( .A(n9853), .ZN(n9851) );
  NAND2_X1 U11732 ( .A1(n14605), .A2(n9752), .ZN(n14510) );
  INV_X1 U11733 ( .A(n14508), .ZN(n10436) );
  OAI21_X1 U11734 ( .B1(n15046), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15220), .ZN(n10127) );
  OAI211_X1 U11735 ( .C1(n14530), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12037), .B(
        n12072), .ZN(n12039) );
  NOR2_X1 U11736 ( .A1(n15104), .A2(n11842), .ZN(n15117) );
  OR2_X1 U11737 ( .A1(n9683), .A2(n15239), .ZN(n9964) );
  AND2_X1 U11738 ( .A1(n9596), .A2(n9764), .ZN(n10387) );
  NAND2_X1 U11739 ( .A1(n15117), .A2(n10453), .ZN(n9965) );
  NAND2_X1 U11740 ( .A1(n15220), .A2(n12088), .ZN(n15155) );
  INV_X1 U11741 ( .A(n15155), .ZN(n10162) );
  NAND2_X1 U11742 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U11743 ( .A1(n15239), .A2(n15469), .ZN(n15202) );
  OR2_X1 U11744 ( .A1(n10177), .A2(n9672), .ZN(n10174) );
  NAND2_X1 U11745 ( .A1(n15249), .A2(n10176), .ZN(n10175) );
  NOR2_X1 U11746 ( .A1(n10049), .A2(n9672), .ZN(n10176) );
  AND2_X1 U11747 ( .A1(n9674), .A2(n10425), .ZN(n10424) );
  INV_X1 U11748 ( .A(n14925), .ZN(n10425) );
  INV_X1 U11749 ( .A(n10158), .ZN(n10157) );
  OR2_X1 U11750 ( .A1(n14000), .A2(n14035), .ZN(n14189) );
  OR2_X1 U11751 ( .A1(n12092), .A2(n15397), .ZN(n15460) );
  INV_X1 U11752 ( .A(n11595), .ZN(n11940) );
  CLKBUF_X1 U11753 ( .A(n12061), .Z(n13428) );
  AND2_X1 U11754 ( .A1(n11937), .A2(n13463), .ZN(n12091) );
  INV_X1 U11755 ( .A(n11593), .ZN(n9831) );
  NAND2_X1 U11756 ( .A1(n13577), .A2(n21501), .ZN(n10283) );
  INV_X1 U11757 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21275) );
  NOR2_X1 U11758 ( .A1(n12132), .A2(n20799), .ZN(n20933) );
  NAND2_X1 U11759 ( .A1(n20799), .A2(n15555), .ZN(n21088) );
  INV_X1 U11760 ( .A(n11743), .ZN(n15555) );
  AND2_X1 U11761 ( .A1(n20803), .A2(n21286), .ZN(n21200) );
  INV_X1 U11762 ( .A(n21087), .ZN(n21232) );
  NOR2_X1 U11763 ( .A1(n21279), .A2(n10062), .ZN(n21425) );
  NOR2_X1 U11764 ( .A1(n20975), .A2(n21121), .ZN(n21378) );
  AND4_X1 U11765 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11547) );
  AND4_X1 U11766 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11525) );
  AND4_X1 U11767 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11527) );
  AND4_X1 U11768 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11526) );
  NAND2_X1 U11769 ( .A1(n20799), .A2(n11743), .ZN(n21372) );
  OAI221_X1 U11770 ( .B1(n14227), .B2(n15575), .C1(n17321), .C2(n15575), .A(
        n21501), .ZN(n20975) );
  AOI21_X1 U11771 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21327), .A(n20975), 
        .ZN(n21439) );
  NAND2_X2 U11772 ( .A1(n11923), .A2(n11922), .ZN(n17305) );
  NAND2_X1 U11773 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  NAND2_X1 U11774 ( .A1(n11918), .A2(n11917), .ZN(n11923) );
  INV_X1 U11775 ( .A(n11919), .ZN(n11920) );
  INV_X1 U11776 ( .A(n21590), .ZN(n17309) );
  OR2_X1 U11777 ( .A1(n13030), .A2(n20550), .ZN(n13100) );
  OR2_X1 U11778 ( .A1(n12649), .A2(n10793), .ZN(n14374) );
  NOR2_X1 U11779 ( .A1(n10349), .A2(n10351), .ZN(n10347) );
  INV_X1 U11780 ( .A(n10498), .ZN(n10351) );
  NOR2_X1 U11781 ( .A1(n10355), .A2(n11351), .ZN(n10354) );
  INV_X1 U11782 ( .A(n10492), .ZN(n10355) );
  NOR2_X1 U11783 ( .A1(n10344), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10343) );
  INV_X1 U11784 ( .A(n10345), .ZN(n10344) );
  OR2_X1 U11785 ( .A1(n11257), .A2(n12689), .ZN(n11419) );
  INV_X1 U11786 ( .A(n14374), .ZN(n13330) );
  AND2_X1 U11787 ( .A1(n10523), .A2(n10521), .ZN(n10520) );
  NOR2_X1 U11788 ( .A1(n10525), .A2(n10522), .ZN(n10521) );
  INV_X1 U11789 ( .A(n12927), .ZN(n10525) );
  INV_X1 U11790 ( .A(n15615), .ZN(n10522) );
  OR2_X1 U11791 ( .A1(n12788), .A2(n12787), .ZN(n14085) );
  NOR2_X1 U11792 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10423) );
  NOR2_X1 U11793 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10422) );
  NOR2_X1 U11794 ( .A1(n15617), .A2(n10419), .ZN(n13094) );
  NAND2_X1 U11795 ( .A1(n10421), .A2(n10420), .ZN(n10419) );
  NOR2_X1 U11796 ( .A1(n15618), .A2(n13096), .ZN(n10420) );
  INV_X1 U11797 ( .A(n15618), .ZN(n10418) );
  NAND2_X1 U11798 ( .A1(n16254), .A2(n16058), .ZN(n16248) );
  OR2_X1 U11799 ( .A1(n16263), .A2(n16057), .ZN(n16058) );
  XNOR2_X1 U11800 ( .A(n16263), .B(n16078), .ZN(n16256) );
  NAND2_X1 U11801 ( .A1(n16256), .A2(n16255), .ZN(n16254) );
  OR2_X1 U11802 ( .A1(n9663), .A2(n12731), .ZN(n12732) );
  NAND2_X1 U11803 ( .A1(n14370), .A2(n20549), .ZN(n13490) );
  AOI21_X1 U11804 ( .B1(n13109), .B2(n16690), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13078) );
  NAND2_X1 U11805 ( .A1(n16429), .A2(n16431), .ZN(n13088) );
  XNOR2_X1 U11806 ( .A(n13077), .B(n13081), .ZN(n13085) );
  NAND2_X1 U11807 ( .A1(n13079), .A2(n16430), .ZN(n13086) );
  NAND2_X1 U11808 ( .A1(n9675), .A2(n15601), .ZN(n15600) );
  NOR2_X1 U11809 ( .A1(n12967), .A2(n10409), .ZN(n12971) );
  NOR2_X1 U11810 ( .A1(n14291), .A2(n14290), .ZN(n15856) );
  NOR2_X1 U11811 ( .A1(n10111), .A2(n16753), .ZN(n16724) );
  AND2_X1 U11812 ( .A1(n11267), .A2(n11422), .ZN(n16462) );
  AND2_X1 U11813 ( .A1(n10526), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10257) );
  NOR2_X1 U11814 ( .A1(n14395), .A2(n9631), .ZN(n15739) );
  NAND2_X1 U11815 ( .A1(n16557), .A2(n12896), .ZN(n16527) );
  AOI21_X1 U11816 ( .B1(n16858), .B2(n17348), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9866) );
  AND2_X1 U11817 ( .A1(n10503), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U11818 ( .A1(n16609), .A2(n10464), .ZN(n9785) );
  NAND2_X1 U11819 ( .A1(n16609), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9789) );
  NAND2_X1 U11820 ( .A1(n16654), .A2(n11142), .ZN(n10461) );
  AND2_X1 U11821 ( .A1(n11145), .A2(n11146), .ZN(n16644) );
  INV_X1 U11822 ( .A(n16654), .ZN(n10200) );
  INV_X1 U11823 ( .A(n10461), .ZN(n10458) );
  INV_X1 U11824 ( .A(n16644), .ZN(n10457) );
  NAND2_X1 U11825 ( .A1(n16666), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16667) );
  NAND2_X1 U11826 ( .A1(n16702), .A2(n11117), .ZN(n16675) );
  NAND2_X1 U11827 ( .A1(n9797), .A2(n16703), .ZN(n16702) );
  CLKBUF_X1 U11828 ( .A(n12679), .Z(n12680) );
  OR2_X1 U11829 ( .A1(n9663), .A2(n12690), .ZN(n12692) );
  OR2_X1 U11830 ( .A1(n9623), .A2(n19745), .ZN(n13478) );
  OR2_X1 U11831 ( .A1(n20508), .A2(n20517), .ZN(n20168) );
  OR2_X1 U11832 ( .A1(n13455), .A2(n13454), .ZN(n13745) );
  OR2_X1 U11833 ( .A1(n13742), .A2(n13741), .ZN(n10229) );
  AND2_X1 U11834 ( .A1(n20358), .A2(n19948), .ZN(n19846) );
  INV_X1 U11835 ( .A(n11053), .ZN(n19841) );
  INV_X1 U11836 ( .A(n20543), .ZN(n19948) );
  AND2_X1 U11837 ( .A1(n19839), .A2(n20508), .ZN(n17045) );
  AND2_X1 U11838 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20199) );
  AND2_X2 U11839 ( .A1(n14022), .A2(n10980), .ZN(n11060) );
  AND3_X1 U11840 ( .A1(n20169), .A2(n20508), .A3(n20494), .ZN(n20492) );
  NOR2_X1 U11842 ( .A1(n20169), .A2(n20168), .ZN(n20209) );
  AND2_X1 U11843 ( .A1(n20230), .A2(n20508), .ZN(n20270) );
  NAND2_X1 U11844 ( .A1(n9931), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9930) );
  NAND2_X1 U11845 ( .A1(n9929), .A2(n14341), .ZN(n9928) );
  AND2_X1 U11846 ( .A1(n19844), .A2(n20508), .ZN(n20354) );
  NAND2_X1 U11847 ( .A1(n17016), .A2(n20559), .ZN(n17018) );
  INV_X1 U11848 ( .A(n20361), .ZN(n20265) );
  OR2_X1 U11849 ( .A1(n20349), .A2(n20348), .ZN(n20360) );
  NAND2_X1 U11850 ( .A1(n13836), .A2(n13835), .ZN(n19516) );
  NOR2_X1 U11851 ( .A1(n17472), .A2(n17471), .ZN(n17470) );
  NAND2_X1 U11852 ( .A1(n10768), .A2(n17774), .ZN(n17468) );
  NOR2_X1 U11853 ( .A1(n18524), .A2(n17504), .ZN(n17505) );
  NOR2_X1 U11854 ( .A1(n10301), .A2(n10589), .ZN(n17613) );
  XNOR2_X1 U11855 ( .A(n10585), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10590) );
  AND2_X1 U11856 ( .A1(n9619), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10309) );
  NOR2_X1 U11857 ( .A1(n18575), .A2(n10298), .ZN(n10297) );
  NAND2_X1 U11858 ( .A1(n10305), .A2(n9638), .ZN(n18609) );
  NAND2_X1 U11859 ( .A1(n9880), .A2(n18734), .ZN(n14179) );
  NAND2_X1 U11860 ( .A1(n18733), .A2(n9879), .ZN(n9880) );
  NOR2_X1 U11861 ( .A1(n14180), .A2(n19015), .ZN(n9879) );
  INV_X1 U11862 ( .A(n18807), .ZN(n18776) );
  OAI211_X1 U11863 ( .C1(n10383), .C2(n10019), .A(n9621), .B(n10017), .ZN(
        n10016) );
  NOR2_X1 U11864 ( .A1(n10383), .A2(n14442), .ZN(n14444) );
  AND2_X1 U11865 ( .A1(n14433), .A2(n10382), .ZN(n10381) );
  NAND2_X1 U11866 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U11867 ( .A1(n18642), .A2(n14428), .ZN(n14429) );
  NAND2_X1 U11868 ( .A1(n18644), .A2(n14427), .ZN(n14428) );
  NAND2_X1 U11869 ( .A1(n13974), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14125) );
  NAND2_X1 U11870 ( .A1(n9884), .A2(n18771), .ZN(n13946) );
  INV_X1 U11871 ( .A(n13937), .ZN(n13943) );
  NAND2_X1 U11872 ( .A1(n10730), .A2(n19681), .ZN(n10364) );
  OR2_X1 U11873 ( .A1(n19514), .A2(n14474), .ZN(n14475) );
  INV_X1 U11874 ( .A(n20662), .ZN(n14927) );
  AND2_X1 U11875 ( .A1(n20662), .A2(n14545), .ZN(n20658) );
  INV_X1 U11876 ( .A(n20786), .ZN(n20731) );
  AND2_X2 U11877 ( .A1(n20574), .A2(n12623), .ZN(n20732) );
  INV_X1 U11878 ( .A(n20732), .ZN(n15169) );
  NAND2_X1 U11879 ( .A1(n12621), .A2(n9585), .ZN(n20797) );
  XNOR2_X1 U11880 ( .A(n9823), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12631) );
  NAND2_X1 U11881 ( .A1(n9824), .A2(n9698), .ZN(n9823) );
  INV_X1 U11882 ( .A(n14492), .ZN(n9824) );
  XNOR2_X1 U11883 ( .A(n10051), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15045) );
  NAND2_X1 U11884 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  NAND2_X1 U11885 ( .A1(n11852), .A2(n10050), .ZN(n10053) );
  INV_X1 U11886 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21327) );
  NOR2_X1 U11887 ( .A1(n20799), .A2(n10129), .ZN(n21233) );
  INV_X1 U11888 ( .A(n12132), .ZN(n10129) );
  NAND2_X1 U11889 ( .A1(n20933), .A2(n21232), .ZN(n20978) );
  OR2_X1 U11890 ( .A1(n17301), .A2(n21501), .ZN(n20568) );
  OAI21_X1 U11891 ( .B1(n13112), .B2(n13111), .A(n13110), .ZN(n13113) );
  XNOR2_X1 U11892 ( .A(n11427), .B(n11430), .ZN(n15594) );
  INV_X1 U11893 ( .A(n15954), .ZN(n19760) );
  NAND2_X1 U11894 ( .A1(n13007), .A2(n13006), .ZN(n19734) );
  NAND2_X1 U11895 ( .A1(n19748), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19767) );
  XNOR2_X1 U11896 ( .A(n15587), .B(n12927), .ZN(n16211) );
  OR2_X1 U11897 ( .A1(n9675), .A2(n15616), .ZN(n16748) );
  OR2_X1 U11898 ( .A1(n16287), .A2(n12699), .ZN(n16301) );
  XNOR2_X1 U11899 ( .A(n16426), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13130) );
  XNOR2_X1 U11900 ( .A(n10192), .B(n16508), .ZN(n16820) );
  AOI21_X1 U11901 ( .B1(n16505), .B2(n16504), .A(n16503), .ZN(n10192) );
  AND2_X1 U11902 ( .A1(n9784), .A2(n9785), .ZN(n16907) );
  INV_X1 U11903 ( .A(n16722), .ZN(n16704) );
  INV_X1 U11904 ( .A(n16697), .ZN(n16717) );
  NAND2_X1 U11905 ( .A1(n19708), .A2(n11239), .ZN(n16700) );
  INV_X1 U11906 ( .A(n16700), .ZN(n16714) );
  NAND2_X1 U11907 ( .A1(n10897), .A2(n16235), .ZN(n16722) );
  NAND3_X1 U11908 ( .A1(n10087), .A2(n10085), .A3(n10082), .ZN(n13132) );
  OAI21_X1 U11909 ( .B1(n11434), .B2(n10084), .A(n10083), .ZN(n10082) );
  OR2_X1 U11910 ( .A1(n16429), .A2(n10088), .ZN(n10087) );
  NAND2_X1 U11911 ( .A1(n16737), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10185) );
  NOR2_X1 U11912 ( .A1(n10184), .A2(n16730), .ZN(n10123) );
  AOI21_X1 U11913 ( .B1(n9979), .B2(n17346), .A(n9978), .ZN(n9977) );
  OR2_X1 U11914 ( .A1(n16735), .A2(n16736), .ZN(n9978) );
  XNOR2_X1 U11915 ( .A(n16427), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16740) );
  NAND2_X1 U11916 ( .A1(n16443), .A2(n10275), .ZN(n10273) );
  OAI21_X1 U11917 ( .B1(n16443), .B2(n10274), .A(n10270), .ZN(n10269) );
  OAI21_X1 U11918 ( .B1(n16748), .B2(n17330), .A(n9924), .ZN(n9923) );
  NOR2_X1 U11919 ( .A1(n9925), .A2(n16743), .ZN(n9924) );
  INV_X1 U11920 ( .A(n16744), .ZN(n9925) );
  INV_X1 U11921 ( .A(n17340), .ZN(n17327) );
  AND2_X1 U11922 ( .A1(n16759), .A2(n13122), .ZN(n16746) );
  XNOR2_X1 U11923 ( .A(n16441), .B(n9808), .ZN(n16751) );
  XNOR2_X1 U11924 ( .A(n16440), .B(n16745), .ZN(n9808) );
  NOR2_X1 U11925 ( .A1(n16452), .A2(n9811), .ZN(n16749) );
  AND2_X1 U11926 ( .A1(n16457), .A2(n16745), .ZN(n9811) );
  XNOR2_X1 U11927 ( .A(n16476), .B(n16475), .ZN(n16778) );
  NAND2_X1 U11928 ( .A1(n10014), .A2(n16511), .ZN(n16816) );
  NAND2_X1 U11929 ( .A1(n10258), .A2(n16809), .ZN(n10014) );
  NOR2_X1 U11930 ( .A1(n16817), .A2(n10013), .ZN(n10012) );
  AND2_X1 U11931 ( .A1(n16818), .A2(n17346), .ZN(n10013) );
  OAI21_X1 U11932 ( .B1(n16513), .B2(n16514), .A(n16530), .ZN(n16518) );
  NAND2_X1 U11933 ( .A1(n16527), .A2(n16825), .ZN(n9862) );
  NAND2_X1 U11934 ( .A1(n16557), .A2(n9653), .ZN(n16830) );
  XNOR2_X1 U11935 ( .A(n16513), .B(n16531), .ZN(n16842) );
  NAND2_X1 U11936 ( .A1(n10488), .A2(n10486), .ZN(n16538) );
  NAND2_X1 U11937 ( .A1(n10480), .A2(n10489), .ZN(n10488) );
  AOI21_X1 U11938 ( .B1(n16849), .B2(n10009), .A(n16861), .ZN(n10008) );
  NOR2_X1 U11939 ( .A1(n16845), .A2(n10197), .ZN(n10009) );
  AOI21_X1 U11940 ( .B1(n16858), .B2(n17348), .A(n9777), .ZN(n10006) );
  NAND2_X1 U11941 ( .A1(n10007), .A2(n16849), .ZN(n16867) );
  NAND2_X1 U11942 ( .A1(n16846), .A2(n16845), .ZN(n10007) );
  AOI21_X1 U11943 ( .B1(n10480), .B2(n10490), .A(n12905), .ZN(n16547) );
  AND2_X1 U11944 ( .A1(n10370), .A2(n9864), .ZN(n9863) );
  NAND2_X1 U11945 ( .A1(n9866), .A2(n9867), .ZN(n9864) );
  NOR2_X1 U11946 ( .A1(n10372), .A2(n10371), .ZN(n10370) );
  INV_X1 U11947 ( .A(n16865), .ZN(n10371) );
  AND2_X1 U11948 ( .A1(n16899), .A2(n12882), .ZN(n16873) );
  NAND2_X1 U11949 ( .A1(n9938), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10462) );
  INV_X1 U11950 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16914) );
  AND2_X1 U11951 ( .A1(n10368), .A2(n11347), .ZN(n16600) );
  NAND2_X1 U11952 ( .A1(n9917), .A2(n9915), .ZN(n17337) );
  AND2_X1 U11953 ( .A1(n16850), .A2(n9759), .ZN(n9915) );
  AND2_X2 U11954 ( .A1(n10978), .A2(n10960), .ZN(n15946) );
  INV_X1 U11955 ( .A(n10259), .ZN(n10959) );
  INV_X1 U11956 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20521) );
  INV_X1 U11957 ( .A(n20494), .ZN(n20517) );
  INV_X1 U11958 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20512) );
  INV_X1 U11959 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20505) );
  OAI21_X1 U11960 ( .B1(n13425), .B2(n13735), .A(n13420), .ZN(n16993) );
  NOR2_X1 U11961 ( .A1(n20543), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13419) );
  NAND2_X1 U11962 ( .A1(n19559), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17445) );
  NOR2_X2 U11963 ( .A1(n19660), .A2(n17785), .ZN(n17716) );
  INV_X1 U11964 ( .A(n17716), .ZN(n17801) );
  NOR2_X2 U11965 ( .A1(n10763), .A2(n10761), .ZN(n17800) );
  NAND2_X1 U11966 ( .A1(n17966), .A2(n9776), .ZN(n17951) );
  NAND2_X1 U11967 ( .A1(n17951), .A2(n18266), .ZN(n17955) );
  INV_X1 U11968 ( .A(n17961), .ZN(n17966) );
  NOR2_X1 U11969 ( .A1(n10320), .A2(n18038), .ZN(n10318) );
  NOR2_X1 U11970 ( .A1(n17610), .A2(n18110), .ZN(n18073) );
  AND2_X1 U11971 ( .A1(n18272), .A2(n10312), .ZN(n18247) );
  AND2_X1 U11972 ( .A1(n18244), .A2(n9760), .ZN(n10312) );
  NOR2_X1 U11973 ( .A1(n18390), .A2(n18274), .ZN(n18275) );
  NOR2_X1 U11974 ( .A1(n18732), .A2(n18878), .ZN(n10207) );
  INV_X1 U11975 ( .A(n18579), .ZN(n10208) );
  NAND2_X1 U11976 ( .A1(n10210), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10209) );
  INV_X1 U11977 ( .A(n18587), .ZN(n10210) );
  OR2_X1 U11978 ( .A1(n18801), .A2(n18394), .ZN(n18732) );
  NAND2_X1 U11979 ( .A1(n9875), .A2(n9872), .ZN(n18910) );
  AOI21_X1 U11980 ( .B1(n18989), .B2(n18628), .A(n9873), .ZN(n9872) );
  INV_X1 U11981 ( .A(n18921), .ZN(n9875) );
  OAI21_X1 U11982 ( .B1(n17248), .B2(n19062), .A(n9874), .ZN(n9873) );
  NAND2_X1 U11983 ( .A1(n17022), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n9799) );
  INV_X1 U11984 ( .A(n12636), .ZN(n10181) );
  OR2_X1 U11985 ( .A1(n11696), .A2(n11695), .ZN(n11700) );
  INV_X1 U11986 ( .A(n10054), .ZN(n11556) );
  INV_X1 U11987 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9833) );
  AND4_X1 U11988 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n11139) );
  NAND2_X1 U11989 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n9990) );
  NAND2_X1 U11990 ( .A1(n11052), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n9987) );
  NAND2_X1 U11991 ( .A1(n11053), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n9984) );
  NAND2_X1 U11992 ( .A1(n11051), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n9985) );
  AOI22_X1 U11993 ( .A1(n11053), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n20234), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U11994 ( .A1(n9813), .A2(n14022), .ZN(n9812) );
  NOR2_X1 U11995 ( .A1(n10963), .A2(n9814), .ZN(n9813) );
  AND2_X1 U11996 ( .A1(n10739), .A2(n10738), .ZN(n10740) );
  AOI22_X1 U11997 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11470) );
  BUF_X1 U11998 ( .A(n12595), .Z(n12497) );
  CLKBUF_X3 U11999 ( .A(n11613), .Z(n12577) );
  AND2_X1 U12001 ( .A1(n11732), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10285) );
  INV_X1 U12002 ( .A(n11837), .ZN(n9956) );
  XNOR2_X1 U12003 ( .A(n11814), .B(n11813), .ZN(n12188) );
  AND2_X1 U12004 ( .A1(n11770), .A2(n11786), .ZN(n10390) );
  OAI211_X1 U12005 ( .C1(n11734), .C2(n10044), .A(n10041), .B(n10039), .ZN(
        n12162) );
  INV_X1 U12006 ( .A(n11786), .ZN(n10044) );
  NAND2_X1 U12007 ( .A1(n10040), .A2(n11786), .ZN(n10039) );
  NOR2_X1 U12008 ( .A1(n11569), .A2(n21501), .ZN(n10155) );
  AND3_X1 U12009 ( .A1(n9821), .A2(n11555), .A3(n11595), .ZN(n10054) );
  INV_X1 U12010 ( .A(n12068), .ZN(n9821) );
  AOI22_X1 U12011 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11502) );
  BUF_X2 U12012 ( .A(n11467), .Z(n11601) );
  AOI22_X1 U12013 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U12014 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U12015 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U12016 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U12017 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n12578), .ZN(n11462) );
  INV_X1 U12018 ( .A(n11891), .ZN(n11910) );
  NAND2_X1 U12019 ( .A1(n11891), .A2(n11928), .ZN(n11916) );
  AOI22_X1 U12020 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U12021 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10878) );
  NOR2_X1 U12022 ( .A1(n10240), .A2(n10236), .ZN(n10235) );
  INV_X1 U12023 ( .A(n10242), .ZN(n10236) );
  NOR2_X1 U12024 ( .A1(n10245), .A2(n10241), .ZN(n10240) );
  NAND2_X1 U12025 ( .A1(n10246), .A2(n10248), .ZN(n10243) );
  INV_X1 U12026 ( .A(n16236), .ZN(n10249) );
  INV_X1 U12027 ( .A(n16492), .ZN(n10090) );
  INV_X1 U12028 ( .A(n10485), .ZN(n10484) );
  OR2_X1 U12029 ( .A1(n15767), .A2(n11143), .ZN(n11401) );
  NOR2_X1 U12030 ( .A1(n16690), .A2(n10030), .ZN(n10029) );
  INV_X1 U12031 ( .A(n11098), .ZN(n10030) );
  NAND2_X1 U12032 ( .A1(n11003), .A2(n16235), .ZN(n9935) );
  OAI21_X1 U12033 ( .B1(n11221), .B2(n10136), .A(n10135), .ZN(n10134) );
  NAND2_X1 U12034 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10135) );
  NOR2_X1 U12035 ( .A1(n9997), .A2(n9994), .ZN(n10936) );
  NAND2_X1 U12036 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NOR2_X1 U12037 ( .A1(n13038), .A2(n11249), .ZN(n9995) );
  NAND2_X1 U12038 ( .A1(n9705), .A2(n9640), .ZN(n10940) );
  NOR2_X1 U12039 ( .A1(n11246), .A2(n19875), .ZN(n10917) );
  AND2_X1 U12040 ( .A1(n12655), .A2(n10916), .ZN(n12869) );
  NAND2_X1 U12041 ( .A1(n9912), .A2(n9691), .ZN(n9911) );
  OAI21_X1 U12042 ( .B1(n10446), .B2(n9692), .A(n9913), .ZN(n9912) );
  INV_X1 U12043 ( .A(n12642), .ZN(n9913) );
  AND3_X1 U12044 ( .A1(n10812), .A2(n10811), .A3(n14341), .ZN(n10813) );
  NAND2_X1 U12045 ( .A1(n14106), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10812) );
  AND2_X1 U12046 ( .A1(n20295), .A2(n20260), .ZN(n17013) );
  NAND2_X1 U12047 ( .A1(n13329), .A2(n12663), .ZN(n10190) );
  AND2_X1 U12048 ( .A1(n10188), .A2(n12876), .ZN(n10187) );
  INV_X1 U12049 ( .A(n10189), .ZN(n10188) );
  OAI21_X1 U12050 ( .B1(n12657), .B2(n12647), .A(n9801), .ZN(n10189) );
  INV_X1 U12051 ( .A(n9996), .ZN(n9801) );
  INV_X1 U12052 ( .A(n18747), .ZN(n10375) );
  AND2_X1 U12053 ( .A1(n17752), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10742) );
  INV_X1 U12054 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12528) );
  NOR2_X1 U12055 ( .A1(n10535), .A2(n10536), .ZN(n10534) );
  INV_X1 U12056 ( .A(n14691), .ZN(n10535) );
  INV_X1 U12057 ( .A(n12590), .ZN(n12616) );
  AND2_X1 U12058 ( .A1(n12314), .A2(n10529), .ZN(n10528) );
  NOR2_X1 U12059 ( .A1(n14590), .A2(n10438), .ZN(n10437) );
  INV_X1 U12060 ( .A(n14606), .ZN(n10438) );
  INV_X1 U12061 ( .A(n11848), .ZN(n9827) );
  NOR2_X1 U12062 ( .A1(n10453), .A2(n10455), .ZN(n10452) );
  AND2_X1 U12063 ( .A1(n15067), .A2(n9765), .ZN(n9829) );
  INV_X1 U12064 ( .A(n14733), .ZN(n10429) );
  AND2_X1 U12065 ( .A1(n12001), .A2(n12000), .ZN(n14804) );
  NAND2_X1 U12066 ( .A1(n15239), .A2(n11835), .ZN(n15200) );
  INV_X1 U12067 ( .A(n11833), .ZN(n10178) );
  OR2_X1 U12068 ( .A1(n11804), .A2(n11803), .ZN(n11815) );
  INV_X1 U12069 ( .A(n11742), .ZN(n10451) );
  AND3_X1 U12070 ( .A1(n11660), .A2(n11659), .A3(n11658), .ZN(n11662) );
  AND2_X1 U12071 ( .A1(n11713), .A2(n20809), .ZN(n11683) );
  NAND2_X1 U12072 ( .A1(n11550), .A2(n10046), .ZN(n13580) );
  NOR2_X1 U12073 ( .A1(n11930), .A2(n14545), .ZN(n10046) );
  AND2_X2 U12074 ( .A1(n11673), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13590) );
  NAND2_X1 U12075 ( .A1(n10061), .A2(n20967), .ZN(n10060) );
  NAND2_X1 U12076 ( .A1(n13680), .A2(n9636), .ZN(n10059) );
  AOI22_X1 U12077 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11492) );
  AND2_X2 U12078 ( .A1(n13594), .A2(n15563), .ZN(n11610) );
  INV_X1 U12079 ( .A(n9587), .ZN(n20800) );
  NAND2_X1 U12080 ( .A1(n11862), .A2(n11861), .ZN(n11919) );
  OR2_X1 U12081 ( .A1(n11916), .A2(n11919), .ZN(n11917) );
  INV_X1 U12082 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14056) );
  XNOR2_X1 U12083 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10894) );
  AND2_X1 U12084 ( .A1(n10786), .A2(n10785), .ZN(n12644) );
  INV_X1 U12085 ( .A(n13038), .ZN(n12645) );
  NOR2_X1 U12086 ( .A1(n10346), .A2(n11260), .ZN(n10345) );
  INV_X1 U12087 ( .A(n10495), .ZN(n10346) );
  NOR2_X1 U12088 ( .A1(n11381), .A2(n10496), .ZN(n10495) );
  AND2_X1 U12089 ( .A1(n11302), .A2(n11335), .ZN(n10337) );
  INV_X1 U12090 ( .A(n14019), .ZN(n10232) );
  NAND2_X1 U12091 ( .A1(n10938), .A2(n9968), .ZN(n9787) );
  INV_X1 U12092 ( .A(n13038), .ZN(n9800) );
  NAND2_X1 U12093 ( .A1(n14010), .A2(n14011), .ZN(n10233) );
  AND2_X1 U12094 ( .A1(n15603), .A2(n15591), .ZN(n10421) );
  AND2_X1 U12095 ( .A1(n15982), .A2(n14096), .ZN(n10396) );
  NOR2_X1 U12096 ( .A1(n15981), .A2(n15980), .ZN(n15982) );
  AND2_X1 U12097 ( .A1(n14417), .A2(n15741), .ZN(n10415) );
  NAND2_X2 U12098 ( .A1(n10898), .A2(n11246), .ZN(n12655) );
  INV_X1 U12099 ( .A(n19875), .ZN(n10898) );
  NOR2_X1 U12100 ( .A1(n12980), .A2(n10412), .ZN(n10411) );
  INV_X1 U12101 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U12102 ( .A1(n10408), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10407) );
  INV_X1 U12103 ( .A(n10409), .ZN(n10408) );
  NAND2_X1 U12104 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10409) );
  NOR2_X1 U12105 ( .A1(n16619), .A2(n10402), .ZN(n10401) );
  INV_X1 U12106 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10402) );
  AND2_X1 U12107 ( .A1(n13288), .A2(n12701), .ZN(n11104) );
  OR2_X1 U12108 ( .A1(n12701), .A2(n12689), .ZN(n11250) );
  INV_X1 U12109 ( .A(n16430), .ZN(n10089) );
  OAI21_X1 U12110 ( .B1(n10472), .B2(n10471), .A(n10473), .ZN(n10470) );
  INV_X1 U12111 ( .A(n16442), .ZN(n10473) );
  INV_X1 U12112 ( .A(n10470), .ZN(n10469) );
  AND2_X1 U12113 ( .A1(n11413), .A2(n16462), .ZN(n10474) );
  INV_X1 U12114 ( .A(n15657), .ZN(n10518) );
  AND2_X1 U12115 ( .A1(n15687), .A2(n15675), .ZN(n10519) );
  AND2_X1 U12116 ( .A1(n15665), .A2(n16690), .ZN(n11276) );
  NOR2_X1 U12117 ( .A1(n12897), .A2(n13117), .ZN(n10110) );
  AND2_X1 U12118 ( .A1(n15684), .A2(n16690), .ZN(n16471) );
  OR2_X1 U12119 ( .A1(n15701), .A2(n11143), .ZN(n11411) );
  INV_X1 U12120 ( .A(n11409), .ZN(n11410) );
  OAI21_X1 U12121 ( .B1(n11408), .B2(n11407), .A(n11406), .ZN(n11409) );
  NOR2_X1 U12122 ( .A1(n11148), .A2(n16930), .ZN(n10526) );
  AND2_X1 U12123 ( .A1(n10478), .A2(n10034), .ZN(n10033) );
  NAND2_X1 U12124 ( .A1(n10038), .A2(n10036), .ZN(n10034) );
  NOR2_X1 U12125 ( .A1(n10484), .A2(n10479), .ZN(n10478) );
  INV_X1 U12126 ( .A(n16569), .ZN(n10479) );
  INV_X1 U12127 ( .A(n10036), .ZN(n10035) );
  INV_X1 U12128 ( .A(n10489), .ZN(n10483) );
  OR2_X1 U12129 ( .A1(n11401), .A2(n16861), .ZN(n12909) );
  NOR2_X1 U12130 ( .A1(n12633), .A2(n16930), .ZN(n10503) );
  OR2_X1 U12131 ( .A1(n15823), .A2(n11143), .ZN(n12901) );
  NAND2_X1 U12132 ( .A1(n10000), .A2(n11324), .ZN(n9780) );
  NAND2_X1 U12133 ( .A1(n10095), .A2(n10094), .ZN(n10000) );
  NAND2_X1 U12134 ( .A1(n10131), .A2(n11109), .ZN(n11115) );
  OAI211_X1 U12135 ( .C1(n14334), .C2(n10938), .A(n9939), .B(n10146), .ZN(
        n10145) );
  OR2_X1 U12136 ( .A1(n11002), .A2(n11001), .ZN(n12718) );
  AND2_X1 U12137 ( .A1(n14112), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14110) );
  AND2_X1 U12138 ( .A1(n20169), .A2(n20517), .ZN(n19839) );
  AOI22_X1 U12139 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U12140 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10829) );
  NOR2_X1 U12141 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U12142 ( .A1(n17484), .A2(n17943), .ZN(n10768) );
  INV_X1 U12143 ( .A(n18590), .ZN(n10292) );
  INV_X1 U12144 ( .A(n14192), .ZN(n10316) );
  NAND2_X1 U12145 ( .A1(n10610), .A2(n13609), .ZN(n18060) );
  INV_X1 U12146 ( .A(n19127), .ZN(n13620) );
  INV_X1 U12147 ( .A(n10586), .ZN(n10305) );
  XNOR2_X1 U12148 ( .A(n14204), .B(n14198), .ZN(n13955) );
  NOR2_X1 U12149 ( .A1(n17450), .A2(n13650), .ZN(n13614) );
  XNOR2_X1 U12150 ( .A(n13939), .B(n14204), .ZN(n13936) );
  OR2_X1 U12151 ( .A1(n13936), .A2(n19073), .ZN(n13937) );
  NAND2_X1 U12152 ( .A1(n14198), .A2(n14214), .ZN(n13939) );
  NOR3_X1 U12153 ( .A1(n13624), .A2(n13832), .A3(n13658), .ZN(n14193) );
  OAI21_X1 U12154 ( .B1(n13614), .B2(n19551), .A(n13830), .ZN(n18414) );
  INV_X1 U12155 ( .A(n10625), .ZN(n9894) );
  INV_X1 U12156 ( .A(n10626), .ZN(n9891) );
  AOI21_X1 U12157 ( .B1(n13906), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9893), .ZN(n9892) );
  AOI21_X1 U12158 ( .B1(n17751), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10203), .ZN(n10681) );
  AND2_X1 U12159 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10203) );
  NOR2_X1 U12160 ( .A1(n19553), .A2(n19567), .ZN(n19094) );
  NAND2_X1 U12161 ( .A1(n10595), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17266) );
  NOR2_X1 U12162 ( .A1(n19122), .A2(n17260), .ZN(n10213) );
  OR2_X1 U12163 ( .A1(n11929), .A2(n11562), .ZN(n13317) );
  NAND2_X1 U12164 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12026) );
  OR2_X1 U12165 ( .A1(n21588), .A2(n14232), .ZN(n20594) );
  NAND2_X1 U12166 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12040) );
  AND2_X1 U12167 ( .A1(n12388), .A2(n12387), .ZN(n14701) );
  AND2_X1 U12168 ( .A1(n11989), .A2(n11988), .ZN(n14846) );
  OAI211_X1 U12169 ( .C1(n14530), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11986), .B(
        n12072), .ZN(n11989) );
  OR2_X1 U12170 ( .A1(n15009), .A2(n13189), .ZN(n13705) );
  NOR2_X1 U12171 ( .A1(n10539), .A2(n10541), .ZN(n10538) );
  NAND2_X1 U12172 ( .A1(n10540), .A2(n14604), .ZN(n10539) );
  INV_X1 U12173 ( .A(n14577), .ZN(n10540) );
  NOR2_X1 U12174 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  OR2_X1 U12175 ( .A1(n12487), .A2(n15091), .ZN(n12489) );
  OR2_X1 U12176 ( .A1(n12489), .A2(n12488), .ZN(n12529) );
  AND2_X1 U12177 ( .A1(n12440), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12441) );
  AND2_X1 U12178 ( .A1(n9673), .A2(n10071), .ZN(n10070) );
  INV_X1 U12179 ( .A(n14646), .ZN(n10071) );
  INV_X1 U12180 ( .A(n12407), .ZN(n12408) );
  OR2_X1 U12181 ( .A1(n12389), .A2(n21627), .ZN(n12407) );
  OR2_X1 U12182 ( .A1(n12366), .A2(n12365), .ZN(n12369) );
  AND2_X1 U12183 ( .A1(n12281), .A2(n12280), .ZN(n12330) );
  AND4_X1 U12184 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n14841) );
  INV_X1 U12185 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U12186 ( .A1(n12182), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12208) );
  INV_X1 U12187 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U12188 ( .A1(n12132), .A2(n11928), .ZN(n11741) );
  OR2_X1 U12189 ( .A1(n14527), .A2(n12056), .ZN(n14529) );
  INV_X1 U12190 ( .A(n15069), .ZN(n9852) );
  AND2_X1 U12191 ( .A1(n10453), .A2(n15298), .ZN(n10050) );
  INV_X1 U12192 ( .A(n15299), .ZN(n10449) );
  AND2_X1 U12193 ( .A1(n12054), .A2(n12053), .ZN(n14508) );
  NAND2_X1 U12194 ( .A1(n14605), .A2(n10437), .ZN(n14592) );
  NAND2_X1 U12195 ( .A1(n14605), .A2(n14606), .ZN(n14608) );
  AND2_X1 U12196 ( .A1(n14659), .A2(n9743), .ZN(n14641) );
  INV_X1 U12197 ( .A(n14642), .ZN(n10433) );
  NAND2_X1 U12198 ( .A1(n9849), .A2(n9848), .ZN(n12036) );
  NAND2_X1 U12199 ( .A1(n12072), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U12200 ( .A1(n14659), .A2(n10434), .ZN(n14647) );
  NAND2_X1 U12201 ( .A1(n12032), .A2(n9842), .ZN(n12034) );
  NAND2_X1 U12202 ( .A1(n14659), .A2(n14660), .ZN(n14662) );
  NAND2_X1 U12203 ( .A1(n9846), .A2(n9845), .ZN(n12023) );
  NAND2_X1 U12204 ( .A1(n12072), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U12205 ( .A1(n12025), .A2(n12024), .ZN(n14703) );
  INV_X1 U12206 ( .A(n14705), .ZN(n12024) );
  INV_X1 U12207 ( .A(n14706), .ZN(n12025) );
  NAND2_X1 U12208 ( .A1(n12018), .A2(n9840), .ZN(n12021) );
  AND2_X1 U12209 ( .A1(n12009), .A2(n9735), .ZN(n14735) );
  AND2_X1 U12210 ( .A1(n12013), .A2(n12012), .ZN(n14751) );
  NAND2_X1 U12211 ( .A1(n12010), .A2(n9838), .ZN(n12013) );
  NAND2_X1 U12212 ( .A1(n12009), .A2(n9728), .ZN(n14749) );
  AND2_X1 U12213 ( .A1(n10427), .A2(n14783), .ZN(n10426) );
  NAND2_X1 U12214 ( .A1(n11991), .A2(n11990), .ZN(n14844) );
  NOR2_X1 U12215 ( .A1(n10049), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U12216 ( .A1(n15258), .A2(n15257), .ZN(n11823) );
  AND2_X1 U12217 ( .A1(n15272), .A2(n11782), .ZN(n10159) );
  INV_X1 U12218 ( .A(n11784), .ZN(n15274) );
  INV_X1 U12219 ( .A(n14002), .ZN(n11959) );
  INV_X1 U12220 ( .A(n14001), .ZN(n11958) );
  NAND2_X1 U12221 ( .A1(n12106), .A2(n11928), .ZN(n11708) );
  NAND2_X1 U12222 ( .A1(n10392), .A2(n10167), .ZN(n10166) );
  INV_X1 U12223 ( .A(n11928), .ZN(n13725) );
  OR2_X1 U12224 ( .A1(n11939), .A2(n12065), .ZN(n13314) );
  CLKBUF_X1 U12225 ( .A(n11995), .Z(n14531) );
  NAND2_X1 U12226 ( .A1(n9844), .A2(n11933), .ZN(n12077) );
  AOI21_X1 U12227 ( .B1(n12056), .B2(n11573), .A(n12064), .ZN(n9844) );
  AND2_X1 U12228 ( .A1(n12107), .A2(n13684), .ZN(n9822) );
  NAND2_X1 U12229 ( .A1(n11644), .A2(n11643), .ZN(n11655) );
  OAI211_X1 U12230 ( .C1(n11647), .C2(n11562), .A(n11646), .B(n11645), .ZN(
        n11654) );
  AND2_X1 U12231 ( .A1(n10393), .A2(n11609), .ZN(n10391) );
  NOR2_X1 U12232 ( .A1(n13317), .A2(n13777), .ZN(n13682) );
  NAND2_X1 U12233 ( .A1(n10055), .A2(n11575), .ZN(n13581) );
  AND2_X1 U12234 ( .A1(n13572), .A2(n13571), .ZN(n17284) );
  NOR2_X1 U12235 ( .A1(n15549), .A2(n20800), .ZN(n21117) );
  AND2_X1 U12236 ( .A1(n15549), .A2(n9587), .ZN(n21194) );
  NOR2_X1 U12237 ( .A1(n15549), .A2(n9587), .ZN(n21324) );
  NAND2_X1 U12238 ( .A1(n15549), .A2(n20800), .ZN(n21087) );
  AND2_X1 U12239 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20803), .ZN(n20846) );
  OR2_X1 U12240 ( .A1(n21372), .A2(n21371), .ZN(n21381) );
  INV_X1 U12241 ( .A(n21372), .ZN(n21434) );
  NOR2_X1 U12242 ( .A1(n11872), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21580) );
  NAND2_X1 U12243 ( .A1(n13038), .A2(n12641), .ZN(n10891) );
  OR2_X1 U12244 ( .A1(n11105), .A2(n13038), .ZN(n10892) );
  AND2_X1 U12245 ( .A1(n10790), .A2(n10789), .ZN(n12649) );
  OR2_X1 U12246 ( .A1(n10788), .A2(n10787), .ZN(n10790) );
  AND2_X1 U12247 ( .A1(n17317), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10787) );
  OAI21_X1 U12248 ( .B1(n13036), .B2(n10556), .A(n13035), .ZN(n13076) );
  NAND2_X1 U12249 ( .A1(n11263), .A2(n9753), .ZN(n11417) );
  AOI21_X1 U12250 ( .B1(n19753), .B2(n15726), .A(n10398), .ZN(n10397) );
  NOR2_X1 U12251 ( .A1(n10494), .A2(n10493), .ZN(n10492) );
  INV_X1 U12252 ( .A(n11358), .ZN(n10493) );
  INV_X1 U12253 ( .A(n10563), .ZN(n10494) );
  NAND2_X1 U12254 ( .A1(n11372), .A2(n10495), .ZN(n11383) );
  NAND2_X1 U12255 ( .A1(n12954), .A2(n9629), .ZN(n12961) );
  AND2_X1 U12256 ( .A1(n11376), .A2(n11375), .ZN(n13276) );
  INV_X1 U12257 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n15864) );
  NOR2_X1 U12258 ( .A1(n10342), .A2(n10341), .ZN(n10336) );
  INV_X1 U12259 ( .A(n15965), .ZN(n15912) );
  AND2_X1 U12260 ( .A1(n13105), .A2(n13104), .ZN(n15955) );
  INV_X1 U12261 ( .A(n9595), .ZN(n16120) );
  INV_X1 U12262 ( .A(n10223), .ZN(n10222) );
  OAI21_X1 U12263 ( .B1(n14010), .B2(n10231), .A(n10226), .ZN(n10223) );
  AND2_X1 U12264 ( .A1(n14089), .A2(n10227), .ZN(n10226) );
  NAND2_X1 U12265 ( .A1(n10230), .A2(n13735), .ZN(n10227) );
  NAND2_X1 U12266 ( .A1(n10233), .A2(n14016), .ZN(n14018) );
  AND2_X1 U12267 ( .A1(n14088), .A2(n14037), .ZN(n14020) );
  NAND2_X1 U12268 ( .A1(n10233), .A2(n10230), .ZN(n14088) );
  OAI21_X1 U12269 ( .B1(n10228), .B2(n14008), .A(n14007), .ZN(n14090) );
  INV_X1 U12270 ( .A(n10229), .ZN(n10228) );
  NAND2_X1 U12271 ( .A1(n10957), .A2(n10956), .ZN(n10976) );
  AND2_X1 U12272 ( .A1(n16116), .A2(n16115), .ZN(n16234) );
  NAND2_X1 U12273 ( .A1(n10244), .A2(n10248), .ZN(n16233) );
  NAND2_X1 U12274 ( .A1(n16247), .A2(n16079), .ZN(n10244) );
  AND2_X1 U12275 ( .A1(n16014), .A2(n16025), .ZN(n10394) );
  AND2_X1 U12276 ( .A1(n14095), .A2(n9734), .ZN(n16274) );
  AND2_X1 U12277 ( .A1(n12856), .A2(n12855), .ZN(n15721) );
  CLKBUF_X1 U12278 ( .A(n12858), .Z(n15723) );
  NAND2_X1 U12279 ( .A1(n14095), .A2(n10396), .ZN(n16279) );
  INV_X1 U12280 ( .A(n12655), .ZN(n13527) );
  AND2_X1 U12281 ( .A1(n12850), .A2(n12849), .ZN(n14324) );
  CLKBUF_X1 U12282 ( .A(n14322), .Z(n14323) );
  AND2_X1 U12283 ( .A1(n10413), .A2(n10118), .ZN(n10117) );
  INV_X1 U12284 ( .A(n14050), .ZN(n10118) );
  AND3_X1 U12285 ( .A1(n12821), .A2(n12820), .A3(n12819), .ZN(n13063) );
  AND3_X1 U12286 ( .A1(n12806), .A2(n12805), .A3(n12804), .ZN(n13759) );
  AND2_X1 U12287 ( .A1(n13551), .A2(n10416), .ZN(n13552) );
  AND3_X1 U12288 ( .A1(n12751), .A2(n12750), .A3(n12749), .ZN(n13553) );
  AND3_X1 U12289 ( .A1(n12765), .A2(n12764), .A3(n12763), .ZN(n13556) );
  AND3_X1 U12290 ( .A1(n12730), .A2(n12729), .A3(n12728), .ZN(n15885) );
  AND2_X1 U12291 ( .A1(n19768), .A2(n13531), .ZN(n14326) );
  AND2_X1 U12292 ( .A1(n19768), .A2(n13529), .ZN(n16408) );
  NOR2_X1 U12293 ( .A1(n13329), .A2(n19706), .ZN(n13487) );
  NAND2_X1 U12294 ( .A1(n10404), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10403) );
  NOR2_X1 U12295 ( .A1(n12996), .A2(n10405), .ZN(n10404) );
  INV_X1 U12296 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10405) );
  AND2_X1 U12297 ( .A1(n12916), .A2(n10410), .ZN(n12989) );
  AND2_X1 U12298 ( .A1(n9649), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U12299 ( .A1(n12916), .A2(n9649), .ZN(n12986) );
  INV_X1 U12300 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U12301 ( .A1(n12916), .A2(n10411), .ZN(n12983) );
  INV_X1 U12302 ( .A(n12964), .ZN(n11241) );
  NAND2_X1 U12303 ( .A1(n10514), .A2(n13279), .ZN(n10513) );
  INV_X1 U12304 ( .A(n10516), .ZN(n10514) );
  INV_X1 U12305 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16619) );
  AND2_X1 U12306 ( .A1(n11166), .A2(n11151), .ZN(n9976) );
  NAND2_X1 U12307 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10400), .ZN(
        n12950) );
  AND4_X1 U12308 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10400) );
  AND2_X1 U12309 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U12310 ( .A1(n13081), .A2(n13078), .ZN(n13082) );
  NAND2_X1 U12311 ( .A1(n13086), .A2(n13081), .ZN(n13083) );
  NOR2_X1 U12312 ( .A1(n13123), .A2(n13163), .ZN(n10106) );
  NAND2_X1 U12313 ( .A1(n13098), .A2(n13097), .ZN(n13127) );
  NAND2_X1 U12314 ( .A1(n13095), .A2(n13096), .ZN(n13097) );
  OR2_X1 U12315 ( .A1(n11434), .A2(n10089), .ZN(n10088) );
  NAND2_X1 U12316 ( .A1(n11434), .A2(n16430), .ZN(n10083) );
  NOR2_X1 U12317 ( .A1(n16431), .A2(n10089), .ZN(n10084) );
  NOR2_X1 U12318 ( .A1(n16731), .A2(n17340), .ZN(n10184) );
  INV_X1 U12319 ( .A(n16739), .ZN(n9979) );
  INV_X1 U12320 ( .A(n16443), .ZN(n10268) );
  NAND2_X1 U12321 ( .A1(n10277), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10276) );
  INV_X1 U12322 ( .A(n16440), .ZN(n10277) );
  NAND2_X1 U12323 ( .A1(n16443), .A2(n10271), .ZN(n10270) );
  NAND2_X1 U12324 ( .A1(n10275), .A2(n10272), .ZN(n10271) );
  INV_X1 U12325 ( .A(n10276), .ZN(n10272) );
  OR2_X1 U12326 ( .A1(n15627), .A2(n11143), .ZN(n16440) );
  NAND2_X1 U12327 ( .A1(n13144), .A2(n13145), .ZN(n15633) );
  INV_X1 U12328 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U12329 ( .A1(n13120), .A2(n9632), .ZN(n16772) );
  INV_X1 U12330 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21670) );
  NAND2_X1 U12331 ( .A1(n16873), .A2(n10110), .ZN(n16781) );
  OR2_X1 U12332 ( .A1(n16937), .A2(n10441), .ZN(n16800) );
  OR2_X1 U12333 ( .A1(n10442), .A2(n16850), .ZN(n10441) );
  AND2_X1 U12334 ( .A1(n15688), .A2(n15687), .ZN(n15674) );
  OR2_X1 U12335 ( .A1(n11411), .A2(n16798), .ZN(n16493) );
  NAND2_X1 U12336 ( .A1(n13120), .A2(n13119), .ZN(n16812) );
  NAND2_X1 U12337 ( .A1(n16873), .A2(n12896), .ZN(n16824) );
  NOR2_X1 U12338 ( .A1(n9973), .A2(n12673), .ZN(n9972) );
  INV_X1 U12339 ( .A(n9974), .ZN(n9973) );
  OR3_X1 U12340 ( .A1(n15751), .A2(n11143), .A3(n16526), .ZN(n16529) );
  NAND2_X1 U12341 ( .A1(n10509), .A2(n10510), .ZN(n15756) );
  INV_X1 U12342 ( .A(n14395), .ZN(n10509) );
  OR2_X1 U12343 ( .A1(n9706), .A2(n12907), .ZN(n10486) );
  NOR2_X1 U12344 ( .A1(n12904), .A2(n10491), .ZN(n10490) );
  INV_X1 U12345 ( .A(n16558), .ZN(n10491) );
  NOR2_X1 U12346 ( .A1(n16866), .A2(n17330), .ZN(n10372) );
  OR2_X1 U12347 ( .A1(n16937), .A2(n10442), .ZN(n16847) );
  NAND2_X1 U12348 ( .A1(n13051), .A2(n10037), .ZN(n10032) );
  NAND2_X1 U12349 ( .A1(n10445), .A2(n12893), .ZN(n10444) );
  INV_X1 U12350 ( .A(n12891), .ZN(n10445) );
  NAND2_X1 U12351 ( .A1(n9616), .A2(n16630), .ZN(n10262) );
  NAND2_X1 U12352 ( .A1(n10264), .A2(n9616), .ZN(n10261) );
  NOR2_X1 U12353 ( .A1(n16943), .A2(n16973), .ZN(n10112) );
  AND3_X1 U12354 ( .A1(n12791), .A2(n12790), .A3(n12789), .ZN(n13639) );
  INV_X1 U12355 ( .A(n15848), .ZN(n10515) );
  OAI211_X1 U12356 ( .C1(n10081), .C2(n11322), .A(n11290), .B(n11289), .ZN(
        n16680) );
  NAND2_X1 U12357 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  INV_X1 U12358 ( .A(n15900), .ZN(n10119) );
  XNOR2_X1 U12359 ( .A(n11115), .B(n11114), .ZN(n9797) );
  NAND2_X1 U12360 ( .A1(n10958), .A2(n10259), .ZN(n10978) );
  AND2_X1 U12361 ( .A1(n16235), .A2(n11291), .ZN(n13288) );
  NAND2_X1 U12362 ( .A1(n13472), .A2(n13471), .ZN(n13474) );
  AND3_X1 U12363 ( .A1(n12880), .A2(n12879), .A3(n12878), .ZN(n14350) );
  CLKBUF_X1 U12364 ( .A(n12675), .Z(n12676) );
  NAND2_X1 U12365 ( .A1(n10908), .A2(n19856), .ZN(n10255) );
  AND2_X1 U12366 ( .A1(n19839), .A2(n20103), .ZN(n19892) );
  AND2_X1 U12367 ( .A1(n20169), .A2(n20509), .ZN(n19947) );
  AND2_X1 U12368 ( .A1(n20230), .A2(n20103), .ZN(n20135) );
  NAND2_X1 U12369 ( .A1(n10869), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10870) );
  NAND2_X1 U12370 ( .A1(n10864), .A2(n14341), .ZN(n10871) );
  INV_X1 U12371 ( .A(n12867), .ZN(n19856) );
  NAND2_X1 U12372 ( .A1(n10505), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U12373 ( .A1(n10507), .A2(n14341), .ZN(n10506) );
  AND2_X1 U12374 ( .A1(n20361), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19880) );
  NOR2_X2 U12375 ( .A1(n14325), .A2(n17028), .ZN(n19884) );
  NOR2_X2 U12376 ( .A1(n17029), .A2(n17028), .ZN(n19883) );
  NAND2_X1 U12377 ( .A1(n14387), .A2(n20559), .ZN(n20551) );
  NOR2_X1 U12378 ( .A1(n13335), .A2(n13334), .ZN(n14377) );
  NOR2_X1 U12379 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14382) );
  INV_X1 U12380 ( .A(n19694), .ZN(n19684) );
  NAND2_X1 U12381 ( .A1(n17748), .A2(n17493), .ZN(n10300) );
  NOR2_X1 U12383 ( .A1(n17481), .A2(n17483), .ZN(n17482) );
  OAI21_X1 U12384 ( .B1(n17555), .B2(n10291), .A(n10290), .ZN(n17544) );
  NAND2_X1 U12385 ( .A1(n10294), .A2(n10292), .ZN(n10291) );
  NAND2_X1 U12386 ( .A1(n10301), .A2(n10294), .ZN(n10290) );
  INV_X1 U12387 ( .A(n18580), .ZN(n10294) );
  NAND2_X1 U12388 ( .A1(n17557), .A2(n18005), .ZN(n17556) );
  NAND2_X1 U12389 ( .A1(n10293), .A2(n10292), .ZN(n10295) );
  INV_X1 U12390 ( .A(n17555), .ZN(n10293) );
  NAND2_X1 U12391 ( .A1(n17704), .A2(n17695), .ZN(n17680) );
  NOR2_X1 U12392 ( .A1(n18422), .A2(n10358), .ZN(n10357) );
  NOR2_X1 U12393 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10613) );
  OR2_X1 U12394 ( .A1(n13934), .A2(n13933), .ZN(n14168) );
  OR2_X1 U12395 ( .A1(n13858), .A2(n13857), .ZN(n13970) );
  OAI21_X1 U12396 ( .B1(n9603), .B2(n17885), .A(n9701), .ZN(n13881) );
  NOR2_X1 U12397 ( .A1(n18473), .A2(n18414), .ZN(n18442) );
  INV_X1 U12398 ( .A(n18473), .ZN(n18474) );
  NAND2_X1 U12399 ( .A1(n14477), .A2(n9648), .ZN(n17081) );
  NAND2_X1 U12400 ( .A1(n18597), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18574) );
  INV_X1 U12401 ( .A(n18650), .ZN(n10306) );
  AND2_X1 U12402 ( .A1(n10571), .A2(n10308), .ZN(n10307) );
  INV_X1 U12403 ( .A(n17627), .ZN(n10308) );
  AND2_X1 U12404 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18942), .ZN(
        n17065) );
  NAND2_X1 U12405 ( .A1(n10305), .A2(n10307), .ZN(n18648) );
  INV_X1 U12406 ( .A(n17638), .ZN(n18700) );
  NOR2_X1 U12407 ( .A1(n10586), .A2(n17627), .ZN(n18701) );
  NAND2_X1 U12408 ( .A1(n10289), .A2(n9639), .ZN(n17126) );
  INV_X1 U12409 ( .A(n17745), .ZN(n10289) );
  AND2_X1 U12410 ( .A1(n18828), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10028) );
  INV_X1 U12411 ( .A(n18861), .ZN(n9874) );
  NAND2_X1 U12412 ( .A1(n9883), .A2(n9695), .ZN(n18697) );
  NOR2_X1 U12413 ( .A1(n18717), .A2(n18969), .ZN(n18944) );
  AND2_X1 U12414 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17249), .ZN(
        n18941) );
  INV_X1 U12415 ( .A(n18697), .ZN(n18985) );
  NAND2_X1 U12416 ( .A1(n18739), .A2(n10021), .ZN(n17130) );
  INV_X1 U12417 ( .A(n14164), .ZN(n10022) );
  NAND2_X1 U12418 ( .A1(n9878), .A2(n9876), .ZN(n18733) );
  INV_X1 U12419 ( .A(n14178), .ZN(n9877) );
  XNOR2_X1 U12420 ( .A(n14174), .B(n14175), .ZN(n18751) );
  NOR2_X1 U12421 ( .A1(n18751), .A2(n19026), .ZN(n18750) );
  NOR2_X1 U12422 ( .A1(n13946), .A2(n13947), .ZN(n14171) );
  AND2_X1 U12423 ( .A1(n9943), .A2(n9710), .ZN(n18772) );
  NAND2_X1 U12424 ( .A1(n18772), .A2(n18773), .ZN(n18771) );
  OAI21_X1 U12425 ( .B1(n18784), .B2(n10378), .A(n10376), .ZN(n18766) );
  INV_X1 U12426 ( .A(n13607), .ZN(n10363) );
  NOR2_X1 U12427 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19533) );
  INV_X1 U12428 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19528) );
  NOR2_X1 U12429 ( .A1(n10732), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19339) );
  OR2_X1 U12430 ( .A1(n10619), .A2(n10618), .ZN(n19111) );
  NOR2_X1 U12431 ( .A1(n19099), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19461) );
  NOR2_X1 U12432 ( .A1(n19102), .A2(n10212), .ZN(n19551) );
  AOI211_X1 U12433 ( .C1(n19679), .C2(n19681), .A(n19677), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19550) );
  NAND2_X1 U12434 ( .A1(n13198), .A2(n13197), .ZN(n13199) );
  AND4_X1 U12435 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n21524), .ZN(
        n13197) );
  NAND2_X1 U12436 ( .A1(n13230), .A2(n13229), .ZN(n13231) );
  AND4_X1 U12437 ( .A1(n13228), .A2(n13227), .A3(n13226), .A4(n21626), .ZN(
        n13229) );
  NOR2_X1 U12438 ( .A1(n12056), .A2(n9837), .ZN(n14554) );
  NAND2_X1 U12439 ( .A1(n14226), .A2(n14225), .ZN(n21588) );
  INV_X1 U12440 ( .A(n20603), .ZN(n20620) );
  AND2_X1 U12441 ( .A1(n14250), .A2(n14238), .ZN(n20647) );
  INV_X1 U12442 ( .A(n20611), .ZN(n20655) );
  INV_X1 U12443 ( .A(n20629), .ZN(n20641) );
  NAND2_X1 U12444 ( .A1(n13646), .A2(n13645), .ZN(n13644) );
  XNOR2_X1 U12445 ( .A(n10432), .B(n13458), .ZN(n13646) );
  AND2_X1 U12446 ( .A1(n13464), .A2(n13463), .ZN(n20662) );
  OR2_X1 U12447 ( .A1(n13460), .A2(n14530), .ZN(n13461) );
  INV_X1 U12448 ( .A(n20658), .ZN(n14933) );
  INV_X1 U12449 ( .A(n15014), .ZN(n15005) );
  NAND2_X1 U12450 ( .A1(n15036), .A2(n13200), .ZN(n15003) );
  INV_X1 U12451 ( .A(n15001), .ZN(n15016) );
  AND2_X1 U12452 ( .A1(n13570), .A2(n13183), .ZN(n13184) );
  OR2_X1 U12453 ( .A1(n13187), .A2(n14545), .ZN(n13188) );
  AND2_X1 U12454 ( .A1(n15003), .A2(n13705), .ZN(n15037) );
  INV_X1 U12455 ( .A(n20695), .ZN(n13432) );
  NOR2_X2 U12456 ( .A1(n20728), .A2(n13777), .ZN(n20713) );
  AND2_X1 U12457 ( .A1(n13772), .A2(n17309), .ZN(n13773) );
  XNOR2_X1 U12458 ( .A(n14224), .B(n14223), .ZN(n14503) );
  INV_X1 U12459 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21627) );
  INV_X1 U12460 ( .A(n20797), .ZN(n20737) );
  NAND2_X1 U12461 ( .A1(n9851), .A2(n9684), .ZN(n14493) );
  XNOR2_X1 U12462 ( .A(n9857), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15312) );
  OAI21_X1 U12463 ( .B1(n11852), .B2(n15239), .A(n9858), .ZN(n9857) );
  NAND2_X1 U12464 ( .A1(n15060), .A2(n15239), .ZN(n9858) );
  NAND2_X1 U12465 ( .A1(n15089), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10128) );
  NAND2_X1 U12466 ( .A1(n10453), .A2(n11844), .ZN(n9962) );
  NAND2_X1 U12467 ( .A1(n15126), .A2(n11844), .ZN(n15125) );
  NAND2_X1 U12468 ( .A1(n9964), .A2(n9965), .ZN(n15126) );
  NAND2_X1 U12469 ( .A1(n10388), .A2(n9596), .ZN(n15141) );
  NAND2_X1 U12470 ( .A1(n10164), .A2(n10161), .ZN(n15156) );
  NAND2_X1 U12471 ( .A1(n15162), .A2(n10162), .ZN(n10161) );
  NAND2_X1 U12472 ( .A1(n15164), .A2(n15155), .ZN(n10164) );
  AND2_X1 U12473 ( .A1(n15185), .A2(n11834), .ZN(n10066) );
  NAND2_X1 U12474 ( .A1(n15541), .A2(n9674), .ZN(n14926) );
  AND2_X1 U12475 ( .A1(n12091), .A2(n13565), .ZN(n20770) );
  OR2_X1 U12476 ( .A1(n20770), .A2(n15510), .ZN(n20782) );
  INV_X1 U12477 ( .A(n9585), .ZN(n21433) );
  INV_X1 U12478 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21623) );
  OR2_X1 U12479 ( .A1(n17305), .A2(n21282), .ZN(n13696) );
  INV_X1 U12480 ( .A(n13696), .ZN(n15575) );
  NOR2_X1 U12481 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15570) );
  OAI211_X1 U12482 ( .C1(n20968), .C2(n21503), .A(n21200), .B(n20806), .ZN(
        n20851) );
  AND2_X1 U12483 ( .A1(n20858), .A2(n20857), .ZN(n20888) );
  AND2_X1 U12484 ( .A1(n20970), .A2(n20969), .ZN(n21000) );
  OAI21_X1 U12485 ( .B1(n20977), .B2(n20976), .A(n21378), .ZN(n21003) );
  AND2_X1 U12486 ( .A1(n21009), .A2(n21008), .ZN(n21038) );
  OAI21_X1 U12487 ( .B1(n21015), .B2(n21014), .A(n21439), .ZN(n21041) );
  OR2_X1 U12488 ( .A1(n21088), .A2(n21087), .ZN(n21125) );
  AND2_X1 U12489 ( .A1(n21123), .A2(n21122), .ZN(n21151) );
  AND2_X1 U12490 ( .A1(n21239), .A2(n21238), .ZN(n21267) );
  INV_X1 U12491 ( .A(n21447), .ZN(n21293) );
  INV_X1 U12492 ( .A(n21454), .ZN(n21297) );
  INV_X1 U12493 ( .A(n21461), .ZN(n21301) );
  INV_X1 U12494 ( .A(n21468), .ZN(n21305) );
  INV_X1 U12495 ( .A(n21482), .ZN(n21313) );
  OR2_X1 U12496 ( .A1(n21372), .A2(n21274), .ZN(n21336) );
  OAI22_X1 U12497 ( .A1(n21288), .A2(n21287), .B1(n21286), .B2(n21285), .ZN(
        n21318) );
  INV_X1 U12498 ( .A(n21491), .ZN(n21319) );
  AND2_X1 U12499 ( .A1(n21330), .A2(n21329), .ZN(n21358) );
  NAND2_X1 U12500 ( .A1(n11562), .A2(n20846), .ZN(n21429) );
  OR2_X1 U12501 ( .A1(n20975), .A2(n20807), .ZN(n21430) );
  NAND2_X1 U12502 ( .A1(n21581), .A2(n20846), .ZN(n21446) );
  OR2_X1 U12503 ( .A1(n20975), .A2(n20816), .ZN(n21447) );
  NAND2_X1 U12504 ( .A1(n20819), .A2(n20846), .ZN(n21453) );
  OR2_X1 U12505 ( .A1(n20975), .A2(n20821), .ZN(n21454) );
  NAND2_X1 U12506 ( .A1(n20824), .A2(n20846), .ZN(n21460) );
  OR2_X1 U12507 ( .A1(n20975), .A2(n20826), .ZN(n21461) );
  NAND2_X1 U12508 ( .A1(n20829), .A2(n20846), .ZN(n21467) );
  OR2_X1 U12509 ( .A1(n20975), .A2(n20831), .ZN(n21468) );
  NAND2_X1 U12510 ( .A1(n20834), .A2(n20846), .ZN(n21474) );
  OR2_X1 U12511 ( .A1(n20975), .A2(n20836), .ZN(n21475) );
  OR2_X1 U12512 ( .A1(n20975), .A2(n20841), .ZN(n21482) );
  OR2_X1 U12513 ( .A1(n21372), .A2(n21087), .ZN(n21498) );
  NAND2_X1 U12514 ( .A1(n11551), .A2(n20846), .ZN(n21488) );
  OR2_X1 U12515 ( .A1(n20975), .A2(n20849), .ZN(n21491) );
  AND2_X1 U12516 ( .A1(n21428), .A2(n21427), .ZN(n21490) );
  NAND2_X1 U12517 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21590) );
  INV_X1 U12518 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21503) );
  INV_X1 U12519 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21500) );
  INV_X1 U12520 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21282) );
  INV_X1 U12521 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21524) );
  INV_X1 U12522 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20356) );
  NAND2_X1 U12523 ( .A1(n13034), .A2(n11265), .ZN(n15641) );
  NAND2_X1 U12524 ( .A1(n11264), .A2(n10555), .ZN(n11265) );
  AND2_X1 U12525 ( .A1(n11350), .A2(n9669), .ZN(n19742) );
  NAND2_X1 U12526 ( .A1(n11359), .A2(n10354), .ZN(n11348) );
  INV_X1 U12527 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16660) );
  OR3_X1 U12528 ( .A1(n20545), .A2(n19745), .A3(n13041), .ZN(n19748) );
  INV_X1 U12529 ( .A(n19767), .ZN(n15951) );
  XNOR2_X1 U12530 ( .A(n12934), .B(n12933), .ZN(n13162) );
  AOI21_X1 U12531 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12931), .ZN(n12933) );
  OR2_X1 U12532 ( .A1(n12844), .A2(n12843), .ZN(n14401) );
  OR2_X1 U12533 ( .A1(n12831), .A2(n12830), .ZN(n14317) );
  OR2_X1 U12534 ( .A1(n12818), .A2(n12817), .ZN(n14318) );
  OR2_X1 U12535 ( .A1(n12747), .A2(n12746), .ZN(n16304) );
  NOR2_X1 U12536 ( .A1(n14274), .A2(n14273), .ZN(n16291) );
  INV_X1 U12537 ( .A(n16301), .ZN(n16311) );
  INV_X1 U12538 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15939) );
  XNOR2_X1 U12539 ( .A(n13094), .B(n13029), .ZN(n14552) );
  AND2_X1 U12540 ( .A1(n16398), .A2(n19770), .ZN(n16424) );
  INV_X1 U12541 ( .A(n19770), .ZN(n19786) );
  INV_X1 U12542 ( .A(n16421), .ZN(n19794) );
  INV_X1 U12543 ( .A(n16398), .ZN(n19790) );
  OR2_X1 U12544 ( .A1(n16408), .A2(n14326), .ZN(n16421) );
  INV_X1 U12545 ( .A(n13536), .ZN(n19795) );
  NAND2_X1 U12546 ( .A1(n19828), .A2(n13537), .ZN(n19798) );
  INV_X1 U12547 ( .A(n19798), .ZN(n19826) );
  NAND2_X1 U12548 ( .A1(n13306), .A2(n13488), .ZN(n19834) );
  NOR2_X1 U12549 ( .A1(n16722), .A2(n10100), .ZN(n10099) );
  INV_X1 U12550 ( .A(n10104), .ZN(n10100) );
  NAND2_X1 U12551 ( .A1(n13088), .A2(n13089), .ZN(n10333) );
  NOR2_X1 U12552 ( .A1(n13084), .A2(n16707), .ZN(n10102) );
  INV_X1 U12553 ( .A(n16682), .ZN(n16719) );
  NAND2_X1 U12554 ( .A1(n16452), .A2(n9658), .ZN(n10101) );
  NAND2_X1 U12555 ( .A1(n16427), .A2(n13081), .ZN(n10098) );
  NAND2_X1 U12556 ( .A1(n10105), .A2(n13081), .ZN(n10104) );
  INV_X1 U12557 ( .A(n10106), .ZN(n10105) );
  OR2_X1 U12558 ( .A1(n9622), .A2(n15631), .ZN(n16752) );
  NAND2_X1 U12559 ( .A1(n10327), .A2(n16457), .ZN(n16768) );
  NAND2_X1 U12560 ( .A1(n10500), .A2(n10499), .ZN(n12923) );
  NAND2_X1 U12561 ( .A1(n10258), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10499) );
  NAND2_X1 U12562 ( .A1(n16557), .A2(n10501), .ZN(n10500) );
  AND2_X1 U12563 ( .A1(n10258), .A2(n9653), .ZN(n10501) );
  XNOR2_X1 U12564 ( .A(n10476), .B(n10547), .ZN(n12924) );
  NAND2_X1 U12565 ( .A1(n16505), .A2(n12912), .ZN(n10476) );
  INV_X1 U12566 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16875) );
  INV_X1 U12567 ( .A(n16556), .ZN(n16859) );
  AND2_X1 U12568 ( .A1(n16974), .A2(n9770), .ZN(n16899) );
  NOR2_X1 U12569 ( .A1(n16937), .A2(n10444), .ZN(n16902) );
  NAND2_X1 U12570 ( .A1(n16609), .A2(n9773), .ZN(n16588) );
  INV_X1 U12571 ( .A(n9785), .ZN(n16601) );
  NAND2_X1 U12572 ( .A1(n10456), .A2(n10460), .ZN(n16645) );
  NAND2_X1 U12573 ( .A1(n16653), .A2(n10461), .ZN(n10456) );
  NOR2_X1 U12574 ( .A1(n10457), .A2(n10151), .ZN(n10152) );
  AND2_X1 U12575 ( .A1(n10458), .A2(n10460), .ZN(n10151) );
  NAND2_X1 U12576 ( .A1(n16974), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16962) );
  NAND2_X1 U12577 ( .A1(n9967), .A2(n11118), .ZN(n10324) );
  INV_X1 U12578 ( .A(n16675), .ZN(n9967) );
  AND2_X1 U12579 ( .A1(n9917), .A2(n9914), .ZN(n16980) );
  AND2_X1 U12580 ( .A1(n16850), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9914) );
  NOR3_X1 U12581 ( .A1(n13286), .A2(n12887), .A3(n13252), .ZN(n17355) );
  CLKBUF_X1 U12582 ( .A(n14010), .Z(n17345) );
  INV_X1 U12583 ( .A(n16844), .ZN(n9916) );
  INV_X1 U12584 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20531) );
  OR2_X1 U12585 ( .A1(n16993), .A2(n13423), .ZN(n20526) );
  AND2_X1 U12586 ( .A1(n13421), .A2(n13422), .ZN(n13423) );
  INV_X1 U12587 ( .A(n20168), .ZN(n20509) );
  NAND2_X1 U12588 ( .A1(n13244), .A2(n12717), .ZN(n15916) );
  INV_X1 U12589 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17317) );
  NAND2_X1 U12590 ( .A1(n13745), .A2(n13456), .ZN(n20494) );
  NAND2_X1 U12591 ( .A1(n14007), .A2(n10229), .ZN(n14009) );
  INV_X1 U12592 ( .A(n14008), .ZN(n13746) );
  AND2_X1 U12593 ( .A1(n14370), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17016) );
  INV_X1 U12594 ( .A(n17002), .ZN(n17010) );
  OAI21_X1 U12595 ( .B1(n11053), .B2(n20552), .A(n20501), .ZN(n19845) );
  OAI21_X1 U12596 ( .B1(n19843), .B2(n20552), .A(n19842), .ZN(n19882) );
  NAND2_X1 U12597 ( .A1(n17045), .A2(n20269), .ZN(n20041) );
  NAND2_X1 U12598 ( .A1(n17040), .A2(n17039), .ZN(n20037) );
  AND2_X1 U12599 ( .A1(n20050), .A2(n20361), .ZN(n20061) );
  INV_X1 U12600 ( .A(n20061), .ZN(n20073) );
  INV_X1 U12601 ( .A(n20041), .ZN(n20072) );
  OAI21_X1 U12602 ( .B1(n20079), .B2(n20171), .A(n20051), .ZN(n20071) );
  OAI21_X1 U12603 ( .B1(n20078), .B2(n20543), .A(n20077), .ZN(n20098) );
  NOR2_X1 U12604 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20141), .ZN(
        n20127) );
  NAND2_X1 U12605 ( .A1(n20135), .A2(n20269), .ZN(n20172) );
  OAI21_X1 U12606 ( .B1(n20202), .B2(n20171), .A(n20170), .ZN(n20193) );
  OAI21_X1 U12607 ( .B1(n20201), .B2(n20543), .A(n20200), .ZN(n20225) );
  INV_X1 U12608 ( .A(n20240), .ZN(n21755) );
  AOI21_X1 U12609 ( .B1(n20552), .B2(n20235), .A(n20237), .ZN(n21752) );
  INV_X1 U12610 ( .A(n20369), .ZN(n20315) );
  INV_X1 U12611 ( .A(n20296), .ZN(n20352) );
  OAI22_X1 U12612 ( .A1(n19851), .A2(n19873), .B1(n21618), .B2(n19871), .ZN(
        n20369) );
  INV_X1 U12613 ( .A(n20311), .ZN(n20367) );
  INV_X1 U12614 ( .A(n20316), .ZN(n21750) );
  INV_X1 U12615 ( .A(n20325), .ZN(n20383) );
  INV_X1 U12616 ( .A(n20330), .ZN(n20389) );
  AND2_X1 U12617 ( .A1(n19880), .A2(n19875), .ZN(n20395) );
  AND2_X1 U12618 ( .A1(n20354), .A2(n20269), .ZN(n20406) );
  AOI22_X1 U12619 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19883), .ZN(n20411) );
  INV_X1 U12620 ( .A(n20340), .ZN(n20401) );
  AND2_X1 U12621 ( .A1(n20360), .A2(n20351), .ZN(n20404) );
  INV_X1 U12622 ( .A(n20493), .ZN(n17050) );
  NAND2_X1 U12623 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20547) );
  AND3_X1 U12624 ( .A1(n20413), .A2(n20477), .A3(n20414), .ZN(n20560) );
  INV_X1 U12625 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20431) );
  NAND2_X1 U12626 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20413), .ZN(n20566) );
  NOR2_X1 U12627 ( .A1(n9898), .A2(n9897), .ZN(n17450) );
  INV_X1 U12628 ( .A(n13629), .ZN(n9898) );
  NOR2_X1 U12629 ( .A1(n17517), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17503) );
  INV_X1 U12630 ( .A(n10303), .ZN(n17492) );
  NOR2_X1 U12631 ( .A1(n17539), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17524) );
  NAND2_X1 U12632 ( .A1(n17524), .A2(n17518), .ZN(n17517) );
  NAND2_X1 U12633 ( .A1(n17545), .A2(n17936), .ZN(n17539) );
  NOR2_X1 U12634 ( .A1(n13258), .A2(n10301), .ZN(n17555) );
  INV_X1 U12635 ( .A(n10295), .ZN(n17554) );
  NOR2_X1 U12636 ( .A1(n17568), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17557) );
  NAND2_X1 U12637 ( .A1(n17579), .A2(n18038), .ZN(n17568) );
  NAND2_X1 U12638 ( .A1(n17748), .A2(n18571), .ZN(n10591) );
  NOR2_X1 U12639 ( .A1(n17589), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17579) );
  NOR2_X1 U12640 ( .A1(n17644), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17621) );
  NAND2_X1 U12641 ( .A1(n17621), .A2(n21713), .ZN(n17617) );
  NOR2_X1 U12642 ( .A1(n17669), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17649) );
  NAND2_X1 U12643 ( .A1(n17649), .A2(n18113), .ZN(n17644) );
  NAND2_X1 U12644 ( .A1(n17723), .A2(n17719), .ZN(n17718) );
  INV_X1 U12645 ( .A(n17774), .ZN(n17805) );
  NOR2_X1 U12646 ( .A1(n17737), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17723) );
  AND3_X1 U12647 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n17778) );
  INV_X1 U12648 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n9869) );
  OR2_X1 U12649 ( .A1(n19695), .A2(n10759), .ZN(n17812) );
  INV_X1 U12650 ( .A(n19131), .ZN(n17935) );
  AND2_X1 U12651 ( .A1(n17955), .A2(n10311), .ZN(n17945) );
  NAND2_X1 U12652 ( .A1(n18269), .A2(n17937), .ZN(n10311) );
  NOR2_X1 U12653 ( .A1(n17936), .A2(n17967), .ZN(n17971) );
  AND2_X1 U12654 ( .A1(n18073), .A2(n10317), .ZN(n17972) );
  AND2_X1 U12655 ( .A1(n9651), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n10317) );
  INV_X1 U12656 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18075) );
  NAND2_X1 U12657 ( .A1(n18073), .A2(n17935), .ZN(n18074) );
  AND2_X1 U12658 ( .A1(n9652), .A2(n9614), .ZN(n10321) );
  NOR2_X1 U12659 ( .A1(n18200), .A2(n17695), .ZN(n10322) );
  NAND2_X1 U12660 ( .A1(n18243), .A2(n9652), .ZN(n18183) );
  NAND2_X1 U12661 ( .A1(n18243), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n18197) );
  AND2_X1 U12662 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18247), .ZN(n18243) );
  NOR2_X1 U12663 ( .A1(n17259), .A2(n9738), .ZN(n18272) );
  INV_X1 U12664 ( .A(n18284), .ZN(n18279) );
  AND2_X1 U12665 ( .A1(n18304), .A2(n10356), .ZN(n18290) );
  AND2_X1 U12666 ( .A1(n9654), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U12667 ( .A1(n18304), .A2(n9654), .ZN(n18296) );
  INV_X1 U12668 ( .A(n18308), .ZN(n18304) );
  NAND2_X1 U12669 ( .A1(n18304), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18303) );
  NOR2_X1 U12670 ( .A1(n18313), .A2(n19131), .ZN(n18309) );
  NAND2_X1 U12671 ( .A1(n18309), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18308) );
  NOR2_X1 U12672 ( .A1(n18352), .A2(n10361), .ZN(n18314) );
  INV_X1 U12673 ( .A(n18318), .ZN(n10362) );
  NAND2_X1 U12674 ( .A1(n18314), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18313) );
  INV_X1 U12675 ( .A(n18319), .ZN(n18382) );
  NAND2_X1 U12676 ( .A1(n18356), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18352) );
  NOR2_X1 U12677 ( .A1(n18361), .A2(n18522), .ZN(n18356) );
  INV_X1 U12678 ( .A(n18408), .ZN(n18357) );
  AND2_X1 U12679 ( .A1(n18383), .A2(n19675), .ZN(n10360) );
  INV_X1 U12680 ( .A(n14168), .ZN(n18401) );
  INV_X1 U12681 ( .A(n13970), .ZN(n18404) );
  INV_X1 U12682 ( .A(n18389), .ZN(n18410) );
  NAND2_X1 U12683 ( .A1(n14203), .A2(n17935), .ZN(n18319) );
  INV_X1 U12684 ( .A(n18413), .ZN(n18378) );
  INV_X1 U12685 ( .A(n18521), .ZN(n18513) );
  INV_X1 U12686 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18522) );
  NAND2_X1 U12687 ( .A1(n18474), .A2(n19551), .ZN(n18521) );
  CLKBUF_X1 U12688 ( .A(n18512), .Z(n18518) );
  NOR2_X1 U12689 ( .A1(n18518), .A2(n19681), .ZN(n18519) );
  NAND2_X1 U12690 ( .A1(n18566), .A2(n9944), .ZN(n17067) );
  AND2_X1 U12691 ( .A1(n17233), .A2(n9945), .ZN(n9944) );
  AND2_X1 U12692 ( .A1(n17189), .A2(n17188), .ZN(n9945) );
  AND2_X1 U12693 ( .A1(n18597), .A2(n9747), .ZN(n18523) );
  INV_X1 U12694 ( .A(n18535), .ZN(n10296) );
  INV_X1 U12695 ( .A(n18566), .ZN(n18555) );
  NOR2_X1 U12696 ( .A1(n18609), .A2(n18610), .ZN(n18597) );
  NOR2_X1 U12697 ( .A1(n10304), .A2(n10586), .ZN(n18631) );
  NAND2_X1 U12698 ( .A1(n10307), .A2(n10306), .ZN(n10304) );
  AOI21_X1 U12699 ( .B1(n18927), .B2(n18812), .A(n10201), .ZN(n18656) );
  NOR2_X1 U12700 ( .A1(n18696), .A2(n18929), .ZN(n10201) );
  INV_X1 U12701 ( .A(n18730), .ZN(n18706) );
  INV_X1 U12702 ( .A(n18696), .ZN(n18698) );
  INV_X1 U12703 ( .A(n9883), .ZN(n14447) );
  INV_X1 U12704 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18753) );
  NOR2_X2 U12705 ( .A1(n19184), .A2(n19205), .ZN(n17078) );
  INV_X1 U12706 ( .A(n17078), .ZN(n19136) );
  INV_X1 U12707 ( .A(n18813), .ZN(n18803) );
  INV_X1 U12708 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19559) );
  NAND2_X1 U12709 ( .A1(n14444), .A2(n14443), .ZN(n10020) );
  INV_X1 U12710 ( .A(n18987), .ZN(n18961) );
  NAND2_X1 U12711 ( .A1(n10379), .A2(n10381), .ZN(n18552) );
  AND2_X1 U12712 ( .A1(n18626), .A2(n18828), .ZN(n18558) );
  NAND2_X1 U12713 ( .A1(n18873), .A2(n19070), .ZN(n18921) );
  NAND2_X1 U12714 ( .A1(n9886), .A2(n19061), .ZN(n18920) );
  OAI21_X1 U12715 ( .B1(n13657), .B2(n13606), .A(n13656), .ZN(n18971) );
  INV_X1 U12716 ( .A(n13608), .ZN(n13606) );
  OR2_X1 U12717 ( .A1(n17250), .A2(n18941), .ZN(n18973) );
  NAND2_X1 U12718 ( .A1(n17130), .A2(n18664), .ZN(n17167) );
  INV_X1 U12719 ( .A(n19007), .ZN(n18956) );
  NAND2_X1 U12720 ( .A1(n18748), .A2(n18747), .ZN(n18746) );
  NAND2_X1 U12721 ( .A1(n14125), .A2(n14124), .ZN(n18748) );
  INV_X1 U12722 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19026) );
  INV_X1 U12723 ( .A(n19072), .ZN(n19042) );
  INV_X1 U12724 ( .A(n9943), .ZN(n18781) );
  NOR2_X1 U12725 ( .A1(n9887), .A2(n19102), .ZN(n9885) );
  OR2_X1 U12726 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  AND2_X1 U12727 ( .A1(n19519), .A2(n19070), .ZN(n19079) );
  NAND3_X1 U12728 ( .A1(n19692), .A2(n19660), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19205) );
  INV_X1 U12729 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19095) );
  INV_X1 U12730 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19541) );
  INV_X1 U12731 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17752) );
  NAND2_X1 U12732 ( .A1(n19132), .A2(n19106), .ZN(n19477) );
  NAND2_X1 U12733 ( .A1(n19132), .A2(n19111), .ZN(n19483) );
  NAND2_X1 U12734 ( .A1(n19132), .A2(n19122), .ZN(n19495) );
  NAND2_X1 U12735 ( .A1(n19132), .A2(n19127), .ZN(n19501) );
  NAND2_X1 U12736 ( .A1(n19132), .A2(n19131), .ZN(n19511) );
  AND2_X1 U12737 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19562), .ZN(n19675) );
  NOR2_X1 U12738 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19685) );
  NOR2_X1 U12739 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19660), .ZN(
        n19553) );
  INV_X1 U12740 ( .A(n17445), .ZN(n19562) );
  AOI21_X1 U12741 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19685), .ZN(n19567) );
  INV_X1 U12742 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19660) );
  INV_X1 U12743 ( .A(n19682), .ZN(n19677) );
  INV_X1 U12744 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21578) );
  NOR2_X2 U12745 ( .A1(n17404), .A2(n17361), .ZN(n17401) );
  OAI211_X1 U12746 ( .C1(n15304), .C2(n20574), .A(n10069), .B(n10068), .ZN(
        P1_U2971) );
  AOI21_X1 U12747 ( .B1(n15172), .B2(n15057), .A(n15056), .ZN(n10069) );
  OR2_X1 U12748 ( .A1(n12102), .A2(n12101), .ZN(n12103) );
  AND2_X1 U12749 ( .A1(n13216), .A2(n13215), .ZN(n13217) );
  OAI21_X1 U12750 ( .B1(n12132), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n9585), 
        .ZN(n15560) );
  NOR2_X1 U12751 ( .A1(n13114), .A2(n13113), .ZN(n13115) );
  AOI211_X1 U12752 ( .C1(n19750), .C2(n15594), .A(n15593), .B(n15592), .ZN(
        n15599) );
  AOI21_X1 U12753 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16287), .A(n16212), .ZN(
        n16213) );
  NOR2_X1 U12754 ( .A1(n11244), .A2(n11243), .ZN(n11436) );
  NAND2_X1 U12755 ( .A1(n13132), .A2(n16713), .ZN(n11435) );
  OAI21_X1 U12756 ( .B1(n16742), .B2(n16707), .A(n16449), .ZN(P2_U2986) );
  NAND2_X1 U12757 ( .A1(n16749), .A2(n16704), .ZN(n9810) );
  OAI21_X1 U12758 ( .B1(n16820), .B2(n16707), .A(n10137), .ZN(P2_U2993) );
  INV_X1 U12759 ( .A(n10138), .ZN(n10137) );
  OAI21_X1 U12760 ( .B1(n16816), .B2(n16722), .A(n10139), .ZN(n10138) );
  AOI21_X1 U12761 ( .B1(n16818), .B2(n16719), .A(n16512), .ZN(n10139) );
  INV_X1 U12762 ( .A(n9791), .ZN(n9790) );
  OAI21_X1 U12763 ( .B1(n16918), .B2(n16707), .A(n16607), .ZN(n9791) );
  NAND2_X1 U12764 ( .A1(n16732), .A2(n17351), .ZN(n10186) );
  NOR2_X1 U12765 ( .A1(n16729), .A2(n10122), .ZN(n10183) );
  AOI211_X1 U12766 ( .C1(n16728), .C2(n16727), .A(n16726), .B(n16725), .ZN(
        n16729) );
  NAND2_X1 U12767 ( .A1(n16737), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10109) );
  AOI21_X1 U12768 ( .B1(n16749), .B2(n16984), .A(n9921), .ZN(n16750) );
  OAI21_X1 U12769 ( .B1(n16746), .B2(n16745), .A(n9922), .ZN(n9921) );
  AOI21_X1 U12770 ( .B1(n16747), .B2(n17327), .A(n9923), .ZN(n9922) );
  OAI21_X1 U12771 ( .B1(n13159), .B2(n16988), .A(n13150), .ZN(n13151) );
  AOI21_X1 U12772 ( .B1(n16778), .B2(n17351), .A(n9947), .ZN(n9966) );
  INV_X1 U12773 ( .A(n16779), .ZN(n9947) );
  INV_X1 U12774 ( .A(n10011), .ZN(n16819) );
  NAND2_X1 U12775 ( .A1(n16831), .A2(n9782), .ZN(P2_U3027) );
  INV_X1 U12776 ( .A(n9783), .ZN(n9782) );
  OAI21_X1 U12777 ( .B1(n16833), .B2(n16988), .A(n16832), .ZN(n9783) );
  AOI211_X1 U12778 ( .C1(n16842), .C2(n17351), .A(n16841), .B(n16840), .ZN(
        n16843) );
  AOI21_X1 U12779 ( .B1(n16556), .B2(n10006), .A(n10003), .ZN(n10002) );
  NAND2_X1 U12780 ( .A1(n16846), .A2(n10008), .ZN(n10001) );
  NAND2_X1 U12781 ( .A1(n16862), .A2(n17351), .ZN(n10373) );
  NAND2_X1 U12782 ( .A1(n16867), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10374) );
  OAI21_X1 U12783 ( .B1(n16587), .B2(n16988), .A(n13068), .ZN(n13069) );
  NAND2_X1 U12784 ( .A1(n9784), .A2(n9680), .ZN(n16917) );
  AND2_X1 U12785 ( .A1(n16974), .A2(n9656), .ZN(n16915) );
  OR2_X1 U12786 ( .A1(n10772), .A2(n10771), .ZN(n10773) );
  OR2_X1 U12787 ( .A1(n17801), .A2(n17478), .ZN(n10288) );
  INV_X1 U12788 ( .A(n17955), .ZN(n17949) );
  NAND2_X1 U12789 ( .A1(n18073), .A2(n9651), .ZN(n18006) );
  NAND2_X1 U12790 ( .A1(n10211), .A2(n9685), .ZN(P3_U2808) );
  NAND2_X1 U12791 ( .A1(n18578), .A2(n18872), .ZN(n10211) );
  AOI21_X1 U12792 ( .B1(n18730), .B2(n18580), .A(n10207), .ZN(n10206) );
  OAI21_X1 U12793 ( .B1(n18910), .B2(n9871), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18914) );
  NOR2_X1 U12794 ( .A1(n19062), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9871) );
  NAND2_X1 U12795 ( .A1(n17361), .A2(U214), .ZN(U212) );
  AND3_X1 U12796 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U12797 ( .A1(n14296), .A2(n9972), .ZN(n9615) );
  CLKBUF_X3 U12798 ( .A(n11634), .Z(n12491) );
  AND2_X1 U12799 ( .A1(n16615), .A2(n16627), .ZN(n9616) );
  NAND2_X1 U12800 ( .A1(n10531), .A2(n10534), .ZN(n14677) );
  AND2_X1 U12801 ( .A1(n15688), .A2(n9730), .ZN(n9617) );
  AND2_X1 U12802 ( .A1(n12717), .A2(n12722), .ZN(n9618) );
  NAND2_X1 U12803 ( .A1(n9980), .A2(n9762), .ZN(n16427) );
  OR2_X1 U12804 ( .A1(n19753), .A2(n19734), .ZN(n10546) );
  INV_X1 U12805 ( .A(n10546), .ZN(n15952) );
  AND2_X1 U12806 ( .A1(n9648), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9619) );
  OR2_X1 U12807 ( .A1(n18663), .A2(n14470), .ZN(n9620) );
  OR2_X1 U12808 ( .A1(n9620), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9621) );
  INV_X1 U12809 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18113) );
  AND2_X1 U12810 ( .A1(n15688), .A2(n9732), .ZN(n9622) );
  AND2_X1 U12811 ( .A1(n11422), .A2(n16459), .ZN(n9624) );
  AND2_X1 U12812 ( .A1(n16612), .A2(n16616), .ZN(n9625) );
  INV_X2 U12813 ( .A(n10590), .ZN(n10301) );
  CLKBUF_X3 U12814 ( .A(n11628), .Z(n12596) );
  NAND2_X1 U12815 ( .A1(n12350), .A2(n9673), .ZN(n14645) );
  NAND2_X1 U12816 ( .A1(n11372), .A2(n10345), .ZN(n9626) );
  AND4_X1 U12817 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n9627) );
  OR2_X1 U12818 ( .A1(n10340), .A2(n10342), .ZN(n9628) );
  NAND2_X1 U12819 ( .A1(n11609), .A2(n21581), .ZN(n10173) );
  AND2_X1 U12820 ( .A1(n10401), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9629) );
  AND2_X1 U12821 ( .A1(n12860), .A2(n9733), .ZN(n15691) );
  AND2_X1 U12822 ( .A1(n12808), .A2(n9681), .ZN(n13062) );
  NAND2_X1 U12823 ( .A1(n13680), .A2(n13679), .ZN(n13573) );
  NAND2_X1 U12824 ( .A1(n14095), .A2(n14096), .ZN(n15967) );
  AND2_X1 U12825 ( .A1(n11841), .A2(n15150), .ZN(n9630) );
  NAND2_X1 U12826 ( .A1(n14296), .A2(n14396), .ZN(n14395) );
  INV_X1 U12827 ( .A(n9938), .ZN(n16568) );
  NAND2_X1 U12828 ( .A1(n9980), .A2(n10503), .ZN(n9938) );
  OR2_X1 U12829 ( .A1(n10511), .A2(n15738), .ZN(n9631) );
  INV_X1 U12830 ( .A(n19879), .ZN(n12699) );
  AND2_X1 U12831 ( .A1(n13119), .A2(n16782), .ZN(n9632) );
  NAND2_X1 U12832 ( .A1(n12350), .A2(n12349), .ZN(n14722) );
  AND4_X1 U12833 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n9633) );
  AND4_X1 U12834 ( .A1(n11007), .A2(n11010), .A3(n11012), .A4(n11006), .ZN(
        n9634) );
  AND3_X1 U12835 ( .A1(n10986), .A2(n10987), .A3(n10972), .ZN(n9635) );
  CLKBUF_X2 U12836 ( .A(n11725), .Z(n11690) );
  NAND2_X1 U12837 ( .A1(n11878), .A2(n11573), .ZN(n13182) );
  INV_X1 U12838 ( .A(n13182), .ZN(n9837) );
  AND2_X1 U12839 ( .A1(n13679), .A2(n10062), .ZN(n9636) );
  OR2_X2 U12840 ( .A1(n15726), .A2(n10398), .ZN(n9637) );
  AND2_X1 U12841 ( .A1(n10307), .A2(n9696), .ZN(n9638) );
  AND2_X1 U12842 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U12843 ( .A1(n9969), .A2(n12869), .ZN(n9640) );
  AND2_X1 U12844 ( .A1(n10472), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9641) );
  NAND2_X1 U12845 ( .A1(n15688), .A2(n9729), .ZN(n13142) );
  AND2_X1 U12846 ( .A1(n10297), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9642) );
  OR2_X1 U12847 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9643) );
  AND2_X1 U12848 ( .A1(n10303), .A2(n10302), .ZN(n9644) );
  AND3_X1 U12849 ( .A1(n12726), .A2(n12725), .A3(n12724), .ZN(n15900) );
  AND2_X1 U12850 ( .A1(n9629), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9645) );
  AND2_X1 U12851 ( .A1(n11152), .A2(n11151), .ZN(n9646) );
  INV_X1 U12852 ( .A(n10212), .ZN(n9897) );
  INV_X1 U12853 ( .A(n10397), .ZN(n15727) );
  AND2_X1 U12854 ( .A1(n18073), .A2(n9750), .ZN(n9647) );
  AND2_X1 U12855 ( .A1(n10572), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9648) );
  AND2_X1 U12856 ( .A1(n12973), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12917) );
  NAND2_X1 U12857 ( .A1(n10515), .A2(n11175), .ZN(n15831) );
  AND2_X1 U12858 ( .A1(n10411), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9649) );
  AND2_X1 U12859 ( .A1(n11991), .A2(n9736), .ZN(n14803) );
  AND2_X1 U12860 ( .A1(n14477), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10573) );
  INV_X1 U12861 ( .A(n19034), .ZN(n19062) );
  AND2_X1 U12862 ( .A1(n11252), .A2(n9935), .ZN(n9650) );
  AND2_X2 U12863 ( .A1(n13652), .A2(n10609), .ZN(n17751) );
  AND2_X1 U12864 ( .A1(n9750), .A2(n10318), .ZN(n9651) );
  AND2_X1 U12865 ( .A1(n10322), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n9652) );
  INV_X1 U12866 ( .A(n13906), .ZN(n10620) );
  AND2_X1 U12867 ( .A1(n12896), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9653) );
  AND2_X1 U12868 ( .A1(n10357), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9654) );
  AND2_X1 U12869 ( .A1(n10110), .A2(n9766), .ZN(n9655) );
  AND2_X1 U12870 ( .A1(n10112), .A2(n9768), .ZN(n9656) );
  AND2_X1 U12871 ( .A1(n16782), .A2(n9767), .ZN(n9657) );
  AND2_X1 U12872 ( .A1(n10106), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9658) );
  INV_X1 U12873 ( .A(n10205), .ZN(n19519) );
  NAND2_X1 U12874 ( .A1(n9886), .A2(n9885), .ZN(n10205) );
  AND2_X2 U12875 ( .A1(n10889), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11091) );
  AND2_X2 U12876 ( .A1(n10876), .A2(n14341), .ZN(n10990) );
  INV_X1 U12877 ( .A(n13880), .ZN(n10621) );
  OR2_X1 U12878 ( .A1(n18645), .A2(n18628), .ZN(n9659) );
  NAND2_X1 U12879 ( .A1(n12871), .A2(n10923), .ZN(n10932) );
  AND2_X2 U12880 ( .A1(n16196), .A2(n14341), .ZN(n11044) );
  OR2_X1 U12881 ( .A1(n14603), .A2(n10541), .ZN(n9660) );
  AND2_X1 U12882 ( .A1(n12214), .A2(n10529), .ZN(n14765) );
  AND2_X1 U12883 ( .A1(n10199), .A2(n10919), .ZN(n12681) );
  NAND2_X2 U12884 ( .A1(n11581), .A2(n11562), .ZN(n11947) );
  XOR2_X1 U12885 ( .A(n11151), .B(n10952), .Z(n9661) );
  NAND2_X1 U12886 ( .A1(n9957), .A2(n9960), .ZN(n15104) );
  NAND2_X1 U12887 ( .A1(n12151), .A2(n12150), .ZN(n14099) );
  NAND2_X1 U12888 ( .A1(n11359), .A2(n11358), .ZN(n11354) );
  NOR2_X1 U12889 ( .A1(n12949), .A2(n16660), .ZN(n12952) );
  NAND2_X1 U12890 ( .A1(n15688), .A2(n10519), .ZN(n15655) );
  NOR2_X1 U12891 ( .A1(n14722), .A2(n14723), .ZN(n14700) );
  AND2_X1 U12892 ( .A1(n12350), .A2(n10070), .ZN(n14633) );
  AND2_X1 U12893 ( .A1(n12350), .A2(n10072), .ZN(n14657) );
  AND2_X1 U12894 ( .A1(n12214), .A2(n10528), .ZN(n14746) );
  NAND2_X1 U12895 ( .A1(n16671), .A2(n16670), .ZN(n16610) );
  NAND2_X1 U12896 ( .A1(n12860), .A2(n12859), .ZN(n13011) );
  NOR2_X1 U12897 ( .A1(n16937), .A2(n12891), .ZN(n9662) );
  NAND2_X1 U12898 ( .A1(n12954), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12956) );
  NAND2_X1 U12899 ( .A1(n11372), .A2(n11369), .ZN(n11368) );
  INV_X1 U12900 ( .A(n10339), .ZN(n11326) );
  NAND2_X1 U12901 ( .A1(n12688), .A2(n11246), .ZN(n9663) );
  INV_X1 U12902 ( .A(n10359), .ZN(n14203) );
  NAND2_X1 U12903 ( .A1(n14196), .A2(n19675), .ZN(n10359) );
  AND2_X1 U12904 ( .A1(n18304), .A2(n10357), .ZN(n9664) );
  OR2_X1 U12905 ( .A1(n9631), .A2(n10508), .ZN(n9665) );
  NOR2_X1 U12906 ( .A1(n12946), .A2(n16699), .ZN(n12945) );
  INV_X1 U12907 ( .A(n10173), .ZN(n10172) );
  INV_X1 U12908 ( .A(n10275), .ZN(n10274) );
  NAND2_X1 U12909 ( .A1(n16440), .A2(n16745), .ZN(n10275) );
  AND2_X1 U12910 ( .A1(n10150), .A2(n10149), .ZN(n9666) );
  AND3_X1 U12911 ( .A1(n9969), .A2(n12655), .A3(n10130), .ZN(n9667) );
  NOR2_X1 U12912 ( .A1(n14722), .A2(n10536), .ZN(n14690) );
  NAND2_X1 U12913 ( .A1(n12214), .A2(n12213), .ZN(n14840) );
  AND4_X1 U12914 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n9668) );
  INV_X2 U12915 ( .A(n11555), .ZN(n14545) );
  NAND2_X1 U12916 ( .A1(n14322), .A2(n10415), .ZN(n15720) );
  NAND2_X1 U12917 ( .A1(n14507), .A2(n9660), .ZN(n15055) );
  NAND2_X1 U12918 ( .A1(n11359), .A2(n10352), .ZN(n9669) );
  AND2_X1 U12919 ( .A1(n9623), .A2(n12881), .ZN(n13236) );
  INV_X1 U12920 ( .A(n16858), .ZN(n9867) );
  NAND2_X1 U12921 ( .A1(n12954), .A2(n10401), .ZN(n9670) );
  OR2_X1 U12922 ( .A1(n16738), .A2(n17340), .ZN(n9671) );
  AND2_X1 U12923 ( .A1(n15239), .A2(n15503), .ZN(n9672) );
  AND2_X1 U12924 ( .A1(n10072), .A2(n14658), .ZN(n9673) );
  AND2_X1 U12925 ( .A1(n11973), .A2(n15540), .ZN(n9674) );
  NOR2_X1 U12926 ( .A1(n13058), .A2(n14295), .ZN(n14296) );
  AND2_X1 U12927 ( .A1(n15688), .A2(n9970), .ZN(n9675) );
  AND2_X1 U12928 ( .A1(n12952), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12954) );
  INV_X1 U12929 ( .A(n15220), .ZN(n10453) );
  AND2_X1 U12930 ( .A1(n11256), .A2(n11335), .ZN(n9676) );
  AND4_X1 U12931 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n9677) );
  AND2_X1 U12932 ( .A1(n14604), .A2(n10075), .ZN(n9678) );
  INV_X1 U12933 ( .A(n11831), .ZN(n10049) );
  OAI21_X1 U12934 ( .B1(n17505), .B2(n10301), .A(n10300), .ZN(n17481) );
  AND3_X1 U12935 ( .A1(n10627), .A2(n9892), .A3(n9891), .ZN(n9679) );
  AND2_X1 U12936 ( .A1(n9785), .A2(n16984), .ZN(n9680) );
  NAND2_X1 U12937 ( .A1(n11301), .A2(n9688), .ZN(n11257) );
  AND2_X1 U12938 ( .A1(n12807), .A2(n10414), .ZN(n9681) );
  AND3_X1 U12939 ( .A1(n10908), .A2(n19856), .A3(n20550), .ZN(n9682) );
  NAND2_X1 U12940 ( .A1(n10388), .A2(n10387), .ZN(n9683) );
  INV_X1 U12941 ( .A(n10278), .ZN(n15228) );
  NAND2_X1 U12942 ( .A1(n11370), .A2(n11419), .ZN(n11372) );
  AND2_X1 U12943 ( .A1(n15069), .A2(n12100), .ZN(n9684) );
  AND3_X1 U12944 ( .A1(n10209), .A2(n10208), .A3(n10206), .ZN(n9685) );
  AND2_X1 U12945 ( .A1(n18243), .A2(n10321), .ZN(n9686) );
  AND2_X1 U12946 ( .A1(n13727), .A2(n10169), .ZN(n9687) );
  INV_X1 U12947 ( .A(n15140), .ZN(n9958) );
  AND3_X1 U12948 ( .A1(n10337), .A2(n10338), .A3(n11327), .ZN(n9688) );
  INV_X1 U12949 ( .A(n20799), .ZN(n21012) );
  AND3_X1 U12950 ( .A1(n10971), .A2(n11003), .A3(n10970), .ZN(n9689) );
  INV_X1 U12951 ( .A(n14100), .ZN(n12150) );
  AND2_X1 U12953 ( .A1(n10448), .A2(n13208), .ZN(n9690) );
  AND2_X1 U12954 ( .A1(n15602), .A2(n15603), .ZN(n15590) );
  OR2_X1 U12955 ( .A1(n12643), .A2(n12645), .ZN(n9691) );
  NAND2_X1 U12956 ( .A1(n16629), .A2(n16630), .ZN(n16611) );
  INV_X1 U12957 ( .A(n14722), .ZN(n10531) );
  INV_X1 U12958 ( .A(n10329), .ZN(n16709) );
  AND3_X1 U12959 ( .A1(n12640), .A2(n12639), .A3(n12638), .ZN(n9692) );
  AND2_X1 U12960 ( .A1(n10454), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9693) );
  AND4_X1 U12961 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n9694) );
  OR2_X1 U12962 ( .A1(n14446), .A2(n14445), .ZN(n9695) );
  AND2_X1 U12963 ( .A1(n10306), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9696) );
  INV_X1 U12964 ( .A(n14855), .ZN(n12214) );
  AND2_X1 U12965 ( .A1(n11120), .A2(n9906), .ZN(n9697) );
  OR2_X1 U12966 ( .A1(n9853), .A2(n9852), .ZN(n9698) );
  AND2_X1 U12967 ( .A1(n9942), .A2(n10029), .ZN(n9699) );
  NOR2_X1 U12968 ( .A1(n14395), .A2(n15770), .ZN(n15754) );
  NAND2_X1 U12969 ( .A1(n19856), .A2(n14366), .ZN(n9700) );
  AND2_X1 U12970 ( .A1(n14322), .A2(n14417), .ZN(n14418) );
  INV_X1 U12971 ( .A(n10511), .ZN(n10510) );
  NAND2_X1 U12972 ( .A1(n10512), .A2(n11201), .ZN(n10511) );
  INV_X1 U12973 ( .A(n13679), .ZN(n10061) );
  AND2_X1 U12974 ( .A1(n18807), .A2(n18704), .ZN(n18573) );
  AND2_X1 U12975 ( .A1(n10386), .A2(n10385), .ZN(n9701) );
  INV_X1 U12976 ( .A(n9902), .ZN(n16426) );
  NAND2_X1 U12977 ( .A1(n10392), .A2(n11609), .ZN(n9702) );
  INV_X1 U12978 ( .A(n10460), .ZN(n10459) );
  NAND2_X1 U12979 ( .A1(n10200), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U12980 ( .A1(n14142), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12981 ( .A1(n9671), .A2(n9977), .ZN(n9704) );
  NOR2_X1 U12982 ( .A1(n14618), .A2(n14619), .ZN(n14602) );
  AND2_X1 U12983 ( .A1(n10221), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9705) );
  AND2_X1 U12984 ( .A1(n16548), .A2(n16559), .ZN(n9706) );
  INV_X1 U12985 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16699) );
  OR2_X1 U12986 ( .A1(n13727), .A2(n10169), .ZN(n9707) );
  INV_X1 U12987 ( .A(n10038), .ZN(n10037) );
  NAND2_X1 U12988 ( .A1(n13054), .A2(n12903), .ZN(n10038) );
  AND2_X1 U12989 ( .A1(n14641), .A2(n14620), .ZN(n14605) );
  INV_X1 U12990 ( .A(n10264), .ZN(n10263) );
  NAND2_X1 U12991 ( .A1(n9625), .A2(n10265), .ZN(n10264) );
  NAND2_X1 U12992 ( .A1(n11317), .A2(n17338), .ZN(n11118) );
  INV_X1 U12993 ( .A(n11118), .ZN(n16676) );
  AND3_X1 U12994 ( .A1(n11013), .A2(n11008), .A3(n11011), .ZN(n9708) );
  OR2_X1 U12995 ( .A1(n10701), .A2(n10700), .ZN(n19106) );
  INV_X1 U12996 ( .A(n19106), .ZN(n10214) );
  NAND2_X1 U12997 ( .A1(n19131), .A2(n19111), .ZN(n13624) );
  INV_X1 U12998 ( .A(n13624), .ZN(n10216) );
  AND2_X1 U12999 ( .A1(n20549), .A2(n9700), .ZN(n9709) );
  OR2_X1 U13000 ( .A1(n21734), .A2(n13944), .ZN(n9710) );
  AND3_X1 U13001 ( .A1(n12662), .A2(n10190), .A3(n10187), .ZN(n9711) );
  NAND2_X1 U13002 ( .A1(n10468), .A2(n10466), .ZN(n16429) );
  OR2_X1 U13003 ( .A1(n15186), .A2(n15190), .ZN(n9712) );
  AND2_X1 U13004 ( .A1(n10805), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9713) );
  AND2_X1 U13005 ( .A1(n11387), .A2(n9625), .ZN(n9714) );
  AND2_X1 U13006 ( .A1(n10416), .A2(n12792), .ZN(n9715) );
  NOR2_X1 U13007 ( .A1(n16455), .A2(n16456), .ZN(n9716) );
  AND2_X1 U13008 ( .A1(n10352), .A2(n15712), .ZN(n9717) );
  NOR2_X1 U13009 ( .A1(n10453), .A2(n10449), .ZN(n10448) );
  AND2_X1 U13010 ( .A1(n11555), .A2(n12068), .ZN(n12107) );
  AND2_X1 U13011 ( .A1(n9676), .A2(n10497), .ZN(n9718) );
  AND2_X1 U13012 ( .A1(n15185), .A2(n15188), .ZN(n9854) );
  AND2_X1 U13013 ( .A1(n10909), .A2(n12867), .ZN(n9719) );
  NOR2_X1 U13014 ( .A1(n13085), .A2(n13078), .ZN(n9720) );
  AND2_X1 U13015 ( .A1(n9865), .A2(n9863), .ZN(n9721) );
  NAND2_X1 U13016 ( .A1(n16723), .A2(n17346), .ZN(n9722) );
  AND3_X1 U13017 ( .A1(n12847), .A2(n12846), .A3(n12845), .ZN(n14050) );
  OR2_X1 U13018 ( .A1(n10169), .A2(n10172), .ZN(n9723) );
  INV_X1 U13019 ( .A(n13084), .ZN(n10332) );
  OR2_X1 U13020 ( .A1(n17468), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9724) );
  INV_X1 U13021 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9820) );
  INV_X1 U13022 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20501) );
  INV_X1 U13023 ( .A(n11808), .ZN(n10280) );
  OR2_X1 U13024 ( .A1(n11551), .A2(n21503), .ZN(n10549) );
  INV_X1 U13025 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10732) );
  INV_X2 U13026 ( .A(n16308), .ZN(n16287) );
  INV_X1 U13027 ( .A(n17330), .ZN(n17346) );
  INV_X1 U13028 ( .A(n10202), .ZN(n18801) );
  INV_X1 U13029 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11578) );
  INV_X1 U13030 ( .A(n13024), .ZN(n12854) );
  INV_X2 U13031 ( .A(n13024), .ZN(n13026) );
  NAND2_X1 U13032 ( .A1(n12736), .A2(n12735), .ZN(n13551) );
  NAND2_X1 U13033 ( .A1(n13551), .A2(n13550), .ZN(n13549) );
  INV_X1 U13034 ( .A(n20967), .ZN(n10062) );
  NOR2_X1 U13035 ( .A1(n15848), .A2(n10513), .ZN(n13057) );
  INV_X1 U13036 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13037 ( .A1(n12808), .A2(n12807), .ZN(n13061) );
  NOR2_X1 U13038 ( .A1(n12967), .A2(n16562), .ZN(n12968) );
  NOR2_X1 U13039 ( .A1(n14703), .A2(n14692), .ZN(n14680) );
  AND2_X1 U13040 ( .A1(n15541), .A2(n10424), .ZN(n14879) );
  NAND2_X1 U13041 ( .A1(n12009), .A2(n12008), .ZN(n14748) );
  AND2_X1 U13042 ( .A1(n18597), .A2(n10297), .ZN(n9725) );
  NAND2_X1 U13043 ( .A1(n12161), .A2(n12160), .ZN(n14875) );
  NAND2_X1 U13044 ( .A1(n9618), .A2(n13244), .ZN(n15899) );
  OR2_X1 U13045 ( .A1(n12967), .A2(n10407), .ZN(n9726) );
  NAND2_X1 U13046 ( .A1(n12916), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12977) );
  AND2_X1 U13047 ( .A1(n16974), .A2(n10112), .ZN(n9727) );
  AND2_X1 U13048 ( .A1(n12008), .A2(n10430), .ZN(n9728) );
  AND2_X1 U13049 ( .A1(n10519), .A2(n10518), .ZN(n9729) );
  AND2_X1 U13050 ( .A1(n9729), .A2(n9971), .ZN(n9730) );
  NOR2_X1 U13051 ( .A1(n15848), .A2(n10516), .ZN(n13278) );
  AND2_X1 U13052 ( .A1(n11991), .A2(n10427), .ZN(n14782) );
  AND2_X1 U13053 ( .A1(n10249), .A2(n10248), .ZN(n9731) );
  NAND2_X1 U13054 ( .A1(n12808), .A2(n10413), .ZN(n14024) );
  AND2_X1 U13055 ( .A1(n11295), .A2(n11307), .ZN(n11301) );
  INV_X1 U13056 ( .A(n11301), .ZN(n10340) );
  AND2_X1 U13057 ( .A1(n9730), .A2(n15630), .ZN(n9732) );
  NAND2_X1 U13058 ( .A1(n13996), .A2(n12131), .ZN(n14032) );
  AND2_X1 U13059 ( .A1(n12917), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12916) );
  AND2_X1 U13060 ( .A1(n14680), .A2(n14681), .ZN(n14659) );
  AND2_X1 U13061 ( .A1(n12859), .A2(n10116), .ZN(n9733) );
  AND2_X1 U13062 ( .A1(n14879), .A2(n14880), .ZN(n14864) );
  AND2_X1 U13063 ( .A1(n10396), .A2(n10250), .ZN(n9734) );
  AND2_X1 U13064 ( .A1(n9728), .A2(n10429), .ZN(n9735) );
  AND2_X1 U13065 ( .A1(n12954), .A2(n9645), .ZN(n12962) );
  NAND2_X1 U13066 ( .A1(n15541), .A2(n15540), .ZN(n14931) );
  INV_X1 U13067 ( .A(n11369), .ZN(n10496) );
  AND2_X1 U13068 ( .A1(n16978), .A2(n12888), .ZN(n16967) );
  INV_X1 U13069 ( .A(n16630), .ZN(n10266) );
  NAND2_X1 U13070 ( .A1(n10395), .A2(n16014), .ZN(n16260) );
  NAND2_X1 U13071 ( .A1(n18597), .A2(n9642), .ZN(n10577) );
  INV_X1 U13072 ( .A(n11327), .ZN(n10341) );
  AND2_X1 U13073 ( .A1(n10428), .A2(n11990), .ZN(n9736) );
  NAND2_X1 U13074 ( .A1(n20559), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13735) );
  OR2_X1 U13075 ( .A1(n10714), .A2(n10713), .ZN(n19102) );
  INV_X1 U13076 ( .A(n19102), .ZN(n19681) );
  NAND2_X1 U13077 ( .A1(n11769), .A2(n21584), .ZN(n9737) );
  OR2_X1 U13078 ( .A1(n17261), .A2(n17260), .ZN(n9738) );
  AND2_X1 U13079 ( .A1(n10421), .A2(n10418), .ZN(n9739) );
  AND2_X1 U13080 ( .A1(n9734), .A2(n16271), .ZN(n9740) );
  INV_X1 U13081 ( .A(n10198), .ZN(n10197) );
  NAND2_X1 U13082 ( .A1(n16850), .A2(n16851), .ZN(n10198) );
  INV_X1 U13083 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17478) );
  INV_X1 U13084 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12960) );
  AND2_X1 U13085 ( .A1(n11038), .A2(n9650), .ZN(n9741) );
  NAND2_X1 U13086 ( .A1(n14296), .A2(n9974), .ZN(n12672) );
  INV_X1 U13087 ( .A(n10349), .ZN(n10348) );
  OR2_X1 U13088 ( .A1(n11274), .A2(n10350), .ZN(n10349) );
  INV_X1 U13089 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20559) );
  INV_X1 U13090 ( .A(n14732), .ZN(n12349) );
  AND2_X1 U13091 ( .A1(n12348), .A2(n12347), .ZN(n14732) );
  INV_X1 U13092 ( .A(n10231), .ZN(n10230) );
  NAND2_X1 U13093 ( .A1(n14016), .A2(n10232), .ZN(n10231) );
  OR2_X1 U13094 ( .A1(n11050), .A2(n11049), .ZN(n11252) );
  INV_X1 U13095 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16562) );
  INV_X1 U13096 ( .A(n11277), .ZN(n10350) );
  AND2_X1 U13097 ( .A1(n13040), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17055) );
  AND2_X1 U13098 ( .A1(n10523), .A2(n15615), .ZN(n9742) );
  AND2_X1 U13099 ( .A1(n10434), .A2(n10433), .ZN(n9743) );
  AND2_X1 U13100 ( .A1(n10528), .A2(n14747), .ZN(n9744) );
  AND2_X1 U13101 ( .A1(n9733), .A2(n15692), .ZN(n9745) );
  AND2_X1 U13102 ( .A1(n10120), .A2(n9739), .ZN(n9746) );
  AND2_X1 U13103 ( .A1(n9642), .A2(n10296), .ZN(n9747) );
  AND2_X1 U13104 ( .A1(n9735), .A2(n14724), .ZN(n9748) );
  AND2_X1 U13105 ( .A1(n10415), .A2(n12857), .ZN(n9749) );
  INV_X1 U13106 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15663) );
  INV_X1 U13107 ( .A(n18184), .ZN(n18270) );
  INV_X1 U13108 ( .A(n18270), .ZN(n18266) );
  INV_X1 U13109 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10298) );
  INV_X1 U13110 ( .A(n19513), .ZN(n10204) );
  INV_X1 U13111 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10797) );
  INV_X1 U13112 ( .A(n17493), .ZN(n10302) );
  INV_X1 U13113 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10497) );
  NOR2_X2 U13114 ( .A1(n19708), .A2(n16235), .ZN(n16713) );
  INV_X1 U13115 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10299) );
  INV_X1 U13116 ( .A(n17215), .ZN(n18394) );
  AND2_X1 U13117 ( .A1(n17935), .A2(n10319), .ZN(n9750) );
  NOR3_X1 U13118 ( .A1(n12993), .A2(n12992), .A3(n12996), .ZN(n12997) );
  OR2_X1 U13119 ( .A1(n12993), .A2(n12992), .ZN(n9751) );
  NOR2_X1 U13120 ( .A1(n12993), .A2(n10403), .ZN(n13000) );
  AND2_X1 U13121 ( .A1(n18523), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14477) );
  INV_X1 U13122 ( .A(n10612), .ZN(n13651) );
  INV_X1 U13123 ( .A(n16520), .ZN(n10398) );
  AND2_X1 U13124 ( .A1(n10437), .A2(n10436), .ZN(n9752) );
  INV_X1 U13125 ( .A(n18663), .ZN(n18644) );
  AND2_X1 U13126 ( .A1(n10498), .A2(n16240), .ZN(n9753) );
  AND2_X1 U13127 ( .A1(n18243), .A2(n10322), .ZN(n9754) );
  NAND2_X1 U13128 ( .A1(n13014), .A2(n13013), .ZN(n9755) );
  OR2_X1 U13129 ( .A1(n14426), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9756) );
  AND2_X1 U13130 ( .A1(n14477), .A2(n9619), .ZN(n9757) );
  AND2_X1 U13131 ( .A1(n10295), .A2(n17748), .ZN(n9758) );
  AND2_X1 U13132 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9759) );
  AND2_X1 U13133 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n9760) );
  INV_X2 U13134 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21501) );
  NAND2_X2 U13135 ( .A1(n19702), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20477) );
  INV_X1 U13136 ( .A(n19075), .ZN(n19022) );
  NAND2_X1 U13137 ( .A1(n10608), .A2(n13609), .ZN(n9761) );
  NOR2_X1 U13138 ( .A1(n17126), .A2(n18753), .ZN(n17149) );
  INV_X1 U13139 ( .A(n18790), .ZN(n9899) );
  INV_X1 U13140 ( .A(n20796), .ZN(n20798) );
  AND3_X1 U13141 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17724) );
  INV_X1 U13142 ( .A(n15067), .ZN(n10455) );
  AND2_X1 U13143 ( .A1(n10526), .A2(n10561), .ZN(n9762) );
  OR2_X1 U13144 ( .A1(n11851), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9763) );
  NAND2_X1 U13145 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17745) );
  AND2_X1 U13146 ( .A1(n11843), .A2(n11842), .ZN(n9764) );
  AND3_X1 U13147 ( .A1(n11847), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9765) );
  AND2_X1 U13148 ( .A1(n16782), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U13149 ( .A1(n16450), .A2(n16451), .ZN(n9767) );
  AND2_X1 U13150 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9768) );
  INV_X1 U13151 ( .A(n11426), .ZN(n10471) );
  AND2_X1 U13152 ( .A1(n10526), .A2(n9657), .ZN(n9769) );
  AND2_X1 U13153 ( .A1(n9656), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U13154 ( .A1(n9764), .A2(n10389), .ZN(n9771) );
  AND2_X1 U13155 ( .A1(n9762), .A2(n9903), .ZN(n9772) );
  INV_X1 U13156 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17338) );
  INV_X1 U13157 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18431) );
  INV_X1 U13158 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n9868) );
  INV_X1 U13159 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10136) );
  INV_X1 U13160 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n9870) );
  AND2_X1 U13161 ( .A1(n10464), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9773) );
  INV_X1 U13162 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17756) );
  INV_X1 U13163 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10358) );
  NOR2_X1 U13164 ( .A1(n16914), .A2(n16919), .ZN(n10464) );
  AND2_X1 U13165 ( .A1(n10326), .A2(n16782), .ZN(n9774) );
  AND2_X1 U13166 ( .A1(n16525), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9775) );
  AND2_X1 U13167 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n9776) );
  INV_X1 U13168 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16861) );
  INV_X1 U13169 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9814) );
  NAND2_X1 U13170 ( .A1(n16861), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9777) );
  OAI211_X1 U13171 ( .C1(n16733), .C2(n17348), .A(n10186), .B(n10183), .ZN(
        P2_U3017) );
  OAI21_X1 U13172 ( .B1(n16816), .B2(n17348), .A(n10012), .ZN(n10011) );
  INV_X1 U13173 ( .A(n17348), .ZN(n16984) );
  INV_X1 U13174 ( .A(n21466), .ZN(n9778) );
  INV_X1 U13175 ( .A(n9778), .ZN(n9779) );
  AOI22_X2 U13176 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9584), .B1(DATAI_27_), 
        .B2(n9613), .ZN(n21399) );
  INV_X1 U13177 ( .A(n19061), .ZN(n9887) );
  NAND4_X1 U13178 ( .A1(n9781), .A2(n11120), .A3(n11112), .A4(n11118), .ZN(
        n9794) );
  INV_X1 U13179 ( .A(n11114), .ZN(n11116) );
  NAND3_X2 U13180 ( .A1(n9689), .A2(n9635), .A3(n9861), .ZN(n9932) );
  NAND2_X1 U13181 ( .A1(n9980), .A2(n10502), .ZN(n16567) );
  NAND2_X1 U13182 ( .A1(n9787), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10915) );
  NAND2_X1 U13183 ( .A1(n9787), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10934) );
  AOI21_X1 U13184 ( .B1(n9787), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10949), .ZN(n10952) );
  NAND2_X1 U13185 ( .A1(n16667), .A2(n9788), .ZN(n16653) );
  OAI21_X1 U13186 ( .B1(n16609), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n9789), .ZN(n16929) );
  NAND2_X1 U13187 ( .A1(n16608), .A2(n9790), .ZN(P2_U3003) );
  NAND2_X1 U13188 ( .A1(n9792), .A2(n11113), .ZN(n16666) );
  NAND4_X1 U13189 ( .A1(n10140), .A2(n11119), .A3(n9794), .A4(n9793), .ZN(
        n9792) );
  NAND3_X1 U13190 ( .A1(n11110), .A2(n9927), .A3(n10141), .ZN(n9793) );
  AOI22_X1 U13191 ( .A1(n11053), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n20234), .ZN(n11078) );
  AND2_X4 U13192 ( .A1(n9666), .A2(n9796), .ZN(n9980) );
  OAI21_X1 U13193 ( .B1(n16703), .B2(n9797), .A(n16702), .ZN(n16985) );
  NAND2_X1 U13194 ( .A1(n20234), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10964) );
  NAND2_X1 U13195 ( .A1(n20234), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9798) );
  NOR2_X2 U13196 ( .A1(n14022), .A2(n10963), .ZN(n20234) );
  NAND2_X1 U13197 ( .A1(n9934), .A2(n11038), .ZN(n11099) );
  AND2_X2 U13198 ( .A1(n10912), .A2(n12867), .ZN(n9996) );
  NAND2_X1 U13199 ( .A1(n13154), .A2(n16984), .ZN(n13153) );
  INV_X2 U13200 ( .A(n10911), .ZN(n12660) );
  AND3_X4 U13201 ( .A1(n14348), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16202) );
  NAND4_X1 U13202 ( .A1(n9713), .A2(n10808), .A3(n10806), .A4(n10807), .ZN(
        n9804) );
  NAND2_X1 U13203 ( .A1(n10802), .A2(n10800), .ZN(n9805) );
  NAND3_X1 U13204 ( .A1(n10801), .A2(n10803), .A3(n14341), .ZN(n9806) );
  NAND3_X1 U13205 ( .A1(n9810), .A2(n9716), .A3(n9807), .ZN(P2_U2987) );
  OR2_X1 U13206 ( .A1(n16751), .A2(n16707), .ZN(n9807) );
  NOR2_X2 U13207 ( .A1(n14010), .A2(n10963), .ZN(n17022) );
  INV_X2 U13208 ( .A(n10962), .ZN(n14010) );
  NAND3_X1 U13209 ( .A1(n11325), .A2(n11324), .A3(n9817), .ZN(n9816) );
  NOR2_X1 U13210 ( .A1(n11322), .A2(n16690), .ZN(n9817) );
  OAI21_X1 U13211 ( .B1(n10465), .B2(n10090), .A(n13138), .ZN(n9818) );
  INV_X1 U13212 ( .A(n11347), .ZN(n9819) );
  AND2_X2 U13213 ( .A1(n14060), .A2(n13594), .ZN(n11611) );
  NOR2_X4 U13214 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14060) );
  NOR2_X2 U13215 ( .A1(n20819), .A2(n20824), .ZN(n13684) );
  AND2_X2 U13216 ( .A1(n11852), .A2(n10195), .ZN(n14492) );
  NAND3_X1 U13217 ( .A1(n9957), .A2(n9960), .A3(n9765), .ZN(n9825) );
  NAND3_X1 U13218 ( .A1(n9957), .A2(n9960), .A3(n9829), .ZN(n9828) );
  NAND3_X2 U13219 ( .A1(n11672), .A2(n21501), .A3(n20854), .ZN(n10392) );
  NAND2_X1 U13220 ( .A1(n11593), .A2(n11594), .ZN(n20854) );
  NAND2_X2 U13221 ( .A1(n9831), .A2(n10124), .ZN(n11672) );
  NAND2_X4 U13222 ( .A1(n11814), .A2(n11826), .ZN(n15239) );
  OAI21_X1 U13223 ( .B1(n13577), .B2(n10286), .A(n9836), .ZN(n9835) );
  XNOR2_X1 U13224 ( .A(n11733), .B(n9836), .ZN(n12106) );
  NAND3_X1 U13225 ( .A1(n9952), .A2(n15154), .A3(n15149), .ZN(n10388) );
  OR2_X2 U13226 ( .A1(n15283), .A2(n10451), .ZN(n10160) );
  NAND2_X2 U13227 ( .A1(n15291), .A2(n10153), .ZN(n20776) );
  NAND2_X1 U13228 ( .A1(n20550), .A2(n10916), .ZN(n10920) );
  XNOR2_X2 U13229 ( .A(n11100), .B(n12723), .ZN(n11114) );
  NAND3_X2 U13230 ( .A1(n9934), .A2(n9933), .A3(n9932), .ZN(n11100) );
  NOR2_X1 U13231 ( .A1(n19875), .A2(n20559), .ZN(n13421) );
  NAND2_X1 U13232 ( .A1(n19875), .A2(n12656), .ZN(n9999) );
  NAND2_X1 U13233 ( .A1(n11246), .A2(n19875), .ZN(n10909) );
  NAND2_X4 U13234 ( .A1(n9928), .A2(n9930), .ZN(n19875) );
  NAND3_X1 U13235 ( .A1(n9862), .A2(n16830), .A3(n16984), .ZN(n16831) );
  NAND3_X1 U13236 ( .A1(n9862), .A2(n16830), .A3(n16704), .ZN(n16522) );
  NAND3_X1 U13237 ( .A1(n9721), .A2(n10374), .A3(n10373), .ZN(P2_U3030) );
  NAND2_X1 U13238 ( .A1(n16556), .A2(n9866), .ZN(n9865) );
  NOR2_X1 U13239 ( .A1(n18750), .A2(n14176), .ZN(n9881) );
  NOR2_X1 U13240 ( .A1(n14176), .A2(n9877), .ZN(n9876) );
  INV_X1 U13241 ( .A(n18750), .ZN(n9878) );
  OR2_X1 U13242 ( .A1(n9881), .A2(n14178), .ZN(n18734) );
  INV_X1 U13243 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9882) );
  INV_X2 U13244 ( .A(n9889), .ZN(n17260) );
  OR2_X2 U13245 ( .A1(n10633), .A2(n9890), .ZN(n9889) );
  INV_X1 U13246 ( .A(n10731), .ZN(n10365) );
  OR2_X2 U13247 ( .A1(n18730), .A2(n18573), .ZN(n18813) );
  AND2_X2 U13248 ( .A1(n18817), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18730) );
  INV_X1 U13249 ( .A(n11100), .ZN(n10094) );
  NAND3_X1 U13250 ( .A1(n9998), .A2(n12685), .A3(n9901), .ZN(n9997) );
  NAND2_X1 U13251 ( .A1(n9980), .A2(n9772), .ZN(n9902) );
  INV_X1 U13252 ( .A(n13130), .ZN(n13131) );
  NAND2_X1 U13253 ( .A1(n9982), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9904) );
  NAND2_X1 U13254 ( .A1(n9981), .A2(n14341), .ZN(n9905) );
  NAND2_X1 U13255 ( .A1(n16676), .A2(n11119), .ZN(n9906) );
  NAND4_X1 U13256 ( .A1(n10878), .A2(n10879), .A3(n10880), .A4(n10877), .ZN(
        n9908) );
  NAND4_X1 U13257 ( .A1(n10875), .A2(n10874), .A3(n10872), .A4(n10873), .ZN(
        n9909) );
  NAND2_X1 U13258 ( .A1(n16844), .A2(n12885), .ZN(n9919) );
  AND3_X1 U13259 ( .A1(n9719), .A2(n10908), .A3(n9926), .ZN(n12865) );
  NAND4_X1 U13260 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n9929) );
  NAND4_X1 U13261 ( .A1(n10843), .A2(n10845), .A3(n10844), .A4(n10842), .ZN(
        n9931) );
  OAI21_X1 U13262 ( .B1(n9936), .B2(n16722), .A(n16537), .ZN(P2_U2996) );
  OAI21_X1 U13263 ( .B1(n9936), .B2(n17348), .A(n16843), .ZN(P2_U3028) );
  NAND2_X1 U13264 ( .A1(n16528), .A2(n16527), .ZN(n9936) );
  OAI21_X1 U13265 ( .B1(n16458), .B2(n9937), .A(n13161), .ZN(P2_U2989) );
  NAND2_X1 U13266 ( .A1(n13154), .A2(n16704), .ZN(n9937) );
  NAND3_X1 U13267 ( .A1(n9968), .A2(n10938), .A3(n10146), .ZN(n9941) );
  NAND2_X1 U13268 ( .A1(n9633), .A2(n9694), .ZN(n9942) );
  NOR2_X1 U13269 ( .A1(n18794), .A2(n13943), .ZN(n18783) );
  AND2_X2 U13270 ( .A1(n18724), .A2(n17065), .ZN(n18637) );
  NAND2_X1 U13271 ( .A1(n16494), .A2(n16492), .ZN(n13136) );
  NAND3_X1 U13272 ( .A1(n10465), .A2(n9946), .A3(n11410), .ZN(n16494) );
  NAND3_X1 U13273 ( .A1(n9714), .A2(n16670), .A3(n16671), .ZN(n9946) );
  XNOR2_X2 U13274 ( .A(n11577), .B(n11667), .ZN(n11594) );
  NAND2_X1 U13275 ( .A1(n15258), .A2(n9950), .ZN(n9948) );
  INV_X1 U13276 ( .A(n15149), .ZN(n9949) );
  NAND2_X2 U13277 ( .A1(n9949), .A2(n9596), .ZN(n9960) );
  NAND2_X1 U13278 ( .A1(n15153), .A2(n11839), .ZN(n9959) );
  OAI21_X1 U13279 ( .B1(n16780), .B2(n17348), .A(n9966), .ZN(P2_U3022) );
  INV_X1 U13280 ( .A(n10256), .ZN(n10253) );
  NAND2_X1 U13281 ( .A1(n9969), .A2(n10912), .ZN(n10901) );
  NAND3_X1 U13282 ( .A1(n9996), .A2(n12870), .A3(n9969), .ZN(n12873) );
  NAND3_X1 U13283 ( .A1(n11152), .A2(n11162), .A3(n9976), .ZN(n14291) );
  NAND2_X1 U13284 ( .A1(n9646), .A2(n11162), .ZN(n14209) );
  NAND2_X1 U13285 ( .A1(n9980), .A2(n10526), .ZN(n10258) );
  NAND2_X1 U13286 ( .A1(n9980), .A2(n9769), .ZN(n16457) );
  OAI21_X1 U13287 ( .B1(n9980), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16626), .ZN(n16941) );
  NAND2_X1 U13288 ( .A1(n9980), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16626) );
  NAND4_X1 U13289 ( .A1(n10827), .A2(n10826), .A3(n10829), .A4(n10828), .ZN(
        n9981) );
  NAND4_X1 U13290 ( .A1(n10832), .A2(n10833), .A3(n10831), .A4(n10830), .ZN(
        n9982) );
  NAND2_X1 U13291 ( .A1(n11054), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n9986) );
  NAND3_X1 U13292 ( .A1(n16860), .A2(n10002), .A3(n10001), .ZN(P2_U3029) );
  INV_X1 U13293 ( .A(n10016), .ZN(n10015) );
  OAI21_X1 U13294 ( .B1(n14442), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10018), .ZN(n10017) );
  MUX2_X1 U13295 ( .A(n17060), .B(n18663), .S(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n10018) );
  OR2_X1 U13296 ( .A1(n14442), .A2(n9620), .ZN(n10019) );
  NOR2_X1 U13297 ( .A1(n17061), .A2(n18644), .ZN(n14442) );
  INV_X1 U13298 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U13299 ( .A1(n10027), .A2(n13974), .ZN(n10024) );
  INV_X1 U13300 ( .A(n10026), .ZN(n10025) );
  NOR2_X1 U13301 ( .A1(n10375), .A2(n21719), .ZN(n10027) );
  XNOR2_X2 U13302 ( .A(n14123), .B(n14121), .ZN(n13974) );
  AND3_X2 U13303 ( .A1(n18626), .A2(n10028), .A3(n14435), .ZN(n18542) );
  NAND3_X1 U13304 ( .A1(n10379), .A2(n14434), .A3(n10381), .ZN(n14435) );
  NAND2_X2 U13305 ( .A1(n18556), .A2(n9659), .ZN(n18626) );
  INV_X1 U13306 ( .A(n11229), .ZN(n11157) );
  NAND3_X1 U13307 ( .A1(n11734), .A2(n11743), .A3(n10042), .ZN(n10041) );
  NAND2_X1 U13308 ( .A1(n10045), .A2(n9737), .ZN(n11784) );
  OR2_X2 U13309 ( .A1(n13580), .A2(n12015), .ZN(n13176) );
  NAND3_X1 U13310 ( .A1(n10196), .A2(n15069), .A3(n10448), .ZN(n10052) );
  AND2_X1 U13311 ( .A1(n11928), .A2(n10054), .ZN(n12083) );
  NAND2_X1 U13312 ( .A1(n10055), .A2(n11561), .ZN(n11929) );
  NAND2_X2 U13313 ( .A1(n11672), .A2(n11671), .ZN(n13680) );
  NAND2_X1 U13314 ( .A1(n10057), .A2(n11672), .ZN(n10056) );
  NOR2_X2 U13315 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U13316 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11481) );
  AND2_X1 U13317 ( .A1(n15185), .A2(n10063), .ZN(n15153) );
  XNOR2_X1 U13318 ( .A(n15203), .B(n10066), .ZN(n15458) );
  OAI21_X1 U13319 ( .B1(n15312), .B2(n20574), .A(n15066), .ZN(P1_U2972) );
  NAND3_X1 U13320 ( .A1(n11743), .A2(n11734), .A3(n10390), .ZN(n11801) );
  OR2_X1 U13321 ( .A1(n15055), .A2(n20797), .ZN(n10068) );
  NAND2_X1 U13322 ( .A1(n10073), .A2(n12151), .ZN(n14855) );
  NAND2_X1 U13323 ( .A1(n10929), .A2(n10928), .ZN(n10930) );
  NAND2_X2 U13324 ( .A1(n10193), .A2(n10943), .ZN(n10077) );
  AOI21_X4 U13325 ( .B1(n11576), .B2(n11942), .A(n21501), .ZN(n11667) );
  NAND2_X1 U13326 ( .A1(n10477), .A2(n10481), .ZN(n16513) );
  INV_X1 U13327 ( .A(n14437), .ZN(n18526) );
  NAND2_X1 U13328 ( .A1(n18526), .A2(n18818), .ZN(n18525) );
  NAND2_X1 U13329 ( .A1(n10904), .A2(n10917), .ZN(n10911) );
  OR2_X2 U13330 ( .A1(n15743), .A2(n16534), .ZN(n15726) );
  NOR2_X2 U13331 ( .A1(n15895), .A2(n16696), .ZN(n15882) );
  NOR2_X2 U13332 ( .A1(n15786), .A2(n10543), .ZN(n15771) );
  NOR2_X2 U13333 ( .A1(n13268), .A2(n16606), .ZN(n15817) );
  NOR2_X2 U13334 ( .A1(n15858), .A2(n15860), .ZN(n15841) );
  NAND2_X1 U13335 ( .A1(n12982), .A2(n16498), .ZN(n15678) );
  NAND2_X1 U13336 ( .A1(n13004), .A2(n16435), .ZN(n13091) );
  NAND2_X1 U13337 ( .A1(n12995), .A2(n16465), .ZN(n15620) );
  NAND2_X1 U13338 ( .A1(n13002), .A2(n16445), .ZN(n15595) );
  NAND2_X1 U13339 ( .A1(n12988), .A2(n16480), .ZN(n15645) );
  NAND2_X1 U13340 ( .A1(n10399), .A2(n19733), .ZN(n15709) );
  NAND2_X1 U13341 ( .A1(n10194), .A2(n10930), .ZN(n10193) );
  INV_X1 U13342 ( .A(n16820), .ZN(n10252) );
  NAND2_X1 U13343 ( .A1(n10252), .A2(n17351), .ZN(n10251) );
  OAI21_X1 U13344 ( .B1(n10451), .B2(n15282), .A(n11780), .ZN(n10125) );
  NAND2_X1 U13345 ( .A1(n11681), .A2(n11680), .ZN(n10282) );
  XNOR2_X2 U13346 ( .A(n10077), .B(n10953), .ZN(n10975) );
  NAND3_X1 U13347 ( .A1(n13133), .A2(n13135), .A3(n13134), .ZN(P2_U3016) );
  NAND4_X1 U13348 ( .A1(n10931), .A2(n10545), .A3(n12654), .A4(n14385), .ZN(
        n10078) );
  XNOR2_X2 U13349 ( .A(n11150), .B(n9661), .ZN(n10962) );
  NAND2_X1 U13350 ( .A1(n16429), .A2(n10086), .ZN(n10085) );
  AND2_X1 U13351 ( .A1(n11434), .A2(n16431), .ZN(n10086) );
  NAND2_X1 U13352 ( .A1(n10260), .A2(n16492), .ZN(n10092) );
  NOR2_X1 U13353 ( .A1(n14105), .A2(n10093), .ZN(n14347) );
  NOR2_X1 U13354 ( .A1(n10182), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12688) );
  AND2_X1 U13355 ( .A1(n9996), .A2(n10130), .ZN(n12872) );
  AND2_X2 U13356 ( .A1(n10930), .A2(n10943), .ZN(n10958) );
  INV_X1 U13357 ( .A(n13088), .ZN(n10096) );
  NAND2_X1 U13358 ( .A1(n10096), .A2(n9720), .ZN(n10103) );
  NAND3_X1 U13359 ( .A1(n10097), .A2(n13090), .A3(n10107), .ZN(P2_U2983) );
  NAND3_X1 U13360 ( .A1(n10103), .A2(n10102), .A3(n10333), .ZN(n10097) );
  NAND3_X1 U13361 ( .A1(n10101), .A2(n10104), .A3(n10098), .ZN(n13175) );
  NAND3_X1 U13362 ( .A1(n10101), .A2(n10099), .A3(n10098), .ZN(n10107) );
  AND3_X2 U13363 ( .A1(n10103), .A2(n10333), .A3(n10332), .ZN(n13172) );
  INV_X1 U13364 ( .A(n10111), .ZN(n16757) );
  NAND3_X1 U13365 ( .A1(n12671), .A2(n13490), .A3(n12653), .ZN(n10113) );
  NAND2_X1 U13366 ( .A1(n12860), .A2(n9745), .ZN(n15673) );
  INV_X1 U13367 ( .A(n15673), .ZN(n13015) );
  NAND2_X1 U13368 ( .A1(n12808), .A2(n10117), .ZN(n14049) );
  INV_X2 U13369 ( .A(n13270), .ZN(n12808) );
  NAND3_X1 U13370 ( .A1(n9618), .A2(n10119), .A3(n13244), .ZN(n15884) );
  NAND2_X1 U13371 ( .A1(n13144), .A2(n10120), .ZN(n15617) );
  NAND2_X1 U13372 ( .A1(n13144), .A2(n9746), .ZN(n13095) );
  NAND3_X1 U13373 ( .A1(n10185), .A2(n10123), .A3(n9722), .ZN(n10122) );
  NAND2_X1 U13374 ( .A1(n20930), .A2(n10124), .ZN(n21235) );
  INV_X1 U13375 ( .A(n10125), .ZN(n10279) );
  OAI21_X1 U13376 ( .B1(n10450), .B2(n10125), .A(n11785), .ZN(n15266) );
  AND2_X1 U13377 ( .A1(n10127), .A2(n9643), .ZN(n10126) );
  NAND2_X2 U13378 ( .A1(n15058), .A2(n15107), .ZN(n15046) );
  NOR2_X2 U13379 ( .A1(n10256), .A2(n10255), .ZN(n12864) );
  NAND3_X1 U13380 ( .A1(n11101), .A2(n16708), .A3(n11100), .ZN(n10131) );
  NAND2_X1 U13381 ( .A1(n16676), .A2(n10141), .ZN(n10140) );
  NAND2_X1 U13382 ( .A1(n10143), .A2(n10148), .ZN(n10147) );
  NAND3_X1 U13383 ( .A1(n10143), .A2(n10142), .A3(n10148), .ZN(n10948) );
  NAND2_X1 U13384 ( .A1(n10147), .A2(n10145), .ZN(n10144) );
  NAND3_X1 U13385 ( .A1(n11146), .A2(n10458), .A3(n10460), .ZN(n10149) );
  NAND2_X1 U13386 ( .A1(n10457), .A2(n11146), .ZN(n10150) );
  OAI21_X1 U13387 ( .B1(n16653), .B2(n10459), .A(n10152), .ZN(n16646) );
  NOR2_X1 U13388 ( .A1(n15291), .A2(n10153), .ZN(n20771) );
  NAND2_X1 U13389 ( .A1(n11568), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U13390 ( .A1(n10154), .A2(n11571), .ZN(n11577) );
  NAND2_X1 U13391 ( .A1(n11568), .A2(n10155), .ZN(n10154) );
  NAND3_X1 U13392 ( .A1(n10279), .A2(n10160), .A3(n11808), .ZN(n10156) );
  INV_X1 U13393 ( .A(n10160), .ZN(n10450) );
  OAI21_X1 U13394 ( .B1(n11785), .B2(n10280), .A(n11810), .ZN(n10158) );
  INV_X1 U13395 ( .A(n13727), .ZN(n10170) );
  NOR2_X1 U13396 ( .A1(n13727), .A2(n9723), .ZN(n10165) );
  NAND2_X1 U13397 ( .A1(n10179), .A2(n10177), .ZN(n10278) );
  NAND2_X1 U13398 ( .A1(n10182), .A2(n20501), .ZN(n13024) );
  NAND2_X1 U13399 ( .A1(n10182), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12693) );
  NAND2_X1 U13400 ( .A1(n10182), .A2(n12867), .ZN(n10905) );
  AOI21_X1 U13401 ( .B1(n10916), .B2(n10893), .A(n10181), .ZN(n10180) );
  NAND2_X2 U13402 ( .A1(n10283), .A2(n11732), .ZN(n11743) );
  NAND2_X1 U13403 ( .A1(n10191), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16629) );
  OAI21_X1 U13404 ( .B1(n10191), .B2(n10266), .A(n10263), .ZN(n10369) );
  OAI21_X1 U13405 ( .B1(n10191), .B2(n10262), .A(n10261), .ZN(n11347) );
  NAND2_X1 U13406 ( .A1(n10955), .A2(n10954), .ZN(n10194) );
  NAND2_X1 U13407 ( .A1(n10955), .A2(n10954), .ZN(n10259) );
  INV_X1 U13408 ( .A(n10917), .ZN(n10903) );
  NAND2_X1 U13409 ( .A1(n10916), .A2(n10917), .ZN(n10918) );
  NAND2_X2 U13410 ( .A1(n10202), .A2(n18394), .ZN(n18696) );
  NOR2_X2 U13411 ( .A1(n17451), .A2(n19681), .ZN(n10202) );
  NAND3_X1 U13412 ( .A1(n10216), .A2(n10728), .A3(n10213), .ZN(n10212) );
  NAND2_X1 U13413 ( .A1(n10903), .A2(n10909), .ZN(n12657) );
  NAND2_X1 U13414 ( .A1(n10903), .A2(n10217), .ZN(n10900) );
  NAND2_X1 U13415 ( .A1(n14008), .A2(n14007), .ZN(n10224) );
  INV_X1 U13416 ( .A(n14007), .ZN(n10225) );
  NAND2_X1 U13417 ( .A1(n16247), .A2(n10235), .ZN(n10234) );
  OAI211_X1 U13418 ( .C1(n16247), .C2(n10248), .A(n10246), .B(n10239), .ZN(
        n16232) );
  NAND2_X1 U13419 ( .A1(n16247), .A2(n10245), .ZN(n10239) );
  INV_X1 U13420 ( .A(n10246), .ZN(n10241) );
  AND2_X1 U13421 ( .A1(n16243), .A2(n16234), .ZN(n10242) );
  NOR2_X1 U13422 ( .A1(n10247), .A2(n16119), .ZN(n10245) );
  NAND2_X1 U13423 ( .A1(n10247), .A2(n16119), .ZN(n10246) );
  INV_X1 U13424 ( .A(n16079), .ZN(n10247) );
  INV_X1 U13425 ( .A(n16119), .ZN(n10248) );
  NAND2_X1 U13426 ( .A1(n16819), .A2(n10251), .ZN(P2_U3025) );
  NAND2_X1 U13427 ( .A1(n10254), .A2(n12654), .ZN(n12679) );
  NAND2_X1 U13428 ( .A1(n12660), .A2(n17030), .ZN(n10254) );
  NAND2_X1 U13429 ( .A1(n10976), .A2(n10259), .ZN(n13425) );
  AND2_X2 U13430 ( .A1(n10985), .A2(n14010), .ZN(n20139) );
  OAI211_X1 U13431 ( .C1(n16441), .C2(n10273), .A(n10267), .B(n10269), .ZN(
        n16742) );
  NAND3_X1 U13432 ( .A1(n16441), .A2(n10268), .A3(n10276), .ZN(n10267) );
  INV_X1 U13433 ( .A(n11733), .ZN(n10281) );
  NAND3_X1 U13434 ( .A1(n17476), .A2(n17477), .A3(n10288), .ZN(P3_U2642) );
  OR2_X1 U13435 ( .A1(n17505), .A2(n10301), .ZN(n10303) );
  NAND2_X1 U13436 ( .A1(n14477), .A2(n10309), .ZN(n10585) );
  INV_X1 U13437 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10310) );
  INV_X1 U13438 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U13439 ( .A1(n12875), .A2(n19860), .ZN(n10323) );
  OAI21_X1 U13440 ( .B1(n10324), .B2(n16678), .A(n16677), .ZN(n17332) );
  INV_X1 U13441 ( .A(n16511), .ZN(n10325) );
  NAND2_X1 U13442 ( .A1(n10328), .A2(n16758), .ZN(n10327) );
  INV_X1 U13443 ( .A(n10328), .ZN(n16458) );
  NAND2_X1 U13444 ( .A1(n11101), .A2(n11100), .ZN(n10329) );
  NAND4_X1 U13445 ( .A1(n10851), .A2(n10853), .A3(n10852), .A4(n10854), .ZN(
        n10334) );
  NAND4_X1 U13446 ( .A1(n10856), .A2(n10858), .A3(n10857), .A4(n10859), .ZN(
        n10335) );
  NAND2_X1 U13447 ( .A1(n11301), .A2(n10336), .ZN(n10339) );
  NAND2_X1 U13448 ( .A1(n11301), .A2(n11302), .ZN(n11282) );
  NAND2_X1 U13449 ( .A1(n11372), .A2(n10343), .ZN(n11364) );
  AND2_X1 U13450 ( .A1(n11356), .A2(n10348), .ZN(n11263) );
  NAND2_X1 U13451 ( .A1(n11356), .A2(n10347), .ZN(n11264) );
  NAND2_X1 U13452 ( .A1(n11356), .A2(n11277), .ZN(n11273) );
  NAND2_X1 U13453 ( .A1(n11359), .A2(n9717), .ZN(n11278) );
  NAND2_X1 U13454 ( .A1(n11359), .A2(n10492), .ZN(n11353) );
  NAND2_X1 U13455 ( .A1(n14196), .A2(n10360), .ZN(n18390) );
  NAND3_X1 U13456 ( .A1(n10362), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .ZN(n10361) );
  NAND3_X1 U13457 ( .A1(n16670), .A2(n9625), .A3(n16671), .ZN(n10368) );
  NAND2_X1 U13458 ( .A1(n13965), .A2(n21734), .ZN(n10377) );
  INV_X1 U13459 ( .A(n13965), .ZN(n10378) );
  NAND2_X1 U13460 ( .A1(n18786), .A2(n13965), .ZN(n18768) );
  NAND2_X1 U13461 ( .A1(n18784), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18786) );
  NAND2_X2 U13462 ( .A1(n18766), .A2(n13968), .ZN(n14123) );
  OR2_X1 U13463 ( .A1(n17247), .A2(n18644), .ZN(n10379) );
  NAND2_X1 U13464 ( .A1(n17247), .A2(n14430), .ZN(n10380) );
  AND2_X1 U13465 ( .A1(n14470), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10384) );
  NAND3_X1 U13466 ( .A1(n10598), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A3(
        n13654), .ZN(n10385) );
  NAND3_X1 U13467 ( .A1(n13654), .A2(n10597), .A3(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10386) );
  INV_X1 U13468 ( .A(n10567), .ZN(n10393) );
  NAND3_X1 U13469 ( .A1(n11814), .A2(n12152), .A3(n11928), .ZN(n11807) );
  NAND2_X1 U13470 ( .A1(n19753), .A2(n9637), .ZN(n10399) );
  NAND3_X1 U13471 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U13472 ( .A1(n14322), .A2(n9749), .ZN(n12858) );
  NAND2_X1 U13473 ( .A1(n13551), .A2(n9715), .ZN(n13270) );
  NOR2_X1 U13474 ( .A1(n15617), .A2(n15618), .ZN(n15602) );
  NAND2_X1 U13475 ( .A1(n11991), .A2(n10426), .ZN(n14762) );
  NAND2_X1 U13476 ( .A1(n12009), .A2(n9748), .ZN(n14706) );
  NAND2_X1 U13477 ( .A1(n10432), .A2(n10431), .ZN(n14002) );
  NAND2_X1 U13478 ( .A1(n15281), .A2(n11742), .ZN(n15271) );
  NAND2_X1 U13479 ( .A1(n15283), .A2(n15282), .ZN(n15281) );
  NAND2_X1 U13480 ( .A1(n11846), .A2(n15220), .ZN(n15107) );
  NAND2_X1 U13481 ( .A1(n11846), .A2(n10452), .ZN(n10454) );
  NAND2_X1 U13482 ( .A1(n10463), .A2(n10462), .ZN(n16579) );
  NAND3_X1 U13483 ( .A1(n9938), .A2(n16609), .A3(n9773), .ZN(n10463) );
  NAND2_X1 U13484 ( .A1(n10475), .A2(n12915), .ZN(P2_U3026) );
  NAND2_X1 U13485 ( .A1(n12924), .A2(n17351), .ZN(n10475) );
  NAND2_X1 U13486 ( .A1(n11326), .A2(n9676), .ZN(n11329) );
  NAND2_X1 U13487 ( .A1(n11263), .A2(n11268), .ZN(n15644) );
  INV_X1 U13488 ( .A(n11263), .ZN(n11270) );
  NAND2_X4 U13489 ( .A1(n10506), .A2(n10504), .ZN(n19879) );
  NAND4_X1 U13490 ( .A1(n10835), .A2(n10836), .A3(n10834), .A4(n10837), .ZN(
        n10505) );
  NAND4_X1 U13491 ( .A1(n10841), .A2(n10839), .A3(n10838), .A4(n10840), .ZN(
        n10507) );
  AND2_X1 U13492 ( .A1(n9622), .A2(n9742), .ZN(n15587) );
  NAND2_X1 U13493 ( .A1(n9622), .A2(n10520), .ZN(n12934) );
  AND2_X2 U13494 ( .A1(n13590), .A2(n10527), .ZN(n11724) );
  NAND2_X1 U13495 ( .A1(n11672), .A2(n20854), .ZN(n14245) );
  NAND2_X1 U13496 ( .A1(n12214), .A2(n9744), .ZN(n14731) );
  NOR2_X1 U13497 ( .A1(n14603), .A2(n14589), .ZN(n14588) );
  NAND2_X1 U13498 ( .A1(n9623), .A2(n12678), .ZN(n17330) );
  NAND2_X1 U13499 ( .A1(n9623), .A2(n20536), .ZN(n17348) );
  NAND2_X1 U13500 ( .A1(n11414), .A2(n11415), .ZN(n11424) );
  OR2_X1 U13501 ( .A1(n14020), .A2(n14090), .ZN(n14021) );
  NAND2_X1 U13502 ( .A1(n14090), .A2(n14020), .ZN(n14038) );
  OAI21_X1 U13503 ( .B1(n16211), .B2(n15945), .A(n13099), .ZN(n13114) );
  INV_X1 U13504 ( .A(n12950), .ZN(n11240) );
  NAND2_X1 U13505 ( .A1(n13131), .A2(n16984), .ZN(n13134) );
  INV_X1 U13506 ( .A(n12858), .ZN(n12860) );
  AOI21_X1 U13507 ( .B1(n16713), .B2(n16732), .A(n16436), .ZN(n16437) );
  NAND2_X1 U13508 ( .A1(n13132), .A2(n17351), .ZN(n13133) );
  NAND2_X1 U13509 ( .A1(n11950), .A2(n11947), .ZN(n11995) );
  NOR2_X1 U13510 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  NAND2_X1 U13511 ( .A1(n13034), .A2(n19868), .ZN(n13035) );
  CLKBUF_X1 U13512 ( .A(n13270), .Z(n13758) );
  AOI22_X1 U13513 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10837) );
  AOI21_X1 U13514 ( .B1(n10876), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n10810), .ZN(n10814) );
  OR2_X1 U13515 ( .A1(n11115), .A2(n11116), .ZN(n11117) );
  AND3_X1 U13516 ( .A1(n19879), .A2(n11246), .A3(n12656), .ZN(n10910) );
  AOI22_X1 U13517 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13518 ( .A1(n12114), .A2(n12115), .ZN(n15549) );
  NOR2_X1 U13519 ( .A1(n15587), .A2(n15586), .ZN(n16723) );
  OAI21_X1 U13520 ( .B1(n14552), .B2(n15954), .A(n13045), .ZN(n13046) );
  AND2_X1 U13521 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10855) );
  AND2_X1 U13522 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10825) );
  AND2_X1 U13523 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10810) );
  AND2_X1 U13524 ( .A1(n11932), .A2(n11931), .ZN(n12073) );
  NAND2_X1 U13525 ( .A1(n12196), .A2(n12195), .ZN(n14876) );
  AOI21_X1 U13526 ( .B1(n14888), .B2(n20756), .A(n14542), .ZN(n14543) );
  INV_X1 U13527 ( .A(n14101), .ZN(n12151) );
  CLKBUF_X1 U13528 ( .A(n12106), .Z(n20799) );
  NOR2_X1 U13529 ( .A1(n12969), .A2(n12968), .ZN(n10543) );
  OR2_X1 U13530 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10544) );
  OR2_X1 U13531 ( .A1(n19559), .A2(n19570), .ZN(n19676) );
  INV_X1 U13532 ( .A(n17616), .ZN(n17591) );
  INV_X1 U13533 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19619) );
  AND2_X1 U13534 ( .A1(n16502), .A2(n12913), .ZN(n10547) );
  AND3_X1 U13535 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U13536 ( .A1(n11950), .A2(n11944), .ZN(n10550) );
  AND2_X1 U13537 ( .A1(n14510), .A2(n14509), .ZN(n10551) );
  AND3_X1 U13538 ( .A1(n10888), .A2(n10887), .A3(n10886), .ZN(n10552) );
  AND2_X1 U13539 ( .A1(n11249), .A2(n15939), .ZN(n10553) );
  AND3_X1 U13540 ( .A1(n16235), .A2(n12867), .A3(n19868), .ZN(n10554) );
  INV_X1 U13541 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n21618) );
  INV_X1 U13542 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16669) );
  INV_X1 U13543 ( .A(n19647), .ZN(n19690) );
  INV_X1 U13544 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11842) );
  INV_X1 U13545 ( .A(n14325), .ZN(n17029) );
  AND2_X1 U13546 ( .A1(n12689), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10555) );
  OR2_X1 U13547 ( .A1(n19868), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10556) );
  OR2_X1 U13548 ( .A1(n19868), .A2(n11247), .ZN(n10557) );
  OR2_X1 U13549 ( .A1(n16848), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10558) );
  INV_X1 U13550 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11843) );
  INV_X1 U13551 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11142) );
  OR2_X1 U13552 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10559) );
  INV_X1 U13553 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19614) );
  INV_X1 U13554 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19616) );
  INV_X1 U13555 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13273) );
  NAND2_X2 U13556 ( .A1(n21511), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21577) );
  AND2_X1 U13557 ( .A1(n15016), .A2(BUF1_REG_30__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13558 ( .A1(n15036), .A2(n13188), .ZN(n15038) );
  INV_X1 U13559 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11850) );
  AND3_X1 U13560 ( .A1(n11149), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16451), .ZN(n10561) );
  INV_X2 U13561 ( .A(U214), .ZN(n17404) );
  AND2_X1 U13562 ( .A1(n13240), .A2(n13425), .ZN(n10562) );
  OR2_X1 U13563 ( .A1(n19868), .A2(n11261), .ZN(n10563) );
  INV_X1 U13564 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19657) );
  INV_X1 U13565 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11251) );
  AND2_X1 U13566 ( .A1(n19647), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19589) );
  INV_X1 U13567 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13342) );
  INV_X2 U13568 ( .A(n13950), .ZN(n19075) );
  INV_X1 U13569 ( .A(n15754), .ZN(n15755) );
  NAND2_X2 U13570 ( .A1(n20662), .A2(n11551), .ZN(n14935) );
  INV_X1 U13571 ( .A(n13186), .ZN(n15009) );
  INV_X2 U13572 ( .A(n15009), .ZN(n15036) );
  AOI21_X1 U13573 ( .B1(n13185), .B2(n13184), .A(n20568), .ZN(n13186) );
  AND3_X1 U13574 ( .A1(n21275), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10565) );
  AND2_X1 U13575 ( .A1(n12710), .A2(n12691), .ZN(n10566) );
  INV_X1 U13576 ( .A(n12697), .ZN(n13025) );
  NAND2_X1 U13577 ( .A1(n13291), .A2(n13292), .ZN(n12705) );
  NAND2_X1 U13578 ( .A1(n11666), .A2(n11665), .ZN(n10567) );
  AND4_X1 U13579 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n10568) );
  AND4_X1 U13580 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n10569) );
  INV_X1 U13581 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U13582 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10854) );
  INV_X1 U13583 ( .A(n11880), .ZN(n11867) );
  XNOR2_X1 U13584 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11865) );
  INV_X1 U13585 ( .A(n14857), .ZN(n12213) );
  OR2_X1 U13586 ( .A1(n11753), .A2(n11752), .ZN(n11774) );
  INV_X1 U13587 ( .A(n11333), .ZN(n11256) );
  NAND2_X1 U13588 ( .A1(n11158), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10951) );
  INV_X1 U13589 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12992) );
  INV_X1 U13590 ( .A(n15849), .ZN(n11175) );
  AOI21_X1 U13591 ( .B1(n12655), .B2(n12647), .A(n12699), .ZN(n10899) );
  NOR2_X1 U13592 ( .A1(n11930), .A2(n11573), .ZN(n11549) );
  OR2_X1 U13593 ( .A1(n11860), .A2(n11859), .ZN(n11862) );
  NOR2_X1 U13594 ( .A1(n12240), .A2(n14848), .ZN(n12241) );
  AND2_X1 U13595 ( .A1(n11798), .A2(n11797), .ZN(n11800) );
  AOI22_X1 U13596 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11464) );
  OR2_X1 U13597 ( .A1(n11796), .A2(n11795), .ZN(n11816) );
  INV_X1 U13598 ( .A(n11700), .ZN(n11736) );
  NAND2_X1 U13599 ( .A1(n11557), .A2(n11556), .ZN(n11559) );
  INV_X1 U13600 ( .A(n16267), .ZN(n16014) );
  NAND2_X1 U13601 ( .A1(n16235), .A2(n12718), .ZN(n11003) );
  INV_X1 U13602 ( .A(n15915), .ZN(n12722) );
  INV_X1 U13603 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13740) );
  INV_X1 U13604 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14427) );
  INV_X1 U13605 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10594) );
  OR4_X1 U13606 ( .A1(n11909), .A2(n11902), .A3(n11877), .A4(n11890), .ZN(
        n11871) );
  OR2_X1 U13607 ( .A1(n12522), .A2(n12521), .ZN(n12545) );
  OR2_X1 U13608 ( .A1(n11950), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11951) );
  AND2_X1 U13609 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12569) );
  INV_X1 U13610 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12488) );
  AND2_X1 U13611 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12280) );
  AND2_X1 U13612 ( .A1(n12241), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12281) );
  INV_X1 U13613 ( .A(n13998), .ZN(n12129) );
  INV_X1 U13614 ( .A(n11818), .ZN(n11827) );
  INV_X1 U13615 ( .A(n11683), .ZN(n11684) );
  NAND2_X1 U13616 ( .A1(n11240), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12949) );
  INV_X1 U13617 ( .A(n12862), .ZN(n12859) );
  INV_X1 U13618 ( .A(n11253), .ZN(n12731) );
  INV_X1 U13619 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16532) );
  OAI21_X1 U13620 ( .B1(n19868), .B2(n10553), .A(n11250), .ZN(n11296) );
  NOR2_X1 U13621 ( .A1(n11143), .A2(n16727), .ZN(n11429) );
  AND2_X1 U13622 ( .A1(n13017), .A2(n13016), .ZN(n15659) );
  INV_X1 U13623 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21702) );
  INV_X1 U13624 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n21601) );
  INV_X1 U13625 ( .A(n17106), .ZN(n10572) );
  AOI21_X1 U13626 ( .B1(n10748), .B2(n10747), .A(n10746), .ZN(n10753) );
  INV_X1 U13627 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17882) );
  INV_X1 U13628 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21664) );
  INV_X1 U13629 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14436) );
  INV_X1 U13630 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17843) );
  INV_X1 U13631 ( .A(n14545), .ZN(n11551) );
  NAND2_X1 U13632 ( .A1(n20594), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14244) );
  INV_X1 U13633 ( .A(n14763), .ZN(n12008) );
  OR2_X1 U13634 ( .A1(n17305), .A2(n13178), .ZN(n13185) );
  NAND2_X1 U13635 ( .A1(n12569), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14221) );
  NAND2_X1 U13636 ( .A1(n12408), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12439) );
  AND2_X1 U13637 ( .A1(n12105), .A2(n12239), .ZN(n14793) );
  NAND2_X1 U13638 ( .A1(n12142), .A2(n12141), .ZN(n14033) );
  INV_X1 U13639 ( .A(n14932), .ZN(n11973) );
  INV_X1 U13640 ( .A(n21235), .ZN(n21424) );
  INV_X1 U13641 ( .A(n20975), .ZN(n20803) );
  INV_X1 U13642 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21276) );
  AND2_X1 U13643 ( .A1(n13022), .A2(n13021), .ZN(n15618) );
  AND2_X1 U13644 ( .A1(n16040), .A2(n16039), .ZN(n16077) );
  INV_X1 U13645 ( .A(n15721), .ZN(n12857) );
  NAND2_X1 U13646 ( .A1(n13083), .A2(n13082), .ZN(n13084) );
  AND2_X1 U13647 ( .A1(n11421), .A2(n13147), .ZN(n16460) );
  INV_X1 U13648 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21729) );
  NOR2_X1 U13649 ( .A1(n10902), .A2(n10909), .ZN(n10906) );
  AND2_X1 U13650 ( .A1(n12681), .A2(n10554), .ZN(n14372) );
  NAND2_X1 U13651 ( .A1(n14039), .A2(n20501), .ZN(n14015) );
  INV_X1 U13652 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17687) );
  INV_X1 U13653 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n21633) );
  INV_X1 U13654 ( .A(n10588), .ZN(n10571) );
  OR2_X1 U13655 ( .A1(n9659), .A2(n18624), .ZN(n18603) );
  OR2_X1 U13656 ( .A1(n18227), .A2(n10638), .ZN(n10639) );
  NAND2_X1 U13657 ( .A1(n11552), .A2(n11551), .ZN(n12061) );
  INV_X1 U13658 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14848) );
  NOR2_X1 U13659 ( .A1(n14244), .A2(n11573), .ZN(n14250) );
  OR2_X1 U13660 ( .A1(n20593), .A2(n21571), .ZN(n20637) );
  INV_X1 U13661 ( .A(n12107), .ZN(n13189) );
  NAND2_X1 U13662 ( .A1(n12530), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12567) );
  NAND2_X1 U13663 ( .A1(n12441), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12487) );
  NAND2_X1 U13664 ( .A1(n12330), .A2(n12329), .ZN(n12366) );
  AND3_X1 U13665 ( .A1(n12212), .A2(n12211), .A3(n12210), .ZN(n14857) );
  AND2_X1 U13666 ( .A1(n12039), .A2(n12038), .ZN(n14642) );
  AND2_X1 U13667 ( .A1(n12030), .A2(n12029), .ZN(n14681) );
  OR2_X1 U13668 ( .A1(n20766), .A2(n15486), .ZN(n15516) );
  AOI21_X1 U13669 ( .B1(n15220), .B2(n15152), .A(n15229), .ZN(n15187) );
  AND2_X1 U13670 ( .A1(n12084), .A2(n12083), .ZN(n13565) );
  INV_X1 U13671 ( .A(n20770), .ZN(n20744) );
  INV_X1 U13672 ( .A(n14245), .ZN(n21375) );
  OR2_X1 U13673 ( .A1(n21327), .A2(n20855), .ZN(n20887) );
  AND2_X1 U13674 ( .A1(n20934), .A2(n21432), .ZN(n20938) );
  AND2_X1 U13675 ( .A1(n21084), .A2(n21083), .ZN(n21111) );
  AND2_X1 U13676 ( .A1(n21160), .A2(n21159), .ZN(n21187) );
  INV_X1 U13677 ( .A(n21283), .ZN(n21316) );
  AND2_X1 U13678 ( .A1(n21368), .A2(n21367), .ZN(n21416) );
  NAND2_X1 U13679 ( .A1(n20839), .A2(n20846), .ZN(n21481) );
  NAND2_X1 U13680 ( .A1(n10920), .A2(n13038), .ZN(n12868) );
  AOI21_X1 U13681 ( .B1(n13076), .B2(n19750), .A(n13044), .ZN(n13045) );
  INV_X1 U13682 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15677) );
  INV_X1 U13683 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15733) );
  INV_X1 U13684 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16573) );
  INV_X1 U13685 ( .A(n19748), .ZN(n19737) );
  INV_X1 U13686 ( .A(n17339), .ZN(n19745) );
  AND2_X1 U13687 ( .A1(n13010), .A2(n13009), .ZN(n15706) );
  INV_X1 U13688 ( .A(n16409), .ZN(n16392) );
  NAND2_X2 U13689 ( .A1(n13231), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n14325)
         );
  INV_X1 U13690 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16798) );
  AND2_X1 U13691 ( .A1(n16876), .A2(n10558), .ZN(n16849) );
  INV_X1 U13692 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16703) );
  AOI21_X1 U13693 ( .B1(n14015), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13419), .ZN(n13420) );
  INV_X1 U13694 ( .A(n20508), .ZN(n20103) );
  NAND2_X1 U13695 ( .A1(n20501), .A2(n20552), .ZN(n20543) );
  AND2_X1 U13696 ( .A1(n20552), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20262) );
  NAND2_X1 U13697 ( .A1(n20514), .A2(n20361), .ZN(n17028) );
  AND2_X1 U13698 ( .A1(n16992), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13040) );
  OR2_X1 U13699 ( .A1(n17801), .A2(n14481), .ZN(n11440) );
  INV_X1 U13700 ( .A(n10765), .ZN(n10756) );
  INV_X1 U13701 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18054) );
  AOI21_X1 U13702 ( .B1(n13619), .B2(n13618), .A(n13836), .ZN(n19513) );
  INV_X1 U13703 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18084) );
  AND2_X1 U13704 ( .A1(n18929), .A2(n14460), .ZN(n17237) );
  INV_X1 U13705 ( .A(n17623), .ZN(n18703) );
  AND2_X1 U13706 ( .A1(n18673), .A2(n18944), .ZN(n18942) );
  NOR2_X1 U13707 ( .A1(n13605), .A2(n13604), .ZN(n13656) );
  INV_X1 U13708 ( .A(n18664), .ZN(n18988) );
  NAND2_X1 U13709 ( .A1(n19684), .A2(n14193), .ZN(n19061) );
  NOR2_X1 U13710 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19094), .ZN(n19387) );
  INV_X1 U13711 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19872) );
  NOR2_X1 U13712 ( .A1(n19660), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19409) );
  NAND2_X1 U13713 ( .A1(n20594), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14235) );
  AND2_X1 U13714 ( .A1(n20594), .A2(n14713), .ZN(n20629) );
  INV_X1 U13715 ( .A(n14935), .ZN(n20659) );
  INV_X1 U13716 ( .A(n15038), .ZN(n14997) );
  OR2_X1 U13717 ( .A1(n14929), .A2(n14922), .ZN(n14924) );
  INV_X1 U13718 ( .A(n20742), .ZN(n15172) );
  OR2_X1 U13719 ( .A1(n17305), .A2(n13314), .ZN(n17295) );
  INV_X1 U13720 ( .A(n20574), .ZN(n20738) );
  INV_X1 U13721 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13208) );
  INV_X1 U13722 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15330) );
  AND2_X1 U13723 ( .A1(n15462), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15445) );
  INV_X1 U13724 ( .A(n20784), .ZN(n20760) );
  AND2_X1 U13725 ( .A1(n12091), .A2(n12063), .ZN(n20756) );
  NAND2_X1 U13726 ( .A1(n13573), .A2(n13681), .ZN(n21279) );
  OAI22_X1 U13727 ( .A1(n20812), .A2(n20811), .B1(n21202), .B2(n20810), .ZN(
        n20850) );
  OAI22_X1 U13728 ( .A1(n20900), .A2(n20899), .B1(n21202), .B2(n21051), .ZN(
        n20923) );
  OAI22_X1 U13729 ( .A1(n20939), .A2(n20938), .B1(n21503), .B2(n20937), .ZN(
        n20962) );
  INV_X1 U13730 ( .A(n20978), .ZN(n21002) );
  INV_X1 U13731 ( .A(n21075), .ZN(n21040) );
  OAI22_X1 U13732 ( .A1(n21053), .A2(n21052), .B1(n21051), .B2(n21286), .ZN(
        n21077) );
  OAI21_X1 U13733 ( .B1(n21086), .B2(n10565), .A(n21439), .ZN(n21114) );
  INV_X1 U13734 ( .A(n21125), .ZN(n21153) );
  OAI211_X1 U13735 ( .C1(n21129), .C2(n21282), .A(n21200), .B(n21128), .ZN(
        n21154) );
  INV_X1 U13736 ( .A(n21231), .ZN(n21189) );
  OAI22_X1 U13737 ( .A1(n21204), .A2(n21203), .B1(n21202), .B2(n21364), .ZN(
        n21227) );
  OAI21_X1 U13738 ( .B1(n21244), .B2(n21243), .A(n21439), .ZN(n21270) );
  INV_X1 U13739 ( .A(n21430), .ZN(n21289) );
  INV_X1 U13740 ( .A(n21475), .ZN(n21309) );
  INV_X1 U13741 ( .A(n21336), .ZN(n21360) );
  OAI211_X1 U13742 ( .C1(n21380), .C2(n21379), .A(n21378), .B(n21377), .ZN(
        n21419) );
  INV_X1 U13743 ( .A(n21381), .ZN(n21494) );
  NAND2_X1 U13744 ( .A1(n21500), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17301) );
  INV_X1 U13745 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21511) );
  INV_X1 U13746 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21520) );
  INV_X1 U13747 ( .A(n17055), .ZN(n19706) );
  INV_X1 U13748 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16602) );
  INV_X1 U13749 ( .A(n19750), .ZN(n15941) );
  AND2_X1 U13750 ( .A1(n20545), .A2(n13039), .ZN(n19750) );
  AND2_X1 U13751 ( .A1(n20545), .A2(n12935), .ZN(n19761) );
  OR2_X1 U13752 ( .A1(n12802), .A2(n12801), .ZN(n14096) );
  OR2_X1 U13753 ( .A1(n12762), .A2(n12761), .ZN(n16313) );
  INV_X1 U13754 ( .A(n13028), .ZN(n13029) );
  AND2_X1 U13755 ( .A1(n14326), .A2(n14325), .ZN(n16409) );
  OR2_X1 U13756 ( .A1(n16003), .A2(n16002), .ZN(n16271) );
  AND2_X1 U13757 ( .A1(n14326), .A2(n17029), .ZN(n16395) );
  NAND2_X1 U13758 ( .A1(n13523), .A2(n17055), .ZN(n13526) );
  INV_X1 U13759 ( .A(n19768), .ZN(n19785) );
  INV_X1 U13760 ( .A(n13537), .ZN(n20548) );
  INV_X1 U13761 ( .A(n13343), .ZN(n19830) );
  INV_X2 U13762 ( .A(n19834), .ZN(n19836) );
  OAI21_X1 U13763 ( .B1(n13159), .B2(n16707), .A(n13158), .ZN(n13160) );
  AND2_X1 U13764 ( .A1(n15857), .A2(n15848), .ZN(n16650) );
  INV_X1 U13765 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16745) );
  AND2_X1 U13766 ( .A1(n15725), .A2(n12672), .ZN(n16829) );
  INV_X1 U13767 ( .A(n16988), .ZN(n17351) );
  NAND2_X1 U13768 ( .A1(n9623), .A2(n12684), .ZN(n17340) );
  NOR2_X1 U13769 ( .A1(n20543), .A2(n20356), .ZN(n20514) );
  INV_X1 U13770 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16992) );
  NOR2_X1 U13771 ( .A1(n19888), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19881) );
  OR3_X1 U13772 ( .A1(n19921), .A2(n20265), .A3(n19920), .ZN(n19940) );
  OAI21_X1 U13773 ( .B1(n19956), .B2(n19955), .A(n19954), .ZN(n19980) );
  OAI21_X1 U13774 ( .B1(n17044), .B2(n17043), .A(n17042), .ZN(n20036) );
  NAND2_X1 U13775 ( .A1(n17018), .A2(n17017), .ZN(n20361) );
  AND2_X1 U13776 ( .A1(n20199), .A2(n20076), .ZN(n20110) );
  NAND2_X1 U13777 ( .A1(n20112), .A2(n20111), .ZN(n20129) );
  OAI21_X1 U13778 ( .B1(n20142), .B2(n20141), .A(n20140), .ZN(n20164) );
  INV_X1 U13779 ( .A(n20172), .ZN(n20194) );
  INV_X1 U13780 ( .A(n20205), .ZN(n20224) );
  INV_X1 U13781 ( .A(n20388), .ZN(n20281) );
  OAI21_X1 U13782 ( .B1(n20308), .B2(n20307), .A(n20306), .ZN(n20343) );
  INV_X1 U13783 ( .A(n20526), .ZN(n20269) );
  INV_X1 U13784 ( .A(n20320), .ZN(n20377) );
  INV_X1 U13785 ( .A(n19734), .ZN(n19757) );
  AND2_X1 U13786 ( .A1(n20522), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17356) );
  INV_X1 U13787 ( .A(n20566), .ZN(n19702) );
  INV_X1 U13788 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20428) );
  NAND2_X1 U13789 ( .A1(n19675), .A2(n19516), .ZN(n18473) );
  AND2_X1 U13790 ( .A1(n11441), .A2(n11440), .ZN(n11442) );
  INV_X1 U13791 ( .A(n17594), .ZN(n17592) );
  NAND2_X1 U13792 ( .A1(n10592), .A2(n10591), .ZN(n13259) );
  INV_X1 U13793 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21713) );
  INV_X1 U13794 ( .A(n17812), .ZN(n17785) );
  INV_X1 U13795 ( .A(n19566), .ZN(n17781) );
  INV_X1 U13796 ( .A(n17806), .ZN(n17796) );
  INV_X1 U13797 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17936) );
  NAND2_X1 U13798 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17972), .ZN(n17967) );
  INV_X1 U13799 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18257) );
  INV_X1 U13800 ( .A(n18320), .ZN(n18350) );
  OAI211_X1 U13801 ( .C1(n19682), .C2(n19681), .A(n9897), .B(n18474), .ZN(
        n18512) );
  NAND2_X1 U13802 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17106) );
  OR2_X1 U13803 ( .A1(n14157), .A2(n14156), .ZN(n17215) );
  INV_X1 U13804 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17144) );
  NOR2_X1 U13805 ( .A1(n19559), .A2(n19680), .ZN(n18790) );
  AND2_X1 U13806 ( .A1(n14455), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18828) );
  INV_X1 U13807 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18969) );
  AND2_X1 U13808 ( .A1(n19693), .A2(n10757), .ZN(n13950) );
  AND2_X1 U13809 ( .A1(n19074), .A2(n17215), .ZN(n19007) );
  INV_X1 U13810 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21719) );
  AND2_X1 U13811 ( .A1(n19070), .A2(n17216), .ZN(n19074) );
  AND2_X1 U13812 ( .A1(n13845), .A2(n19675), .ZN(n19070) );
  INV_X1 U13813 ( .A(n19387), .ZN(n19184) );
  INV_X1 U13814 ( .A(n19456), .ZN(n19155) );
  INV_X1 U13815 ( .A(n19512), .ZN(n19178) );
  INV_X1 U13816 ( .A(n19162), .ZN(n19201) );
  INV_X1 U13817 ( .A(n19159), .ZN(n19223) );
  INV_X1 U13818 ( .A(n19249), .ZN(n19266) );
  AND2_X1 U13819 ( .A1(n19560), .A2(n19319), .ZN(n19289) );
  INV_X1 U13820 ( .A(n19274), .ZN(n19313) );
  NOR2_X1 U13821 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19528), .ZN(
        n19316) );
  INV_X1 U13822 ( .A(n19362), .ZN(n19364) );
  INV_X1 U13823 ( .A(n19363), .ZN(n19404) );
  INV_X1 U13824 ( .A(n19384), .ZN(n19426) );
  AND2_X1 U13825 ( .A1(n19560), .A2(n19436), .ZN(n19451) );
  INV_X1 U13826 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19692) );
  NOR3_X1 U13827 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19589), .A3(n19572), 
        .ZN(n13830) );
  INV_X1 U13828 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21652) );
  NAND2_X2 U13829 ( .A1(n13199), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20796)
         );
  INV_X1 U13830 ( .A(U212), .ZN(n17403) );
  OR3_X1 U13831 ( .A1(n17305), .A2(n13428), .A3(n20568), .ZN(n14226) );
  INV_X1 U13832 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21373) );
  INV_X1 U13833 ( .A(n20647), .ZN(n20615) );
  OR2_X1 U13834 ( .A1(n13705), .A2(n20798), .ZN(n15014) );
  OR2_X1 U13835 ( .A1(n13705), .A2(n20796), .ZN(n15001) );
  INV_X1 U13836 ( .A(n15226), .ZN(n15029) );
  INV_X1 U13837 ( .A(n14973), .ZN(n20849) );
  INV_X1 U13838 ( .A(n14006), .ZN(n20821) );
  OR2_X1 U13839 ( .A1(n13432), .A2(n20688), .ZN(n20667) );
  OR2_X1 U13840 ( .A1(n20695), .A2(n11573), .ZN(n20663) );
  OR2_X1 U13841 ( .A1(n13431), .A2(n17305), .ZN(n20695) );
  NOR2_X1 U13842 ( .A1(n14226), .A2(n13773), .ZN(n13800) );
  INV_X1 U13843 ( .A(n20723), .ZN(n13804) );
  NAND2_X2 U13844 ( .A1(n15169), .A2(n13729), .ZN(n20742) );
  OR2_X2 U13845 ( .A1(n17295), .A2(n20568), .ZN(n20574) );
  INV_X1 U13846 ( .A(n20756), .ZN(n20788) );
  INV_X1 U13847 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20780) );
  NAND2_X2 U13848 ( .A1(n12091), .A2(n11943), .ZN(n20784) );
  AOI21_X1 U13849 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21501), .A(n13575), 
        .ZN(n13698) );
  NAND2_X1 U13850 ( .A1(n20933), .A2(n21117), .ZN(n20880) );
  NAND2_X1 U13851 ( .A1(n20933), .A2(n21324), .ZN(n20927) );
  NAND2_X1 U13852 ( .A1(n20933), .A2(n21194), .ZN(n20966) );
  OR2_X1 U13853 ( .A1(n21088), .A2(n21274), .ZN(n21044) );
  OR2_X1 U13854 ( .A1(n21088), .A2(n21006), .ZN(n21075) );
  OR2_X1 U13855 ( .A1(n21088), .A2(n21371), .ZN(n21109) );
  NAND2_X1 U13856 ( .A1(n21233), .A2(n21117), .ZN(n21193) );
  NAND2_X1 U13857 ( .A1(n21233), .A2(n21324), .ZN(n21231) );
  NAND2_X1 U13858 ( .A1(n21233), .A2(n21194), .ZN(n21273) );
  NAND2_X1 U13859 ( .A1(n21233), .A2(n21232), .ZN(n21323) );
  NAND2_X1 U13860 ( .A1(n21434), .A2(n21324), .ZN(n21422) );
  NOR2_X1 U13861 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21587) );
  INV_X1 U13862 ( .A(n21569), .ZN(n21505) );
  INV_X1 U13863 ( .A(n21577), .ZN(n21579) );
  OR2_X1 U13864 ( .A1(n21520), .A2(n21577), .ZN(n21543) );
  NAND2_X1 U13865 ( .A1(n15959), .A2(n13100), .ZN(n20545) );
  NAND2_X1 U13866 ( .A1(n10896), .A2(n17055), .ZN(n19708) );
  NOR2_X1 U13867 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  NAND2_X1 U13868 ( .A1(n19835), .A2(n13033), .ZN(n15954) );
  INV_X1 U13869 ( .A(n19761), .ZN(n15945) );
  NAND2_X1 U13870 ( .A1(n13487), .A2(n13330), .ZN(n15959) );
  AND2_X1 U13871 ( .A1(n13424), .A2(n17055), .ZN(n16308) );
  NAND2_X1 U13872 ( .A1(n12699), .A2(n19768), .ZN(n19770) );
  NAND2_X1 U13873 ( .A1(n19768), .A2(n13527), .ZN(n16398) );
  NAND2_X1 U13874 ( .A1(n13526), .A2(n13525), .ZN(n19768) );
  AND2_X1 U13875 ( .A1(n13372), .A2(n13371), .ZN(n19863) );
  OR2_X1 U13876 ( .A1(n19828), .A2(n13492), .ZN(n13536) );
  OR2_X1 U13877 ( .A1(n13735), .A2(n16992), .ZN(n13537) );
  NAND2_X1 U13878 ( .A1(n13491), .A2(n20560), .ZN(n19828) );
  INV_X1 U13879 ( .A(n19835), .ZN(n13488) );
  OR2_X1 U13880 ( .A1(n13306), .A2(n16235), .ZN(n13343) );
  INV_X1 U13881 ( .A(n16713), .ZN(n16707) );
  INV_X1 U13882 ( .A(n13151), .ZN(n13152) );
  INV_X1 U13883 ( .A(n13069), .ZN(n13070) );
  NAND2_X1 U13884 ( .A1(n9623), .A2(n20537), .ZN(n16988) );
  INV_X1 U13885 ( .A(n10797), .ZN(n17004) );
  NAND2_X1 U13886 ( .A1(n19892), .A2(n20526), .ZN(n19898) );
  NAND2_X1 U13887 ( .A1(n19892), .A2(n20269), .ZN(n19943) );
  NAND2_X1 U13888 ( .A1(n19947), .A2(n20269), .ZN(n19978) );
  NAND2_X1 U13889 ( .A1(n19947), .A2(n20526), .ZN(n19984) );
  INV_X1 U13890 ( .A(n20037), .ZN(n20022) );
  NAND2_X1 U13891 ( .A1(n17045), .A2(n20526), .ZN(n20040) );
  NAND2_X1 U13892 ( .A1(n20492), .A2(n20526), .ZN(n20102) );
  AOI22_X1 U13893 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19883), .ZN(n21759) );
  NAND2_X1 U13894 ( .A1(n20209), .A2(n20526), .ZN(n20229) );
  INV_X1 U13895 ( .A(n20397), .ZN(n20256) );
  AOI22_X1 U13896 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19883), .ZN(n20400) );
  INV_X1 U13897 ( .A(n20491), .ZN(n20412) );
  INV_X1 U13898 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20429) );
  INV_X1 U13899 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20459) );
  INV_X1 U13900 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19680) );
  NAND2_X1 U13901 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  INV_X1 U13902 ( .A(n17573), .ZN(n17585) );
  INV_X1 U13903 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17744) );
  INV_X1 U13904 ( .A(n17800), .ZN(n17768) );
  INV_X1 U13905 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18005) );
  NAND2_X1 U13906 ( .A1(n19131), .A2(n18272), .ZN(n18184) );
  INV_X1 U13907 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18265) );
  AND2_X1 U13908 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18369), .ZN(n18372) );
  NOR2_X1 U13909 ( .A1(n14140), .A2(n14139), .ZN(n18397) );
  NOR2_X1 U13910 ( .A1(n18273), .A2(n18319), .ZN(n18407) );
  INV_X1 U13911 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18429) );
  NAND2_X1 U13912 ( .A1(n18442), .A2(n9889), .ZN(n18440) );
  INV_X1 U13913 ( .A(n18442), .ZN(n18471) );
  INV_X1 U13914 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19096) );
  INV_X1 U13915 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19107) );
  INV_X1 U13916 ( .A(n18519), .ZN(n18515) );
  INV_X1 U13917 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18862) );
  INV_X1 U13918 ( .A(n19070), .ZN(n19080) );
  INV_X1 U13919 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19010) );
  NAND2_X1 U13920 ( .A1(n19080), .A2(n19075), .ZN(n19072) );
  INV_X1 U13921 ( .A(n19079), .ZN(n19021) );
  INV_X1 U13922 ( .A(n17280), .ZN(n13720) );
  NAND2_X1 U13923 ( .A1(n13636), .A2(n13635), .ZN(n17280) );
  NAND2_X1 U13924 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19228), .ZN(
        n19249) );
  INV_X1 U13925 ( .A(n19358), .ZN(n19294) );
  NAND2_X1 U13926 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19410), .ZN(
        n19432) );
  INV_X1 U13927 ( .A(n19504), .ZN(n19431) );
  NAND2_X1 U13928 ( .A1(n19132), .A2(n9889), .ZN(n19465) );
  NAND2_X1 U13929 ( .A1(n19132), .A2(n19117), .ZN(n19489) );
  NAND4_X1 U13930 ( .A1(n19692), .A2(n19657), .A3(n19680), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n19566) );
  INV_X1 U13931 ( .A(n19656), .ZN(n19571) );
  NAND2_X1 U13932 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19682) );
  INV_X1 U13933 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19601) );
  INV_X1 U13934 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19626) );
  NOR2_X1 U13935 ( .A1(n14325), .A2(n13232), .ZN(n17361) );
  INV_X1 U13936 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19133) );
  INV_X1 U13937 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19124) );
  INV_X1 U13938 ( .A(n17401), .ZN(n17406) );
  INV_X1 U13939 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n21626) );
  OAI21_X1 U13940 ( .B1(n15045), .B2(n20784), .A(n13217), .ZN(P1_U3002) );
  OR4_X1 U13941 ( .A1(n13285), .A2(n13284), .A3(n13283), .A4(n13282), .ZN(
        P2_U2844) );
  OR4_X1 U13942 ( .A1(n13257), .A2(n13256), .A3(n13255), .A4(n13254), .ZN(
        P2_U3044) );
  OR4_X1 U13943 ( .A1(n13266), .A2(n13265), .A3(n13264), .A4(n13263), .ZN(
        P3_U2651) );
  NAND2_X1 U13944 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17163) );
  NOR2_X1 U13945 ( .A1(n17163), .A2(n17687), .ZN(n17626) );
  NAND2_X1 U13946 ( .A1(n17149), .A2(n17626), .ZN(n10586) );
  NAND2_X1 U13947 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17627) );
  NAND2_X1 U13948 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17638) );
  NAND2_X1 U13949 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18650) );
  NAND2_X1 U13950 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18610) );
  NAND2_X1 U13951 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18575) );
  NAND2_X1 U13952 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18535) );
  XNOR2_X1 U13953 ( .A(n10310), .B(n9757), .ZN(n17071) );
  AOI21_X1 U13954 ( .B1(n17081), .B2(n17478), .A(n9757), .ZN(n17472) );
  INV_X1 U13955 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21668) );
  INV_X1 U13956 ( .A(n10573), .ZN(n10576) );
  NOR2_X1 U13957 ( .A1(n21668), .A2(n10576), .ZN(n10574) );
  OR2_X1 U13958 ( .A1(n10574), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10575) );
  AND2_X1 U13959 ( .A1(n17081), .A2(n10575), .ZN(n17483) );
  OAI22_X1 U13960 ( .A1(n21668), .A2(n10573), .B1(n10576), .B2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17493) );
  INV_X1 U13961 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10578) );
  INV_X1 U13962 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18816) );
  NOR2_X1 U13963 ( .A1(n18816), .A2(n10577), .ZN(n10581) );
  INV_X1 U13964 ( .A(n10581), .ZN(n10580) );
  OR2_X1 U13965 ( .A1(n18535), .A2(n10580), .ZN(n17095) );
  AOI21_X1 U13966 ( .B1(n10578), .B2(n17095), .A(n10573), .ZN(n18524) );
  INV_X1 U13967 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18550) );
  NOR2_X1 U13968 ( .A1(n18550), .A2(n10580), .ZN(n10579) );
  OAI21_X1 U13969 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n10579), .A(
        n17095), .ZN(n18537) );
  INV_X1 U13970 ( .A(n18537), .ZN(n17514) );
  AOI21_X1 U13971 ( .B1(n18550), .B2(n10580), .A(n10579), .ZN(n18546) );
  NAND2_X1 U13972 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9725), .ZN(
        n18534) );
  AOI21_X1 U13973 ( .B1(n10299), .B2(n18534), .A(n10581), .ZN(n18560) );
  INV_X1 U13974 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18577) );
  NAND2_X1 U13975 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18597), .ZN(
        n18571) );
  NOR2_X1 U13976 ( .A1(n10298), .A2(n18571), .ZN(n10584) );
  NAND2_X1 U13977 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10584), .ZN(
        n10583) );
  INV_X1 U13978 ( .A(n18534), .ZN(n10582) );
  AOI21_X1 U13979 ( .B1(n18577), .B2(n10583), .A(n10582), .ZN(n18580) );
  XOR2_X1 U13980 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n10584), .Z(
        n18590) );
  AOI21_X1 U13981 ( .B1(n10298), .B2(n18571), .A(n10584), .ZN(n18599) );
  NOR2_X1 U13982 ( .A1(n18816), .A2(n10586), .ZN(n17150) );
  INV_X1 U13983 ( .A(n17150), .ZN(n10587) );
  NOR2_X1 U13984 ( .A1(n17627), .A2(n10587), .ZN(n17623) );
  NOR2_X1 U13985 ( .A1(n10588), .A2(n18703), .ZN(n18647) );
  NAND2_X1 U13986 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18647), .ZN(
        n17611) );
  INV_X1 U13987 ( .A(n17611), .ZN(n17603) );
  INV_X1 U13988 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17803) );
  AND2_X1 U13989 ( .A1(n17603), .A2(n17803), .ZN(n10589) );
  INV_X1 U13990 ( .A(n17613), .ZN(n10592) );
  NOR2_X1 U13991 ( .A1(n18599), .A2(n13259), .ZN(n13258) );
  NOR2_X1 U13992 ( .A1(n17544), .A2(n10301), .ZN(n17536) );
  NOR2_X1 U13993 ( .A1(n18560), .A2(n17536), .ZN(n17535) );
  NOR2_X1 U13994 ( .A1(n17535), .A2(n10301), .ZN(n17529) );
  NOR2_X1 U13995 ( .A1(n18546), .A2(n17529), .ZN(n17528) );
  NOR2_X1 U13996 ( .A1(n17528), .A2(n10301), .ZN(n17513) );
  NOR2_X1 U13997 ( .A1(n17514), .A2(n17513), .ZN(n17512) );
  NOR2_X1 U13998 ( .A1(n17512), .A2(n10301), .ZN(n17504) );
  NOR2_X1 U13999 ( .A1(n17482), .A2(n10301), .ZN(n17471) );
  NOR2_X1 U14000 ( .A1(n17470), .A2(n10301), .ZN(n11437) );
  OAI21_X1 U14001 ( .B1(n17071), .B2(n11437), .A(n17781), .ZN(n10593) );
  AOI21_X1 U14002 ( .B1(n17071), .B2(n11437), .A(n10593), .ZN(n10774) );
  NAND3_X1 U14003 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(P3_REIP_REG_24__SCAN_IN), .ZN(n10766) );
  INV_X1 U14004 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19631) );
  INV_X1 U14005 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19628) );
  INV_X1 U14006 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U14007 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U14008 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10605) );
  INV_X1 U14009 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U14010 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U14011 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10599) );
  OAI211_X1 U14012 ( .C1(n9603), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        n10602) );
  INV_X1 U14013 ( .A(n10602), .ZN(n10604) );
  INV_X1 U14014 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17896) );
  OR2_X1 U14015 ( .A1(n18227), .A2(n17896), .ZN(n10603) );
  NAND4_X1 U14016 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10619) );
  INV_X1 U14017 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U14018 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10617) );
  AND2_X2 U14019 ( .A1(n13609), .A2(n10609), .ZN(n13869) );
  AOI22_X1 U14020 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10616) );
  INV_X4 U14021 ( .A(n18060), .ZN(n18234) );
  AOI22_X1 U14022 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10615) );
  AND2_X4 U14023 ( .A1(n13651), .A2(n10613), .ZN(n18235) );
  AOI22_X1 U14024 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10614) );
  NAND4_X1 U14025 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10618) );
  INV_X1 U14026 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10628) );
  INV_X1 U14027 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U14028 ( .A1(n18095), .A2(n10622), .B1(n13880), .B2(n18084), .ZN(
        n10626) );
  INV_X1 U14029 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10624) );
  INV_X1 U14030 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10623) );
  OAI22_X1 U14031 ( .A1(n9588), .A2(n10624), .B1(n18123), .B2(n10623), .ZN(
        n10625) );
  INV_X4 U14032 ( .A(n18125), .ZN(n18232) );
  AOI22_X1 U14033 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U14034 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U14035 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U14036 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U14037 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10629) );
  NAND4_X1 U14038 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10633) );
  AOI22_X1 U14039 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U14040 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n18205), .ZN(n10641) );
  INV_X1 U14041 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U14042 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10635) );
  NAND2_X1 U14043 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10634) );
  OAI211_X1 U14044 ( .C1(n9603), .C2(n10636), .A(n10635), .B(n10634), .ZN(
        n10637) );
  INV_X1 U14045 ( .A(n10637), .ZN(n10640) );
  INV_X1 U14046 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10638) );
  NAND4_X1 U14047 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10648) );
  AOI22_X1 U14048 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U14049 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U14050 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U14051 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U14052 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10647) );
  AOI22_X1 U14053 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U14054 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10655) );
  INV_X1 U14055 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18013) );
  NAND2_X1 U14056 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10650) );
  NAND2_X1 U14057 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10649) );
  OAI211_X1 U14058 ( .C1(n9602), .C2(n18013), .A(n10650), .B(n10649), .ZN(
        n10651) );
  INV_X1 U14059 ( .A(n10651), .ZN(n10654) );
  INV_X1 U14060 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10652) );
  OR2_X1 U14061 ( .A1(n18227), .A2(n10652), .ZN(n10653) );
  NAND4_X1 U14062 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        n10662) );
  AOI22_X1 U14063 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U14064 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U14065 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U14066 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10657) );
  NAND4_X1 U14067 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10661) );
  AOI22_X1 U14068 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U14069 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10668) );
  INV_X1 U14070 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17995) );
  NAND2_X1 U14071 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U14072 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10663) );
  OAI211_X1 U14073 ( .C1(n9603), .C2(n17995), .A(n10664), .B(n10663), .ZN(
        n10665) );
  INV_X1 U14074 ( .A(n10665), .ZN(n10667) );
  OR2_X1 U14075 ( .A1(n18227), .A2(n21633), .ZN(n10666) );
  NAND4_X1 U14076 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10675) );
  AOI22_X1 U14077 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U14078 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U14079 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U14080 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U14081 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  AOI22_X1 U14082 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10682) );
  INV_X1 U14083 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18126) );
  NAND2_X1 U14084 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10677) );
  NAND2_X1 U14085 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10676) );
  OAI211_X1 U14086 ( .C1(n9602), .C2(n18126), .A(n10677), .B(n10676), .ZN(
        n10678) );
  INV_X1 U14087 ( .A(n10678), .ZN(n10680) );
  INV_X1 U14088 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18124) );
  OR2_X1 U14089 ( .A1(n18227), .A2(n18124), .ZN(n10679) );
  NAND4_X1 U14090 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n10688) );
  AOI22_X1 U14091 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U14092 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U14093 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U14094 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10683) );
  NAND4_X1 U14095 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10687) );
  NAND2_X1 U14096 ( .A1(n19122), .A2(n19127), .ZN(n10720) );
  NOR4_X2 U14097 ( .A1(n19111), .A2(n10727), .A3(n19117), .A4(n10720), .ZN(
        n10729) );
  AOI22_X1 U14098 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U14099 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10694) );
  INV_X1 U14100 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U14101 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10690) );
  NAND2_X1 U14102 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10689) );
  OAI211_X1 U14103 ( .C1(n9602), .C2(n18041), .A(n10690), .B(n10689), .ZN(
        n10691) );
  INV_X1 U14104 ( .A(n10691), .ZN(n10693) );
  OR2_X1 U14105 ( .A1(n18227), .A2(n17843), .ZN(n10692) );
  NAND4_X1 U14106 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10701) );
  AOI22_X1 U14107 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U14108 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U14109 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U14110 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10696) );
  NAND4_X1 U14111 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10700) );
  NAND2_X1 U14112 ( .A1(n19122), .A2(n10214), .ZN(n13832) );
  INV_X1 U14113 ( .A(n13832), .ZN(n10716) );
  NAND2_X1 U14114 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10703) );
  NAND2_X1 U14115 ( .A1(n18205), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10702) );
  OAI211_X1 U14116 ( .C1(n17882), .C2(n18227), .A(n10703), .B(n10702), .ZN(
        n10704) );
  INV_X1 U14117 ( .A(n10704), .ZN(n10708) );
  AOI22_X1 U14118 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13906), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U14119 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U14120 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10705) );
  NAND4_X1 U14121 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10714) );
  AOI22_X1 U14122 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14134), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U14123 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U14124 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U14125 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U14126 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  NOR2_X1 U14127 ( .A1(n17260), .A2(n19102), .ZN(n13648) );
  NAND2_X1 U14128 ( .A1(n14199), .A2(n19131), .ZN(n10715) );
  NAND2_X1 U14129 ( .A1(n13648), .A2(n10715), .ZN(n13631) );
  OAI21_X1 U14130 ( .B1(n10716), .B2(n10728), .A(n13631), .ZN(n10724) );
  INV_X1 U14131 ( .A(n19111), .ZN(n10725) );
  INV_X1 U14132 ( .A(n19117), .ZN(n10718) );
  INV_X1 U14133 ( .A(n14199), .ZN(n10717) );
  AOI22_X1 U14134 ( .A1(n10725), .A2(n10727), .B1(n10718), .B2(n10717), .ZN(
        n10723) );
  NAND2_X1 U14135 ( .A1(n19102), .A2(n17260), .ZN(n13650) );
  NAND2_X1 U14136 ( .A1(n10214), .A2(n13650), .ZN(n13625) );
  AOI21_X1 U14137 ( .B1(n19131), .B2(n10720), .A(n10718), .ZN(n10719) );
  AOI21_X1 U14138 ( .B1(n10720), .B2(n13625), .A(n10719), .ZN(n10722) );
  NOR2_X1 U14139 ( .A1(n19106), .A2(n10720), .ZN(n13833) );
  OAI21_X1 U14140 ( .B1(n10728), .B2(n13833), .A(n17260), .ZN(n10721) );
  NAND3_X1 U14141 ( .A1(n10723), .A2(n10722), .A3(n10721), .ZN(n13623) );
  NAND2_X1 U14142 ( .A1(n10729), .A2(n13603), .ZN(n13607) );
  NAND2_X1 U14143 ( .A1(n10725), .A2(n10214), .ZN(n13657) );
  INV_X1 U14144 ( .A(n13657), .ZN(n10726) );
  NOR2_X1 U14145 ( .A1(n13620), .A2(n19122), .ZN(n13626) );
  NAND2_X1 U14146 ( .A1(n10726), .A2(n13626), .ZN(n14192) );
  NOR2_X1 U14147 ( .A1(n10727), .A2(n14192), .ZN(n10730) );
  NAND2_X1 U14148 ( .A1(n10729), .A2(n19106), .ZN(n13629) );
  MUX2_X1 U14149 ( .A(n19095), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10737) );
  MUX2_X1 U14150 ( .A(n10732), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13617) );
  NAND2_X1 U14151 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19528), .ZN(
        n13615) );
  INV_X1 U14152 ( .A(n13615), .ZN(n10733) );
  NAND2_X1 U14153 ( .A1(n13617), .A2(n10733), .ZN(n10735) );
  NAND2_X1 U14154 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10732), .ZN(
        n10734) );
  NAND2_X1 U14155 ( .A1(n10735), .A2(n10734), .ZN(n10736) );
  NAND2_X1 U14156 ( .A1(n10736), .A2(n10737), .ZN(n10739) );
  OAI21_X1 U14157 ( .B1(n10737), .B2(n10736), .A(n10739), .ZN(n10750) );
  NAND2_X1 U14158 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19095), .ZN(
        n10738) );
  AOI21_X1 U14159 ( .B1(n10740), .B2(n19524), .A(n10742), .ZN(n10748) );
  OR2_X1 U14160 ( .A1(n10748), .A2(n19541), .ZN(n10744) );
  INV_X1 U14161 ( .A(n10740), .ZN(n10741) );
  NAND2_X1 U14162 ( .A1(n10741), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U14163 ( .A1(n10745), .A2(n10742), .ZN(n10743) );
  NAND2_X1 U14164 ( .A1(n10745), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10747) );
  NOR2_X1 U14165 ( .A1(n17752), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10746) );
  INV_X1 U14166 ( .A(n13617), .ZN(n10751) );
  XNOR2_X1 U14167 ( .A(n10751), .B(n13615), .ZN(n10752) );
  NAND2_X1 U14168 ( .A1(n10753), .A2(n10752), .ZN(n13835) );
  NOR2_X4 U14169 ( .A1(n19517), .A2(n18473), .ZN(n19695) );
  NOR2_X4 U14170 ( .A1(n21652), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19647) );
  NOR2_X1 U14171 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19572) );
  INV_X1 U14172 ( .A(n13830), .ZN(n19679) );
  INV_X1 U14173 ( .A(n19550), .ZN(n10754) );
  OR2_X2 U14174 ( .A1(n10763), .A2(n10754), .ZN(n17806) );
  INV_X1 U14175 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19608) );
  INV_X1 U14176 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19593) );
  NAND2_X1 U14177 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17795) );
  NOR2_X1 U14178 ( .A1(n19593), .A2(n17795), .ZN(n17755) );
  NAND2_X1 U14179 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n17712) );
  INV_X1 U14180 ( .A(n17712), .ZN(n10755) );
  NAND4_X1 U14181 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n17755), .A4(n10755), .ZN(n17703) );
  NOR2_X1 U14182 ( .A1(n19601), .A2(n17703), .ZN(n17678) );
  NAND4_X1 U14183 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17678), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17650) );
  NOR2_X1 U14184 ( .A1(n19608), .A2(n17650), .ZN(n17637) );
  NAND2_X1 U14185 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17637), .ZN(n10764) );
  NOR2_X2 U14186 ( .A1(n19613), .A2(n17634), .ZN(n17616) );
  NAND3_X1 U14187 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n10765) );
  INV_X1 U14188 ( .A(n17551), .ZN(n17563) );
  INV_X1 U14189 ( .A(n17531), .ZN(n17501) );
  NOR2_X2 U14190 ( .A1(n10766), .A2(n17501), .ZN(n17480) );
  NAND4_X1 U14191 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17480), .ZN(n11438) );
  INV_X1 U14192 ( .A(n19409), .ZN(n19560) );
  NOR2_X1 U14193 ( .A1(n17445), .A2(n19560), .ZN(n19555) );
  INV_X1 U14194 ( .A(n19555), .ZN(n10758) );
  NOR2_X1 U14195 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19693) );
  NOR2_X1 U14196 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n10757) );
  NAND3_X1 U14197 ( .A1(n10758), .A2(n19075), .A3(n19566), .ZN(n10759) );
  OAI22_X1 U14198 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n11438), .B1(n10310), 
        .B2(n17801), .ZN(n10772) );
  AND2_X1 U14199 ( .A1(n19102), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n10760) );
  OR2_X1 U14200 ( .A1(n19550), .A2(n10760), .ZN(n10761) );
  NAND2_X1 U14201 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19102), .ZN(n10762) );
  AOI211_X4 U14202 ( .C1(n19680), .C2(n19682), .A(n10763), .B(n10762), .ZN(
        n17774) );
  NAND2_X1 U14203 ( .A1(n17778), .A2(n18257), .ZN(n17773) );
  NAND2_X1 U14204 ( .A1(n17754), .A2(n17744), .ZN(n17737) );
  INV_X1 U14205 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17719) );
  INV_X1 U14206 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17695) );
  INV_X1 U14207 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17670) );
  NAND2_X1 U14208 ( .A1(n17679), .A2(n17670), .ZN(n17669) );
  NAND2_X1 U14209 ( .A1(n17601), .A2(n18075), .ZN(n17589) );
  INV_X1 U14210 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18038) );
  INV_X1 U14211 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17518) );
  INV_X1 U14212 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17497) );
  NAND2_X1 U14213 ( .A1(n17503), .A2(n17497), .ZN(n17496) );
  INV_X1 U14214 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17943) );
  NOR2_X1 U14215 ( .A1(n17805), .A2(n10768), .ZN(n11439) );
  OAI21_X1 U14216 ( .B1(n17800), .B2(n11439), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n10770) );
  NOR3_X1 U14217 ( .A1(n17785), .A2(n19613), .A3(n10764), .ZN(n17635) );
  NAND4_X1 U14218 ( .A1(n17635), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n17564) );
  NOR2_X1 U14219 ( .A1(n17564), .A2(n10765), .ZN(n13260) );
  NAND4_X1 U14220 ( .A1(n13260), .A2(P3_REIP_REG_23__SCAN_IN), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n17519) );
  NOR2_X1 U14221 ( .A1(n17519), .A2(n10766), .ZN(n17479) );
  INV_X1 U14222 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19644) );
  NAND2_X1 U14223 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17487) );
  NOR2_X1 U14224 ( .A1(n19644), .A2(n17487), .ZN(n10767) );
  NAND2_X1 U14225 ( .A1(n17812), .A2(n17806), .ZN(n17594) );
  AOI21_X1 U14226 ( .B1(n17479), .B2(n10767), .A(n17592), .ZN(n17467) );
  NAND2_X1 U14227 ( .A1(n17467), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10769) );
  NAND3_X1 U14228 ( .A1(n10770), .A2(n10769), .A3(n9724), .ZN(n10771) );
  OR2_X1 U14229 ( .A1(n10774), .A2(n10773), .ZN(P3_U2641) );
  NAND2_X1 U14230 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20531), .ZN(
        n10791) );
  OAI21_X1 U14231 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20531), .A(
        n10791), .ZN(n10893) );
  INV_X1 U14232 ( .A(n10791), .ZN(n10775) );
  NAND2_X1 U14233 ( .A1(n10894), .A2(n10775), .ZN(n10777) );
  NAND2_X1 U14234 ( .A1(n20521), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U14235 ( .A1(n10777), .A2(n10776), .ZN(n10781) );
  NAND2_X1 U14236 ( .A1(n10781), .A2(n10780), .ZN(n10779) );
  NAND2_X1 U14237 ( .A1(n20512), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10778) );
  NAND2_X1 U14238 ( .A1(n10779), .A2(n10778), .ZN(n10784) );
  XNOR2_X1 U14239 ( .A(n10784), .B(n10783), .ZN(n12642) );
  XNOR2_X1 U14240 ( .A(n10781), .B(n10780), .ZN(n12641) );
  NOR2_X1 U14241 ( .A1(n14341), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10782) );
  NOR2_X1 U14242 ( .A1(n17317), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10785) );
  INV_X1 U14243 ( .A(n10792), .ZN(n10794) );
  INV_X1 U14244 ( .A(n10786), .ZN(n10788) );
  NAND2_X1 U14245 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13342), .ZN(
        n10789) );
  XNOR2_X1 U14246 ( .A(n10894), .B(n10791), .ZN(n12636) );
  AND2_X1 U14247 ( .A1(n12636), .A2(n10792), .ZN(n10793) );
  OAI21_X1 U14248 ( .B1(n10893), .B2(n10794), .A(n13330), .ZN(n10796) );
  AND2_X2 U14249 ( .A1(n16202), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15993) );
  INV_X1 U14250 ( .A(n15993), .ZN(n10795) );
  NOR2_X1 U14251 ( .A1(n14110), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13338) );
  AOI21_X1 U14252 ( .B1(n10795), .B2(n13338), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n20524) );
  MUX2_X1 U14253 ( .A(n10796), .B(n20524), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20538) );
  INV_X2 U14254 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14334) );
  AND3_X4 U14255 ( .A1(n10797), .A2(n14334), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U14256 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10803) );
  INV_X1 U14257 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U14258 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U14259 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U14260 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U14261 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U14262 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16197), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U14263 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U14264 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U14265 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U14266 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U14267 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10811) );
  NAND4_X1 U14268 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n10824) );
  NAND2_X1 U14269 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10817) );
  NAND2_X1 U14270 ( .A1(n10817), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10818) );
  AOI21_X1 U14271 ( .B1(n10876), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n10818), .ZN(n10822) );
  AOI22_X1 U14272 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U14273 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U14274 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U14275 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  AOI22_X1 U14276 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10828) );
  AOI21_X1 U14277 ( .B1(n10876), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n10825), .ZN(n10827) );
  AOI22_X1 U14278 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U14279 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U14280 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U14281 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U14282 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U14283 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U14284 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U14285 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U14286 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U14287 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U14288 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U14289 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U14290 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U14291 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U14292 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U14293 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U14294 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U14295 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U14296 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U14297 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U14298 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U14299 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U14300 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10857) );
  AOI21_X1 U14301 ( .B1(n10876), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n10855), .ZN(n10856) );
  AOI22_X1 U14302 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U14303 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U14304 ( .A1(n16026), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U14305 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U14306 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10864) );
  AOI22_X1 U14307 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U14308 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U14309 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U14310 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10865) );
  NAND4_X1 U14311 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10869) );
  AOI22_X1 U14312 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14106), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U14313 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U14314 ( .A1(n10876), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14315 ( .A1(n16086), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U14316 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10876), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U14317 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U14318 ( .A1(n14363), .A2(n12645), .ZN(n12914) );
  AOI22_X1 U14319 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n16041), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10885) );
  AND2_X2 U14320 ( .A1(n14106), .A2(n14341), .ZN(n14107) );
  AOI22_X1 U14321 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11026), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U14322 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10990), .B1(
        n11125), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10883) );
  AND2_X2 U14323 ( .A1(n10881), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11039) );
  AOI22_X1 U14324 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10882) );
  AND2_X2 U14325 ( .A1(n10809), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12756) );
  AOI22_X1 U14326 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10888) );
  AND2_X2 U14327 ( .A1(n16202), .A2(n14341), .ZN(n11069) );
  AOI22_X1 U14328 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11069), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U14329 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U14330 ( .A1(n16048), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14409), .ZN(n10890) );
  NAND2_X1 U14331 ( .A1(n10892), .A2(n10891), .ZN(n11245) );
  INV_X1 U14332 ( .A(n10893), .ZN(n12637) );
  NAND2_X1 U14333 ( .A1(n10894), .A2(n12637), .ZN(n12635) );
  NAND2_X1 U14334 ( .A1(n11245), .A2(n12635), .ZN(n10895) );
  NOR2_X1 U14335 ( .A1(n12644), .A2(n12642), .ZN(n12643) );
  AOI21_X1 U14336 ( .B1(n10895), .B2(n12643), .A(n12649), .ZN(n20534) );
  NAND2_X1 U14337 ( .A1(n20534), .A2(n20536), .ZN(n12667) );
  OAI21_X1 U14338 ( .B1(n20538), .B2(n12914), .A(n12667), .ZN(n10896) );
  INV_X1 U14339 ( .A(n19708), .ZN(n10897) );
  INV_X1 U14340 ( .A(n12656), .ZN(n12647) );
  INV_X1 U14341 ( .A(n10902), .ZN(n10904) );
  OAI21_X1 U14342 ( .B1(n10906), .B2(n10905), .A(n10911), .ZN(n12682) );
  INV_X1 U14343 ( .A(n12656), .ZN(n10907) );
  NAND2_X1 U14344 ( .A1(n10907), .A2(n19879), .ZN(n10921) );
  NAND2_X1 U14345 ( .A1(n10921), .A2(n9999), .ZN(n10908) );
  INV_X2 U14346 ( .A(n17030), .ZN(n20550) );
  INV_X1 U14347 ( .A(n12679), .ZN(n14364) );
  NAND2_X1 U14348 ( .A1(n19879), .A2(n19875), .ZN(n13530) );
  NOR2_X1 U14349 ( .A1(n13530), .A2(n11246), .ZN(n10913) );
  NAND2_X1 U14350 ( .A1(n14364), .A2(n10545), .ZN(n12675) );
  AOI22_X1 U14351 ( .A1(n12675), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n14382), .ZN(n10914) );
  NAND2_X1 U14352 ( .A1(n10915), .A2(n10914), .ZN(n10928) );
  INV_X1 U14353 ( .A(n10928), .ZN(n10926) );
  NAND2_X1 U14354 ( .A1(n10918), .A2(n10912), .ZN(n10919) );
  INV_X1 U14355 ( .A(n10921), .ZN(n10922) );
  NAND2_X1 U14356 ( .A1(n12660), .A2(n20557), .ZN(n14385) );
  NAND2_X1 U14357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U14358 ( .A1(n10926), .A2(n10927), .ZN(n10943) );
  INV_X1 U14359 ( .A(n10927), .ZN(n10929) );
  NAND2_X1 U14360 ( .A1(n10931), .A2(n10932), .ZN(n14335) );
  AOI22_X1 U14361 ( .A1(n14335), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14382), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U14362 ( .A1(n10934), .A2(n10933), .ZN(n10954) );
  INV_X1 U14363 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19722) );
  INV_X1 U14364 ( .A(n14382), .ZN(n20544) );
  NAND2_X1 U14365 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10935) );
  OAI211_X1 U14366 ( .C1(n10950), .C2(n19722), .A(n20544), .B(n10935), .ZN(
        n10937) );
  INV_X1 U14367 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11249) );
  NOR2_X1 U14368 ( .A1(n10937), .A2(n10936), .ZN(n10939) );
  NAND2_X1 U14369 ( .A1(n11158), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10941) );
  OAI21_X1 U14370 ( .B1(n20512), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16992), 
        .ZN(n10944) );
  NAND2_X1 U14371 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10946) );
  OR2_X1 U14372 ( .A1(n10950), .A2(n20431), .ZN(n10945) );
  OAI211_X1 U14373 ( .C1(n11229), .C2(n11247), .A(n10946), .B(n10945), .ZN(
        n10947) );
  NOR2_X1 U14374 ( .A1(n20544), .A2(n20505), .ZN(n10949) );
  INV_X1 U14375 ( .A(n10954), .ZN(n10957) );
  INV_X1 U14376 ( .A(n10955), .ZN(n10956) );
  NAND2_X1 U14377 ( .A1(n10975), .A2(n13425), .ZN(n10966) );
  INV_X1 U14378 ( .A(n10966), .ZN(n10961) );
  INV_X1 U14379 ( .A(n10958), .ZN(n10974) );
  NAND2_X1 U14380 ( .A1(n10974), .A2(n10959), .ZN(n10960) );
  BUF_X4 U14381 ( .A(n10962), .Z(n14022) );
  INV_X2 U14382 ( .A(n10975), .ZN(n13240) );
  INV_X1 U14383 ( .A(n15946), .ZN(n10965) );
  NOR2_X2 U14384 ( .A1(n10967), .A2(n14010), .ZN(n11051) );
  OR2_X2 U14385 ( .A1(n10966), .A2(n15946), .ZN(n10968) );
  NOR2_X2 U14386 ( .A1(n14022), .A2(n10968), .ZN(n11052) );
  AOI22_X1 U14387 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11051), .B1(
        n11052), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10972) );
  NOR2_X2 U14388 ( .A1(n10967), .A2(n14022), .ZN(n11077) );
  NOR2_X2 U14389 ( .A1(n14010), .A2(n10968), .ZN(n11055) );
  AOI22_X1 U14390 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11055), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U14391 ( .A1(n10562), .A2(n15946), .ZN(n10969) );
  NOR2_X2 U14392 ( .A1(n10969), .A2(n14010), .ZN(n11053) );
  NOR2_X2 U14393 ( .A1(n14022), .A2(n10969), .ZN(n11054) );
  AOI22_X1 U14394 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11053), .B1(
        n11054), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10970) );
  INV_X1 U14395 ( .A(n13425), .ZN(n15962) );
  AND2_X1 U14396 ( .A1(n15962), .A2(n10974), .ZN(n10979) );
  AND2_X1 U14397 ( .A1(n13240), .A2(n10979), .ZN(n10985) );
  BUF_X1 U14398 ( .A(n10975), .Z(n14333) );
  INV_X1 U14399 ( .A(n10976), .ZN(n10977) );
  NOR2_X1 U14400 ( .A1(n10978), .A2(n10977), .ZN(n10981) );
  AND2_X1 U14401 ( .A1(n14333), .A2(n10981), .ZN(n10980) );
  AOI22_X1 U14402 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11059), .B1(
        n11060), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10989) );
  AND2_X1 U14403 ( .A1(n14333), .A2(n10979), .ZN(n10984) );
  AOI22_X1 U14404 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11082), .B1(
        n20349), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10988) );
  AND2_X1 U14405 ( .A1(n13240), .A2(n10981), .ZN(n10982) );
  INV_X1 U14406 ( .A(n10982), .ZN(n10983) );
  NOR2_X1 U14407 ( .A1(n14022), .A2(n10983), .ZN(n11058) );
  AOI22_X1 U14408 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11057), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U14409 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20261), .B1(
        n20139), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14410 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16041), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14411 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14107), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U14412 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10990), .B1(
        n11125), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U14413 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11069), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10991) );
  NAND4_X1 U14414 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n11002) );
  AOI22_X1 U14415 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14416 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14417 ( .A1(n15993), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14418 ( .A1(n11091), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14409), .ZN(n10997) );
  NAND4_X1 U14419 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11001) );
  AOI22_X1 U14420 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17022), .B1(
        n11051), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11005) );
  AOI21_X1 U14421 ( .B1(n11058), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n16235), .ZN(n11004) );
  AND2_X1 U14422 ( .A1(n11005), .A2(n11004), .ZN(n11009) );
  AOI22_X1 U14423 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11055), .B1(
        n11052), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14424 ( .A1(n11054), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11007) );
  AOI22_X1 U14425 ( .A1(n11077), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n20139), .ZN(n11013) );
  AOI22_X1 U14426 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11057), .B1(
        n20349), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14427 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11082), .B1(
        n11059), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U14428 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11060), .B1(
        n20261), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14107), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14430 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16041), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14431 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10990), .B1(
        n11125), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14432 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11044), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11014) );
  NAND4_X1 U14433 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11025) );
  NAND2_X1 U14434 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14435 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11018) );
  AND2_X1 U14436 ( .A1(n11019), .A2(n11018), .ZN(n11023) );
  AOI22_X1 U14437 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14438 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14439 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n14409), .ZN(n11020) );
  NAND4_X1 U14440 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11024) );
  AOI22_X1 U14441 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16041), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14442 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14107), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10990), .B1(
        n11125), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14444 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11027) );
  NAND4_X1 U14445 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11036) );
  AOI22_X1 U14446 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14409), .ZN(n11034) );
  AOI22_X1 U14447 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14448 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14449 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9589), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U14450 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11035) );
  INV_X1 U14451 ( .A(n11104), .ZN(n11037) );
  INV_X1 U14452 ( .A(n11105), .ZN(n12709) );
  NAND2_X1 U14453 ( .A1(n11037), .A2(n12709), .ZN(n11038) );
  AOI22_X1 U14454 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n16041), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U14455 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11026), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U14456 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U14457 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U14458 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n11050) );
  AOI22_X1 U14459 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14409), .ZN(n11048) );
  AOI22_X1 U14460 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11069), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U14461 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14462 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n16048), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11045) );
  NAND4_X1 U14463 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11049) );
  AOI22_X1 U14464 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n11057), .B1(
        n20204), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14465 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11082), .B1(
        n20349), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11059), .B1(
        n11060), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14467 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20261), .B1(
        n20139), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14468 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n16041), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14469 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n14107), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14471 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U14472 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11075) );
  AOI22_X1 U14473 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n14409), .ZN(n11073) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n11091), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14475 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14476 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n11069), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11070) );
  NAND4_X1 U14477 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11074) );
  NOR2_X1 U14478 ( .A1(n11075), .A2(n11074), .ZN(n12727) );
  NAND2_X1 U14479 ( .A1(n12727), .A2(n16235), .ZN(n11076) );
  AOI22_X1 U14480 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11077), .B1(
        n11052), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14481 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11051), .B1(
        n11055), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n17022), .B1(
        n11054), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11082), .B1(
        n20204), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14484 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11057), .B1(
        n20349), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11059), .B1(
        n11060), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20261), .B1(
        n20139), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11026), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14489 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14490 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11087) );
  NAND4_X1 U14491 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11097) );
  AOI22_X1 U14492 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14409), .ZN(n11095) );
  AOI22_X1 U14493 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14494 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n16048), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11092) );
  NAND4_X1 U14496 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n11096) );
  NAND2_X1 U14497 ( .A1(n12731), .A2(n16235), .ZN(n11098) );
  INV_X1 U14498 ( .A(n11252), .ZN(n12723) );
  NAND2_X1 U14499 ( .A1(n11114), .A2(n16703), .ZN(n11112) );
  INV_X1 U14500 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13237) );
  INV_X1 U14501 ( .A(n11291), .ZN(n12690) );
  XNOR2_X1 U14502 ( .A(n12690), .B(n12701), .ZN(n11102) );
  INV_X1 U14503 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13287) );
  NOR2_X1 U14504 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  NAND2_X1 U14505 ( .A1(n11102), .A2(n13289), .ZN(n11103) );
  XOR2_X1 U14506 ( .A(n11102), .B(n13289), .Z(n13361) );
  NAND2_X1 U14507 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13361), .ZN(
        n13360) );
  NAND2_X1 U14508 ( .A1(n11103), .A2(n13360), .ZN(n11106) );
  XNOR2_X1 U14509 ( .A(n13237), .B(n11106), .ZN(n13251) );
  XNOR2_X1 U14510 ( .A(n11105), .B(n11104), .ZN(n13250) );
  NAND2_X1 U14511 ( .A1(n13251), .A2(n13250), .ZN(n13249) );
  NAND2_X1 U14512 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11106), .ZN(
        n11107) );
  NAND2_X1 U14513 ( .A1(n13249), .A2(n11107), .ZN(n11108) );
  INV_X1 U14514 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17354) );
  XNOR2_X1 U14515 ( .A(n11108), .B(n17354), .ZN(n16708) );
  NAND2_X1 U14516 ( .A1(n11108), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14517 ( .A1(n11112), .A2(n11115), .ZN(n11110) );
  INV_X1 U14518 ( .A(n11115), .ZN(n11111) );
  INV_X1 U14519 ( .A(n11119), .ZN(n16678) );
  NAND2_X1 U14520 ( .A1(n16678), .A2(n11324), .ZN(n11113) );
  NAND2_X1 U14521 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14522 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14523 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14409), .ZN(
        n11122) );
  NAND2_X1 U14524 ( .A1(n11091), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14525 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14526 ( .A1(n15993), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U14527 ( .A1(n11125), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14528 ( .A1(n10990), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14529 ( .A1(n16042), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14530 ( .A1(n11026), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14531 ( .A1(n16041), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14532 ( .A1(n14107), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14533 ( .A1(n11044), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14534 ( .A1(n16048), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14535 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14536 ( .A1(n10996), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11134) );
  NAND4_X1 U14537 ( .A1(n11141), .A2(n11140), .A3(n11139), .A4(n11138), .ZN(
        n11254) );
  INV_X1 U14538 ( .A(n11254), .ZN(n11143) );
  OAI21_X1 U14539 ( .B1(n11144), .B2(n11143), .A(n21729), .ZN(n11145) );
  NAND2_X1 U14540 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16524) );
  NAND2_X1 U14541 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11147) );
  NOR2_X1 U14542 ( .A1(n16524), .A2(n11147), .ZN(n12896) );
  NAND2_X1 U14543 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U14544 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16885) );
  NOR2_X1 U14545 ( .A1(n12892), .A2(n16885), .ZN(n12632) );
  AND2_X1 U14546 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13118) );
  NAND4_X1 U14547 ( .A1(n12896), .A2(n12632), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n13118), .ZN(n11148) );
  NAND2_X1 U14548 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16769) );
  NAND2_X1 U14549 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16753) );
  NOR2_X1 U14550 ( .A1(n16769), .A2(n16753), .ZN(n11149) );
  AND2_X1 U14551 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16451) );
  NAND2_X1 U14552 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13123) );
  INV_X1 U14553 ( .A(n11150), .ZN(n11152) );
  INV_X1 U14554 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U14555 ( .A1(n12928), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U14556 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11153) );
  OAI211_X1 U14557 ( .C1(n11229), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11156) );
  AOI21_X1 U14558 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11156), .ZN(n14208) );
  INV_X1 U14559 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n15902) );
  INV_X1 U14560 ( .A(n11158), .ZN(n11235) );
  OR2_X1 U14561 ( .A1(n11235), .A2(n16703), .ZN(n11160) );
  AOI22_X1 U14562 ( .A1(n12928), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11159) );
  OAI211_X1 U14563 ( .C1(n12930), .C2(n15902), .A(n11160), .B(n11159), .ZN(
        n14044) );
  INV_X1 U14564 ( .A(n14044), .ZN(n11161) );
  NOR2_X1 U14565 ( .A1(n14208), .A2(n11161), .ZN(n11162) );
  INV_X1 U14566 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U14567 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11164) );
  INV_X1 U14568 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20438) );
  OR2_X1 U14569 ( .A1(n11221), .A2(n20438), .ZN(n11163) );
  OAI211_X1 U14570 ( .C1(n11229), .C2(n14280), .A(n11164), .B(n11163), .ZN(
        n11165) );
  AOI21_X1 U14571 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11165), .ZN(n14278) );
  INV_X1 U14572 ( .A(n14278), .ZN(n11166) );
  INV_X1 U14573 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U14574 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11168) );
  INV_X1 U14575 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20440) );
  OR2_X1 U14576 ( .A1(n11221), .A2(n20440), .ZN(n11167) );
  OAI211_X1 U14577 ( .C1(n11229), .C2(n11255), .A(n11168), .B(n11167), .ZN(
        n11169) );
  AOI21_X1 U14578 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11169), .ZN(n14290) );
  OR2_X1 U14579 ( .A1(n11235), .A2(n21729), .ZN(n11171) );
  AOI22_X1 U14580 ( .A1(n12928), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11170) );
  OAI211_X1 U14581 ( .C1(n11229), .C2(n15864), .A(n11171), .B(n11170), .ZN(
        n15855) );
  NAND2_X1 U14582 ( .A1(n15856), .A2(n15855), .ZN(n15848) );
  NAND2_X1 U14583 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11173) );
  INV_X1 U14584 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20444) );
  OR2_X1 U14585 ( .A1(n11221), .A2(n20444), .ZN(n11172) );
  OAI211_X1 U14586 ( .C1(n12930), .C2(n10497), .A(n11173), .B(n11172), .ZN(
        n11174) );
  AOI21_X1 U14587 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11174), .ZN(n15849) );
  INV_X1 U14588 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n16299) );
  NAND2_X1 U14589 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11177) );
  INV_X1 U14590 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20446) );
  OR2_X1 U14591 ( .A1(n11221), .A2(n20446), .ZN(n11176) );
  OAI211_X1 U14592 ( .C1(n11229), .C2(n16299), .A(n11177), .B(n11176), .ZN(
        n11178) );
  AOI21_X1 U14593 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11178), .ZN(n15832) );
  OR2_X1 U14594 ( .A1(n11235), .A2(n16914), .ZN(n11180) );
  AOI22_X1 U14595 ( .A1(n12928), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11179) );
  OAI211_X1 U14596 ( .C1(n11229), .C2(n13273), .A(n11180), .B(n11179), .ZN(
        n13279) );
  INV_X1 U14597 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14598 ( .A1(n12928), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14599 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11181) );
  OAI211_X1 U14600 ( .C1(n12930), .C2(n11258), .A(n11182), .B(n11181), .ZN(
        n11183) );
  AOI21_X1 U14601 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11183), .ZN(n13060) );
  INV_X1 U14602 ( .A(n13060), .ZN(n11187) );
  INV_X1 U14603 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11186) );
  INV_X1 U14604 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16901) );
  OR2_X1 U14605 ( .A1(n11235), .A2(n16901), .ZN(n11185) );
  AOI22_X1 U14606 ( .A1(n12928), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11184) );
  OAI211_X1 U14607 ( .C1(n12930), .C2(n11186), .A(n11185), .B(n11184), .ZN(
        n14080) );
  AND2_X1 U14608 ( .A1(n11187), .A2(n14080), .ZN(n11188) );
  NAND2_X1 U14609 ( .A1(n13057), .A2(n11188), .ZN(n13058) );
  INV_X1 U14610 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U14611 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11190) );
  INV_X1 U14612 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20453) );
  OR2_X1 U14613 ( .A1(n11221), .A2(n20453), .ZN(n11189) );
  OAI211_X1 U14614 ( .C1(n12930), .C2(n15793), .A(n11190), .B(n11189), .ZN(
        n11191) );
  AOI21_X1 U14615 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11191), .ZN(n14295) );
  INV_X1 U14616 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11377) );
  OR2_X1 U14617 ( .A1(n11235), .A2(n16875), .ZN(n11193) );
  AOI22_X1 U14618 ( .A1(n12928), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11192) );
  OAI211_X1 U14619 ( .C1(n12930), .C2(n11377), .A(n11193), .B(n11192), .ZN(
        n14396) );
  INV_X1 U14620 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n16288) );
  NAND2_X1 U14621 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11195) );
  INV_X1 U14622 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20457) );
  OR2_X1 U14623 ( .A1(n11221), .A2(n20457), .ZN(n11194) );
  OAI211_X1 U14624 ( .C1(n12930), .C2(n16288), .A(n11195), .B(n11194), .ZN(
        n11196) );
  AOI21_X1 U14625 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11196), .ZN(n15770) );
  INV_X1 U14626 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U14627 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11198) );
  OR2_X1 U14628 ( .A1(n11221), .A2(n20459), .ZN(n11197) );
  OAI211_X1 U14629 ( .C1(n12930), .C2(n11199), .A(n11198), .B(n11197), .ZN(
        n11200) );
  AOI21_X1 U14630 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11200), .ZN(n15758) );
  INV_X1 U14631 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14632 ( .A1(n12928), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U14633 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11202) );
  OAI211_X1 U14634 ( .C1(n11229), .C2(n11261), .A(n11203), .B(n11202), .ZN(
        n11204) );
  AOI21_X1 U14635 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11204), .ZN(n15738) );
  INV_X1 U14636 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15729) );
  INV_X1 U14637 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16825) );
  OR2_X1 U14638 ( .A1(n11235), .A2(n16825), .ZN(n11206) );
  AOI22_X1 U14639 ( .A1(n12928), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11205) );
  OAI211_X1 U14640 ( .C1(n11229), .C2(n15729), .A(n11206), .B(n11205), .ZN(
        n15724) );
  INV_X1 U14641 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14642 ( .A1(n12928), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14643 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11207) );
  OAI211_X1 U14644 ( .C1(n12930), .C2(n11209), .A(n11208), .B(n11207), .ZN(
        n11210) );
  AOI21_X1 U14645 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11210), .ZN(n12673) );
  INV_X1 U14646 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15712) );
  NAND2_X1 U14647 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11212) );
  INV_X1 U14648 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20464) );
  OR2_X1 U14649 ( .A1(n11221), .A2(n20464), .ZN(n11211) );
  OAI211_X1 U14650 ( .C1(n12930), .C2(n15712), .A(n11212), .B(n11211), .ZN(
        n11213) );
  AOI21_X1 U14651 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11213), .ZN(n15705) );
  NOR2_X2 U14652 ( .A1(n9615), .A2(n15705), .ZN(n15688) );
  INV_X1 U14653 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15697) );
  OR2_X1 U14654 ( .A1(n11235), .A2(n16798), .ZN(n11215) );
  AOI22_X1 U14655 ( .A1(n12928), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11214) );
  OAI211_X1 U14656 ( .C1(n15697), .C2(n12930), .A(n11215), .B(n11214), .ZN(
        n15687) );
  INV_X1 U14657 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11262) );
  OR2_X1 U14658 ( .A1(n11235), .A2(n21670), .ZN(n11217) );
  AOI22_X1 U14659 ( .A1(n12928), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11216) );
  OAI211_X1 U14660 ( .C1(n11262), .C2(n11229), .A(n11217), .B(n11216), .ZN(
        n15675) );
  INV_X1 U14661 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U14662 ( .A1(n12928), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U14663 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11218) );
  OAI211_X1 U14664 ( .C1(n12930), .C2(n11268), .A(n11219), .B(n11218), .ZN(
        n11220) );
  AOI21_X1 U14665 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11220), .ZN(n15657) );
  INV_X1 U14666 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n21691) );
  NAND2_X1 U14667 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11223) );
  INV_X1 U14668 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20471) );
  OR2_X1 U14669 ( .A1(n11221), .A2(n20471), .ZN(n11222) );
  OAI211_X1 U14670 ( .C1(n12930), .C2(n21691), .A(n11223), .B(n11222), .ZN(
        n11224) );
  AOI21_X1 U14671 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11224), .ZN(n13143) );
  INV_X1 U14672 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16240) );
  INV_X1 U14673 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16758) );
  OR2_X1 U14674 ( .A1(n11235), .A2(n16758), .ZN(n11226) );
  AOI22_X1 U14675 ( .A1(n12928), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11225) );
  OAI211_X1 U14676 ( .C1(n16240), .C2(n11229), .A(n11226), .B(n11225), .ZN(
        n15630) );
  INV_X1 U14677 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15623) );
  OR2_X1 U14678 ( .A1(n11235), .A2(n16745), .ZN(n11228) );
  AOI22_X1 U14679 ( .A1(n12928), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11227) );
  OAI211_X1 U14680 ( .C1(n15623), .C2(n12930), .A(n11228), .B(n11227), .ZN(
        n15615) );
  INV_X1 U14681 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16728) );
  AOI22_X1 U14682 ( .A1(n12928), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11231) );
  NAND2_X1 U14683 ( .A1(n11157), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11230) );
  OAI211_X1 U14684 ( .C1(n11235), .C2(n16728), .A(n11231), .B(n11230), .ZN(
        n15601) );
  INV_X1 U14685 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14686 ( .A1(n12928), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11232) );
  OAI21_X1 U14687 ( .B1(n12930), .B2(n11233), .A(n11232), .ZN(n11234) );
  AOI21_X1 U14688 ( .B1(n12932), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11234), .ZN(n15583) );
  INV_X1 U14689 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11238) );
  INV_X1 U14690 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13163) );
  OR2_X1 U14691 ( .A1(n11235), .A2(n13163), .ZN(n11237) );
  AOI22_X1 U14692 ( .A1(n12928), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11236) );
  OAI211_X1 U14693 ( .C1(n11238), .C2(n12930), .A(n11237), .B(n11236), .ZN(
        n12927) );
  NAND2_X1 U14694 ( .A1(n16992), .A2(n20501), .ZN(n20493) );
  NAND2_X1 U14695 ( .A1(n20493), .A2(n20543), .ZN(n20515) );
  NAND2_X1 U14696 ( .A1(n20515), .A2(n20559), .ZN(n11239) );
  AND2_X1 U14697 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20516) );
  NOR2_X1 U14698 ( .A1(n16211), .A2(n16682), .ZN(n11244) );
  NAND2_X1 U14699 ( .A1(n12962), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12964) );
  NAND2_X1 U14700 ( .A1(n12989), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12993) );
  NAND2_X1 U14701 ( .A1(n13000), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12937) );
  INV_X1 U14702 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13107) );
  XNOR2_X1 U14703 ( .A(n12937), .B(n13107), .ZN(n13092) );
  NAND2_X1 U14704 ( .A1(n20356), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U14705 ( .A1(n13735), .A2(n13005), .ZN(n13675) );
  NAND2_X2 U14706 ( .A1(n17050), .A2(n13006), .ZN(n17339) );
  NAND2_X1 U14707 ( .A1(n19745), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U14708 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11242) );
  OAI211_X1 U14709 ( .C1(n13092), .C2(n16717), .A(n13126), .B(n11242), .ZN(
        n11243) );
  INV_X1 U14710 ( .A(n11245), .ZN(n11248) );
  OAI21_X1 U14711 ( .B1(n11248), .B2(n12689), .A(n10557), .ZN(n11297) );
  MUX2_X1 U14712 ( .A(n12718), .B(n11251), .S(n12689), .Z(n11307) );
  MUX2_X1 U14713 ( .A(n11252), .B(n15902), .S(n12689), .Z(n11302) );
  MUX2_X1 U14714 ( .A(n12727), .B(P2_EBX_REG_5__SCAN_IN), .S(n12689), .Z(
        n11283) );
  MUX2_X1 U14715 ( .A(n11253), .B(n14280), .S(n12689), .Z(n11327) );
  MUX2_X1 U14716 ( .A(n11255), .B(n11254), .S(n19868), .Z(n11335) );
  NOR2_X1 U14717 ( .A1(n19868), .A2(n15864), .ZN(n11333) );
  NAND2_X1 U14718 ( .A1(n11373), .A2(n13273), .ZN(n11370) );
  NAND2_X1 U14719 ( .A1(n12689), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11369) );
  NOR2_X1 U14720 ( .A1(n19868), .A2(n11258), .ZN(n11381) );
  NOR2_X1 U14721 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n11259) );
  NOR2_X1 U14722 ( .A1(n19868), .A2(n11259), .ZN(n11260) );
  NAND2_X1 U14723 ( .A1(n12689), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11358) );
  NOR2_X1 U14724 ( .A1(n19868), .A2(n15729), .ZN(n11351) );
  NAND2_X1 U14725 ( .A1(n11278), .A2(n11419), .ZN(n11356) );
  NAND2_X1 U14726 ( .A1(n12689), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11277) );
  NOR2_X1 U14727 ( .A1(n19868), .A2(n11262), .ZN(n11274) );
  INV_X1 U14728 ( .A(n11414), .ZN(n13034) );
  OAI21_X1 U14729 ( .B1(n15641), .B2(n11143), .A(n16758), .ZN(n11267) );
  NAND2_X1 U14730 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11266) );
  NOR2_X1 U14731 ( .A1(n19868), .A2(n11268), .ZN(n11269) );
  INV_X1 U14732 ( .A(n11419), .ZN(n11361) );
  AOI21_X1 U14733 ( .B1(n11270), .B2(n11269), .A(n11361), .ZN(n11271) );
  AND2_X1 U14734 ( .A1(n11271), .A2(n15644), .ZN(n15665) );
  INV_X1 U14735 ( .A(n11276), .ZN(n11272) );
  INV_X1 U14736 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U14737 ( .A1(n11272), .A2(n13121), .ZN(n16473) );
  INV_X1 U14738 ( .A(n11274), .ZN(n11275) );
  XNOR2_X1 U14739 ( .A(n11273), .B(n11275), .ZN(n15684) );
  INV_X1 U14740 ( .A(n16471), .ZN(n16472) );
  NAND2_X1 U14741 ( .A1(n16472), .A2(n21670), .ZN(n13137) );
  AND2_X1 U14742 ( .A1(n16473), .A2(n13137), .ZN(n11413) );
  NAND2_X1 U14743 ( .A1(n11276), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16474) );
  NAND2_X1 U14744 ( .A1(n11278), .A2(n10350), .ZN(n11279) );
  NAND2_X1 U14745 ( .A1(n11273), .A2(n11279), .ZN(n15701) );
  NAND2_X1 U14746 ( .A1(n16493), .A2(n21670), .ZN(n11280) );
  NAND2_X1 U14747 ( .A1(n11280), .A2(n16471), .ZN(n11281) );
  AND2_X1 U14748 ( .A1(n16474), .A2(n11281), .ZN(n13138) );
  NAND2_X1 U14749 ( .A1(n11282), .A2(n11283), .ZN(n11284) );
  NAND2_X1 U14750 ( .A1(n9628), .A2(n11284), .ZN(n15890) );
  AND2_X1 U14751 ( .A1(n15890), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14752 ( .A1(n11322), .A2(n11287), .ZN(n11290) );
  OAI21_X1 U14753 ( .B1(n11143), .B2(n17338), .A(n15890), .ZN(n11288) );
  OAI21_X1 U14754 ( .B1(n15890), .B2(n17338), .A(n11288), .ZN(n11289) );
  MUX2_X1 U14755 ( .A(n11291), .B(n12637), .S(n13038), .Z(n11292) );
  MUX2_X1 U14756 ( .A(n11292), .B(P2_EBX_REG_0__SCAN_IN), .S(n12689), .Z(
        n15957) );
  NAND2_X1 U14757 ( .A1(n15957), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13358) );
  NAND3_X1 U14758 ( .A1(n12689), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U14759 ( .A1(n11296), .A2(n11293), .ZN(n15940) );
  NOR2_X1 U14760 ( .A1(n13358), .A2(n15940), .ZN(n11294) );
  NAND2_X1 U14761 ( .A1(n13358), .A2(n15940), .ZN(n13357) );
  OAI21_X1 U14762 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11294), .A(
        n13357), .ZN(n13767) );
  INV_X1 U14763 ( .A(n11295), .ZN(n11309) );
  NAND2_X1 U14764 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  NAND2_X1 U14765 ( .A1(n11309), .A2(n11298), .ZN(n15929) );
  XNOR2_X1 U14766 ( .A(n15929), .B(n13237), .ZN(n13766) );
  OR2_X1 U14767 ( .A1(n13767), .A2(n13766), .ZN(n13245) );
  INV_X1 U14768 ( .A(n15929), .ZN(n11299) );
  NAND2_X1 U14769 ( .A1(n11299), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11300) );
  NAND2_X1 U14770 ( .A1(n13245), .A2(n11300), .ZN(n16710) );
  INV_X1 U14771 ( .A(n11302), .ZN(n11303) );
  NAND2_X1 U14772 ( .A1(n10340), .A2(n11303), .ZN(n11304) );
  NAND2_X1 U14773 ( .A1(n11282), .A2(n11304), .ZN(n16693) );
  NAND2_X1 U14774 ( .A1(n16693), .A2(n16703), .ZN(n11311) );
  OAI21_X1 U14775 ( .B1(n16710), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11311), .ZN(n11306) );
  NOR2_X1 U14776 ( .A1(n11306), .A2(n16690), .ZN(n11305) );
  NAND2_X1 U14777 ( .A1(n16709), .A2(n11305), .ZN(n11316) );
  INV_X1 U14778 ( .A(n11306), .ZN(n11314) );
  INV_X1 U14779 ( .A(n11307), .ZN(n11308) );
  NAND2_X1 U14780 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  AND2_X1 U14781 ( .A1(n11310), .A2(n10340), .ZN(n16688) );
  NAND3_X1 U14782 ( .A1(n16710), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11311), .ZN(n11312) );
  OAI21_X1 U14783 ( .B1(n16703), .B2(n16693), .A(n11312), .ZN(n11313) );
  AOI21_X1 U14784 ( .B1(n11314), .B2(n16688), .A(n11313), .ZN(n11315) );
  NAND2_X1 U14785 ( .A1(n11316), .A2(n11315), .ZN(n16679) );
  NAND2_X1 U14786 ( .A1(n16680), .A2(n16679), .ZN(n11321) );
  NAND2_X1 U14787 ( .A1(n11317), .A2(n15890), .ZN(n11319) );
  AOI21_X1 U14788 ( .B1(n15890), .B2(n16690), .A(n17338), .ZN(n11318) );
  NAND2_X1 U14789 ( .A1(n11319), .A2(n11318), .ZN(n11320) );
  NAND2_X1 U14790 ( .A1(n11321), .A2(n11320), .ZN(n16670) );
  INV_X1 U14791 ( .A(n11323), .ZN(n11325) );
  NAND2_X1 U14792 ( .A1(n9628), .A2(n10341), .ZN(n11328) );
  AND2_X1 U14793 ( .A1(n10339), .A2(n11328), .ZN(n19751) );
  INV_X1 U14794 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16973) );
  NAND2_X1 U14795 ( .A1(n12689), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11330) );
  MUX2_X1 U14796 ( .A(n12689), .B(n11330), .S(n11329), .Z(n11332) );
  INV_X1 U14797 ( .A(n11331), .ZN(n11337) );
  NAND2_X1 U14798 ( .A1(n11332), .A2(n11337), .ZN(n15847) );
  INV_X1 U14799 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16930) );
  OAI21_X1 U14800 ( .B1(n15847), .B2(n11143), .A(n16930), .ZN(n16628) );
  NAND2_X1 U14801 ( .A1(n11257), .A2(n11333), .ZN(n11334) );
  AND2_X1 U14802 ( .A1(n11329), .A2(n11334), .ZN(n15863) );
  NAND2_X1 U14803 ( .A1(n15863), .A2(n16690), .ZN(n11341) );
  NAND2_X1 U14804 ( .A1(n11341), .A2(n21729), .ZN(n16640) );
  INV_X1 U14805 ( .A(n11335), .ZN(n11336) );
  XNOR2_X1 U14806 ( .A(n10339), .B(n11336), .ZN(n11343) );
  NAND2_X1 U14807 ( .A1(n11343), .A2(n11142), .ZN(n16657) );
  AND2_X1 U14808 ( .A1(n16640), .A2(n16657), .ZN(n16631) );
  AND2_X1 U14809 ( .A1(n16628), .A2(n16631), .ZN(n16612) );
  NAND2_X1 U14810 ( .A1(n12689), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11338) );
  MUX2_X1 U14811 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11338), .S(n11337), .Z(
        n11339) );
  NAND2_X1 U14812 ( .A1(n11339), .A2(n11419), .ZN(n15837) );
  OR2_X1 U14813 ( .A1(n15837), .A2(n11143), .ZN(n11340) );
  INV_X1 U14814 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16919) );
  NAND2_X1 U14815 ( .A1(n11340), .A2(n16919), .ZN(n16616) );
  INV_X1 U14816 ( .A(n11341), .ZN(n11342) );
  NAND2_X1 U14817 ( .A1(n11342), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16641) );
  INV_X1 U14818 ( .A(n11343), .ZN(n15879) );
  NAND2_X1 U14819 ( .A1(n15879), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16656) );
  AND2_X1 U14820 ( .A1(n16641), .A2(n16656), .ZN(n16630) );
  NAND2_X1 U14821 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11344) );
  OR2_X1 U14822 ( .A1(n15837), .A2(n11344), .ZN(n16615) );
  INV_X1 U14823 ( .A(n15847), .ZN(n11346) );
  AND2_X1 U14824 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U14825 ( .A1(n11346), .A2(n11345), .ZN(n16627) );
  NAND2_X1 U14826 ( .A1(n12689), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U14827 ( .A(n12689), .B(n11349), .S(n11348), .Z(n11350) );
  NAND2_X1 U14828 ( .A1(n19742), .A2(n16690), .ZN(n11403) );
  INV_X1 U14829 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U14830 ( .A1(n11403), .A2(n12883), .ZN(n12913) );
  INV_X1 U14831 ( .A(n11351), .ZN(n11352) );
  XNOR2_X1 U14832 ( .A(n11353), .B(n11352), .ZN(n15735) );
  NAND2_X1 U14833 ( .A1(n15735), .A2(n16690), .ZN(n11392) );
  NAND2_X1 U14834 ( .A1(n11392), .A2(n16825), .ZN(n16515) );
  XNOR2_X1 U14835 ( .A(n11354), .B(n10563), .ZN(n11393) );
  NAND2_X1 U14836 ( .A1(n11393), .A2(n16690), .ZN(n11355) );
  INV_X1 U14837 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16526) );
  NAND2_X1 U14838 ( .A1(n11355), .A2(n16526), .ZN(n16530) );
  AND2_X1 U14839 ( .A1(n16515), .A2(n16530), .ZN(n12912) );
  AND2_X1 U14840 ( .A1(n12913), .A2(n12912), .ZN(n16504) );
  AND3_X1 U14841 ( .A1(n9669), .A2(n12689), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n11357) );
  OR2_X1 U14842 ( .A1(n11357), .A2(n11356), .ZN(n15716) );
  INV_X1 U14843 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16809) );
  OAI21_X1 U14844 ( .B1(n15716), .B2(n11143), .A(n16809), .ZN(n16507) );
  OR2_X1 U14845 ( .A1(n11359), .A2(n11358), .ZN(n11360) );
  NAND2_X1 U14846 ( .A1(n11354), .A2(n11360), .ZN(n15767) );
  NAND2_X1 U14847 ( .A1(n11401), .A2(n16861), .ZN(n12908) );
  NOR2_X1 U14848 ( .A1(n19868), .A2(n16288), .ZN(n11362) );
  AOI21_X1 U14849 ( .B1(n9626), .B2(n11362), .A(n11361), .ZN(n11363) );
  NAND2_X1 U14850 ( .A1(n11364), .A2(n11363), .ZN(n15778) );
  XNOR2_X1 U14851 ( .A(n11394), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16548) );
  NAND2_X1 U14852 ( .A1(n12689), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11365) );
  MUX2_X1 U14853 ( .A(n12689), .B(n11365), .S(n11383), .Z(n11366) );
  OR2_X1 U14854 ( .A1(n11383), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11379) );
  AND2_X1 U14855 ( .A1(n11366), .A2(n11379), .ZN(n15792) );
  NAND2_X1 U14856 ( .A1(n15792), .A2(n16690), .ZN(n11398) );
  INV_X1 U14857 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U14858 ( .A1(n11398), .A2(n11367), .ZN(n16569) );
  NAND2_X1 U14859 ( .A1(n11370), .A2(n10496), .ZN(n11371) );
  NAND2_X1 U14860 ( .A1(n11368), .A2(n11371), .ZN(n15823) );
  NAND2_X1 U14861 ( .A1(n12901), .A2(n16901), .ZN(n13052) );
  INV_X1 U14862 ( .A(n11372), .ZN(n11376) );
  INV_X1 U14863 ( .A(n11373), .ZN(n11374) );
  NAND3_X1 U14864 ( .A1(n11374), .A2(n12689), .A3(P2_EBX_REG_11__SCAN_IN), 
        .ZN(n11375) );
  NAND2_X1 U14865 ( .A1(n13276), .A2(n16690), .ZN(n11388) );
  NAND2_X1 U14866 ( .A1(n11388), .A2(n16914), .ZN(n16597) );
  AND2_X1 U14867 ( .A1(n13052), .A2(n16597), .ZN(n12903) );
  NOR2_X1 U14868 ( .A1(n19868), .A2(n11377), .ZN(n11378) );
  NAND2_X1 U14869 ( .A1(n11379), .A2(n11378), .ZN(n11380) );
  NAND2_X1 U14870 ( .A1(n11380), .A2(n9626), .ZN(n15784) );
  OAI21_X1 U14871 ( .B1(n15784), .B2(n11143), .A(n16875), .ZN(n16559) );
  NAND2_X1 U14872 ( .A1(n11368), .A2(n11381), .ZN(n11382) );
  NAND2_X1 U14873 ( .A1(n11383), .A2(n11382), .ZN(n15811) );
  OR2_X1 U14874 ( .A1(n15811), .A2(n11143), .ZN(n11384) );
  INV_X1 U14875 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13050) );
  NAND2_X1 U14876 ( .A1(n11384), .A2(n13050), .ZN(n13054) );
  AND4_X1 U14877 ( .A1(n16569), .A2(n12903), .A3(n16559), .A4(n13054), .ZN(
        n11385) );
  AND3_X1 U14878 ( .A1(n12908), .A2(n16548), .A3(n11385), .ZN(n11386) );
  AND3_X1 U14879 ( .A1(n16504), .A2(n16507), .A3(n11386), .ZN(n11387) );
  INV_X1 U14880 ( .A(n11387), .ZN(n11408) );
  XNOR2_X1 U14881 ( .A(n12901), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16590) );
  INV_X1 U14882 ( .A(n11388), .ZN(n11389) );
  NAND2_X1 U14883 ( .A1(n11389), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16598) );
  AND2_X1 U14884 ( .A1(n16590), .A2(n16598), .ZN(n11407) );
  INV_X1 U14885 ( .A(n15716), .ZN(n11391) );
  AND2_X1 U14886 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U14887 ( .A1(n11391), .A2(n11390), .ZN(n16506) );
  OR2_X1 U14888 ( .A1(n11392), .A2(n16825), .ZN(n16516) );
  INV_X1 U14889 ( .A(n11393), .ZN(n15751) );
  AND2_X1 U14890 ( .A1(n16516), .A2(n16529), .ZN(n12910) );
  INV_X1 U14891 ( .A(n11394), .ZN(n11395) );
  NAND2_X1 U14892 ( .A1(n11395), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12906) );
  INV_X1 U14893 ( .A(n15784), .ZN(n11397) );
  AND2_X1 U14894 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11396) );
  NAND2_X1 U14895 ( .A1(n11397), .A2(n11396), .ZN(n16558) );
  INV_X1 U14896 ( .A(n11398), .ZN(n11399) );
  NAND2_X1 U14897 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16570) );
  NAND2_X1 U14898 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11400) );
  OR2_X1 U14899 ( .A1(n15811), .A2(n11400), .ZN(n13053) );
  AND4_X1 U14900 ( .A1(n12906), .A2(n16558), .A3(n16570), .A4(n13053), .ZN(
        n11402) );
  AND2_X1 U14901 ( .A1(n11402), .A2(n12909), .ZN(n11405) );
  INV_X1 U14902 ( .A(n11403), .ZN(n11404) );
  NAND2_X1 U14903 ( .A1(n11404), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16502) );
  AND4_X1 U14904 ( .A1(n16506), .A2(n12910), .A3(n11405), .A4(n16502), .ZN(
        n11406) );
  NAND2_X1 U14905 ( .A1(n11411), .A2(n16798), .ZN(n16492) );
  NAND2_X1 U14906 ( .A1(n12689), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11415) );
  INV_X1 U14907 ( .A(n11415), .ZN(n11416) );
  NAND2_X1 U14908 ( .A1(n11417), .A2(n11416), .ZN(n11418) );
  NAND2_X1 U14909 ( .A1(n11424), .A2(n11418), .ZN(n15627) );
  NAND2_X1 U14910 ( .A1(n11419), .A2(n16690), .ZN(n11421) );
  AOI21_X1 U14911 ( .B1(n16440), .B2(n16745), .A(n16460), .ZN(n11420) );
  OR2_X1 U14912 ( .A1(n11421), .A2(n13147), .ZN(n16459) );
  NOR2_X1 U14913 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11426) );
  INV_X1 U14914 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15605) );
  NOR2_X1 U14915 ( .A1(n19868), .A2(n15605), .ZN(n11423) );
  INV_X1 U14916 ( .A(n11431), .ZN(n11427) );
  NAND2_X1 U14917 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  NAND2_X1 U14918 ( .A1(n11427), .A2(n11425), .ZN(n15608) );
  OR2_X1 U14919 ( .A1(n15608), .A2(n11143), .ZN(n16442) );
  NAND2_X1 U14920 ( .A1(n12689), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U14921 ( .A1(n15594), .A2(n16690), .ZN(n11428) );
  INV_X1 U14922 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16727) );
  NAND2_X1 U14923 ( .A1(n11428), .A2(n16727), .ZN(n16431) );
  NAND2_X1 U14924 ( .A1(n12689), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11432) );
  INV_X1 U14925 ( .A(n13078), .ZN(n13080) );
  AND2_X1 U14926 ( .A1(n16690), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11433) );
  NAND2_X1 U14927 ( .A1(n13109), .A2(n11433), .ZN(n13079) );
  NAND2_X1 U14928 ( .A1(n13080), .A2(n13079), .ZN(n11434) );
  OAI211_X1 U14929 ( .C1(n16722), .C2(n13130), .A(n11436), .B(n11435), .ZN(
        P2_U2984) );
  NOR2_X1 U14930 ( .A1(n10301), .A2(n19566), .ZN(n17788) );
  INV_X1 U14931 ( .A(n17788), .ZN(n17802) );
  NOR3_X1 U14932 ( .A1(n17071), .A2(n11437), .A3(n17802), .ZN(n11446) );
  INV_X1 U14933 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19646) );
  INV_X1 U14934 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19649) );
  AOI221_X1 U14935 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n19646), .C2(n19649), .A(n11438), .ZN(n11445) );
  INV_X1 U14936 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17814) );
  NAND2_X1 U14937 ( .A1(n11439), .A2(n17814), .ZN(n11443) );
  AOI22_X1 U14938 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n17467), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17800), .ZN(n11441) );
  INV_X1 U14939 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14481) );
  OR3_X1 U14940 ( .A1(n11446), .A2(n11445), .A3(n11444), .ZN(P3_U2640) );
  AND2_X2 U14941 ( .A1(n11451), .A2(n13590), .ZN(n11628) );
  AND2_X4 U14942 ( .A1(n13590), .A2(n15563), .ZN(n12538) );
  AOI22_X1 U14943 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14944 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11610), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14945 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11448) );
  AND2_X2 U14946 ( .A1(n13590), .A2(n14060), .ZN(n11719) );
  AND2_X2 U14947 ( .A1(n11452), .A2(n15563), .ZN(n11634) );
  AOI22_X1 U14948 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11457) );
  AND2_X4 U14949 ( .A1(n11451), .A2(n13594), .ZN(n12605) );
  AND2_X2 U14950 ( .A1(n11451), .A2(n11453), .ZN(n11613) );
  AOI22_X1 U14951 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11613), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14952 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11455) );
  AND2_X4 U14953 ( .A1(n14060), .A2(n11453), .ZN(n12409) );
  AND2_X2 U14954 ( .A1(n11453), .A2(n15563), .ZN(n11725) );
  AOI22_X1 U14955 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11454) );
  AND4_X2 U14956 ( .A1(n11457), .A2(n11456), .A3(n11455), .A4(n11454), .ZN(
        n11458) );
  INV_X1 U14957 ( .A(n11554), .ZN(n11478) );
  AOI22_X1 U14958 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14959 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14960 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11613), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14961 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14962 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14963 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11467), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14964 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11468) );
  NAND4_X1 U14965 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11477) );
  AOI22_X1 U14966 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14967 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14968 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14969 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14970 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11476) );
  AOI21_X2 U14971 ( .B1(n11478), .B2(n12068), .A(n14545), .ZN(n11932) );
  AOI22_X1 U14972 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14973 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14974 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14975 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14976 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14977 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U14978 ( .A1(n11932), .A2(n11940), .ZN(n11587) );
  INV_X1 U14979 ( .A(n11587), .ZN(n11489) );
  INV_X1 U14980 ( .A(n13187), .ZN(n11488) );
  NAND2_X1 U14981 ( .A1(n11489), .A2(n11488), .ZN(n11589) );
  NAND2_X1 U14982 ( .A1(n11589), .A2(n11588), .ZN(n11548) );
  AOI22_X1 U14983 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14984 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14985 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14986 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14987 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14988 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14989 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14990 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9600), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14991 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14992 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14993 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11611), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14994 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14995 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11634), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14996 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11725), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14997 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11511) );
  NAND2_X1 U14998 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11510) );
  NAND2_X1 U14999 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U15000 ( .A1(n11634), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U15001 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U15002 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U15003 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U15004 ( .A1(n9600), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11512) );
  NAND2_X1 U15005 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11519) );
  NAND2_X1 U15006 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U15007 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U15008 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11516) );
  NAND2_X1 U15009 ( .A1(n11467), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U15010 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U15011 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11521) );
  NAND2_X1 U15012 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11520) );
  NAND4_X4 U15013 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n21581) );
  NAND2_X1 U15014 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U15015 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U15016 ( .A1(n11611), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U15017 ( .A1(n11634), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U15018 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U15019 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U15020 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11533) );
  NAND2_X1 U15021 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U15022 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U15023 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U15024 ( .A1(n9600), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U15025 ( .A1(n9606), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U15026 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11543) );
  NAND2_X1 U15027 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11542) );
  NAND2_X1 U15028 ( .A1(n11725), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11541) );
  NAND2_X1 U15029 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11540) );
  NAND4_X4 U15030 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11562) );
  INV_X2 U15031 ( .A(n11562), .ZN(n11573) );
  NAND2_X1 U15032 ( .A1(n11573), .A2(n21581), .ZN(n14243) );
  INV_X1 U15033 ( .A(n20824), .ZN(n11581) );
  NAND2_X1 U15034 ( .A1(n11995), .A2(n11930), .ZN(n12067) );
  NAND4_X1 U15035 ( .A1(n11548), .A2(n13176), .A3(n14243), .A4(n12067), .ZN(
        n11553) );
  NAND2_X1 U15036 ( .A1(n11550), .A2(n11549), .ZN(n13313) );
  INV_X1 U15037 ( .A(n13313), .ZN(n11552) );
  XNOR2_X1 U15038 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11872) );
  NOR2_X2 U15039 ( .A1(n12061), .A2(n11872), .ZN(n11572) );
  NOR2_X1 U15040 ( .A1(n11553), .A2(n11572), .ZN(n11567) );
  NAND2_X1 U15041 ( .A1(n12069), .A2(n11554), .ZN(n11625) );
  NAND2_X1 U15042 ( .A1(n11625), .A2(n12107), .ZN(n11557) );
  INV_X1 U15043 ( .A(n12065), .ZN(n11561) );
  OAI21_X1 U15044 ( .B1(n13187), .B2(n11573), .A(n13772), .ZN(n11563) );
  NAND2_X1 U15045 ( .A1(n11589), .A2(n11563), .ZN(n11933) );
  NAND2_X1 U15046 ( .A1(n20819), .A2(n11562), .ZN(n11585) );
  OAI21_X1 U15047 ( .B1(n12065), .B2(n11950), .A(n11585), .ZN(n11564) );
  INV_X1 U15048 ( .A(n11564), .ZN(n11565) );
  OAI21_X1 U15049 ( .B1(n11580), .B2(n13684), .A(n11573), .ZN(n11566) );
  NAND4_X1 U15050 ( .A1(n11567), .A2(n11929), .A3(n13582), .A4(n11566), .ZN(
        n11568) );
  NAND2_X1 U15051 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11677) );
  OAI21_X1 U15052 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11677), .ZN(n21198) );
  NAND2_X1 U15053 ( .A1(n17301), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11668) );
  OAI21_X1 U15054 ( .B1(n12622), .B2(n21198), .A(n11668), .ZN(n11570) );
  INV_X1 U15055 ( .A(n11570), .ZN(n11571) );
  INV_X1 U15056 ( .A(n11572), .ZN(n11574) );
  NOR2_X1 U15057 ( .A1(n12065), .A2(n13182), .ZN(n11575) );
  AND2_X2 U15058 ( .A1(n13581), .A2(n13176), .ZN(n11942) );
  INV_X1 U15059 ( .A(n17301), .ZN(n11579) );
  MUX2_X1 U15060 ( .A(n11579), .B(n12622), .S(n21327), .Z(n11642) );
  OAI21_X2 U15061 ( .B1(n11711), .B2(n11578), .A(n11642), .ZN(n12120) );
  NAND2_X1 U15062 ( .A1(n11580), .A2(n9837), .ZN(n12075) );
  OR2_X1 U15063 ( .A1(n13187), .A2(n11581), .ZN(n11584) );
  NAND2_X1 U15064 ( .A1(n15570), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20571) );
  INV_X1 U15065 ( .A(n20571), .ZN(n11582) );
  NAND2_X1 U15066 ( .A1(n14243), .A2(n11582), .ZN(n11583) );
  AOI21_X1 U15067 ( .B1(n14554), .B2(n11584), .A(n11583), .ZN(n11592) );
  NAND2_X1 U15068 ( .A1(n13684), .A2(n12127), .ZN(n11586) );
  NAND2_X1 U15069 ( .A1(n11586), .A2(n11585), .ZN(n12064) );
  AOI21_X1 U15070 ( .B1(n21584), .B2(n11587), .A(n12064), .ZN(n11591) );
  NAND3_X1 U15071 ( .A1(n11589), .A2(n15567), .A3(n21581), .ZN(n11590) );
  NAND4_X1 U15072 ( .A1(n12075), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n12121) );
  INV_X1 U15073 ( .A(n11717), .ZN(n11608) );
  AOI22_X1 U15074 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U15075 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U15076 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U15077 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U15078 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11607) );
  AOI22_X1 U15079 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U15080 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U15081 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11603) );
  INV_X2 U15082 ( .A(n11633), .ZN(n12512) );
  AOI22_X1 U15083 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U15084 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  NAND2_X1 U15085 ( .A1(n11608), .A2(n11657), .ZN(n11609) );
  INV_X1 U15086 ( .A(n11610), .ZN(n11633) );
  CLKBUF_X3 U15087 ( .A(n11611), .Z(n12511) );
  AOI22_X1 U15088 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U15089 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n12595), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U15090 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12395), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U15091 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U15092 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11623) );
  AOI22_X1 U15093 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12602), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U15094 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12496), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U15095 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U15096 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12449), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U15097 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n11622) );
  NAND2_X1 U15098 ( .A1(n11648), .A2(n11657), .ZN(n11737) );
  OAI21_X1 U15099 ( .B1(n11648), .B2(n11657), .A(n11737), .ZN(n11624) );
  INV_X1 U15100 ( .A(n11624), .ZN(n11626) );
  AOI21_X1 U15101 ( .B1(n11626), .B2(n21584), .A(n11625), .ZN(n11627) );
  AOI22_X1 U15102 ( .A1(n11724), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U15103 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U15104 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U15105 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U15106 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11640) );
  AOI22_X1 U15107 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U15108 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U15109 ( .A1(n11719), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U15110 ( .A1(n11610), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U15111 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  OR2_X2 U15112 ( .A1(n11640), .A2(n11639), .ZN(n11818) );
  MUX2_X1 U15113 ( .A(n11824), .B(n11656), .S(n11648), .Z(n11641) );
  INV_X1 U15114 ( .A(n11641), .ZN(n11644) );
  NAND2_X1 U15115 ( .A1(n11642), .A2(n21501), .ZN(n11643) );
  INV_X1 U15116 ( .A(n11648), .ZN(n11647) );
  NAND2_X1 U15117 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11646) );
  AOI21_X1 U15118 ( .B1(n11940), .B2(n11818), .A(n21501), .ZN(n11645) );
  OR2_X1 U15119 ( .A1(n13772), .A2(n11648), .ZN(n13723) );
  NAND2_X1 U15120 ( .A1(n11573), .A2(n20824), .ZN(n13722) );
  AND2_X1 U15121 ( .A1(n13723), .A2(n13722), .ZN(n11649) );
  NAND2_X1 U15122 ( .A1(n20894), .A2(n11649), .ZN(n11651) );
  INV_X1 U15123 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13749) );
  AOI21_X1 U15124 ( .B1(n11649), .B2(n13725), .A(n13749), .ZN(n11650) );
  NAND2_X1 U15125 ( .A1(n11651), .A2(n11650), .ZN(n13727) );
  NAND2_X1 U15126 ( .A1(n11652), .A2(n10170), .ZN(n11653) );
  INV_X1 U15127 ( .A(n11656), .ZN(n11660) );
  NAND2_X1 U15128 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11659) );
  INV_X1 U15129 ( .A(n11716), .ZN(n11697) );
  NAND2_X1 U15130 ( .A1(n11697), .A2(n11657), .ZN(n11658) );
  NAND2_X1 U15131 ( .A1(n11661), .A2(n11662), .ZN(n11666) );
  INV_X1 U15132 ( .A(n11661), .ZN(n11664) );
  INV_X1 U15133 ( .A(n11662), .ZN(n11663) );
  NAND2_X1 U15134 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  INV_X1 U15135 ( .A(n11667), .ZN(n11670) );
  AND2_X1 U15136 ( .A1(n11668), .A2(n11569), .ZN(n11669) );
  INV_X1 U15137 ( .A(n13680), .ZN(n11681) );
  NAND2_X1 U15138 ( .A1(n17301), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11674) );
  INV_X1 U15139 ( .A(n12622), .ZN(n11713) );
  INV_X1 U15140 ( .A(n11677), .ZN(n11676) );
  NAND2_X1 U15141 ( .A1(n11676), .A2(n21276), .ZN(n20928) );
  NAND2_X1 U15142 ( .A1(n11677), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11678) );
  NAND2_X1 U15143 ( .A1(n20928), .A2(n11678), .ZN(n20809) );
  AOI21_X1 U15144 ( .B1(n11682), .B2(n21501), .A(n11683), .ZN(n11679) );
  INV_X1 U15145 ( .A(n11679), .ZN(n11680) );
  INV_X1 U15146 ( .A(n11682), .ZN(n11685) );
  NAND3_X1 U15147 ( .A1(n10061), .A2(n13680), .A3(n21501), .ZN(n11704) );
  NAND2_X1 U15148 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11699) );
  AOI22_X1 U15149 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U15150 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U15151 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U15152 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U15153 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11696) );
  AOI22_X1 U15154 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U15155 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U15156 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U15157 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U15158 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11695) );
  NAND2_X1 U15159 ( .A1(n11697), .A2(n11700), .ZN(n11698) );
  NAND2_X1 U15160 ( .A1(n11699), .A2(n11698), .ZN(n11702) );
  NOR2_X1 U15161 ( .A1(n11736), .A2(n11717), .ZN(n11701) );
  XNOR2_X1 U15162 ( .A(n11702), .B(n11701), .ZN(n11703) );
  XNOR2_X1 U15163 ( .A(n11737), .B(n11736), .ZN(n11706) );
  INV_X1 U15164 ( .A(n13722), .ZN(n11705) );
  AOI21_X1 U15165 ( .B1(n11706), .B2(n21584), .A(n11705), .ZN(n11707) );
  NAND2_X1 U15166 ( .A1(n11708), .A2(n11707), .ZN(n15291) );
  NAND2_X1 U15167 ( .A1(n11709), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11710) );
  INV_X1 U15168 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20764) );
  NAND2_X1 U15169 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10565), .ZN(
        n21110) );
  NAND2_X1 U15170 ( .A1(n21275), .A2(n21110), .ZN(n11712) );
  NOR3_X1 U15171 ( .A1(n21275), .A2(n21276), .A3(n21195), .ZN(n21441) );
  NAND2_X1 U15172 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21441), .ZN(
        n21489) );
  AOI22_X1 U15173 ( .A1(n11713), .A2(n21120), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17301), .ZN(n11714) );
  AOI22_X1 U15174 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U15175 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U15176 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U15177 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11720) );
  NAND4_X1 U15178 ( .A1(n11723), .A2(n11722), .A3(n11721), .A4(n11720), .ZN(
        n11731) );
  AOI22_X1 U15179 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U15180 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U15181 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U15182 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11726) );
  NAND4_X1 U15183 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11730) );
  AOI22_X1 U15184 ( .A1(n11921), .A2(n11772), .B1(n11891), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11732) );
  INV_X1 U15185 ( .A(n11734), .ZN(n11735) );
  NAND2_X1 U15186 ( .A1(n11737), .A2(n11736), .ZN(n11773) );
  INV_X1 U15187 ( .A(n11772), .ZN(n11738) );
  XNOR2_X1 U15188 ( .A(n11773), .B(n11738), .ZN(n11739) );
  NAND2_X1 U15189 ( .A1(n11739), .A2(n21584), .ZN(n11740) );
  NAND2_X1 U15190 ( .A1(n11741), .A2(n11740), .ZN(n15282) );
  AOI22_X1 U15191 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U15192 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U15193 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U15194 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11744) );
  NAND4_X1 U15195 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11753) );
  AOI22_X1 U15196 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U15197 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U15198 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U15199 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11748) );
  NAND4_X1 U15200 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  NAND2_X1 U15201 ( .A1(n11921), .A2(n11774), .ZN(n11755) );
  NAND2_X1 U15202 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U15203 ( .A1(n11755), .A2(n11754), .ZN(n11770) );
  AOI22_X1 U15204 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U15205 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U15206 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U15207 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U15208 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11765) );
  AOI22_X1 U15209 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11763) );
  INV_X1 U15210 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21701) );
  AOI22_X1 U15211 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U15212 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U15213 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11760) );
  NAND4_X1 U15214 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11764) );
  NAND2_X1 U15215 ( .A1(n11921), .A2(n11802), .ZN(n11767) );
  NAND2_X1 U15216 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U15217 ( .A1(n11767), .A2(n11766), .ZN(n11786) );
  AND2_X1 U15218 ( .A1(n11772), .A2(n11774), .ZN(n11768) );
  NAND2_X1 U15219 ( .A1(n11773), .A2(n11768), .ZN(n11804) );
  XNOR2_X1 U15220 ( .A(n11804), .B(n11802), .ZN(n11769) );
  INV_X1 U15221 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15273) );
  NAND2_X1 U15222 ( .A1(n12149), .A2(n11928), .ZN(n11778) );
  NAND2_X1 U15223 ( .A1(n11773), .A2(n11772), .ZN(n11775) );
  XNOR2_X1 U15224 ( .A(n11775), .B(n11774), .ZN(n11776) );
  NAND2_X1 U15225 ( .A1(n11776), .A2(n21584), .ZN(n11777) );
  NOR2_X1 U15226 ( .A1(n15272), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U15227 ( .A1(n15272), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15228 ( .A1(n11781), .A2(n15273), .ZN(n11783) );
  AND2_X1 U15229 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U15230 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U15231 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U15232 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15233 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11787) );
  NAND4_X1 U15234 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11796) );
  AOI22_X1 U15235 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U15236 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U15237 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U15238 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U15239 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11795) );
  NAND2_X1 U15240 ( .A1(n11921), .A2(n11816), .ZN(n11798) );
  NAND2_X1 U15241 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U15242 ( .A1(n11801), .A2(n11800), .ZN(n12152) );
  INV_X1 U15243 ( .A(n11802), .ZN(n11803) );
  XNOR2_X1 U15244 ( .A(n11815), .B(n11816), .ZN(n11805) );
  NAND2_X1 U15245 ( .A1(n11805), .A2(n21584), .ZN(n11806) );
  INV_X1 U15246 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15534) );
  NAND2_X1 U15247 ( .A1(n15264), .A2(n15534), .ZN(n11808) );
  INV_X1 U15248 ( .A(n15264), .ZN(n11809) );
  NAND2_X1 U15249 ( .A1(n11809), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U15250 ( .A1(n11921), .A2(n11818), .ZN(n11812) );
  NAND2_X1 U15251 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U15252 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  INV_X1 U15253 ( .A(n11815), .ZN(n11817) );
  NAND2_X1 U15254 ( .A1(n11817), .A2(n11816), .ZN(n11828) );
  XNOR2_X1 U15255 ( .A(n11828), .B(n11818), .ZN(n11819) );
  AND2_X1 U15256 ( .A1(n11819), .A2(n21584), .ZN(n11820) );
  AOI21_X1 U15257 ( .B1(n12188), .B2(n11928), .A(n11820), .ZN(n11821) );
  INV_X1 U15258 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U15259 ( .A1(n11821), .A2(n15519), .ZN(n15257) );
  INV_X1 U15260 ( .A(n11821), .ZN(n11822) );
  NAND2_X1 U15261 ( .A1(n11822), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15256) );
  INV_X1 U15262 ( .A(n11824), .ZN(n11825) );
  OR3_X1 U15263 ( .A1(n11828), .A2(n11827), .A3(n13772), .ZN(n11829) );
  INV_X1 U15264 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11830) );
  NAND2_X1 U15265 ( .A1(n15247), .A2(n11830), .ZN(n11831) );
  INV_X1 U15266 ( .A(n15247), .ZN(n11832) );
  NAND2_X1 U15267 ( .A1(n11832), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11833) );
  INV_X1 U15268 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U15269 ( .A1(n15239), .A2(n15453), .ZN(n11834) );
  INV_X1 U15270 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U15271 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11835) );
  INV_X1 U15272 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U15273 ( .A1(n15239), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11836) );
  INV_X1 U15274 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U15275 ( .A1(n15239), .A2(n15177), .ZN(n11837) );
  NAND3_X1 U15276 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U15277 ( .A1(n15239), .A2(n11838), .ZN(n11839) );
  NAND2_X1 U15278 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15188) );
  NOR2_X1 U15279 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U15280 ( .A1(n15198), .A2(n15469), .ZN(n15152) );
  NOR2_X1 U15281 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15424) );
  INV_X1 U15282 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21716) );
  NAND2_X1 U15283 ( .A1(n15424), .A2(n21716), .ZN(n11840) );
  OAI21_X1 U15284 ( .B1(n15152), .B2(n11840), .A(n15220), .ZN(n11841) );
  NAND2_X1 U15285 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15150) );
  INV_X1 U15286 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11845) );
  INV_X1 U15287 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11844) );
  XNOR2_X1 U15288 ( .A(n15239), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15140) );
  NAND2_X1 U15289 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15105) );
  INV_X1 U15290 ( .A(n15105), .ZN(n11847) );
  INV_X1 U15291 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12031) );
  NAND2_X1 U15292 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11848) );
  NAND3_X1 U15293 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15067) );
  NOR2_X1 U15294 ( .A1(n11849), .A2(n15220), .ZN(n15078) );
  INV_X1 U15295 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U15296 ( .A1(n15320), .A2(n15330), .ZN(n11851) );
  NOR2_X1 U15297 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15299) );
  AND2_X1 U15298 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U15299 ( .A1(n15239), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11853) );
  XNOR2_X1 U15300 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U15301 ( .A1(n21327), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U15302 ( .A1(n11868), .A2(n11867), .ZN(n11855) );
  NAND2_X1 U15303 ( .A1(n21195), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U15304 ( .A1(n11855), .A2(n11854), .ZN(n11870) );
  XNOR2_X1 U15305 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U15306 ( .A1(n11870), .A2(n11869), .ZN(n11857) );
  NAND2_X1 U15307 ( .A1(n21276), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15308 ( .A1(n11857), .A2(n11856), .ZN(n11866) );
  NOR2_X1 U15309 ( .A1(n14056), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11858) );
  INV_X1 U15310 ( .A(n11864), .ZN(n11860) );
  INV_X1 U15311 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14063) );
  NOR2_X1 U15312 ( .A1(n14063), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11859) );
  INV_X1 U15313 ( .A(n11863), .ZN(n11861) );
  AND2_X1 U15314 ( .A1(n11864), .A2(n11863), .ZN(n11909) );
  XNOR2_X1 U15315 ( .A(n11866), .B(n11865), .ZN(n11902) );
  XNOR2_X1 U15316 ( .A(n11868), .B(n11867), .ZN(n11877) );
  XNOR2_X1 U15317 ( .A(n11870), .B(n11869), .ZN(n11890) );
  NAND2_X1 U15318 ( .A1(n11919), .A2(n11871), .ZN(n13179) );
  INV_X1 U15319 ( .A(n13179), .ZN(n13316) );
  INV_X1 U15320 ( .A(n21580), .ZN(n15582) );
  AOI21_X1 U15321 ( .B1(n21581), .B2(n15582), .A(n17309), .ZN(n11873) );
  NAND2_X1 U15322 ( .A1(n13316), .A2(n11873), .ZN(n11927) );
  NAND2_X1 U15323 ( .A1(n11921), .A2(n21581), .ZN(n11875) );
  NAND2_X1 U15324 ( .A1(n11478), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U15325 ( .A1(n11875), .A2(n11874), .ZN(n11886) );
  INV_X1 U15326 ( .A(n11886), .ZN(n11876) );
  NAND2_X1 U15327 ( .A1(n11876), .A2(n21581), .ZN(n11908) );
  INV_X1 U15328 ( .A(n11877), .ZN(n11889) );
  NAND2_X1 U15329 ( .A1(n11478), .A2(n11562), .ZN(n11879) );
  NAND2_X1 U15330 ( .A1(n11879), .A2(n13777), .ZN(n11895) );
  OAI21_X1 U15331 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21327), .A(
        n11880), .ZN(n11881) );
  INV_X1 U15332 ( .A(n11881), .ZN(n11882) );
  OAI211_X1 U15333 ( .C1(n12065), .C2(n11573), .A(n11895), .B(n11882), .ZN(
        n11885) );
  NAND2_X1 U15334 ( .A1(n11921), .A2(n11882), .ZN(n11883) );
  NAND2_X1 U15335 ( .A1(n11916), .A2(n11883), .ZN(n11884) );
  OAI211_X1 U15336 ( .C1(n11886), .C2(n11889), .A(n11885), .B(n11884), .ZN(
        n11888) );
  NAND2_X1 U15337 ( .A1(n11886), .A2(n11889), .ZN(n11887) );
  OAI211_X1 U15338 ( .C1(n11908), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        n11894) );
  INV_X1 U15339 ( .A(n11890), .ZN(n11896) );
  NAND2_X1 U15340 ( .A1(n11921), .A2(n11896), .ZN(n11892) );
  OAI211_X1 U15341 ( .C1(n11896), .C2(n11910), .A(n11895), .B(n11892), .ZN(
        n11893) );
  NAND2_X1 U15342 ( .A1(n11894), .A2(n11893), .ZN(n11899) );
  INV_X1 U15343 ( .A(n11895), .ZN(n11897) );
  NAND3_X1 U15344 ( .A1(n11897), .A2(n11896), .A3(n11921), .ZN(n11898) );
  NAND2_X1 U15345 ( .A1(n11899), .A2(n11898), .ZN(n11901) );
  NAND2_X1 U15346 ( .A1(n11910), .A2(n11902), .ZN(n11900) );
  NAND2_X1 U15347 ( .A1(n11901), .A2(n11900), .ZN(n11905) );
  INV_X1 U15348 ( .A(n11916), .ZN(n11903) );
  NAND2_X1 U15349 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  NAND2_X1 U15350 ( .A1(n11905), .A2(n11904), .ZN(n11907) );
  NAND2_X1 U15351 ( .A1(n11910), .A2(n11909), .ZN(n11906) );
  NAND2_X1 U15352 ( .A1(n11907), .A2(n11906), .ZN(n11915) );
  INV_X1 U15353 ( .A(n11908), .ZN(n11913) );
  INV_X1 U15354 ( .A(n11909), .ZN(n11911) );
  NOR2_X1 U15355 ( .A1(n11911), .A2(n11910), .ZN(n11912) );
  AOI22_X1 U15356 ( .A1(n11913), .A2(n11912), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21501), .ZN(n11914) );
  NAND2_X1 U15357 ( .A1(n11915), .A2(n11914), .ZN(n11918) );
  OAI21_X1 U15358 ( .B1(n21581), .B2(n21580), .A(n21590), .ZN(n14239) );
  OAI211_X1 U15359 ( .C1(n13580), .C2(n14239), .A(n11562), .B(n13189), .ZN(
        n11924) );
  INV_X1 U15360 ( .A(n11924), .ZN(n11925) );
  OR2_X1 U15361 ( .A1(n17305), .A2(n11925), .ZN(n11926) );
  MUX2_X1 U15362 ( .A(n11927), .B(n11926), .S(n12069), .Z(n11936) );
  AOI21_X1 U15363 ( .B1(n15567), .B2(n11573), .A(n11930), .ZN(n11938) );
  NAND2_X1 U15364 ( .A1(n13187), .A2(n11940), .ZN(n11931) );
  NAND2_X1 U15365 ( .A1(n11938), .A2(n12073), .ZN(n11939) );
  NAND2_X1 U15366 ( .A1(n13317), .A2(n11939), .ZN(n11934) );
  NAND2_X1 U15367 ( .A1(n11934), .A2(n11933), .ZN(n13568) );
  AOI21_X1 U15368 ( .B1(n17305), .B2(n12083), .A(n13568), .ZN(n11935) );
  NAND2_X1 U15369 ( .A1(n11936), .A2(n11935), .ZN(n11937) );
  NAND2_X1 U15370 ( .A1(n11938), .A2(n9837), .ZN(n13591) );
  OR2_X1 U15371 ( .A1(n12062), .A2(n11940), .ZN(n11941) );
  NAND4_X1 U15372 ( .A1(n11942), .A2(n13591), .A3(n13314), .A4(n11941), .ZN(
        n11943) );
  NAND2_X1 U15373 ( .A1(n11947), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11945) );
  INV_X1 U15374 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11944) );
  NAND2_X1 U15375 ( .A1(n11945), .A2(n10550), .ZN(n13458) );
  INV_X1 U15376 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11946) );
  NAND2_X1 U15377 ( .A1(n13645), .A2(n11946), .ZN(n11949) );
  INV_X1 U15378 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20793) );
  NAND2_X1 U15379 ( .A1(n11947), .A2(n20793), .ZN(n11948) );
  NAND3_X1 U15380 ( .A1(n11949), .A2(n11948), .A3(n11950), .ZN(n11952) );
  NAND2_X1 U15381 ( .A1(n11947), .A2(n20780), .ZN(n11954) );
  INV_X1 U15382 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U15383 ( .A1(n13645), .A2(n11955), .ZN(n11953) );
  NAND3_X1 U15384 ( .A1(n11954), .A2(n11953), .A3(n12072), .ZN(n11957) );
  NAND2_X1 U15385 ( .A1(n12056), .A2(n11955), .ZN(n11956) );
  AND2_X1 U15386 ( .A1(n11957), .A2(n11956), .ZN(n14001) );
  NAND2_X1 U15387 ( .A1(n11959), .A2(n11958), .ZN(n14000) );
  NAND2_X2 U15388 ( .A1(n13645), .A2(n12072), .ZN(n12047) );
  OR2_X1 U15389 ( .A1(n12047), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U15390 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11960) );
  OAI211_X1 U15391 ( .C1(n12015), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12050), .B(
        n11960), .ZN(n11961) );
  NAND2_X1 U15392 ( .A1(n11962), .A2(n11961), .ZN(n14035) );
  NAND2_X1 U15393 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U15394 ( .A1(n12050), .A2(n11963), .ZN(n11966) );
  OR2_X1 U15395 ( .A1(n14530), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n11965) );
  INV_X1 U15396 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15397 ( .A1(n11966), .A2(n11965), .B1(n12056), .B2(n11964), .ZN(
        n14190) );
  OR2_X1 U15398 ( .A1(n12047), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11969) );
  NAND2_X1 U15399 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11967) );
  OAI211_X1 U15400 ( .C1(n14530), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12050), .B(
        n11967), .ZN(n11968) );
  AND2_X1 U15401 ( .A1(n11969), .A2(n11968), .ZN(n15540) );
  NAND2_X1 U15402 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11970) );
  NAND2_X1 U15403 ( .A1(n12050), .A2(n11970), .ZN(n11972) );
  OR2_X1 U15404 ( .A1(n14530), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n11971) );
  INV_X1 U15405 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U15406 ( .A1(n11972), .A2(n11971), .B1(n12056), .B2(n14934), .ZN(
        n14932) );
  OR2_X1 U15407 ( .A1(n12047), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15408 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11974) );
  OAI211_X1 U15409 ( .C1(n14530), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12050), .B(
        n11974), .ZN(n11975) );
  NAND2_X1 U15410 ( .A1(n11976), .A2(n11975), .ZN(n14925) );
  NAND2_X1 U15411 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11977) );
  NAND2_X1 U15412 ( .A1(n12050), .A2(n11977), .ZN(n11979) );
  OR2_X1 U15413 ( .A1(n14530), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U15414 ( .A1(n11979), .A2(n11978), .ZN(n11982) );
  INV_X1 U15415 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U15416 ( .A1(n12056), .A2(n11980), .ZN(n11981) );
  NAND2_X1 U15417 ( .A1(n11982), .A2(n11981), .ZN(n14880) );
  OR2_X1 U15418 ( .A1(n12047), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U15419 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11983) );
  OAI211_X1 U15420 ( .C1(P1_EBX_REG_9__SCAN_IN), .C2(n12015), .A(n11947), .B(
        n11983), .ZN(n11984) );
  AND2_X1 U15421 ( .A1(n11985), .A2(n11984), .ZN(n14865) );
  NAND2_X1 U15422 ( .A1(n14864), .A2(n14865), .ZN(n14843) );
  INV_X1 U15423 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U15424 ( .A1(n11947), .A2(n15493), .ZN(n11986) );
  INV_X1 U15425 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U15426 ( .A1(n12056), .A2(n11987), .ZN(n11988) );
  OR2_X1 U15427 ( .A1(n12047), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U15428 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11992) );
  OAI211_X1 U15429 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n14530), .A(n12050), .B(
        n11992), .ZN(n11993) );
  NAND2_X1 U15430 ( .A1(n11994), .A2(n11993), .ZN(n14830) );
  MUX2_X1 U15431 ( .A(n12047), .B(n12072), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11997) );
  OR2_X1 U15432 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U15433 ( .A1(n11997), .A2(n11996), .ZN(n14805) );
  NAND2_X1 U15434 ( .A1(n12050), .A2(n11998), .ZN(n11999) );
  OAI21_X1 U15435 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n14530), .A(n11999), .ZN(
        n12001) );
  INV_X1 U15436 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U15437 ( .A1(n12056), .A2(n14917), .ZN(n12000) );
  NOR2_X1 U15438 ( .A1(n14805), .A2(n14804), .ZN(n12002) );
  INV_X1 U15439 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U15440 ( .A1(n11947), .A2(n15444), .ZN(n12003) );
  OAI211_X1 U15441 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n14530), .A(n12003), .B(
        n12072), .ZN(n12005) );
  INV_X1 U15442 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U15443 ( .A1(n12056), .A2(n14915), .ZN(n12004) );
  NAND2_X1 U15444 ( .A1(n12005), .A2(n12004), .ZN(n14783) );
  MUX2_X1 U15445 ( .A(n12047), .B(n12072), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12007) );
  OR2_X1 U15446 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U15447 ( .A1(n12007), .A2(n12006), .ZN(n14763) );
  NAND2_X1 U15448 ( .A1(n12050), .A2(n12088), .ZN(n12010) );
  INV_X1 U15449 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U15450 ( .A1(n12056), .A2(n12011), .ZN(n12012) );
  OR2_X1 U15451 ( .A1(n12047), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U15452 ( .A1(n12072), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12014) );
  OAI211_X1 U15453 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n12015), .A(n11947), .B(
        n12014), .ZN(n12016) );
  NAND2_X1 U15454 ( .A1(n12017), .A2(n12016), .ZN(n14733) );
  NAND2_X1 U15455 ( .A1(n12050), .A2(n11843), .ZN(n12018) );
  INV_X1 U15456 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U15457 ( .A1(n12056), .A2(n12019), .ZN(n12020) );
  NAND2_X1 U15458 ( .A1(n12021), .A2(n12020), .ZN(n14724) );
  OR2_X1 U15459 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12022) );
  NAND2_X1 U15460 ( .A1(n12023), .A2(n12022), .ZN(n14705) );
  NAND2_X1 U15461 ( .A1(n11947), .A2(n12026), .ZN(n12028) );
  OR2_X1 U15462 ( .A1(n14530), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12027) );
  INV_X1 U15463 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14908) );
  AOI22_X1 U15464 ( .A1(n12028), .A2(n12027), .B1(n12056), .B2(n14908), .ZN(
        n14692) );
  MUX2_X1 U15465 ( .A(n12047), .B(n12072), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12030) );
  OR2_X1 U15466 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12029) );
  NAND2_X1 U15467 ( .A1(n12050), .A2(n12031), .ZN(n12032) );
  INV_X1 U15468 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14905) );
  NAND2_X1 U15469 ( .A1(n12056), .A2(n14905), .ZN(n12033) );
  NAND2_X1 U15470 ( .A1(n12034), .A2(n12033), .ZN(n14660) );
  OR2_X1 U15471 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U15472 ( .A1(n12036), .A2(n12035), .ZN(n14649) );
  NAND2_X1 U15473 ( .A1(n11947), .A2(n15330), .ZN(n12037) );
  INV_X1 U15474 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21704) );
  NAND2_X1 U15475 ( .A1(n12056), .A2(n21704), .ZN(n12038) );
  OR2_X1 U15476 ( .A1(n12047), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n12042) );
  OAI211_X1 U15477 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14530), .A(n11947), .B(
        n12040), .ZN(n12041) );
  AND2_X1 U15478 ( .A1(n12042), .A2(n12041), .ZN(n14620) );
  INV_X1 U15479 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U15480 ( .A1(n11947), .A2(n15070), .ZN(n12043) );
  OAI211_X1 U15481 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n14530), .A(n12043), .B(
        n12072), .ZN(n12046) );
  INV_X1 U15482 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U15483 ( .A1(n12056), .A2(n12044), .ZN(n12045) );
  NAND2_X1 U15484 ( .A1(n12046), .A2(n12045), .ZN(n14606) );
  MUX2_X1 U15485 ( .A(n12047), .B(n12072), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12049) );
  OR2_X1 U15486 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U15487 ( .A1(n12049), .A2(n12048), .ZN(n14590) );
  INV_X1 U15488 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U15489 ( .A1(n12050), .A2(n15052), .ZN(n12051) );
  OAI211_X1 U15490 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n14530), .A(n12051), .B(
        n12072), .ZN(n12054) );
  INV_X1 U15491 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U15492 ( .A1(n12056), .A2(n12052), .ZN(n12053) );
  OR2_X1 U15493 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12055) );
  OR2_X1 U15494 ( .A1(n14530), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U15495 ( .A1(n12055), .A2(n12057), .ZN(n12058) );
  MUX2_X1 U15496 ( .A(n12058), .B(n12057), .S(n12056), .Z(n13209) );
  OAI22_X1 U15497 ( .A1(n14527), .A2(n12072), .B1(n12058), .B2(n14510), .ZN(
        n12060) );
  AND2_X1 U15498 ( .A1(n14530), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12059) );
  AOI21_X1 U15499 ( .B1(n14531), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12059), .ZN(
        n14526) );
  XNOR2_X1 U15500 ( .A(n12060), .B(n14526), .ZN(n14891) );
  OAI22_X1 U15501 ( .A1(n13428), .A2(n21581), .B1(n20829), .B2(n12062), .ZN(
        n12063) );
  INV_X1 U15502 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12100) );
  NAND2_X1 U15503 ( .A1(n12091), .A2(n13682), .ZN(n15372) );
  INV_X1 U15504 ( .A(n14243), .ZN(n21583) );
  NAND2_X1 U15505 ( .A1(n21583), .A2(n12065), .ZN(n12066) );
  AND2_X1 U15506 ( .A1(n12067), .A2(n12066), .ZN(n12084) );
  OAI21_X1 U15507 ( .B1(n12069), .B2(n20839), .A(n11551), .ZN(n12070) );
  OAI21_X1 U15508 ( .B1(n12070), .B2(n13684), .A(n21581), .ZN(n12071) );
  OAI211_X1 U15509 ( .C1(n12073), .C2(n12072), .A(n12084), .B(n12071), .ZN(
        n12074) );
  INV_X1 U15510 ( .A(n12074), .ZN(n12076) );
  NAND2_X1 U15511 ( .A1(n12076), .A2(n12075), .ZN(n13583) );
  OR2_X1 U15512 ( .A1(n12077), .A2(n13583), .ZN(n12078) );
  NAND2_X1 U15513 ( .A1(n12091), .A2(n12078), .ZN(n15366) );
  NAND2_X2 U15514 ( .A1(n15372), .A2(n15366), .ZN(n15510) );
  NAND2_X1 U15515 ( .A1(n15372), .A2(n13749), .ZN(n20783) );
  NAND2_X1 U15516 ( .A1(n15510), .A2(n20783), .ZN(n20766) );
  AND3_X1 U15517 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15485) );
  AND2_X1 U15518 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12079) );
  AND2_X1 U15519 ( .A1(n15485), .A2(n12079), .ZN(n15477) );
  NAND3_X1 U15520 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U15521 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20745) );
  NOR2_X1 U15522 ( .A1(n12080), .A2(n20745), .ZN(n12081) );
  AND2_X1 U15523 ( .A1(n15477), .A2(n12081), .ZN(n15461) );
  AND2_X1 U15524 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12082) );
  AND2_X1 U15525 ( .A1(n15461), .A2(n12082), .ZN(n15394) );
  INV_X1 U15526 ( .A(n15394), .ZN(n15452) );
  OR2_X1 U15527 ( .A1(n20766), .A2(n15452), .ZN(n12086) );
  NOR2_X1 U15528 ( .A1(n20745), .A2(n15273), .ZN(n12085) );
  NAND2_X1 U15529 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U15530 ( .A1(n20780), .A2(n20767), .ZN(n20743) );
  AND2_X1 U15531 ( .A1(n12085), .A2(n20743), .ZN(n15511) );
  AND3_X1 U15532 ( .A1(n15511), .A2(n15477), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U15533 ( .A1(n20770), .A2(n15445), .ZN(n15368) );
  NAND2_X1 U15534 ( .A1(n12086), .A2(n15368), .ZN(n15388) );
  AND2_X1 U15535 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U15536 ( .A1(n15388), .A2(n12087), .ZN(n15431) );
  NOR3_X1 U15537 ( .A1(n15177), .A2(n21716), .A3(n12088), .ZN(n12093) );
  INV_X1 U15538 ( .A(n12093), .ZN(n15406) );
  NOR2_X1 U15539 ( .A1(n15431), .A2(n15406), .ZN(n15408) );
  AND2_X1 U15540 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U15541 ( .A1(n15408), .A2(n12089), .ZN(n15377) );
  NAND2_X1 U15542 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12096) );
  OR2_X2 U15543 ( .A1(n15358), .A2(n12096), .ZN(n15344) );
  NAND2_X1 U15544 ( .A1(n10455), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12090) );
  NOR2_X1 U15545 ( .A1(n15344), .A2(n12090), .ZN(n13211) );
  NAND3_X1 U15546 ( .A1(n13211), .A2(n15298), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14540) );
  INV_X1 U15547 ( .A(n20782), .ZN(n15518) );
  INV_X1 U15548 ( .A(n15298), .ZN(n13212) );
  NOR2_X1 U15549 ( .A1(n15366), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12092) );
  OR2_X2 U15550 ( .A1(n12622), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20786) );
  NOR2_X1 U15551 ( .A1(n12091), .A2(n20731), .ZN(n15397) );
  NOR2_X1 U15552 ( .A1(n15460), .A2(n20782), .ZN(n12098) );
  INV_X1 U15553 ( .A(n12098), .ZN(n14536) );
  AND4_X1 U15554 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n12093), .ZN(n15370) );
  NAND2_X1 U15555 ( .A1(n15445), .A2(n15370), .ZN(n15371) );
  NAND2_X1 U15556 ( .A1(n15394), .A2(n15370), .ZN(n15375) );
  OAI21_X1 U15557 ( .B1(n15510), .B2(n15371), .A(n15375), .ZN(n12094) );
  NAND3_X1 U15558 ( .A1(n12094), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12095) );
  AOI21_X1 U15559 ( .B1(n12095), .B2(n20782), .A(n15460), .ZN(n15350) );
  NAND2_X1 U15560 ( .A1(n20782), .A2(n12096), .ZN(n12097) );
  AND2_X1 U15561 ( .A1(n15350), .A2(n12097), .ZN(n15332) );
  NAND2_X1 U15562 ( .A1(n20782), .A2(n15067), .ZN(n15322) );
  AND3_X1 U15563 ( .A1(n15332), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15322), .ZN(n15313) );
  NOR2_X1 U15564 ( .A1(n15313), .A2(n12098), .ZN(n15306) );
  AOI21_X1 U15565 ( .B1(n13212), .B2(n14536), .A(n15306), .ZN(n13210) );
  OAI211_X1 U15566 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15518), .A(
        n13210), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14537) );
  INV_X1 U15567 ( .A(n14537), .ZN(n12099) );
  AOI21_X1 U15568 ( .B1(n12100), .B2(n14540), .A(n12099), .ZN(n12102) );
  NAND2_X1 U15569 ( .A1(n20731), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n12626) );
  INV_X1 U15570 ( .A(n12626), .ZN(n12101) );
  AOI21_X1 U15571 ( .B1(n14891), .B2(n20756), .A(n12103), .ZN(n12104) );
  OAI21_X1 U15572 ( .B1(n12631), .B2(n20784), .A(n12104), .ZN(P1_U3001) );
  NAND2_X1 U15573 ( .A1(n12106), .A2(n12105), .ZN(n12112) );
  NAND2_X1 U15574 ( .A1(n12107), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12139) );
  XNOR2_X1 U15575 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15290) );
  AOI21_X1 U15576 ( .B1(n12587), .B2(n15290), .A(n14497), .ZN(n12109) );
  NAND2_X1 U15577 ( .A1(n14498), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12108) );
  OAI211_X1 U15578 ( .C1(n12139), .C2(n11673), .A(n12109), .B(n12108), .ZN(
        n12110) );
  INV_X1 U15579 ( .A(n12110), .ZN(n12111) );
  NAND2_X1 U15580 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  NAND2_X1 U15581 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15582 ( .A1(n12113), .A2(n12131), .ZN(n13999) );
  INV_X1 U15583 ( .A(n13999), .ZN(n12130) );
  NAND2_X1 U15584 ( .A1(n9702), .A2(n10567), .ZN(n12115) );
  NAND2_X1 U15585 ( .A1(n15549), .A2(n12105), .ZN(n12119) );
  INV_X2 U15586 ( .A(n10549), .ZN(n14498) );
  AOI22_X1 U15587 ( .A1(n14498), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21503), .ZN(n12117) );
  INV_X1 U15588 ( .A(n12139), .ZN(n12143) );
  NAND2_X1 U15589 ( .A1(n12143), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12116) );
  AND2_X1 U15590 ( .A1(n12117), .A2(n12116), .ZN(n12118) );
  NAND2_X1 U15591 ( .A1(n12119), .A2(n12118), .ZN(n13643) );
  INV_X1 U15592 ( .A(n12121), .ZN(n12122) );
  XNOR2_X1 U15593 ( .A(n12120), .B(n12122), .ZN(n20930) );
  NAND2_X1 U15594 ( .A1(n20930), .A2(n12105), .ZN(n12126) );
  AOI22_X1 U15595 ( .A1(n14498), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21503), .ZN(n12124) );
  NAND2_X1 U15596 ( .A1(n12143), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12123) );
  AND2_X1 U15597 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  NAND2_X1 U15598 ( .A1(n12126), .A2(n12125), .ZN(n13467) );
  AOI21_X1 U15599 ( .B1(n9587), .B2(n12127), .A(n21503), .ZN(n13466) );
  NAND2_X1 U15600 ( .A1(n13467), .A2(n13466), .ZN(n13465) );
  OR2_X1 U15601 ( .A1(n13467), .A2(n14228), .ZN(n12128) );
  NAND2_X1 U15602 ( .A1(n13465), .A2(n12128), .ZN(n13642) );
  NAND2_X1 U15603 ( .A1(n13643), .A2(n13642), .ZN(n13998) );
  NAND2_X1 U15604 ( .A1(n12130), .A2(n12129), .ZN(n13996) );
  NAND2_X1 U15605 ( .A1(n12132), .A2(n12105), .ZN(n12142) );
  NAND2_X1 U15606 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12134) );
  INV_X1 U15607 ( .A(n12134), .ZN(n12136) );
  NOR2_X1 U15608 ( .A1(n12134), .A2(n12133), .ZN(n12153) );
  INV_X1 U15609 ( .A(n12153), .ZN(n12135) );
  OAI21_X1 U15610 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12136), .A(
        n12135), .ZN(n15285) );
  AOI22_X1 U15611 ( .A1(n12619), .A2(n15285), .B1(n14497), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U15612 ( .A1(n14498), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12137) );
  OAI211_X1 U15613 ( .C1(n12139), .C2(n14056), .A(n12138), .B(n12137), .ZN(
        n12140) );
  INV_X1 U15614 ( .A(n12140), .ZN(n12141) );
  NAND2_X1 U15615 ( .A1(n14032), .A2(n14033), .ZN(n14101) );
  NAND2_X1 U15616 ( .A1(n12143), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12147) );
  INV_X1 U15617 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20656) );
  AOI21_X1 U15618 ( .B1(n20656), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12144) );
  AOI21_X1 U15619 ( .B1(n14498), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12144), .ZN(
        n12146) );
  XNOR2_X1 U15620 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n12153), .ZN(
        n20741) );
  NOR2_X1 U15621 ( .A1(n20741), .A2(n14228), .ZN(n12145) );
  AOI21_X1 U15622 ( .B1(n12147), .B2(n12146), .A(n12145), .ZN(n12148) );
  AOI21_X1 U15623 ( .B1(n12149), .B2(n12105), .A(n12148), .ZN(n14100) );
  NAND2_X1 U15624 ( .A1(n12152), .A2(n12105), .ZN(n12161) );
  NAND2_X1 U15625 ( .A1(n12163), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12166) );
  INV_X1 U15626 ( .A(n12166), .ZN(n12154) );
  NAND2_X1 U15627 ( .A1(n12154), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12190) );
  INV_X1 U15628 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U15629 ( .A1(n12166), .A2(n12155), .ZN(n12156) );
  NAND2_X1 U15630 ( .A1(n12190), .A2(n12156), .ZN(n20623) );
  NAND2_X1 U15631 ( .A1(n20623), .A2(n12619), .ZN(n12158) );
  NAND2_X1 U15632 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12157) );
  NAND2_X1 U15633 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  AOI21_X1 U15634 ( .B1(n14498), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12159), .ZN(
        n12160) );
  NAND2_X1 U15635 ( .A1(n12162), .A2(n12105), .ZN(n12171) );
  INV_X1 U15636 ( .A(n12163), .ZN(n12164) );
  INV_X1 U15637 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20625) );
  NAND2_X1 U15638 ( .A1(n12164), .A2(n20625), .ZN(n12165) );
  NAND2_X1 U15639 ( .A1(n12166), .A2(n12165), .ZN(n20636) );
  NAND2_X1 U15640 ( .A1(n20636), .A2(n12619), .ZN(n12168) );
  NAND2_X1 U15641 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12167) );
  NAND2_X1 U15642 ( .A1(n12168), .A2(n12167), .ZN(n12169) );
  AOI21_X1 U15643 ( .B1(n14498), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12169), .ZN(
        n12170) );
  NAND2_X1 U15644 ( .A1(n12171), .A2(n12170), .ZN(n14217) );
  AOI22_X1 U15645 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12602), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15646 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15647 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15648 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12449), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12172) );
  NAND4_X1 U15649 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n12181) );
  AOI22_X1 U15650 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11718), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15651 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12395), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15652 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15653 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12512), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12176) );
  NAND4_X1 U15654 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12180) );
  OAI21_X1 U15655 ( .B1(n12181), .B2(n12180), .A(n12105), .ZN(n12186) );
  NAND2_X1 U15656 ( .A1(n14498), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12185) );
  NAND2_X1 U15657 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12184) );
  INV_X1 U15658 ( .A(n12190), .ZN(n12182) );
  XNOR2_X1 U15659 ( .A(n12208), .B(n12207), .ZN(n15252) );
  NAND2_X1 U15660 ( .A1(n15252), .A2(n12619), .ZN(n12183) );
  NAND4_X1 U15661 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n14877) );
  NAND3_X1 U15662 ( .A1(n14875), .A2(n14217), .A3(n14877), .ZN(n12187) );
  NAND2_X1 U15663 ( .A1(n12188), .A2(n12105), .ZN(n12196) );
  INV_X1 U15664 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12189) );
  NAND2_X1 U15665 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  NAND2_X1 U15666 ( .A1(n12208), .A2(n12191), .ZN(n20602) );
  NAND2_X1 U15667 ( .A1(n20602), .A2(n12619), .ZN(n12193) );
  NAND2_X1 U15668 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U15669 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  AOI21_X1 U15670 ( .B1(n14498), .B2(P1_EAX_REG_7__SCAN_IN), .A(n12194), .ZN(
        n12195) );
  AOI22_X1 U15671 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15672 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15673 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15674 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15675 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12206) );
  AOI22_X1 U15676 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15677 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15678 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15679 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15680 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12205) );
  OAI21_X1 U15681 ( .B1(n12206), .B2(n12205), .A(n12105), .ZN(n12212) );
  NAND2_X1 U15682 ( .A1(n14498), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12211) );
  OAI21_X1 U15683 ( .B1(n12208), .B2(n12207), .A(n21702), .ZN(n12209) );
  NAND2_X1 U15684 ( .A1(n12209), .A2(n12240), .ZN(n15243) );
  AOI22_X1 U15685 ( .A1(n15243), .A2(n12619), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n14497), .ZN(n12210) );
  AOI22_X1 U15686 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15687 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15688 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15689 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15690 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12224) );
  AOI22_X1 U15691 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15692 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15693 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15694 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15695 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  OAI21_X1 U15696 ( .B1(n12224), .B2(n12223), .A(n12105), .ZN(n12228) );
  NAND2_X1 U15697 ( .A1(n14498), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12227) );
  XNOR2_X1 U15698 ( .A(n12240), .B(n14848), .ZN(n15235) );
  NAND2_X1 U15699 ( .A1(n15235), .A2(n12619), .ZN(n12226) );
  NAND2_X1 U15700 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12225) );
  AOI22_X1 U15701 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15702 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15703 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15704 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15705 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12238) );
  AOI22_X1 U15706 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15707 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15708 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15709 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U15710 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12237) );
  OR2_X1 U15711 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  INV_X1 U15712 ( .A(n14497), .ZN(n12344) );
  INV_X1 U15713 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14826) );
  NAND2_X1 U15714 ( .A1(n14498), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12245) );
  INV_X1 U15715 ( .A(n12281), .ZN(n12273) );
  INV_X1 U15716 ( .A(n12241), .ZN(n12242) );
  NAND2_X1 U15717 ( .A1(n12242), .A2(n14826), .ZN(n12243) );
  NAND2_X1 U15718 ( .A1(n12273), .A2(n12243), .ZN(n15224) );
  NAND2_X1 U15719 ( .A1(n15224), .A2(n12619), .ZN(n12244) );
  OAI211_X1 U15720 ( .C1(n12344), .C2(n14826), .A(n12245), .B(n12244), .ZN(
        n14789) );
  INV_X1 U15721 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12274) );
  OR2_X1 U15722 ( .A1(n12273), .A2(n12274), .ZN(n12247) );
  INV_X1 U15723 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12246) );
  XNOR2_X1 U15724 ( .A(n12247), .B(n12246), .ZN(n15204) );
  NAND2_X1 U15725 ( .A1(n15204), .A2(n12619), .ZN(n12262) );
  AOI22_X1 U15726 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15727 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15728 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15729 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12248) );
  NAND4_X1 U15730 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12257) );
  AOI22_X1 U15731 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15732 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15733 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15734 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15735 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12256) );
  OAI21_X1 U15736 ( .B1(n12257), .B2(n12256), .A(n12105), .ZN(n12260) );
  NAND2_X1 U15737 ( .A1(n14498), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15738 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12258) );
  AND3_X1 U15739 ( .A1(n12260), .A2(n12259), .A3(n12258), .ZN(n12261) );
  NAND2_X1 U15740 ( .A1(n12262), .A2(n12261), .ZN(n14796) );
  AOI22_X1 U15741 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12538), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15742 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15743 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15744 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U15745 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12272) );
  AOI22_X1 U15746 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15747 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15748 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15749 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15750 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12271) );
  NOR2_X1 U15751 ( .A1(n12272), .A2(n12271), .ZN(n12279) );
  INV_X1 U15752 ( .A(n12105), .ZN(n12278) );
  XNOR2_X1 U15753 ( .A(n12273), .B(n12274), .ZN(n15216) );
  NAND2_X1 U15754 ( .A1(n15216), .A2(n12619), .ZN(n12277) );
  NOR2_X1 U15755 ( .A1(n12344), .A2(n12274), .ZN(n12275) );
  AOI21_X1 U15756 ( .B1(n14498), .B2(P1_EAX_REG_12__SCAN_IN), .A(n12275), .ZN(
        n12276) );
  OAI211_X1 U15757 ( .C1(n12279), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        n14794) );
  OAI211_X1 U15758 ( .C1(n14793), .C2(n14789), .A(n14796), .B(n14794), .ZN(
        n12313) );
  NAND2_X1 U15759 ( .A1(n12330), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12283) );
  INV_X1 U15760 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12282) );
  XNOR2_X1 U15761 ( .A(n12283), .B(n12282), .ZN(n15181) );
  INV_X1 U15762 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U15763 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15764 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15765 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15766 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U15767 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12293) );
  AOI22_X1 U15768 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15769 ( .A1(n12497), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15770 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15771 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U15772 ( .A1(n12291), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12292) );
  OAI21_X1 U15773 ( .B1(n12293), .B2(n12292), .A(n12105), .ZN(n12295) );
  NAND2_X1 U15774 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12294) );
  OAI211_X1 U15775 ( .C1(n20669), .C2(n10549), .A(n12295), .B(n12294), .ZN(
        n12296) );
  AOI21_X1 U15776 ( .B1(n15181), .B2(n12619), .A(n12296), .ZN(n14768) );
  INV_X1 U15777 ( .A(n12330), .ZN(n12298) );
  INV_X1 U15778 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12297) );
  XNOR2_X1 U15779 ( .A(n12298), .B(n12297), .ZN(n15194) );
  AOI22_X1 U15780 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15781 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15782 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15783 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12299) );
  NAND4_X1 U15784 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12308) );
  AOI22_X1 U15785 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15786 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15787 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15788 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15789 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12307) );
  OAI21_X1 U15790 ( .B1(n12308), .B2(n12307), .A(n12105), .ZN(n12311) );
  NAND2_X1 U15791 ( .A1(n14498), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15792 ( .A1(n14497), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12309) );
  NAND3_X1 U15793 ( .A1(n12311), .A2(n12310), .A3(n12309), .ZN(n12312) );
  AOI21_X1 U15794 ( .B1(n15194), .B2(n12619), .A(n12312), .ZN(n14777) );
  NOR3_X1 U15795 ( .A1(n12313), .A2(n14768), .A3(n14777), .ZN(n12314) );
  INV_X1 U15796 ( .A(n15567), .ZN(n12315) );
  NAND2_X1 U15797 ( .A1(n12590), .A2(n14228), .ZN(n12434) );
  AOI22_X1 U15798 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15799 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12496), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12320) );
  AOI21_X1 U15800 ( .B1(n12597), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12619), .ZN(n12317) );
  NAND2_X1 U15801 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12316) );
  AND2_X1 U15802 ( .A1(n12317), .A2(n12316), .ZN(n12319) );
  AOI22_X1 U15803 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12318) );
  NAND4_X1 U15804 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n12327) );
  AOI22_X1 U15805 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12602), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15806 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11718), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15807 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15808 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n9607), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12322) );
  NAND4_X1 U15809 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12326) );
  OR2_X1 U15810 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND2_X1 U15811 ( .A1(n12434), .A2(n12328), .ZN(n12332) );
  AOI22_X1 U15812 ( .A1(n14498), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21503), .ZN(n12331) );
  XNOR2_X1 U15813 ( .A(n12366), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15171) );
  AOI22_X1 U15814 ( .A1(n12332), .A2(n12331), .B1(n12619), .B2(n15171), .ZN(
        n14747) );
  INV_X1 U15815 ( .A(n14731), .ZN(n12350) );
  INV_X1 U15816 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15168) );
  OR2_X1 U15817 ( .A1(n12366), .A2(n15168), .ZN(n12333) );
  INV_X1 U15818 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14740) );
  XNOR2_X1 U15819 ( .A(n12333), .B(n14740), .ZN(n15158) );
  NAND2_X1 U15820 ( .A1(n15158), .A2(n12619), .ZN(n12348) );
  AOI22_X1 U15821 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15822 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15823 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15824 ( .A1(n12497), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12334) );
  NAND4_X1 U15825 ( .A1(n12337), .A2(n12336), .A3(n12335), .A4(n12334), .ZN(
        n12343) );
  AOI22_X1 U15826 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12578), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15827 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15828 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15829 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12338) );
  NAND4_X1 U15830 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n12342) );
  OR2_X1 U15831 ( .A1(n12343), .A2(n12342), .ZN(n12346) );
  INV_X1 U15832 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15002) );
  OAI22_X1 U15833 ( .A1(n10549), .A2(n15002), .B1(n14740), .B2(n12344), .ZN(
        n12345) );
  AOI21_X1 U15834 ( .B1(n12616), .B2(n12346), .A(n12345), .ZN(n12347) );
  AOI22_X1 U15835 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15836 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15837 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15838 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12351) );
  NAND4_X1 U15839 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12362) );
  AOI22_X1 U15840 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15841 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15842 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U15843 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12356) );
  NAND2_X1 U15844 ( .A1(n12449), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12355) );
  AND3_X1 U15845 ( .A1(n12356), .A2(n12355), .A3(n14228), .ZN(n12357) );
  NAND4_X1 U15846 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12361) );
  OAI21_X1 U15847 ( .B1(n12362), .B2(n12361), .A(n12434), .ZN(n12364) );
  AOI22_X1 U15848 ( .A1(n14498), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21503), .ZN(n12363) );
  NAND2_X1 U15849 ( .A1(n12364), .A2(n12363), .ZN(n12368) );
  NAND2_X1 U15850 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12365) );
  XNOR2_X1 U15851 ( .A(n12369), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15146) );
  NAND2_X1 U15852 ( .A1(n15146), .A2(n12619), .ZN(n12367) );
  NAND2_X1 U15853 ( .A1(n12368), .A2(n12367), .ZN(n14723) );
  INV_X1 U15854 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15144) );
  INV_X1 U15855 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14714) );
  OAI21_X1 U15856 ( .B1(n12369), .B2(n15144), .A(n14714), .ZN(n12372) );
  NAND2_X1 U15857 ( .A1(n12372), .A2(n12389), .ZN(n15136) );
  OR2_X1 U15858 ( .A1(n15136), .A2(n14228), .ZN(n12388) );
  AOI22_X1 U15859 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15860 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15861 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15862 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15863 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12382) );
  AOI22_X1 U15864 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15865 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15866 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15867 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15868 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12381) );
  NOR2_X1 U15869 ( .A1(n12382), .A2(n12381), .ZN(n12386) );
  NAND2_X1 U15870 ( .A1(n21503), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12383) );
  NAND2_X1 U15871 ( .A1(n14228), .A2(n12383), .ZN(n12384) );
  AOI21_X1 U15872 ( .B1(n14498), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12384), .ZN(
        n12385) );
  OAI21_X1 U15873 ( .B1(n12590), .B2(n12386), .A(n12385), .ZN(n12387) );
  NAND2_X1 U15874 ( .A1(n12389), .A2(n21627), .ZN(n12390) );
  AND2_X1 U15875 ( .A1(n12407), .A2(n12390), .ZN(n15129) );
  AOI22_X1 U15876 ( .A1(n14498), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21503), .ZN(n12406) );
  AOI22_X1 U15877 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15878 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15879 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15880 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12409), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15881 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12404) );
  INV_X1 U15882 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15883 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12395), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12397) );
  AOI21_X1 U15884 ( .B1(n12604), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n12619), .ZN(n12396) );
  OAI211_X1 U15885 ( .C1(n11596), .C2(n12398), .A(n12397), .B(n12396), .ZN(
        n12399) );
  INV_X1 U15886 ( .A(n12399), .ZN(n12402) );
  AOI22_X1 U15887 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15888 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12400) );
  NAND3_X1 U15889 ( .A1(n12402), .A2(n12401), .A3(n12400), .ZN(n12403) );
  OAI21_X1 U15890 ( .B1(n12404), .B2(n12403), .A(n12434), .ZN(n12405) );
  AOI22_X1 U15891 ( .A1(n15129), .A2(n12619), .B1(n12406), .B2(n12405), .ZN(
        n14691) );
  OAI21_X1 U15892 ( .B1(n12408), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n12439), .ZN(n15120) );
  INV_X1 U15893 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14984) );
  AOI22_X1 U15894 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12604), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15895 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15896 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15897 ( .A1(n12409), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12410) );
  NAND4_X1 U15898 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n12410), .ZN(
        n12419) );
  AOI22_X1 U15899 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15900 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15901 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15902 ( .A1(n12449), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15903 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12418) );
  OAI21_X1 U15904 ( .B1(n12419), .B2(n12418), .A(n12616), .ZN(n12421) );
  OAI21_X1 U15905 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21373), .A(
        n21503), .ZN(n12420) );
  OAI211_X1 U15906 ( .C1(n10549), .C2(n14984), .A(n12421), .B(n12420), .ZN(
        n12422) );
  OAI21_X1 U15907 ( .B1(n15120), .B2(n14228), .A(n12422), .ZN(n14678) );
  XNOR2_X1 U15908 ( .A(n12439), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14663) );
  AOI22_X1 U15909 ( .A1(n14498), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21503), .ZN(n12438) );
  AOI22_X1 U15910 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15911 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15912 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15913 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12423) );
  NAND4_X1 U15914 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        n12436) );
  INV_X1 U15915 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15916 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12428) );
  AOI21_X1 U15917 ( .B1(n12604), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12619), .ZN(n12427) );
  OAI211_X1 U15918 ( .C1(n11596), .C2(n12429), .A(n12428), .B(n12427), .ZN(
        n12430) );
  INV_X1 U15919 ( .A(n12430), .ZN(n12433) );
  AOI22_X1 U15920 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12602), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15921 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12431) );
  NAND3_X1 U15922 ( .A1(n12433), .A2(n12432), .A3(n12431), .ZN(n12435) );
  OAI21_X1 U15923 ( .B1(n12436), .B2(n12435), .A(n12434), .ZN(n12437) );
  AOI22_X1 U15924 ( .A1(n14663), .A2(n12619), .B1(n12438), .B2(n12437), .ZN(
        n14658) );
  INV_X1 U15925 ( .A(n12439), .ZN(n12440) );
  INV_X1 U15926 ( .A(n12441), .ZN(n12443) );
  INV_X1 U15927 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15928 ( .A1(n12443), .A2(n12442), .ZN(n12444) );
  NAND2_X1 U15929 ( .A1(n12487), .A2(n12444), .ZN(n15100) );
  AOI22_X1 U15930 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15931 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15932 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15933 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U15934 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12455) );
  AOI22_X1 U15935 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12496), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15936 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12603), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15937 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12395), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15938 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12577), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12450) );
  NAND4_X1 U15939 ( .A1(n12453), .A2(n12452), .A3(n12451), .A4(n12450), .ZN(
        n12454) );
  NOR2_X1 U15940 ( .A1(n12455), .A2(n12454), .ZN(n12483) );
  AOI22_X1 U15941 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15942 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15943 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15944 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15945 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12466) );
  AOI22_X1 U15946 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15947 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15948 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15949 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15950 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12465) );
  NOR2_X1 U15951 ( .A1(n12466), .A2(n12465), .ZN(n12482) );
  XNOR2_X1 U15952 ( .A(n12483), .B(n12482), .ZN(n12469) );
  OAI21_X1 U15953 ( .B1(n21373), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n21503), .ZN(n12468) );
  NAND2_X1 U15954 ( .A1(n14498), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n12467) );
  OAI211_X1 U15955 ( .C1(n12590), .C2(n12469), .A(n12468), .B(n12467), .ZN(
        n12470) );
  OAI21_X1 U15956 ( .B1(n15100), .B2(n14228), .A(n12470), .ZN(n14646) );
  XNOR2_X1 U15957 ( .A(n12487), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15095) );
  INV_X1 U15958 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15091) );
  NOR2_X1 U15959 ( .A1(n15091), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12471) );
  AOI211_X1 U15960 ( .C1(n14498), .C2(P1_EAX_REG_24__SCAN_IN), .A(n12619), .B(
        n12471), .ZN(n12486) );
  AOI22_X1 U15961 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15962 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15963 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15964 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12472) );
  NAND4_X1 U15965 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12481) );
  AOI22_X1 U15966 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15967 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15968 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15969 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15970 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  OR2_X1 U15971 ( .A1(n12481), .A2(n12480), .ZN(n12504) );
  NOR2_X1 U15972 ( .A1(n12483), .A2(n12482), .ZN(n12505) );
  XOR2_X1 U15973 ( .A(n12504), .B(n12505), .Z(n12484) );
  NAND2_X1 U15974 ( .A1(n12484), .A2(n12616), .ZN(n12485) );
  AOI22_X1 U15975 ( .A1(n15095), .A2(n12619), .B1(n12486), .B2(n12485), .ZN(
        n14634) );
  NAND2_X1 U15976 ( .A1(n14633), .A2(n14634), .ZN(n14618) );
  NAND2_X1 U15977 ( .A1(n12489), .A2(n12488), .ZN(n12490) );
  NAND2_X1 U15978 ( .A1(n12529), .A2(n12490), .ZN(n15083) );
  AOI22_X1 U15979 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15980 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15981 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15982 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12492) );
  NAND4_X1 U15983 ( .A1(n12495), .A2(n12494), .A3(n12493), .A4(n12492), .ZN(
        n12503) );
  AOI22_X1 U15984 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12496), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15985 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12497), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15986 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15987 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12498) );
  NAND4_X1 U15988 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n12502) );
  NOR2_X1 U15989 ( .A1(n12503), .A2(n12502), .ZN(n12524) );
  NAND2_X1 U15990 ( .A1(n12505), .A2(n12504), .ZN(n12523) );
  XNOR2_X1 U15991 ( .A(n12524), .B(n12523), .ZN(n12508) );
  AOI21_X1 U15992 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21503), .A(
        n12619), .ZN(n12507) );
  NAND2_X1 U15993 ( .A1(n14498), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12506) );
  OAI211_X1 U15994 ( .C1(n12508), .C2(n12590), .A(n12507), .B(n12506), .ZN(
        n12509) );
  OAI21_X1 U15995 ( .B1(n15083), .B2(n14228), .A(n12509), .ZN(n14619) );
  XNOR2_X1 U15996 ( .A(n12529), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14609) );
  AOI21_X1 U15997 ( .B1(n12528), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12510) );
  AOI21_X1 U15998 ( .B1(n14498), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12510), .ZN(
        n12527) );
  AOI22_X1 U15999 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U16000 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U16001 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U16002 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12513) );
  NAND4_X1 U16003 ( .A1(n12516), .A2(n12515), .A3(n12514), .A4(n12513), .ZN(
        n12522) );
  AOI22_X1 U16004 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11718), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U16005 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U16006 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U16007 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12517) );
  NAND4_X1 U16008 ( .A1(n12520), .A2(n12519), .A3(n12518), .A4(n12517), .ZN(
        n12521) );
  NOR2_X1 U16009 ( .A1(n12524), .A2(n12523), .ZN(n12546) );
  XOR2_X1 U16010 ( .A(n12545), .B(n12546), .Z(n12525) );
  NAND2_X1 U16011 ( .A1(n12525), .A2(n12616), .ZN(n12526) );
  AOI22_X1 U16012 ( .A1(n14609), .A2(n12619), .B1(n12527), .B2(n12526), .ZN(
        n14604) );
  INV_X1 U16013 ( .A(n12530), .ZN(n12532) );
  INV_X1 U16014 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U16015 ( .A1(n12532), .A2(n12531), .ZN(n12533) );
  NAND2_X1 U16016 ( .A1(n12567), .A2(n12533), .ZN(n15063) );
  AOI22_X1 U16017 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U16018 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U16019 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12577), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U16020 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12534) );
  NAND4_X1 U16021 ( .A1(n12537), .A2(n12536), .A3(n12535), .A4(n12534), .ZN(
        n12544) );
  AOI22_X1 U16022 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U16023 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U16024 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U16025 ( .A1(n12538), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12539) );
  NAND4_X1 U16026 ( .A1(n12542), .A2(n12541), .A3(n12540), .A4(n12539), .ZN(
        n12543) );
  NOR2_X1 U16027 ( .A1(n12544), .A2(n12543), .ZN(n12563) );
  NAND2_X1 U16028 ( .A1(n12546), .A2(n12545), .ZN(n12562) );
  XNOR2_X1 U16029 ( .A(n12563), .B(n12562), .ZN(n12549) );
  AOI21_X1 U16030 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21503), .A(
        n12619), .ZN(n12548) );
  NAND2_X1 U16031 ( .A1(n14498), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12547) );
  OAI211_X1 U16032 ( .C1(n12549), .C2(n12590), .A(n12548), .B(n12547), .ZN(
        n12550) );
  OAI21_X1 U16033 ( .B1(n15063), .B2(n14228), .A(n12550), .ZN(n14589) );
  XNOR2_X1 U16034 ( .A(n12567), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15057) );
  INV_X1 U16035 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15054) );
  NOR2_X1 U16036 ( .A1(n15054), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12551) );
  AOI211_X1 U16037 ( .C1(n14498), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12619), .B(
        n12551), .ZN(n12566) );
  AOI22_X1 U16038 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U16039 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U16040 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U16041 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12552) );
  NAND4_X1 U16042 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12561) );
  AOI22_X1 U16043 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U16044 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U16045 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U16046 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U16047 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12560) );
  OR2_X1 U16048 ( .A1(n12561), .A2(n12560), .ZN(n12585) );
  NOR2_X1 U16049 ( .A1(n12563), .A2(n12562), .ZN(n12586) );
  XOR2_X1 U16050 ( .A(n12585), .B(n12586), .Z(n12564) );
  NAND2_X1 U16051 ( .A1(n12564), .A2(n12616), .ZN(n12565) );
  AOI22_X1 U16052 ( .A1(n15057), .A2(n12619), .B1(n12566), .B2(n12565), .ZN(
        n14506) );
  INV_X1 U16053 ( .A(n12567), .ZN(n12568) );
  INV_X1 U16054 ( .A(n12569), .ZN(n12571) );
  INV_X1 U16055 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U16056 ( .A1(n12571), .A2(n12570), .ZN(n12572) );
  NAND2_X1 U16057 ( .A1(n14221), .A2(n12572), .ZN(n15041) );
  AOI22_X1 U16058 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U16059 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U16060 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U16061 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U16062 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12584) );
  AOI22_X1 U16063 ( .A1(n12577), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U16064 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U16065 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U16066 ( .A1(n12578), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12579) );
  NAND4_X1 U16067 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12583) );
  NOR2_X1 U16068 ( .A1(n12584), .A2(n12583), .ZN(n12594) );
  NAND2_X1 U16069 ( .A1(n12586), .A2(n12585), .ZN(n12593) );
  XNOR2_X1 U16070 ( .A(n12594), .B(n12593), .ZN(n12591) );
  AOI21_X1 U16071 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21503), .A(
        n12587), .ZN(n12589) );
  NAND2_X1 U16072 ( .A1(n14498), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12588) );
  OAI211_X1 U16073 ( .C1(n12591), .C2(n12590), .A(n12589), .B(n12588), .ZN(
        n12592) );
  OAI21_X1 U16074 ( .B1(n15041), .B2(n14228), .A(n12592), .ZN(n14577) );
  XNOR2_X1 U16075 ( .A(n14221), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14567) );
  NOR2_X1 U16076 ( .A1(n12594), .A2(n12593), .ZN(n12613) );
  AOI22_X1 U16077 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U16078 ( .A1(n11613), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12449), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U16079 ( .A1(n12596), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U16080 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12597), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12598) );
  NAND4_X1 U16081 ( .A1(n12601), .A2(n12600), .A3(n12599), .A4(n12598), .ZN(
        n12611) );
  AOI22_X1 U16082 ( .A1(n12602), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U16083 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12603), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U16084 ( .A1(n12604), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U16085 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9599), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12606) );
  NAND4_X1 U16086 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12610) );
  NOR2_X1 U16087 ( .A1(n12611), .A2(n12610), .ZN(n12612) );
  XNOR2_X1 U16088 ( .A(n12613), .B(n12612), .ZN(n12617) );
  INV_X1 U16089 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16090 ( .A1(n21503), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12614) );
  OAI211_X1 U16091 ( .C1(n10549), .C2(n13202), .A(n14228), .B(n12614), .ZN(
        n12615) );
  AOI21_X1 U16092 ( .B1(n12617), .B2(n12616), .A(n12615), .ZN(n12618) );
  AOI21_X1 U16093 ( .B1(n14567), .B2(n12619), .A(n12618), .ZN(n14496) );
  INV_X1 U16094 ( .A(n14496), .ZN(n12620) );
  XNOR2_X1 U16095 ( .A(n14576), .B(n12620), .ZN(n14566) );
  NAND3_X1 U16096 ( .A1(n21501), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n17319) );
  INV_X1 U16097 ( .A(n17319), .ZN(n12621) );
  INV_X1 U16098 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12628) );
  NAND2_X1 U16099 ( .A1(n21433), .A2(n12622), .ZN(n21589) );
  NAND2_X1 U16100 ( .A1(n21589), .A2(n21501), .ZN(n12623) );
  NAND2_X1 U16101 ( .A1(n21501), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12625) );
  NAND2_X1 U16102 ( .A1(n21373), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U16103 ( .A1(n12625), .A2(n12624), .ZN(n13729) );
  NAND2_X1 U16104 ( .A1(n14567), .A2(n15172), .ZN(n12627) );
  OAI211_X1 U16105 ( .C1(n12628), .C2(n15169), .A(n12627), .B(n12626), .ZN(
        n12629) );
  AOI21_X1 U16106 ( .B1(n14566), .B2(n20737), .A(n12629), .ZN(n12630) );
  OAI21_X1 U16107 ( .B1(n12631), .B2(n20574), .A(n12630), .ZN(P1_U2969) );
  INV_X1 U16108 ( .A(n12632), .ZN(n12633) );
  INV_X1 U16109 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20413) );
  NOR2_X1 U16110 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20421) );
  INV_X1 U16111 ( .A(n20421), .ZN(n20414) );
  AND2_X1 U16112 ( .A1(n20560), .A2(n20547), .ZN(n14366) );
  INV_X1 U16113 ( .A(n12641), .ZN(n12634) );
  NAND2_X1 U16114 ( .A1(n10130), .A2(n12634), .ZN(n12640) );
  NAND2_X1 U16115 ( .A1(n12645), .A2(n12635), .ZN(n12639) );
  NAND2_X1 U16116 ( .A1(n17030), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13492) );
  AOI21_X1 U16117 ( .B1(n12645), .B2(n12644), .A(n12649), .ZN(n12646) );
  NAND2_X1 U16118 ( .A1(n12652), .A2(n20550), .ZN(n12648) );
  NAND2_X1 U16119 ( .A1(n12648), .A2(n12647), .ZN(n12653) );
  INV_X1 U16120 ( .A(n13492), .ZN(n12650) );
  NAND2_X1 U16121 ( .A1(n14363), .A2(n20549), .ZN(n12669) );
  OAI21_X1 U16122 ( .B1(n13527), .B2(n12656), .A(n12867), .ZN(n12663) );
  NAND2_X1 U16123 ( .A1(n17030), .A2(n19879), .ZN(n12658) );
  OAI211_X1 U16124 ( .C1(n10921), .C2(n20549), .A(n12867), .B(n12658), .ZN(
        n12659) );
  NAND3_X1 U16125 ( .A1(n12660), .A2(n14366), .A3(n13330), .ZN(n12662) );
  NAND2_X1 U16126 ( .A1(n12657), .A2(n19879), .ZN(n12661) );
  NAND2_X1 U16127 ( .A1(n12661), .A2(n20557), .ZN(n12876) );
  MUX2_X1 U16128 ( .A(n12660), .B(n19856), .S(n10916), .Z(n12665) );
  INV_X1 U16129 ( .A(n20547), .ZN(n20553) );
  NOR2_X1 U16130 ( .A1(n14374), .A2(n20553), .ZN(n12664) );
  NAND2_X1 U16131 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  AND3_X1 U16132 ( .A1(n13332), .A2(n12667), .A3(n12666), .ZN(n12668) );
  OAI21_X1 U16133 ( .B1(n20538), .B2(n12669), .A(n12668), .ZN(n12670) );
  INV_X1 U16134 ( .A(n12670), .ZN(n12671) );
  NAND2_X1 U16135 ( .A1(n12672), .A2(n12673), .ZN(n12674) );
  NAND2_X1 U16136 ( .A1(n9615), .A2(n12674), .ZN(n19730) );
  NAND2_X1 U16137 ( .A1(n12676), .A2(n16235), .ZN(n12677) );
  NAND2_X1 U16138 ( .A1(n12677), .A2(n10931), .ZN(n12678) );
  NAND2_X1 U16139 ( .A1(n12680), .A2(n20549), .ZN(n12683) );
  NAND2_X1 U16140 ( .A1(n12681), .A2(n12682), .ZN(n14103) );
  NAND2_X1 U16141 ( .A1(n12683), .A2(n14103), .ZN(n12684) );
  NAND2_X1 U16142 ( .A1(n13027), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12687) );
  NOR2_X1 U16143 ( .A1(n19879), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U16144 ( .A1(n12848), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12686) );
  AND2_X1 U16145 ( .A1(n12687), .A2(n12686), .ZN(n12862) );
  NAND2_X1 U16146 ( .A1(n13527), .A2(n12854), .ZN(n12710) );
  MUX2_X1 U16147 ( .A(n19879), .B(n20531), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12691) );
  NAND2_X1 U16148 ( .A1(n12692), .A2(n10566), .ZN(n13291) );
  NAND2_X1 U16149 ( .A1(n13027), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12696) );
  INV_X1 U16150 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13532) );
  OAI211_X1 U16151 ( .C1(n19879), .C2(n13532), .A(n12693), .B(n20501), .ZN(
        n12694) );
  INV_X1 U16152 ( .A(n12694), .ZN(n12695) );
  NAND2_X1 U16153 ( .A1(n12696), .A2(n12695), .ZN(n13292) );
  AOI22_X1 U16154 ( .A1(n12697), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12854), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12698) );
  XNOR2_X1 U16155 ( .A(n12705), .B(n12706), .ZN(n13472) );
  NOR2_X1 U16156 ( .A1(n13527), .A2(n12699), .ZN(n12700) );
  MUX2_X1 U16157 ( .A(n12700), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n12704) );
  INV_X1 U16158 ( .A(n12701), .ZN(n12702) );
  NOR2_X1 U16159 ( .A1(n9663), .A2(n12702), .ZN(n12703) );
  NOR2_X1 U16160 ( .A1(n12704), .A2(n12703), .ZN(n13471) );
  INV_X1 U16161 ( .A(n12706), .ZN(n12707) );
  NAND2_X1 U16162 ( .A1(n12705), .A2(n12707), .ZN(n12708) );
  NAND2_X1 U16163 ( .A1(n13474), .A2(n12708), .ZN(n12716) );
  OR2_X1 U16164 ( .A1(n9663), .A2(n12709), .ZN(n12711) );
  OAI211_X1 U16165 ( .C1(n20501), .C2(n20512), .A(n12711), .B(n12710), .ZN(
        n12714) );
  XNOR2_X1 U16166 ( .A(n12716), .B(n12714), .ZN(n13242) );
  NAND2_X1 U16167 ( .A1(n13027), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U16168 ( .A1(n12697), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12712) );
  AND2_X1 U16169 ( .A1(n12713), .A2(n12712), .ZN(n13241) );
  INV_X1 U16170 ( .A(n12714), .ZN(n12715) );
  NAND2_X1 U16171 ( .A1(n12716), .A2(n12715), .ZN(n12717) );
  INV_X1 U16172 ( .A(n9663), .ZN(n12803) );
  AOI22_X1 U16173 ( .A1(n12803), .A2(n12718), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n12697), .ZN(n12721) );
  OAI22_X1 U16174 ( .A1(n13024), .A2(n17354), .B1(n20505), .B2(n20501), .ZN(
        n12719) );
  AOI21_X1 U16175 ( .B1(n13027), .B2(P2_REIP_REG_3__SCAN_IN), .A(n12719), .ZN(
        n12720) );
  AND2_X1 U16176 ( .A1(n12721), .A2(n12720), .ZN(n15915) );
  NAND2_X1 U16177 ( .A1(n13027), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U16178 ( .A1(n12697), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12725) );
  OR2_X1 U16179 ( .A1(n9663), .A2(n12723), .ZN(n12724) );
  NAND2_X1 U16180 ( .A1(n13027), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U16182 ( .A1(n12848), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12729) );
  OR2_X1 U16183 ( .A1(n9663), .A2(n12727), .ZN(n12728) );
  OAI21_X2 U16184 ( .B1(n15884), .B2(n15885), .A(n12732), .ZN(n13547) );
  AOI22_X1 U16185 ( .A1(n12848), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12734) );
  OAI21_X1 U16186 ( .B1(n12733), .B2(n20438), .A(n12734), .ZN(n13546) );
  NAND2_X1 U16187 ( .A1(n13547), .A2(n13546), .ZN(n12736) );
  OR2_X1 U16188 ( .A1(n9663), .A2(n11143), .ZN(n12735) );
  AOI22_X1 U16189 ( .A1(n12848), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12737) );
  OAI21_X1 U16190 ( .B1(n12733), .B2(n20440), .A(n12737), .ZN(n13550) );
  NAND2_X1 U16191 ( .A1(n13027), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16192 ( .A1(n12848), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16193 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U16194 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U16195 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U16196 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U16197 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12747) );
  AOI22_X1 U16198 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14409), .ZN(n12745) );
  AOI22_X1 U16199 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U16200 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11044), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U16201 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U16202 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12746) );
  INV_X1 U16203 ( .A(n16304), .ZN(n12748) );
  OR2_X1 U16204 ( .A1(n9663), .A2(n12748), .ZN(n12749) );
  NAND2_X1 U16205 ( .A1(n13027), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16206 ( .A1(n12848), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13026), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U16207 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n16041), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16208 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11026), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U16209 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16210 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11069), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12752) );
  NAND4_X1 U16211 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12762) );
  AOI22_X1 U16212 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n14409), .ZN(n12760) );
  AOI22_X1 U16213 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16214 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U16215 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11044), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U16216 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  INV_X1 U16217 ( .A(n16313), .ZN(n16292) );
  OR2_X1 U16218 ( .A1(n9663), .A2(n16292), .ZN(n12763) );
  INV_X1 U16219 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20447) );
  AOI22_X1 U16220 ( .A1(n12697), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16221 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16222 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16223 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16224 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12767) );
  NAND4_X1 U16225 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12776) );
  AOI22_X1 U16226 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14409), .ZN(n12774) );
  AOI22_X1 U16227 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16228 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11044), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U16229 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12771) );
  NAND4_X1 U16230 ( .A1(n12774), .A2(n12773), .A3(n12772), .A4(n12771), .ZN(
        n12775) );
  OR2_X1 U16231 ( .A1(n12776), .A2(n12775), .ZN(n16294) );
  NAND2_X1 U16232 ( .A1(n12803), .A2(n16294), .ZN(n12777) );
  OAI211_X1 U16233 ( .C1(n12733), .C2(n20447), .A(n12778), .B(n12777), .ZN(
        n13271) );
  NAND2_X1 U16234 ( .A1(n13027), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16235 ( .A1(n12848), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U16236 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16237 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12781) );
  AOI22_X1 U16238 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U16239 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12779) );
  NAND4_X1 U16240 ( .A1(n12782), .A2(n12781), .A3(n12780), .A4(n12779), .ZN(
        n12788) );
  AOI22_X1 U16241 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14409), .ZN(n12786) );
  AOI22_X1 U16242 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U16243 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11044), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16244 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12783) );
  NAND4_X1 U16245 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12787) );
  INV_X1 U16246 ( .A(n14085), .ZN(n16298) );
  OR2_X1 U16247 ( .A1(n9663), .A2(n16298), .ZN(n12789) );
  INV_X1 U16248 ( .A(n13639), .ZN(n13269) );
  AND2_X1 U16249 ( .A1(n13271), .A2(n13269), .ZN(n12792) );
  NAND2_X1 U16250 ( .A1(n13027), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U16251 ( .A1(n12848), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16252 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n16041), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16253 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14107), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U16254 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U16255 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12793) );
  NAND4_X1 U16256 ( .A1(n12796), .A2(n12795), .A3(n12794), .A4(n12793), .ZN(
        n12802) );
  AOI22_X1 U16257 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11069), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U16258 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16259 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11044), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U16260 ( .A1(n11091), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14409), .ZN(n12797) );
  NAND4_X1 U16261 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12801) );
  NAND2_X1 U16262 ( .A1(n12803), .A2(n14096), .ZN(n12804) );
  NAND2_X1 U16263 ( .A1(n13027), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16264 ( .A1(n12848), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U16265 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16266 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U16267 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U16268 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12809) );
  NAND4_X1 U16269 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12809), .ZN(
        n12818) );
  AOI22_X1 U16270 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n14409), .ZN(n12816) );
  AOI22_X1 U16271 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16272 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11044), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16273 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12813) );
  NAND4_X1 U16274 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12817) );
  INV_X1 U16275 ( .A(n14318), .ZN(n14298) );
  OR2_X1 U16276 ( .A1(n9663), .A2(n14298), .ZN(n12819) );
  AOI22_X1 U16277 ( .A1(n12848), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16278 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n16041), .B1(
        n16042), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U16279 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n14107), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U16280 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16281 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12822) );
  NAND4_X1 U16282 ( .A1(n12825), .A2(n12824), .A3(n12823), .A4(n12822), .ZN(
        n12831) );
  AOI22_X1 U16283 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14409), .ZN(n12829) );
  AOI22_X1 U16284 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11069), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U16285 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n9589), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U16286 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11044), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12826) );
  NAND4_X1 U16287 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        n12830) );
  INV_X1 U16288 ( .A(n14317), .ZN(n12832) );
  OR2_X1 U16289 ( .A1(n9663), .A2(n12832), .ZN(n12833) );
  OAI211_X1 U16290 ( .C1(n12733), .C2(n20453), .A(n12834), .B(n12833), .ZN(
        n14025) );
  NAND2_X1 U16291 ( .A1(n13027), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12847) );
  INV_X1 U16292 ( .A(n13025), .ZN(n12848) );
  AOI22_X1 U16293 ( .A1(n12848), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U16294 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U16295 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16296 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16297 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12835) );
  NAND4_X1 U16298 ( .A1(n12838), .A2(n12837), .A3(n12836), .A4(n12835), .ZN(
        n12844) );
  AOI22_X1 U16299 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14409), .ZN(n12842) );
  AOI22_X1 U16300 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U16301 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11044), .B1(
        n16048), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U16302 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12839) );
  NAND4_X1 U16303 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n12843) );
  INV_X1 U16304 ( .A(n14401), .ZN(n14306) );
  OR2_X1 U16305 ( .A1(n9663), .A2(n14306), .ZN(n12845) );
  NAND2_X1 U16306 ( .A1(n13027), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U16307 ( .A1(n12848), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12849) );
  NOR2_X2 U16308 ( .A1(n14049), .A2(n14324), .ZN(n14322) );
  AOI22_X1 U16309 ( .A1(n12848), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U16310 ( .B1(n12733), .B2(n20459), .A(n12851), .ZN(n14417) );
  INV_X1 U16311 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U16312 ( .A1(n12697), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U16313 ( .B1(n12733), .B2(n12853), .A(n12852), .ZN(n15741) );
  NAND2_X1 U16314 ( .A1(n13027), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U16315 ( .A1(n12848), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12855) );
  INV_X1 U16316 ( .A(n13011), .ZN(n12861) );
  AOI21_X1 U16317 ( .B1(n12862), .B2(n15723), .A(n12861), .ZN(n19731) );
  INV_X1 U16318 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n12863) );
  NOR2_X1 U16319 ( .A1(n17339), .A2(n12863), .ZN(n12920) );
  NAND2_X1 U16320 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13484) );
  INV_X1 U16321 ( .A(n13484), .ZN(n13235) );
  NAND2_X1 U16322 ( .A1(n13237), .A2(n13484), .ZN(n12885) );
  OR2_X1 U16323 ( .A1(n12864), .A2(n12865), .ZN(n12866) );
  MUX2_X1 U16324 ( .A(n12867), .B(n12866), .S(n20550), .Z(n12880) );
  INV_X1 U16325 ( .A(n13524), .ZN(n13303) );
  OAI21_X1 U16326 ( .B1(n9996), .B2(n12647), .A(n13303), .ZN(n12874) );
  INV_X1 U16327 ( .A(n12869), .ZN(n12870) );
  NAND2_X1 U16328 ( .A1(n12872), .A2(n12871), .ZN(n13521) );
  AND3_X1 U16329 ( .A1(n12874), .A2(n12873), .A3(n13521), .ZN(n12879) );
  NAND2_X1 U16330 ( .A1(n12875), .A2(n20549), .ZN(n14345) );
  NAND2_X1 U16331 ( .A1(n14345), .A2(n12876), .ZN(n12877) );
  NAND2_X1 U16332 ( .A1(n12877), .A2(n19860), .ZN(n12878) );
  NAND2_X1 U16333 ( .A1(n14350), .A2(n10932), .ZN(n12881) );
  NAND2_X1 U16334 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16943) );
  INV_X1 U16335 ( .A(n16885), .ZN(n13065) );
  NAND2_X1 U16336 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n13065), .ZN(
        n12894) );
  INV_X1 U16337 ( .A(n12894), .ZN(n12882) );
  AOI211_X1 U16338 ( .C1(n12883), .C2(n16825), .A(n13118), .B(n16824), .ZN(
        n12884) );
  AOI211_X1 U16339 ( .C1(n17327), .C2(n19731), .A(n12920), .B(n12884), .ZN(
        n12899) );
  NAND2_X1 U16340 ( .A1(n16974), .A2(n16973), .ZN(n12889) );
  NAND2_X1 U16341 ( .A1(n16850), .A2(n17354), .ZN(n17341) );
  INV_X1 U16342 ( .A(n13478), .ZN(n13286) );
  INV_X1 U16343 ( .A(n13236), .ZN(n16848) );
  AOI21_X1 U16344 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13235), .A(
        n16848), .ZN(n12887) );
  INV_X1 U16345 ( .A(n12885), .ZN(n12886) );
  AND2_X1 U16346 ( .A1(n16844), .A2(n12886), .ZN(n13252) );
  AND2_X1 U16347 ( .A1(n17341), .A2(n17355), .ZN(n16978) );
  OAI21_X1 U16348 ( .B1(n17338), .B2(n16703), .A(n16850), .ZN(n12888) );
  NAND2_X1 U16349 ( .A1(n12889), .A2(n16967), .ZN(n16954) );
  AND2_X1 U16350 ( .A1(n16850), .A2(n16943), .ZN(n12890) );
  AND2_X1 U16351 ( .A1(n16850), .A2(n16930), .ZN(n12891) );
  NAND2_X1 U16352 ( .A1(n16850), .A2(n12892), .ZN(n12893) );
  NAND2_X1 U16353 ( .A1(n16850), .A2(n12894), .ZN(n12895) );
  INV_X1 U16354 ( .A(n12896), .ZN(n12897) );
  INV_X1 U16355 ( .A(n13120), .ZN(n16834) );
  NAND2_X1 U16356 ( .A1(n16834), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12898) );
  OAI211_X1 U16357 ( .C1(n19730), .C2(n17330), .A(n12899), .B(n12898), .ZN(
        n12900) );
  AOI21_X1 U16358 ( .B1(n12923), .B2(n16984), .A(n12900), .ZN(n12915) );
  OAI21_X1 U16359 ( .B1(n12901), .B2(n16901), .A(n13053), .ZN(n12902) );
  INV_X1 U16360 ( .A(n16570), .ZN(n12904) );
  INV_X1 U16361 ( .A(n16559), .ZN(n12905) );
  INV_X1 U16362 ( .A(n12906), .ZN(n12907) );
  NAND2_X1 U16363 ( .A1(n12909), .A2(n12908), .ZN(n16539) );
  INV_X1 U16364 ( .A(n16513), .ZN(n12911) );
  INV_X1 U16365 ( .A(n12914), .ZN(n20537) );
  NOR2_X1 U16366 ( .A1(n12917), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12918) );
  OR2_X1 U16367 ( .A1(n12916), .A2(n12918), .ZN(n19733) );
  NOR2_X1 U16368 ( .A1(n19733), .A2(n16717), .ZN(n12919) );
  AOI211_X1 U16369 ( .C1(n16714), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12920), .B(n12919), .ZN(n12921) );
  OAI21_X1 U16370 ( .B1(n19730), .B2(n16682), .A(n12921), .ZN(n12922) );
  AOI21_X1 U16371 ( .B1(n12923), .B2(n16704), .A(n12922), .ZN(n12926) );
  NAND2_X1 U16372 ( .A1(n12924), .A2(n16713), .ZN(n12925) );
  NAND2_X1 U16373 ( .A1(n12926), .A2(n12925), .ZN(P2_U2994) );
  INV_X1 U16374 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16375 ( .A1(n12928), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12929) );
  OAI21_X1 U16376 ( .B1(n12930), .B2(n13101), .A(n12929), .ZN(n12931) );
  INV_X1 U16377 ( .A(n13162), .ZN(n12936) );
  NAND3_X1 U16378 ( .A1(n12660), .A2(n13330), .A3(n17055), .ZN(n13030) );
  NAND2_X1 U16379 ( .A1(n20547), .A2(n20356), .ZN(n13102) );
  NOR2_X1 U16380 ( .A1(n13038), .A2(n13102), .ZN(n12935) );
  NAND2_X1 U16381 ( .A1(n12936), .A2(n19761), .ZN(n13049) );
  INV_X1 U16382 ( .A(n12937), .ZN(n12938) );
  NAND2_X1 U16383 ( .A1(n12938), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12939) );
  MUX2_X2 U16384 ( .A(n13072), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n19753) );
  MUX2_X1 U16385 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16990) );
  INV_X1 U16386 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12942) );
  MUX2_X1 U16387 ( .A(n12942), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15936) );
  NOR2_X1 U16388 ( .A1(n16990), .A2(n15936), .ZN(n15924) );
  INV_X1 U16389 ( .A(n12940), .ZN(n12944) );
  INV_X1 U16390 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U16391 ( .A1(n12942), .A2(n12941), .ZN(n12943) );
  NAND2_X1 U16392 ( .A1(n12944), .A2(n12943), .ZN(n15926) );
  AND2_X1 U16393 ( .A1(n15924), .A2(n15926), .ZN(n15910) );
  OAI21_X1 U16394 ( .B1(n12940), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12946), .ZN(n16716) );
  NAND2_X1 U16395 ( .A1(n15910), .A2(n16716), .ZN(n15895) );
  AND2_X1 U16396 ( .A1(n12946), .A2(n16699), .ZN(n12947) );
  NOR2_X1 U16397 ( .A1(n12945), .A2(n12947), .ZN(n16696) );
  OR2_X1 U16398 ( .A1(n12945), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12948) );
  NAND2_X1 U16399 ( .A1(n12950), .A2(n12948), .ZN(n16684) );
  NAND2_X1 U16400 ( .A1(n15882), .A2(n16684), .ZN(n19752) );
  NAND2_X1 U16401 ( .A1(n12950), .A2(n16669), .ZN(n12951) );
  AND2_X1 U16402 ( .A1(n12949), .A2(n12951), .ZN(n19755) );
  OR2_X2 U16403 ( .A1(n19752), .A2(n19755), .ZN(n19756) );
  AND2_X1 U16404 ( .A1(n12949), .A2(n16660), .ZN(n12953) );
  NOR2_X1 U16405 ( .A1(n12952), .A2(n12953), .ZN(n16662) );
  OR2_X1 U16406 ( .A1(n19756), .A2(n16662), .ZN(n15858) );
  NOR2_X1 U16407 ( .A1(n12952), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12955) );
  OR2_X1 U16408 ( .A1(n12954), .A2(n12955), .ZN(n16648) );
  INV_X1 U16409 ( .A(n16648), .ZN(n15860) );
  OR2_X1 U16410 ( .A1(n12954), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12957) );
  NAND2_X1 U16411 ( .A1(n12956), .A2(n12957), .ZN(n16634) );
  NAND2_X1 U16412 ( .A1(n15841), .A2(n16634), .ZN(n15827) );
  NAND2_X1 U16413 ( .A1(n12956), .A2(n16619), .ZN(n12958) );
  AND2_X1 U16414 ( .A1(n9670), .A2(n12958), .ZN(n16621) );
  OR2_X1 U16415 ( .A1(n15827), .A2(n16621), .ZN(n13268) );
  NAND2_X1 U16416 ( .A1(n9670), .A2(n16602), .ZN(n12959) );
  AND2_X1 U16417 ( .A1(n12961), .A2(n12959), .ZN(n16606) );
  AND2_X1 U16418 ( .A1(n12961), .A2(n12960), .ZN(n12963) );
  OR2_X1 U16419 ( .A1(n12963), .A2(n12962), .ZN(n16592) );
  AND2_X1 U16420 ( .A1(n15817), .A2(n16592), .ZN(n15804) );
  OR2_X1 U16421 ( .A1(n12962), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12965) );
  NAND2_X1 U16422 ( .A1(n12964), .A2(n12965), .ZN(n16582) );
  NAND2_X1 U16423 ( .A1(n15804), .A2(n16582), .ZN(n15798) );
  NAND2_X1 U16424 ( .A1(n12964), .A2(n16573), .ZN(n12966) );
  AND2_X1 U16425 ( .A1(n12967), .A2(n12966), .ZN(n16575) );
  OR2_X1 U16426 ( .A1(n15798), .A2(n16575), .ZN(n15786) );
  AND2_X1 U16427 ( .A1(n12967), .A2(n16562), .ZN(n12969) );
  NOR2_X1 U16428 ( .A1(n12968), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12970) );
  OR2_X1 U16429 ( .A1(n12971), .A2(n12970), .ZN(n16552) );
  AND2_X1 U16430 ( .A1(n15771), .A2(n16552), .ZN(n15759) );
  OR2_X1 U16431 ( .A1(n12971), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12972) );
  NAND2_X1 U16432 ( .A1(n9726), .A2(n12972), .ZN(n16543) );
  NAND2_X1 U16433 ( .A1(n15759), .A2(n16543), .ZN(n15743) );
  INV_X1 U16434 ( .A(n12973), .ZN(n12975) );
  NAND2_X1 U16435 ( .A1(n9726), .A2(n16532), .ZN(n12974) );
  AND2_X1 U16436 ( .A1(n12975), .A2(n12974), .ZN(n16534) );
  AND2_X1 U16437 ( .A1(n12975), .A2(n15733), .ZN(n12976) );
  OR2_X1 U16438 ( .A1(n12976), .A2(n12917), .ZN(n16520) );
  NAND2_X1 U16439 ( .A1(n15709), .A2(n19753), .ZN(n12979) );
  OR2_X1 U16440 ( .A1(n12916), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12978) );
  NAND2_X1 U16441 ( .A1(n12977), .A2(n12978), .ZN(n16510) );
  NAND2_X1 U16442 ( .A1(n12979), .A2(n16510), .ZN(n15694) );
  NAND2_X1 U16443 ( .A1(n15694), .A2(n19753), .ZN(n12982) );
  NAND2_X1 U16444 ( .A1(n12977), .A2(n12980), .ZN(n12981) );
  NAND2_X1 U16445 ( .A1(n12983), .A2(n12981), .ZN(n16498) );
  NAND2_X1 U16446 ( .A1(n15678), .A2(n19753), .ZN(n12985) );
  NAND2_X1 U16447 ( .A1(n12983), .A2(n15677), .ZN(n12984) );
  NAND2_X1 U16448 ( .A1(n12986), .A2(n12984), .ZN(n16486) );
  NAND2_X1 U16449 ( .A1(n12985), .A2(n16486), .ZN(n15666) );
  NAND2_X1 U16450 ( .A1(n15666), .A2(n19753), .ZN(n12988) );
  AND2_X1 U16451 ( .A1(n12986), .A2(n15663), .ZN(n12987) );
  OR2_X1 U16452 ( .A1(n12987), .A2(n12989), .ZN(n16480) );
  NAND2_X1 U16453 ( .A1(n15645), .A2(n19753), .ZN(n12991) );
  OR2_X1 U16454 ( .A1(n12989), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12990) );
  NAND2_X1 U16455 ( .A1(n12993), .A2(n12990), .ZN(n15646) );
  NAND2_X1 U16456 ( .A1(n12991), .A2(n15646), .ZN(n15635) );
  NAND2_X1 U16457 ( .A1(n15635), .A2(n19753), .ZN(n12995) );
  NAND2_X1 U16458 ( .A1(n12993), .A2(n12992), .ZN(n12994) );
  NAND2_X1 U16459 ( .A1(n9751), .A2(n12994), .ZN(n16465) );
  NAND2_X1 U16460 ( .A1(n15620), .A2(n19753), .ZN(n12999) );
  AND2_X1 U16461 ( .A1(n9751), .A2(n12996), .ZN(n12998) );
  OR2_X1 U16462 ( .A1(n12998), .A2(n12997), .ZN(n16454) );
  NAND2_X1 U16463 ( .A1(n12999), .A2(n16454), .ZN(n15610) );
  NAND2_X1 U16464 ( .A1(n15610), .A2(n19753), .ZN(n13002) );
  NOR2_X1 U16465 ( .A1(n12997), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13001) );
  OR2_X1 U16466 ( .A1(n13000), .A2(n13001), .ZN(n16445) );
  NAND2_X1 U16467 ( .A1(n15595), .A2(n19753), .ZN(n13004) );
  OR2_X1 U16468 ( .A1(n13000), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13003) );
  NAND2_X1 U16469 ( .A1(n12937), .A2(n13003), .ZN(n16435) );
  INV_X1 U16470 ( .A(n13005), .ZN(n13007) );
  NAND2_X1 U16471 ( .A1(n19753), .A2(n19757), .ZN(n15965) );
  NAND2_X1 U16472 ( .A1(n15912), .A2(n13092), .ZN(n13111) );
  NOR2_X1 U16473 ( .A1(n13091), .A2(n13111), .ZN(n13047) );
  NAND2_X1 U16474 ( .A1(n13027), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U16475 ( .A1(n12697), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13009) );
  INV_X1 U16476 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20466) );
  AOI22_X1 U16477 ( .A1(n12848), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13012) );
  OAI21_X1 U16478 ( .B1(n12733), .B2(n20466), .A(n13012), .ZN(n15692) );
  NAND2_X1 U16479 ( .A1(n13027), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16480 ( .A1(n12848), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U16481 ( .A1(n13015), .A2(n9755), .ZN(n15658) );
  NAND2_X1 U16482 ( .A1(n13027), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16483 ( .A1(n12848), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13016) );
  NOR2_X2 U16484 ( .A1(n15658), .A2(n15659), .ZN(n13144) );
  AOI22_X1 U16485 ( .A1(n12848), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13018) );
  OAI21_X1 U16486 ( .B1(n12733), .B2(n20471), .A(n13018), .ZN(n13145) );
  NAND2_X1 U16487 ( .A1(n13027), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16488 ( .A1(n12848), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13019) );
  AND2_X1 U16489 ( .A1(n13020), .A2(n13019), .ZN(n15632) );
  NAND2_X1 U16490 ( .A1(n13027), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16491 ( .A1(n12848), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13021) );
  INV_X1 U16492 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U16493 ( .A1(n12848), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13026), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13023) );
  OAI21_X1 U16494 ( .B1(n12733), .B2(n16444), .A(n13023), .ZN(n15603) );
  INV_X1 U16495 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13518) );
  INV_X1 U16496 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20479) );
  OAI222_X1 U16497 ( .A1(n13518), .A2(n13025), .B1(n20479), .B2(n12733), .C1(
        n13024), .C2(n16727), .ZN(n15591) );
  AOI222_X1 U16498 ( .A1(n13027), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n12848), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n13026), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13096) );
  AOI222_X1 U16499 ( .A1(n13027), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12848), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n13026), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13028) );
  INV_X1 U16500 ( .A(n13030), .ZN(n13031) );
  AND2_X2 U16501 ( .A1(n13031), .A2(n20557), .ZN(n19835) );
  INV_X1 U16502 ( .A(n13102), .ZN(n13032) );
  NAND2_X1 U16503 ( .A1(n20560), .A2(n13032), .ZN(n14386) );
  INV_X1 U16504 ( .A(n14386), .ZN(n13033) );
  NAND2_X1 U16505 ( .A1(n13102), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13037) );
  NOR2_X1 U16506 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NAND2_X1 U16507 ( .A1(n13040), .A2(n20262), .ZN(n14389) );
  NAND2_X1 U16508 ( .A1(n19734), .A2(n14389), .ZN(n13041) );
  INV_X1 U16509 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20483) );
  NAND2_X1 U16510 ( .A1(n15951), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13043) );
  NAND3_X1 U16511 ( .A1(n19835), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n14386), 
        .ZN(n13042) );
  OAI211_X1 U16512 ( .C1(n19748), .C2(n20483), .A(n13043), .B(n13042), .ZN(
        n13044) );
  NAND2_X1 U16513 ( .A1(n13049), .A2(n13048), .ZN(P2_U2824) );
  NAND2_X1 U16514 ( .A1(n16579), .A2(n16984), .ZN(n13071) );
  NAND2_X1 U16515 ( .A1(n13051), .A2(n16597), .ZN(n16591) );
  NAND2_X1 U16516 ( .A1(n16591), .A2(n16590), .ZN(n16589) );
  NAND2_X1 U16517 ( .A1(n16589), .A2(n13052), .ZN(n13056) );
  NAND2_X1 U16518 ( .A1(n13054), .A2(n13053), .ZN(n13055) );
  XNOR2_X1 U16519 ( .A(n13056), .B(n13055), .ZN(n16587) );
  INV_X1 U16520 ( .A(n16899), .ZN(n16886) );
  OAI21_X1 U16521 ( .B1(n16886), .B2(n13065), .A(n16902), .ZN(n16889) );
  NAND2_X1 U16522 ( .A1(n13057), .A2(n14080), .ZN(n14082) );
  INV_X1 U16523 ( .A(n13058), .ZN(n13059) );
  AOI21_X1 U16524 ( .B1(n13060), .B2(n14082), .A(n13059), .ZN(n16584) );
  INV_X1 U16525 ( .A(n16584), .ZN(n15816) );
  NAND2_X1 U16526 ( .A1(n19745), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16581) );
  AOI21_X1 U16527 ( .B1(n13063), .B2(n13061), .A(n13062), .ZN(n15813) );
  NAND2_X1 U16528 ( .A1(n15813), .A2(n17327), .ZN(n13064) );
  OAI211_X1 U16529 ( .C1(n15816), .C2(n17330), .A(n16581), .B(n13064), .ZN(
        n13067) );
  NOR3_X1 U16530 ( .A1(n16886), .A2(n13065), .A3(n16901), .ZN(n13066) );
  AOI211_X1 U16531 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16889), .A(
        n13067), .B(n13066), .ZN(n13068) );
  NAND2_X1 U16532 ( .A1(n13071), .A2(n13070), .ZN(P2_U3033) );
  NOR2_X1 U16533 ( .A1(n17339), .A2(n20483), .ZN(n13164) );
  AOI21_X1 U16534 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13164), .ZN(n13074) );
  NAND2_X1 U16535 ( .A1(n13072), .A2(n16697), .ZN(n13073) );
  OAI211_X1 U16536 ( .C1(n13162), .C2(n16682), .A(n13074), .B(n13073), .ZN(
        n13075) );
  INV_X1 U16537 ( .A(n13075), .ZN(n13090) );
  NAND2_X1 U16538 ( .A1(n13076), .A2(n16690), .ZN(n13077) );
  INV_X1 U16539 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13081) );
  INV_X1 U16540 ( .A(n13085), .ZN(n13087) );
  NOR2_X1 U16541 ( .A1(n13087), .A2(n13086), .ZN(n13089) );
  INV_X1 U16542 ( .A(n13091), .ZN(n13112) );
  AOI21_X1 U16543 ( .B1(n13112), .B2(n19757), .A(n15952), .ZN(n13093) );
  OR2_X1 U16544 ( .A1(n13093), .A2(n13092), .ZN(n13116) );
  INV_X1 U16545 ( .A(n13094), .ZN(n13098) );
  INV_X1 U16546 ( .A(n13127), .ZN(n16321) );
  NAND2_X1 U16547 ( .A1(n16321), .A2(n19760), .ZN(n13099) );
  INV_X1 U16548 ( .A(n13100), .ZN(n13305) );
  AND2_X1 U16549 ( .A1(n13102), .A2(n13101), .ZN(n13103) );
  NAND2_X1 U16550 ( .A1(n13305), .A2(n13103), .ZN(n13105) );
  NAND2_X1 U16551 ( .A1(n19835), .A2(n14386), .ZN(n13104) );
  AOI22_X1 U16552 ( .A1(n19737), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19746), .ZN(n13106) );
  OAI21_X1 U16553 ( .B1(n13107), .B2(n19767), .A(n13106), .ZN(n13108) );
  AOI21_X1 U16554 ( .B1(n13109), .B2(n19750), .A(n13108), .ZN(n13110) );
  NAND2_X1 U16555 ( .A1(n13116), .A2(n13115), .ZN(P2_U2825) );
  NAND2_X1 U16556 ( .A1(n13118), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13117) );
  INV_X1 U16557 ( .A(n16769), .ZN(n16782) );
  INV_X1 U16558 ( .A(n16753), .ZN(n16450) );
  NAND2_X1 U16559 ( .A1(n16724), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16734) );
  NOR2_X1 U16560 ( .A1(n16734), .A2(n13123), .ZN(n13166) );
  INV_X1 U16561 ( .A(n13118), .ZN(n16810) );
  AOI21_X1 U16562 ( .B1(n16850), .B2(n16810), .A(n16809), .ZN(n13119) );
  NAND2_X1 U16563 ( .A1(n16850), .A2(n16753), .ZN(n13122) );
  OAI21_X1 U16564 ( .B1(n13123), .B2(n16745), .A(n16850), .ZN(n13124) );
  NAND3_X1 U16565 ( .A1(n16746), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13124), .ZN(n13167) );
  OAI21_X1 U16566 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13166), .A(
        n13167), .ZN(n13125) );
  OAI211_X1 U16567 ( .C1(n13127), .C2(n17340), .A(n13126), .B(n13125), .ZN(
        n13129) );
  NOR2_X1 U16568 ( .A1(n16211), .A2(n17330), .ZN(n13128) );
  NOR2_X1 U16569 ( .A1(n13129), .A2(n13128), .ZN(n13135) );
  INV_X1 U16570 ( .A(n13137), .ZN(n13139) );
  OAI21_X1 U16571 ( .B1(n13136), .B2(n13139), .A(n13138), .ZN(n13140) );
  NAND2_X1 U16572 ( .A1(n13140), .A2(n16473), .ZN(n16461) );
  INV_X1 U16573 ( .A(n16460), .ZN(n16438) );
  NAND2_X1 U16574 ( .A1(n16438), .A2(n16459), .ZN(n13141) );
  XNOR2_X1 U16575 ( .A(n16461), .B(n13141), .ZN(n13159) );
  AOI21_X1 U16576 ( .B1(n13143), .B2(n13142), .A(n9617), .ZN(n16244) );
  XNOR2_X1 U16577 ( .A(n13144), .B(n13145), .ZN(n16358) );
  NOR2_X1 U16578 ( .A1(n16358), .A2(n17340), .ZN(n13149) );
  NOR2_X1 U16579 ( .A1(n17339), .A2(n20471), .ZN(n13155) );
  AOI21_X1 U16580 ( .B1(n16757), .B2(n13147), .A(n13155), .ZN(n13146) );
  OAI21_X1 U16581 ( .B1(n16759), .B2(n13147), .A(n13146), .ZN(n13148) );
  AOI211_X1 U16582 ( .C1(n16244), .C2(n17346), .A(n13149), .B(n13148), .ZN(
        n13150) );
  OAI21_X1 U16583 ( .B1(n16458), .B2(n13153), .A(n13152), .ZN(P2_U3021) );
  AOI21_X1 U16584 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n13155), .ZN(n13156) );
  OAI21_X1 U16585 ( .B1(n15646), .B2(n16717), .A(n13156), .ZN(n13157) );
  AOI21_X1 U16586 ( .B1(n16244), .B2(n16719), .A(n13157), .ZN(n13158) );
  INV_X1 U16587 ( .A(n13160), .ZN(n13161) );
  NOR2_X1 U16588 ( .A1(n13162), .A2(n17330), .ZN(n13171) );
  NOR2_X1 U16589 ( .A1(n13163), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13165) );
  AOI21_X1 U16590 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(n13169) );
  NAND3_X1 U16591 ( .A1(n13167), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16800), .ZN(n13168) );
  OAI211_X1 U16592 ( .C1(n14552), .C2(n17340), .A(n13169), .B(n13168), .ZN(
        n13170) );
  NOR2_X1 U16593 ( .A1(n13171), .A2(n13170), .ZN(n13174) );
  NAND2_X1 U16594 ( .A1(n13172), .A2(n17351), .ZN(n13173) );
  OAI211_X1 U16595 ( .C1(n13175), .C2(n17348), .A(n13174), .B(n13173), .ZN(
        P2_U3015) );
  OAI21_X1 U16596 ( .B1(n17309), .B2(n13176), .A(n13591), .ZN(n13177) );
  INV_X1 U16597 ( .A(n13177), .ZN(n13178) );
  NOR2_X1 U16598 ( .A1(n21581), .A2(n17309), .ZN(n13180) );
  NAND2_X1 U16599 ( .A1(n13310), .A2(n13180), .ZN(n13570) );
  NAND4_X1 U16600 ( .A1(n13181), .A2(n13684), .A3(n14545), .A4(n20839), .ZN(
        n13460) );
  OR2_X1 U16601 ( .A1(n13460), .A2(n13182), .ZN(n13183) );
  NAND2_X1 U16602 ( .A1(n14566), .A2(n14997), .ZN(n13207) );
  NOR4_X1 U16603 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13193) );
  NOR4_X1 U16604 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13192) );
  NOR4_X1 U16605 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13191) );
  NOR4_X1 U16606 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13190) );
  AND4_X1 U16607 ( .A1(n13193), .A2(n13192), .A3(n13191), .A4(n13190), .ZN(
        n13198) );
  NOR4_X1 U16608 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13196) );
  NOR4_X1 U16609 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13195) );
  NOR4_X1 U16610 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13194) );
  NOR2_X1 U16611 ( .A1(n14545), .A2(n20834), .ZN(n13200) );
  INV_X1 U16612 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14027) );
  NOR2_X1 U16613 ( .A1(n20796), .A2(n14027), .ZN(n13201) );
  AOI21_X1 U16614 ( .B1(DATAI_14_), .B2(n20796), .A(n13201), .ZN(n20711) );
  OAI22_X1 U16615 ( .A1(n15003), .A2(n20711), .B1(n15036), .B2(n13202), .ZN(
        n13203) );
  AOI21_X1 U16616 ( .B1(n15005), .B2(DATAI_30_), .A(n13203), .ZN(n13204) );
  INV_X1 U16617 ( .A(n13204), .ZN(n13205) );
  NOR2_X1 U16618 ( .A1(n13205), .A2(n10560), .ZN(n13206) );
  NAND2_X1 U16619 ( .A1(n13207), .A2(n13206), .ZN(P1_U2874) );
  AOI21_X1 U16620 ( .B1(n13209), .B2(n14510), .A(n14527), .ZN(n14894) );
  NAND2_X1 U16621 ( .A1(n14894), .A2(n20756), .ZN(n13216) );
  INV_X1 U16622 ( .A(n13210), .ZN(n13214) );
  INV_X1 U16623 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14578) );
  NOR2_X1 U16624 ( .A1(n20786), .A2(n14578), .ZN(n15039) );
  INV_X1 U16625 ( .A(n13211), .ZN(n15308) );
  NOR3_X1 U16626 ( .A1(n15308), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13212), .ZN(n13213) );
  AOI211_X1 U16627 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n13214), .A(
        n15039), .B(n13213), .ZN(n13215) );
  NOR2_X1 U16628 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13219) );
  NOR4_X1 U16629 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13218) );
  NAND4_X1 U16630 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13219), .A4(n13218), .ZN(n13232) );
  NOR2_X4 U16631 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13232), .ZN(n17425)
         );
  NOR3_X1 U16632 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21578), .ZN(n13221) );
  NOR4_X1 U16633 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13220) );
  NAND4_X1 U16634 ( .A1(n20798), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13221), .A4(
        n13220), .ZN(U214) );
  NOR4_X1 U16635 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13225) );
  NOR4_X1 U16636 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n13224) );
  NOR4_X1 U16637 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13223) );
  NOR4_X1 U16638 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13222) );
  AND4_X1 U16639 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13230) );
  NOR4_X1 U16640 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n13228) );
  NOR4_X1 U16641 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n13227) );
  NOR4_X1 U16642 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U16643 ( .A1(n16844), .A2(n13235), .ZN(n13234) );
  NAND2_X1 U16644 ( .A1(n13236), .A2(n13484), .ZN(n13233) );
  NAND3_X1 U16645 ( .A1(n13234), .A2(n13233), .A3(n13478), .ZN(n13239) );
  AND2_X1 U16646 ( .A1(n13236), .A2(n13235), .ZN(n13238) );
  MUX2_X1 U16647 ( .A(n13239), .B(n13238), .S(n13237), .Z(n13257) );
  NOR2_X1 U16648 ( .A1(n13240), .A2(n17330), .ZN(n13256) );
  OR2_X1 U16649 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  NAND2_X1 U16650 ( .A1(n13244), .A2(n13243), .ZN(n20510) );
  INV_X1 U16651 ( .A(n20510), .ZN(n13248) );
  INV_X1 U16652 ( .A(n13245), .ZN(n13765) );
  AOI211_X1 U16653 ( .C1(n13767), .C2(n13766), .A(n13765), .B(n16988), .ZN(
        n13246) );
  INV_X1 U16654 ( .A(n13246), .ZN(n13247) );
  OR2_X1 U16655 ( .A1(n17339), .A2(n20431), .ZN(n13763) );
  OAI211_X1 U16656 ( .C1(n17340), .C2(n13248), .A(n13247), .B(n13763), .ZN(
        n13255) );
  OAI21_X1 U16657 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13764) );
  INV_X1 U16658 ( .A(n13252), .ZN(n13253) );
  OAI21_X1 U16659 ( .B1(n13764), .B2(n17348), .A(n13253), .ZN(n13254) );
  AOI211_X1 U16660 ( .C1(n18599), .C2(n13259), .A(n13258), .B(n19566), .ZN(
        n13266) );
  AOI211_X1 U16661 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17568), .A(n17557), .B(
        n17805), .ZN(n13265) );
  OAI22_X1 U16662 ( .A1(n10298), .A2(n17801), .B1(n17768), .B2(n10320), .ZN(
        n13264) );
  NAND2_X1 U16663 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17572) );
  NOR2_X1 U16664 ( .A1(n17572), .A2(n17585), .ZN(n13262) );
  OR2_X1 U16665 ( .A1(n17592), .A2(n13260), .ZN(n17562) );
  INV_X1 U16666 ( .A(n17562), .ZN(n13261) );
  MUX2_X1 U16667 ( .A(n13262), .B(n13261), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n13263) );
  INV_X1 U16668 ( .A(n15817), .ZN(n13267) );
  NAND2_X1 U16669 ( .A1(n15912), .A2(n13267), .ZN(n15818) );
  AOI21_X1 U16670 ( .B1(n16606), .B2(n13268), .A(n15818), .ZN(n13285) );
  AND2_X1 U16671 ( .A1(n13552), .A2(n13269), .ZN(n13272) );
  OAI21_X1 U16672 ( .B1(n13272), .B2(n13271), .A(n13758), .ZN(n16911) );
  OAI21_X1 U16673 ( .B1(n15955), .B2(n13273), .A(n17339), .ZN(n13274) );
  AOI21_X1 U16674 ( .B1(n19737), .B2(P2_REIP_REG_11__SCAN_IN), .A(n13274), 
        .ZN(n13275) );
  OAI21_X1 U16675 ( .B1(n16911), .B2(n15954), .A(n13275), .ZN(n13284) );
  INV_X1 U16676 ( .A(n13276), .ZN(n13277) );
  OAI22_X1 U16677 ( .A1(n13277), .A2(n15941), .B1(n16602), .B2(n19767), .ZN(
        n13283) );
  INV_X1 U16678 ( .A(n16606), .ZN(n13281) );
  NOR2_X1 U16679 ( .A1(n13278), .A2(n13279), .ZN(n13280) );
  OR2_X1 U16680 ( .A1(n13057), .A2(n13280), .ZN(n16603) );
  OAI22_X1 U16681 ( .A1(n10546), .A2(n13281), .B1(n16603), .B2(n15945), .ZN(
        n13282) );
  MUX2_X1 U16682 ( .A(n16850), .B(n13286), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13296) );
  AND2_X1 U16683 ( .A1(n13288), .A2(n13287), .ZN(n13290) );
  OR2_X1 U16684 ( .A1(n13290), .A2(n13289), .ZN(n13678) );
  OAI21_X1 U16685 ( .B1(n13292), .B2(n13291), .A(n12705), .ZN(n15953) );
  OAI22_X1 U16686 ( .A1(n17348), .A2(n13678), .B1(n17340), .B2(n15953), .ZN(
        n13295) );
  OAI21_X1 U16687 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15957), .A(
        n13358), .ZN(n13673) );
  OR2_X1 U16688 ( .A1(n17330), .A2(n13425), .ZN(n13293) );
  OR2_X1 U16689 ( .A1(n17339), .A2(n19722), .ZN(n13672) );
  OAI211_X1 U16690 ( .C1(n16988), .C2(n13673), .A(n13293), .B(n13672), .ZN(
        n13294) );
  OR3_X1 U16691 ( .A1(n13296), .A2(n13295), .A3(n13294), .ZN(P2_U3046) );
  MUX2_X1 U16692 ( .A(n20547), .B(P2_STATEBS16_REG_SCAN_IN), .S(n20559), .Z(
        n13297) );
  AND2_X1 U16693 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20522) );
  INV_X1 U16694 ( .A(n17356), .ZN(n17316) );
  NAND2_X1 U16695 ( .A1(n16992), .A2(n20552), .ZN(n14387) );
  OAI211_X1 U16696 ( .C1(n13297), .C2(P2_STATE2_REG_2__SCAN_IN), .A(n17316), 
        .B(n14387), .ZN(n13298) );
  INV_X1 U16697 ( .A(n13298), .ZN(P2_U3178) );
  NOR2_X1 U16698 ( .A1(n20543), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13300) );
  AOI211_X1 U16699 ( .C1(n15959), .C2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n13300), 
        .B(n13305), .ZN(n13299) );
  INV_X1 U16700 ( .A(n13299), .ZN(P2_U2814) );
  INV_X1 U16701 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19703) );
  NAND2_X1 U16702 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20552), .ZN(n17052) );
  OAI22_X1 U16703 ( .A1(n20545), .A2(n19703), .B1(n17052), .B2(n20493), .ZN(
        P2_U2816) );
  INV_X1 U16704 ( .A(n20545), .ZN(n13302) );
  OAI21_X1 U16705 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13300), .A(n13302), 
        .ZN(n13301) );
  OAI21_X1 U16706 ( .B1(n13303), .B2(n13302), .A(n13301), .ZN(P2_U3612) );
  NAND2_X1 U16707 ( .A1(n13310), .A2(n13463), .ZN(n14225) );
  AND2_X1 U16708 ( .A1(n9585), .A2(n21500), .ZN(n14713) );
  AOI21_X1 U16709 ( .B1(n14225), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14713), 
        .ZN(n13304) );
  NAND2_X1 U16710 ( .A1(n14226), .A2(n13304), .ZN(P1_U2801) );
  NAND2_X1 U16711 ( .A1(n13305), .A2(n20547), .ZN(n13306) );
  INV_X1 U16712 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13309) );
  INV_X1 U16713 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13798) );
  OR2_X1 U16714 ( .A1(n14325), .A2(n13798), .ZN(n13308) );
  NAND2_X1 U16715 ( .A1(n14325), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13307) );
  AND2_X1 U16716 ( .A1(n13308), .A2(n13307), .ZN(n14052) );
  INV_X1 U16717 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19800) );
  OAI222_X1 U16718 ( .A1(n19834), .A2(n13309), .B1(n13343), .B2(n14052), .C1(
        n13488), .C2(n19800), .ZN(P2_U2982) );
  AOI21_X1 U16719 ( .B1(n14530), .B2(n15582), .A(n17309), .ZN(n13563) );
  INV_X1 U16720 ( .A(n17305), .ZN(n13312) );
  INV_X1 U16721 ( .A(n13428), .ZN(n13311) );
  OAI22_X1 U16722 ( .A1(n13312), .A2(n9837), .B1(n13311), .B2(n13310), .ZN(
        n20569) );
  AOI211_X1 U16723 ( .C1(n9837), .C2(n21590), .A(n13563), .B(n20569), .ZN(
        n17292) );
  NOR2_X1 U16724 ( .A1(n17292), .A2(n20568), .ZN(n20576) );
  INV_X1 U16725 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13323) );
  NAND3_X1 U16726 ( .A1(n13314), .A2(n13313), .A3(n13591), .ZN(n13315) );
  MUX2_X1 U16727 ( .A(n13565), .B(n13315), .S(n17305), .Z(n13319) );
  NOR2_X1 U16728 ( .A1(n13317), .A2(n13316), .ZN(n13318) );
  OR2_X1 U16729 ( .A1(n13319), .A2(n13318), .ZN(n13320) );
  NAND2_X1 U16730 ( .A1(n13320), .A2(n11551), .ZN(n17294) );
  INV_X1 U16731 ( .A(n17294), .ZN(n13321) );
  NAND2_X1 U16732 ( .A1(n20576), .A2(n13321), .ZN(n13322) );
  OAI21_X1 U16733 ( .B1(n20576), .B2(n13323), .A(n13322), .ZN(P1_U3484) );
  INV_X1 U16734 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17393) );
  OR2_X1 U16735 ( .A1(n14325), .A2(n17393), .ZN(n13325) );
  NAND2_X1 U16736 ( .A1(n14325), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U16737 ( .A1(n13325), .A2(n13324), .ZN(n16363) );
  INV_X1 U16738 ( .A(n16363), .ZN(n13326) );
  NOR2_X1 U16739 ( .A1(n13343), .A2(n13326), .ZN(n19832) );
  INV_X1 U16740 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n13509) );
  INV_X1 U16741 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13510) );
  OAI22_X1 U16742 ( .A1(n19834), .A2(n13509), .B1(n13510), .B2(n13488), .ZN(
        n13327) );
  OR2_X1 U16743 ( .A1(n19832), .A2(n13327), .ZN(P2_U2960) );
  INV_X1 U16744 ( .A(n14366), .ZN(n13328) );
  OR2_X1 U16745 ( .A1(n13329), .A2(n13328), .ZN(n13333) );
  AND2_X1 U16746 ( .A1(n13524), .A2(n20547), .ZN(n14365) );
  NAND3_X1 U16747 ( .A1(n12680), .A2(n13330), .A3(n14365), .ZN(n13331) );
  OAI211_X1 U16748 ( .C1(n13490), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        n13335) );
  INV_X1 U16749 ( .A(n14103), .ZN(n14371) );
  MUX2_X1 U16750 ( .A(n14371), .B(n14372), .S(n14370), .Z(n13334) );
  OR2_X1 U16751 ( .A1(n14377), .A2(n19706), .ZN(n13337) );
  AOI22_X1 U16752 ( .A1(n17356), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n20559), .ZN(n13336) );
  NAND2_X1 U16753 ( .A1(n13337), .A2(n13336), .ZN(n17002) );
  INV_X1 U16754 ( .A(n13338), .ZN(n13339) );
  AND2_X1 U16755 ( .A1(n10130), .A2(n13339), .ZN(n13340) );
  NAND2_X1 U16756 ( .A1(n12864), .A2(n13340), .ZN(n14367) );
  OR3_X1 U16757 ( .A1(n17010), .A2(n14367), .A3(n20493), .ZN(n13341) );
  OAI21_X1 U16758 ( .B1(n13342), .B2(n17002), .A(n13341), .ZN(P2_U3595) );
  INV_X1 U16759 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19812) );
  INV_X1 U16760 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17391) );
  OR2_X1 U16761 ( .A1(n14325), .A2(n17391), .ZN(n13345) );
  NAND2_X1 U16762 ( .A1(n14325), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13344) );
  NAND2_X1 U16763 ( .A1(n13345), .A2(n13344), .ZN(n16355) );
  NAND2_X1 U16764 ( .A1(n19830), .A2(n16355), .ZN(n13400) );
  NAND2_X1 U16765 ( .A1(n19836), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13346) );
  OAI211_X1 U16766 ( .C1(n19812), .C2(n13488), .A(n13400), .B(n13346), .ZN(
        P2_U2976) );
  INV_X1 U16767 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19806) );
  INV_X1 U16768 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n21639) );
  OR2_X1 U16769 ( .A1(n14325), .A2(n21639), .ZN(n13348) );
  NAND2_X1 U16770 ( .A1(n14325), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U16771 ( .A1(n13348), .A2(n13347), .ZN(n16331) );
  NAND2_X1 U16772 ( .A1(n19830), .A2(n16331), .ZN(n13351) );
  NAND2_X1 U16773 ( .A1(n19836), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13349) );
  OAI211_X1 U16774 ( .C1(n19806), .C2(n13488), .A(n13351), .B(n13349), .ZN(
        P2_U2979) );
  INV_X1 U16775 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U16776 ( .A1(n19836), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13350) );
  OAI211_X1 U16777 ( .C1(n13502), .C2(n13488), .A(n13351), .B(n13350), .ZN(
        P2_U2964) );
  INV_X1 U16778 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19810) );
  INV_X1 U16779 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17389) );
  OR2_X1 U16780 ( .A1(n14325), .A2(n17389), .ZN(n13353) );
  NAND2_X1 U16781 ( .A1(n14325), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U16782 ( .A1(n13353), .A2(n13352), .ZN(n16347) );
  NAND2_X1 U16783 ( .A1(n19830), .A2(n16347), .ZN(n13356) );
  NAND2_X1 U16784 ( .A1(n19836), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13354) );
  OAI211_X1 U16785 ( .C1(n19810), .C2(n13488), .A(n13356), .B(n13354), .ZN(
        P2_U2977) );
  INV_X1 U16786 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U16787 ( .A1(n19836), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13355) );
  OAI211_X1 U16788 ( .C1(n13497), .C2(n13488), .A(n13356), .B(n13355), .ZN(
        P2_U2962) );
  OAI21_X1 U16789 ( .B1(n15940), .B2(n13358), .A(n13357), .ZN(n13359) );
  INV_X1 U16790 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13479) );
  XOR2_X1 U16791 ( .A(n13359), .B(n13479), .Z(n13470) );
  NOR2_X1 U16792 ( .A1(n17339), .A2(n20429), .ZN(n13480) );
  OAI21_X1 U16793 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13361), .A(
        n13360), .ZN(n13477) );
  NOR2_X1 U16794 ( .A1(n16722), .A2(n13477), .ZN(n13362) );
  AOI211_X1 U16795 ( .C1(n16713), .C2(n13470), .A(n13480), .B(n13362), .ZN(
        n13364) );
  MUX2_X1 U16796 ( .A(n16717), .B(n16700), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13363) );
  OAI211_X1 U16797 ( .C1(n15946), .C2(n16682), .A(n13364), .B(n13363), .ZN(
        P2_U3013) );
  AOI22_X1 U16798 ( .A1(n19836), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n19835), .ZN(n13367) );
  INV_X1 U16799 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13783) );
  OR2_X1 U16800 ( .A1(n14325), .A2(n13783), .ZN(n13366) );
  NAND2_X1 U16801 ( .A1(n14325), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13365) );
  NAND2_X1 U16802 ( .A1(n13366), .A2(n13365), .ZN(n16370) );
  NAND2_X1 U16803 ( .A1(n19830), .A2(n16370), .ZN(n13388) );
  NAND2_X1 U16804 ( .A1(n13367), .A2(n13388), .ZN(P2_U2974) );
  AOI22_X1 U16805 ( .A1(n19836), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19835), .ZN(n13370) );
  INV_X1 U16806 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13794) );
  OR2_X1 U16807 ( .A1(n14325), .A2(n13794), .ZN(n13369) );
  NAND2_X1 U16808 ( .A1(n14325), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U16809 ( .A1(n13369), .A2(n13368), .ZN(n19866) );
  NAND2_X1 U16810 ( .A1(n19830), .A2(n19866), .ZN(n13406) );
  NAND2_X1 U16811 ( .A1(n13370), .A2(n13406), .ZN(P2_U2972) );
  AOI22_X1 U16812 ( .A1(n19836), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19835), .ZN(n13374) );
  INV_X1 U16813 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13774) );
  OR2_X1 U16814 ( .A1(n14325), .A2(n13774), .ZN(n13372) );
  NAND2_X1 U16815 ( .A1(n14325), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13371) );
  INV_X1 U16816 ( .A(n19863), .ZN(n13373) );
  NAND2_X1 U16817 ( .A1(n19830), .A2(n13373), .ZN(n13408) );
  NAND2_X1 U16818 ( .A1(n13374), .A2(n13408), .ZN(P2_U2971) );
  AOI22_X1 U16819 ( .A1(n19836), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19835), .ZN(n13377) );
  INV_X1 U16820 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17399) );
  OR2_X1 U16821 ( .A1(n14325), .A2(n17399), .ZN(n13376) );
  NAND2_X1 U16822 ( .A1(n14325), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13375) );
  AND2_X1 U16823 ( .A1(n13376), .A2(n13375), .ZN(n19859) );
  INV_X1 U16824 ( .A(n19859), .ZN(n16400) );
  NAND2_X1 U16825 ( .A1(n19830), .A2(n16400), .ZN(n13410) );
  NAND2_X1 U16826 ( .A1(n13377), .A2(n13410), .ZN(P2_U2970) );
  AOI22_X1 U16827 ( .A1(n19836), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19835), .ZN(n13380) );
  INV_X1 U16828 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13779) );
  OR2_X1 U16829 ( .A1(n14325), .A2(n13779), .ZN(n13379) );
  NAND2_X1 U16830 ( .A1(n14325), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U16831 ( .A1(n13379), .A2(n13378), .ZN(n16407) );
  NAND2_X1 U16832 ( .A1(n19830), .A2(n16407), .ZN(n13412) );
  NAND2_X1 U16833 ( .A1(n13380), .A2(n13412), .ZN(P2_U2969) );
  AOI22_X1 U16834 ( .A1(n19836), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n19835), .ZN(n13384) );
  INV_X1 U16835 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13709) );
  OR2_X1 U16836 ( .A1(n14325), .A2(n13709), .ZN(n13382) );
  NAND2_X1 U16837 ( .A1(n14325), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13381) );
  AND2_X1 U16838 ( .A1(n13382), .A2(n13381), .ZN(n19852) );
  INV_X1 U16839 ( .A(n19852), .ZN(n13383) );
  NAND2_X1 U16840 ( .A1(n19830), .A2(n13383), .ZN(n13402) );
  NAND2_X1 U16841 ( .A1(n13384), .A2(n13402), .ZN(P2_U2968) );
  AOI22_X1 U16842 ( .A1(n19836), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n19835), .ZN(n13387) );
  INV_X1 U16843 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13787) );
  OR2_X1 U16844 ( .A1(n14325), .A2(n13787), .ZN(n13386) );
  NAND2_X1 U16845 ( .A1(n14325), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13385) );
  NAND2_X1 U16846 ( .A1(n13386), .A2(n13385), .ZN(n16377) );
  NAND2_X1 U16847 ( .A1(n19830), .A2(n16377), .ZN(n13404) );
  NAND2_X1 U16848 ( .A1(n13387), .A2(n13404), .ZN(P2_U2973) );
  AOI22_X1 U16849 ( .A1(n19836), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19835), .ZN(n13389) );
  NAND2_X1 U16850 ( .A1(n13389), .A2(n13388), .ZN(P2_U2959) );
  AOI22_X1 U16851 ( .A1(n19836), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19835), .ZN(n13392) );
  INV_X1 U16852 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14936) );
  OR2_X1 U16853 ( .A1(n14325), .A2(n14936), .ZN(n13391) );
  NAND2_X1 U16854 ( .A1(n14325), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13390) );
  NAND2_X1 U16855 ( .A1(n13391), .A2(n13390), .ZN(n16326) );
  NAND2_X1 U16856 ( .A1(n19830), .A2(n16326), .ZN(n13393) );
  NAND2_X1 U16857 ( .A1(n13392), .A2(n13393), .ZN(P2_U2965) );
  AOI22_X1 U16858 ( .A1(n19836), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19835), .ZN(n13394) );
  NAND2_X1 U16859 ( .A1(n13394), .A2(n13393), .ZN(P2_U2980) );
  AOI22_X1 U16860 ( .A1(n19836), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19835), .ZN(n13397) );
  INV_X1 U16861 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14949) );
  OR2_X1 U16862 ( .A1(n14325), .A2(n14949), .ZN(n13396) );
  NAND2_X1 U16863 ( .A1(n14325), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U16864 ( .A1(n13396), .A2(n13395), .ZN(n16340) );
  NAND2_X1 U16865 ( .A1(n19830), .A2(n16340), .ZN(n13398) );
  NAND2_X1 U16866 ( .A1(n13397), .A2(n13398), .ZN(P2_U2963) );
  AOI22_X1 U16867 ( .A1(n19836), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19835), .ZN(n13399) );
  NAND2_X1 U16868 ( .A1(n13399), .A2(n13398), .ZN(P2_U2978) );
  AOI22_X1 U16869 ( .A1(n19836), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19835), .ZN(n13401) );
  NAND2_X1 U16870 ( .A1(n13401), .A2(n13400), .ZN(P2_U2961) );
  AOI22_X1 U16871 ( .A1(n19836), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19835), .ZN(n13403) );
  NAND2_X1 U16872 ( .A1(n13403), .A2(n13402), .ZN(P2_U2953) );
  AOI22_X1 U16873 ( .A1(n19836), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19835), .ZN(n13405) );
  NAND2_X1 U16874 ( .A1(n13405), .A2(n13404), .ZN(P2_U2958) );
  AOI22_X1 U16875 ( .A1(n19836), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19835), .ZN(n13407) );
  NAND2_X1 U16876 ( .A1(n13407), .A2(n13406), .ZN(P2_U2957) );
  AOI22_X1 U16877 ( .A1(n19836), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19835), .ZN(n13409) );
  NAND2_X1 U16878 ( .A1(n13409), .A2(n13408), .ZN(P2_U2956) );
  AOI22_X1 U16879 ( .A1(n19836), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19835), .ZN(n13411) );
  NAND2_X1 U16880 ( .A1(n13411), .A2(n13410), .ZN(P2_U2955) );
  AOI22_X1 U16881 ( .A1(n19836), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19835), .ZN(n13413) );
  NAND2_X1 U16882 ( .A1(n13413), .A2(n13412), .ZN(P2_U2954) );
  AOI22_X1 U16883 ( .A1(n19836), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19835), .ZN(n13416) );
  INV_X1 U16884 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13706) );
  OR2_X1 U16885 ( .A1(n14325), .A2(n13706), .ZN(n13415) );
  NAND2_X1 U16886 ( .A1(n14325), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U16887 ( .A1(n13415), .A2(n13414), .ZN(n17019) );
  NAND2_X1 U16888 ( .A1(n19830), .A2(n17019), .ZN(n13417) );
  NAND2_X1 U16889 ( .A1(n13416), .A2(n13417), .ZN(P2_U2967) );
  AOI22_X1 U16890 ( .A1(n19836), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19835), .ZN(n13418) );
  NAND2_X1 U16891 ( .A1(n13418), .A2(n13417), .ZN(P2_U2952) );
  NAND2_X1 U16892 ( .A1(n19875), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14039) );
  AOI21_X1 U16893 ( .B1(n20549), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16894 ( .B1(n14370), .B2(n14103), .A(n10932), .ZN(n13424) );
  MUX2_X1 U16895 ( .A(n13425), .B(n11249), .S(n16287), .Z(n13426) );
  OAI21_X1 U16896 ( .B1(n20526), .B2(n16301), .A(n13426), .ZN(P2_U2887) );
  NAND2_X1 U16897 ( .A1(n13682), .A2(n21580), .ZN(n13561) );
  NAND2_X1 U16898 ( .A1(n13777), .A2(n21580), .ZN(n13427) );
  NOR2_X1 U16899 ( .A1(n13428), .A2(n13427), .ZN(n17303) );
  INV_X1 U16900 ( .A(n17303), .ZN(n13429) );
  NAND2_X1 U16901 ( .A1(n13561), .A2(n13429), .ZN(n13430) );
  NAND2_X1 U16902 ( .A1(n13430), .A2(n13463), .ZN(n13431) );
  NAND2_X1 U16903 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17321) );
  NOR2_X4 U16904 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17321), .ZN(n20688) );
  INV_X2 U16905 ( .A(n20667), .ZN(n20691) );
  AOI22_X1 U16906 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16907 ( .B1(n13202), .B2(n20663), .A(n13433), .ZN(P1_U2906) );
  INV_X1 U16908 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16909 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U16910 ( .B1(n13435), .B2(n20663), .A(n13434), .ZN(P1_U2910) );
  AOI22_X1 U16911 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U16912 ( .B1(n15002), .B2(n20663), .A(n13436), .ZN(P1_U2919) );
  INV_X1 U16913 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U16914 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U16915 ( .B1(n13438), .B2(n20663), .A(n13437), .ZN(P1_U2918) );
  INV_X1 U16916 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U16917 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13439) );
  OAI21_X1 U16918 ( .B1(n13440), .B2(n20663), .A(n13439), .ZN(P1_U2917) );
  INV_X1 U16919 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U16920 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U16921 ( .B1(n14974), .B2(n20663), .A(n13441), .ZN(P1_U2913) );
  INV_X1 U16922 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U16923 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13442) );
  OAI21_X1 U16924 ( .B1(n13443), .B2(n20663), .A(n13442), .ZN(P1_U2916) );
  AOI22_X1 U16925 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13444) );
  OAI21_X1 U16926 ( .B1(n14984), .B2(n20663), .A(n13444), .ZN(P1_U2915) );
  INV_X1 U16927 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U16928 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13445) );
  OAI21_X1 U16929 ( .B1(n13446), .B2(n20663), .A(n13445), .ZN(P1_U2914) );
  INV_X1 U16930 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13448) );
  AOI22_X1 U16931 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13447) );
  OAI21_X1 U16932 ( .B1(n13448), .B2(n20663), .A(n13447), .ZN(P1_U2908) );
  INV_X1 U16933 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13450) );
  AOI22_X1 U16934 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U16935 ( .B1(n13450), .B2(n20663), .A(n13449), .ZN(P1_U2907) );
  INV_X1 U16936 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U16937 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13451) );
  OAI21_X1 U16938 ( .B1(n13452), .B2(n20663), .A(n13451), .ZN(P1_U2909) );
  NAND2_X1 U16939 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20531), .ZN(
        n20295) );
  NAND2_X1 U16940 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20521), .ZN(
        n20260) );
  NOR2_X1 U16941 ( .A1(n20543), .A2(n17013), .ZN(n19915) );
  AOI21_X1 U16942 ( .B1(n14015), .B2(n17004), .A(n19915), .ZN(n13453) );
  XNOR2_X1 U16943 ( .A(n16993), .B(n13743), .ZN(n13454) );
  NAND2_X1 U16944 ( .A1(n13455), .A2(n13454), .ZN(n13456) );
  MUX2_X1 U16945 ( .A(n15946), .B(n15939), .S(n16287), .Z(n13457) );
  OAI21_X1 U16946 ( .B1(n20517), .B2(n16301), .A(n13457), .ZN(P2_U2886) );
  OR2_X1 U16947 ( .A1(n14531), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13459) );
  NAND2_X1 U16948 ( .A1(n13459), .A2(n13458), .ZN(n14284) );
  NAND2_X1 U16949 ( .A1(n17305), .A2(n13565), .ZN(n13462) );
  NAND2_X1 U16950 ( .A1(n13462), .A2(n13461), .ZN(n13464) );
  OAI21_X1 U16951 ( .B1(n13467), .B2(n13466), .A(n13465), .ZN(n14288) );
  OAI222_X1 U16952 ( .A1(n14284), .A2(n14933), .B1(n11944), .B2(n20662), .C1(
        n14288), .C2(n14935), .ZN(P1_U2872) );
  INV_X1 U16953 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16954 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13468) );
  OAI21_X1 U16955 ( .B1(n13469), .B2(n20663), .A(n13468), .ZN(P1_U2920) );
  INV_X1 U16956 ( .A(n13470), .ZN(n13476) );
  OR2_X1 U16957 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NAND2_X1 U16958 ( .A1(n13474), .A2(n13473), .ZN(n20513) );
  INV_X1 U16959 ( .A(n20513), .ZN(n13475) );
  OAI22_X1 U16960 ( .A1(n13476), .A2(n16988), .B1(n13475), .B2(n17340), .ZN(
        n13483) );
  NOR2_X1 U16961 ( .A1(n15946), .A2(n17330), .ZN(n13482) );
  OAI22_X1 U16962 ( .A1(n13479), .A2(n13478), .B1(n17348), .B2(n13477), .ZN(
        n13481) );
  NOR4_X1 U16963 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        n13486) );
  OAI211_X1 U16964 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16850), .B(n13484), .ZN(n13485) );
  NAND2_X1 U16965 ( .A1(n13486), .A2(n13485), .ZN(P2_U3045) );
  INV_X1 U16966 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13495) );
  INV_X1 U16967 ( .A(n13487), .ZN(n13489) );
  OAI21_X1 U16968 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13491) );
  INV_X1 U16969 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13494) );
  INV_X1 U16970 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13493) );
  OAI222_X1 U16971 ( .A1(n13495), .A2(n19798), .B1(n13536), .B2(n13494), .C1(
        n13537), .C2(n13493), .ZN(P2_U2935) );
  INV_X1 U16972 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13498) );
  INV_X1 U16973 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13496) );
  OAI222_X1 U16974 ( .A1(n13498), .A2(n19798), .B1(n13536), .B2(n13497), .C1(
        n13537), .C2(n13496), .ZN(P2_U2925) );
  INV_X1 U16975 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13500) );
  INV_X1 U16976 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n21621) );
  INV_X1 U16977 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13499) );
  OAI222_X1 U16978 ( .A1(n13500), .A2(n19798), .B1(n13536), .B2(n21621), .C1(
        n13537), .C2(n13499), .ZN(P2_U2930) );
  INV_X1 U16979 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13503) );
  INV_X1 U16980 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13501) );
  OAI222_X1 U16981 ( .A1(n13503), .A2(n19798), .B1(n13536), .B2(n13502), .C1(
        n13537), .C2(n13501), .ZN(P2_U2923) );
  INV_X1 U16982 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n13505) );
  INV_X1 U16983 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n21715) );
  INV_X1 U16984 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n13504) );
  OAI222_X1 U16985 ( .A1(n13505), .A2(n19798), .B1(n13537), .B2(n21715), .C1(
        n13504), .C2(n19828), .ZN(P2_U2943) );
  INV_X1 U16986 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13508) );
  INV_X1 U16987 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13507) );
  INV_X1 U16988 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13506) );
  OAI222_X1 U16989 ( .A1(n13508), .A2(n19798), .B1(n13536), .B2(n13507), .C1(
        n13537), .C2(n13506), .ZN(P2_U2933) );
  INV_X1 U16990 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13511) );
  OAI222_X1 U16991 ( .A1(n13511), .A2(n19798), .B1(n13536), .B2(n13510), .C1(
        n13537), .C2(n13509), .ZN(P2_U2927) );
  INV_X1 U16992 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13514) );
  INV_X1 U16993 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13513) );
  INV_X1 U16994 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13512) );
  OAI222_X1 U16995 ( .A1(n13514), .A2(n19798), .B1(n13536), .B2(n13513), .C1(
        n13537), .C2(n13512), .ZN(P2_U2931) );
  INV_X1 U16996 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13516) );
  INV_X1 U16997 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14421) );
  INV_X1 U16998 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13515) );
  OAI222_X1 U16999 ( .A1(n13516), .A2(n19798), .B1(n13536), .B2(n14421), .C1(
        n13537), .C2(n13515), .ZN(P2_U2934) );
  INV_X1 U17000 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13519) );
  INV_X1 U17001 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n13517) );
  OAI222_X1 U17002 ( .A1(n13519), .A2(n19798), .B1(n13536), .B2(n13518), .C1(
        n13517), .C2(n13537), .ZN(P2_U2922) );
  INV_X1 U17003 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13520) );
  INV_X1 U17004 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n21728) );
  INV_X1 U17005 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n21636) );
  OAI222_X1 U17006 ( .A1(n13536), .A2(n13520), .B1(n19798), .B2(n21728), .C1(
        n13537), .C2(n21636), .ZN(P2_U2932) );
  INV_X1 U17007 ( .A(n15953), .ZN(n13528) );
  NAND2_X1 U17008 ( .A1(n20269), .A2(n13528), .ZN(n19788) );
  NAND2_X1 U17009 ( .A1(n14370), .A2(n14372), .ZN(n13522) );
  NAND2_X1 U17010 ( .A1(n13522), .A2(n13521), .ZN(n13523) );
  NAND3_X1 U17011 ( .A1(n20545), .A2(n20547), .A3(n13524), .ZN(n13525) );
  OAI211_X1 U17012 ( .C1(n20269), .C2(n13528), .A(n19788), .B(n19790), .ZN(
        n13535) );
  INV_X1 U17013 ( .A(n13530), .ZN(n13531) );
  OAI22_X1 U17014 ( .A1(n19770), .A2(n15953), .B1(n13532), .B2(n19768), .ZN(
        n13533) );
  AOI21_X1 U17015 ( .B1(n16421), .B2(n17019), .A(n13533), .ZN(n13534) );
  NAND2_X1 U17016 ( .A1(n13535), .A2(n13534), .ZN(P2_U2919) );
  INV_X1 U17017 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13539) );
  AOI22_X1 U17018 ( .A1(n19795), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n20548), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13538) );
  OAI21_X1 U17019 ( .B1(n19798), .B2(n13539), .A(n13538), .ZN(P2_U2928) );
  INV_X1 U17020 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U17021 ( .A1(n19795), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n20548), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13540) );
  OAI21_X1 U17022 ( .B1(n19798), .B2(n13541), .A(n13540), .ZN(P2_U2926) );
  INV_X1 U17023 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U17024 ( .A1(n19795), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n20548), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13542) );
  OAI21_X1 U17025 ( .B1(n19798), .B2(n13543), .A(n13542), .ZN(P2_U2924) );
  INV_X1 U17026 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U17027 ( .A1(n19795), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n20548), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13544) );
  OAI21_X1 U17028 ( .B1(n19798), .B2(n13545), .A(n13544), .ZN(P2_U2929) );
  INV_X1 U17029 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19816) );
  INV_X1 U17030 ( .A(n16377), .ZN(n19874) );
  XOR2_X1 U17031 ( .A(n13547), .B(n13546), .Z(n19759) );
  INV_X1 U17032 ( .A(n19759), .ZN(n13548) );
  OAI222_X1 U17033 ( .A1(n19768), .A2(n19816), .B1(n19874), .B2(n19794), .C1(
        n13548), .C2(n16424), .ZN(P2_U2913) );
  INV_X1 U17034 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19814) );
  INV_X1 U17035 ( .A(n16370), .ZN(n19878) );
  OAI21_X1 U17036 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n16957) );
  OAI222_X1 U17037 ( .A1(n19768), .A2(n19814), .B1(n19878), .B2(n19794), .C1(
        n16957), .C2(n16424), .ZN(P2_U2912) );
  INV_X1 U17038 ( .A(n13552), .ZN(n13640) );
  OR2_X1 U17039 ( .A1(n13549), .A2(n13556), .ZN(n13558) );
  NAND2_X1 U17040 ( .A1(n13558), .A2(n13553), .ZN(n13554) );
  NAND2_X1 U17041 ( .A1(n13640), .A2(n13554), .ZN(n15843) );
  AOI22_X1 U17042 ( .A1(n16421), .A2(n16355), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19785), .ZN(n13555) );
  OAI21_X1 U17043 ( .B1(n15843), .B2(n16424), .A(n13555), .ZN(P2_U2910) );
  NAND2_X1 U17044 ( .A1(n13549), .A2(n13556), .ZN(n13557) );
  AND2_X1 U17045 ( .A1(n13558), .A2(n13557), .ZN(n16946) );
  INV_X1 U17046 ( .A(n16946), .ZN(n13560) );
  AOI22_X1 U17047 ( .A1(n16421), .A2(n16363), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19785), .ZN(n13559) );
  OAI21_X1 U17048 ( .B1(n13560), .B2(n16424), .A(n13559), .ZN(P2_U2911) );
  NAND2_X1 U17049 ( .A1(n13561), .A2(n13580), .ZN(n13564) );
  INV_X1 U17050 ( .A(n13591), .ZN(n13562) );
  AOI21_X1 U17051 ( .B1(n13564), .B2(n13563), .A(n13562), .ZN(n13566) );
  INV_X1 U17052 ( .A(n13565), .ZN(n13592) );
  MUX2_X1 U17053 ( .A(n13566), .B(n13592), .S(n17305), .Z(n13572) );
  NOR2_X1 U17054 ( .A1(n14243), .A2(n20819), .ZN(n13567) );
  NOR2_X1 U17055 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  AND2_X1 U17056 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  INV_X1 U17057 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20575) );
  NOR2_X1 U17058 ( .A1(n21501), .A2(n17321), .ZN(n14067) );
  INV_X1 U17059 ( .A(n14067), .ZN(n17325) );
  OAI22_X1 U17060 ( .A1(n17284), .A2(n20568), .B1(n20575), .B2(n17325), .ZN(
        n13575) );
  INV_X1 U17061 ( .A(n13698), .ZN(n15578) );
  INV_X1 U17062 ( .A(n13581), .ZN(n14061) );
  OR2_X1 U17063 ( .A1(n13573), .A2(n10062), .ZN(n13574) );
  XNOR2_X1 U17064 ( .A(n13574), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20640) );
  NAND4_X1 U17065 ( .A1(n13575), .A2(n15570), .A3(n14061), .A4(n20640), .ZN(
        n13576) );
  OAI21_X1 U17066 ( .B1(n15578), .B2(n14063), .A(n13576), .ZN(P1_U3468) );
  INV_X1 U17067 ( .A(n13578), .ZN(n13579) );
  NAND4_X1 U17068 ( .A1(n13582), .A2(n13581), .A3(n13580), .A4(n13579), .ZN(
        n13584) );
  NOR2_X1 U17069 ( .A1(n13584), .A2(n13583), .ZN(n13688) );
  INV_X1 U17070 ( .A(n13688), .ZN(n15569) );
  NAND2_X1 U17071 ( .A1(n15563), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13585) );
  NAND2_X1 U17072 ( .A1(n13585), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13586) );
  NAND2_X1 U17073 ( .A1(n11633), .A2(n13586), .ZN(n13599) );
  NAND3_X1 U17074 ( .A1(n13688), .A2(n13684), .A3(n13599), .ZN(n13597) );
  NAND2_X1 U17075 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13587) );
  INV_X1 U17076 ( .A(n13587), .ZN(n13588) );
  MUX2_X1 U17077 ( .A(n13588), .B(n13587), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13589) );
  NAND2_X1 U17078 ( .A1(n13682), .A2(n13589), .ZN(n13596) );
  MUX2_X1 U17079 ( .A(n13590), .B(n14056), .S(n15563), .Z(n13593) );
  NAND2_X1 U17080 ( .A1(n13592), .A2(n13591), .ZN(n13686) );
  OAI21_X1 U17081 ( .B1(n13594), .B2(n13593), .A(n13686), .ZN(n13595) );
  NAND3_X1 U17082 ( .A1(n13597), .A2(n13596), .A3(n13595), .ZN(n13598) );
  AOI21_X1 U17083 ( .B1(n21118), .B2(n15569), .A(n13598), .ZN(n14055) );
  INV_X1 U17084 ( .A(n14055), .ZN(n13600) );
  AOI22_X1 U17085 ( .A1(n13600), .A2(n15570), .B1(n15575), .B2(n13599), .ZN(
        n13602) );
  NAND2_X1 U17086 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13698), .ZN(
        n13601) );
  OAI21_X1 U17087 ( .B1(n13602), .B2(n13698), .A(n13601), .ZN(P1_U3469) );
  NOR3_X1 U17088 ( .A1(n19681), .A2(n10216), .A3(n13614), .ZN(n13605) );
  INV_X1 U17089 ( .A(n13603), .ZN(n13604) );
  NAND2_X1 U17090 ( .A1(n13608), .A2(n13607), .ZN(n19081) );
  OAI21_X1 U17091 ( .B1(n18994), .B2(n9882), .A(n18943), .ZN(n13717) );
  INV_X1 U17092 ( .A(n13717), .ZN(n13611) );
  INV_X1 U17093 ( .A(n13609), .ZN(n13610) );
  INV_X1 U17094 ( .A(n13652), .ZN(n13659) );
  NAND2_X1 U17095 ( .A1(n13610), .A2(n13659), .ZN(n13612) );
  AND2_X1 U17096 ( .A1(n18994), .A2(n14199), .ZN(n17254) );
  OAI22_X1 U17097 ( .A1(n13611), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13612), .B2(n17254), .ZN(n19527) );
  INV_X1 U17098 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14470) );
  INV_X1 U17099 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19053) );
  OAI22_X1 U17100 ( .A1(n14470), .A2(n19053), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13662) );
  INV_X1 U17101 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18884) );
  NOR2_X1 U17102 ( .A1(n19559), .A2(n18884), .ZN(n13664) );
  INV_X1 U17103 ( .A(n13612), .ZN(n17799) );
  AOI222_X1 U17104 ( .A1(n19527), .A2(n19693), .B1(n13662), .B2(n13664), .C1(
        n19553), .C2(n17799), .ZN(n13638) );
  NAND2_X1 U17105 ( .A1(n19516), .A2(n19682), .ZN(n13622) );
  AOI221_X1 U17106 ( .B1(n19681), .B2(n17278), .C1(n10212), .C2(n17278), .A(
        n13622), .ZN(n14195) );
  OAI21_X1 U17107 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19528), .A(
        n13615), .ZN(n13616) );
  INV_X1 U17108 ( .A(n13616), .ZN(n13834) );
  AND2_X1 U17109 ( .A1(n13617), .A2(n13834), .ZN(n13619) );
  NAND2_X1 U17110 ( .A1(n13620), .A2(n19117), .ZN(n13658) );
  NAND2_X1 U17111 ( .A1(n19513), .A2(n14193), .ZN(n13621) );
  OAI21_X1 U17112 ( .B1(n13622), .B2(n18414), .A(n13621), .ZN(n13633) );
  INV_X1 U17113 ( .A(n13623), .ZN(n13628) );
  NOR3_X1 U17114 ( .A1(n13626), .A2(n13625), .A3(n13624), .ZN(n13979) );
  AND2_X1 U17115 ( .A1(n14199), .A2(n19117), .ZN(n13977) );
  INV_X1 U17116 ( .A(n13977), .ZN(n13627) );
  NAND3_X1 U17117 ( .A1(n13628), .A2(n13979), .A3(n13627), .ZN(n13630) );
  NAND2_X1 U17118 ( .A1(n13630), .A2(n13629), .ZN(n13632) );
  NAND2_X1 U17119 ( .A1(n13632), .A2(n13631), .ZN(n13844) );
  OR2_X1 U17120 ( .A1(n13633), .A2(n13844), .ZN(n13634) );
  OR2_X1 U17121 ( .A1(n14195), .A2(n13634), .ZN(n19535) );
  NAND2_X1 U17122 ( .A1(n19535), .A2(n19675), .ZN(n13636) );
  INV_X1 U17123 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17452) );
  NAND3_X1 U17124 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19659)
         );
  OR2_X1 U17125 ( .A1(n17452), .A2(n19659), .ZN(n17267) );
  NAND2_X1 U17126 ( .A1(n19657), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19093) );
  AND2_X1 U17127 ( .A1(n17267), .A2(n19093), .ZN(n13635) );
  NAND2_X1 U17128 ( .A1(n13720), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13637) );
  OAI21_X1 U17129 ( .B1(n13638), .B2(n13720), .A(n13637), .ZN(P3_U3289) );
  XNOR2_X1 U17130 ( .A(n13640), .B(n13639), .ZN(n16924) );
  AOI22_X1 U17131 ( .A1(n16421), .A2(n16347), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19785), .ZN(n13641) );
  OAI21_X1 U17132 ( .B1(n16924), .B2(n16424), .A(n13641), .ZN(P2_U2909) );
  OAI21_X1 U17133 ( .B1(n13643), .B2(n13642), .A(n13998), .ZN(n14255) );
  OAI21_X1 U17134 ( .B1(n13646), .B2(n13645), .A(n13644), .ZN(n14237) );
  AOI22_X1 U17135 ( .A1(n20658), .A2(n14237), .B1(n14927), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13647) );
  OAI21_X1 U17136 ( .B1(n14255), .B2(n14935), .A(n13647), .ZN(P1_U2871) );
  INV_X1 U17137 ( .A(n13648), .ZN(n13649) );
  NAND2_X1 U17138 ( .A1(n13650), .A2(n13649), .ZN(n19694) );
  NAND2_X1 U17139 ( .A1(n13651), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17766) );
  INV_X1 U17140 ( .A(n17766), .ZN(n13653) );
  NOR2_X1 U17141 ( .A1(n13652), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13715) );
  NOR2_X1 U17142 ( .A1(n13653), .A2(n13715), .ZN(n17784) );
  INV_X1 U17143 ( .A(n13654), .ZN(n13655) );
  NAND3_X1 U17144 ( .A1(n13717), .A2(n10612), .A3(n13655), .ZN(n13661) );
  OAI21_X1 U17145 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n13713) );
  NAND3_X1 U17146 ( .A1(n13713), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n13659), .ZN(n13660) );
  OAI211_X1 U17147 ( .C1(n19061), .C2(n17784), .A(n13661), .B(n13660), .ZN(
        n19536) );
  INV_X1 U17148 ( .A(n13662), .ZN(n13663) );
  AOI222_X1 U17149 ( .A1(n19536), .A2(n19693), .B1(n13664), .B2(n13663), .C1(
        n19553), .C2(n17784), .ZN(n13666) );
  NAND2_X1 U17150 ( .A1(n13720), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13665) );
  OAI21_X1 U17151 ( .B1(n13720), .B2(n13666), .A(n13665), .ZN(P3_U3288) );
  INV_X1 U17152 ( .A(n20930), .ZN(n14070) );
  OAI22_X1 U17153 ( .A1(n14070), .A2(n13688), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15567), .ZN(n17282) );
  OAI22_X1 U17154 ( .A1(n13696), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21500), .ZN(n13667) );
  AOI21_X1 U17155 ( .B1(n17282), .B2(n15570), .A(n13667), .ZN(n13670) );
  INV_X1 U17156 ( .A(n13682), .ZN(n13668) );
  NOR2_X1 U17157 ( .A1(n13668), .A2(n11578), .ZN(n17281) );
  AOI22_X1 U17158 ( .A1(n17281), .A2(n15570), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13698), .ZN(n13669) );
  OAI21_X1 U17159 ( .B1(n13670), .B2(n13698), .A(n13669), .ZN(P1_U3474) );
  INV_X1 U17160 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19808) );
  INV_X1 U17161 ( .A(n16340), .ZN(n13671) );
  OAI222_X1 U17162 ( .A1(n16911), .A2(n16424), .B1(n19768), .B2(n19808), .C1(
        n19794), .C2(n13671), .ZN(P2_U2908) );
  OAI21_X1 U17163 ( .B1(n16707), .B2(n13673), .A(n13672), .ZN(n13674) );
  AOI21_X1 U17164 ( .B1(n15962), .B2(n16719), .A(n13674), .ZN(n13677) );
  OAI21_X1 U17165 ( .B1(n16714), .B2(n13675), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13676) );
  OAI211_X1 U17166 ( .C1(n13678), .C2(n16722), .A(n13677), .B(n13676), .ZN(
        P2_U3014) );
  OR2_X1 U17167 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  OR2_X1 U17168 ( .A1(n21279), .A2(n13688), .ZN(n13692) );
  NAND2_X1 U17169 ( .A1(n13682), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13683) );
  NAND2_X1 U17170 ( .A1(n13682), .A2(n11569), .ZN(n15566) );
  MUX2_X1 U17171 ( .A(n13683), .B(n15566), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13690) );
  XNOR2_X1 U17172 ( .A(n15563), .B(n11673), .ZN(n13685) );
  AND2_X1 U17173 ( .A1(n13684), .A2(n13685), .ZN(n13687) );
  INV_X1 U17174 ( .A(n13685), .ZN(n13695) );
  AOI22_X1 U17175 ( .A1(n13688), .A2(n13687), .B1(n13686), .B2(n13695), .ZN(
        n13689) );
  AND2_X1 U17176 ( .A1(n13690), .A2(n13689), .ZN(n13691) );
  NAND2_X1 U17177 ( .A1(n13692), .A2(n13691), .ZN(n14053) );
  NOR2_X1 U17178 ( .A1(n21500), .A2(n13749), .ZN(n15573) );
  INV_X1 U17179 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14535) );
  OAI22_X1 U17180 ( .A1(n14535), .A2(n20793), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15572) );
  INV_X1 U17181 ( .A(n15572), .ZN(n13693) );
  NAND2_X1 U17182 ( .A1(n15573), .A2(n13693), .ZN(n13694) );
  OAI21_X1 U17183 ( .B1(n13696), .B2(n13695), .A(n13694), .ZN(n13697) );
  AOI21_X1 U17184 ( .B1(n14053), .B2(n15570), .A(n13697), .ZN(n13699) );
  MUX2_X1 U17185 ( .A(n13699), .B(n11673), .S(n13698), .Z(n13700) );
  INV_X1 U17186 ( .A(n13700), .ZN(P1_U3472) );
  NOR2_X1 U17187 ( .A1(n17800), .A2(n17774), .ZN(n13704) );
  NAND2_X1 U17188 ( .A1(n17260), .A2(n19695), .ZN(n17783) );
  INV_X1 U17189 ( .A(n19693), .ZN(n17256) );
  NAND3_X1 U17190 ( .A1(n17812), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A3(
        n17256), .ZN(n13701) );
  OAI21_X1 U17191 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17783), .A(
        n13701), .ZN(n13702) );
  AOI21_X1 U17192 ( .B1(n17594), .B2(P3_REIP_REG_0__SCAN_IN), .A(n13702), .ZN(
        n13703) );
  OAI21_X1 U17193 ( .B1(n13704), .B2(n9868), .A(n13703), .ZN(P3_U2671) );
  OR2_X1 U17194 ( .A1(n20796), .A2(n13706), .ZN(n13708) );
  NAND2_X1 U17195 ( .A1(n20796), .A2(DATAI_0_), .ZN(n13707) );
  NAND2_X1 U17196 ( .A1(n13708), .A2(n13707), .ZN(n15010) );
  INV_X1 U17197 ( .A(n15010), .ZN(n20807) );
  INV_X1 U17198 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20696) );
  OAI222_X1 U17199 ( .A1(n15038), .A2(n14288), .B1(n15037), .B2(n20807), .C1(
        n15036), .C2(n20696), .ZN(P1_U2904) );
  OR2_X1 U17200 ( .A1(n20796), .A2(n13709), .ZN(n13711) );
  NAND2_X1 U17201 ( .A1(n20796), .A2(DATAI_1_), .ZN(n13710) );
  NAND2_X1 U17202 ( .A1(n13711), .A2(n13710), .ZN(n13803) );
  INV_X1 U17203 ( .A(n13803), .ZN(n20816) );
  INV_X1 U17204 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20693) );
  OAI222_X1 U17205 ( .A1(n15038), .A2(n14255), .B1(n15037), .B2(n20816), .C1(
        n13186), .C2(n20693), .ZN(P1_U2903) );
  NOR2_X1 U17206 ( .A1(n18943), .A2(n13651), .ZN(n13712) );
  AOI211_X1 U17207 ( .C1(n13713), .C2(n17766), .A(n13715), .B(n13712), .ZN(
        n19522) );
  NOR2_X1 U17208 ( .A1(n19522), .A2(n17256), .ZN(n13714) );
  AOI211_X1 U17209 ( .C1(n19553), .C2(n17766), .A(n13714), .B(n13720), .ZN(
        n13721) );
  INV_X1 U17210 ( .A(n13715), .ZN(n13716) );
  AOI22_X1 U17211 ( .A1(n13717), .A2(n13651), .B1(n9887), .B2(n13716), .ZN(
        n19523) );
  NOR3_X1 U17212 ( .A1(n19523), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n17256), .ZN(n13718) );
  AOI21_X1 U17213 ( .B1(n19553), .B2(n9601), .A(n13718), .ZN(n13719) );
  OAI22_X1 U17214 ( .A1(n13721), .A2(n19524), .B1(n13720), .B2(n13719), .ZN(
        P3_U3285) );
  AND3_X1 U17215 ( .A1(n13723), .A2(n13722), .A3(n13749), .ZN(n13724) );
  OAI21_X1 U17216 ( .B1(n9587), .B2(n13725), .A(n13724), .ZN(n13726) );
  NAND2_X1 U17217 ( .A1(n13727), .A2(n13726), .ZN(n13756) );
  INV_X1 U17218 ( .A(n13756), .ZN(n13733) );
  INV_X1 U17219 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13728) );
  NOR2_X1 U17220 ( .A1(n20786), .A2(n13728), .ZN(n13752) );
  INV_X1 U17221 ( .A(n13729), .ZN(n13731) );
  INV_X1 U17222 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13730) );
  AOI21_X1 U17223 ( .B1(n15169), .B2(n13731), .A(n13730), .ZN(n13732) );
  AOI211_X1 U17224 ( .C1(n13733), .C2(n20738), .A(n13752), .B(n13732), .ZN(
        n13734) );
  OAI21_X1 U17225 ( .B1(n20797), .B2(n14288), .A(n13734), .ZN(P1_U2999) );
  INV_X1 U17226 ( .A(n13735), .ZN(n14011) );
  NAND2_X1 U17227 ( .A1(n14333), .A2(n14011), .ZN(n13739) );
  NAND2_X1 U17228 ( .A1(n20199), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14013) );
  INV_X1 U17229 ( .A(n20199), .ZN(n19944) );
  NAND2_X1 U17230 ( .A1(n19944), .A2(n20512), .ZN(n13736) );
  NAND2_X1 U17231 ( .A1(n14013), .A2(n13736), .ZN(n17014) );
  NOR2_X1 U17232 ( .A1(n17014), .A2(n20543), .ZN(n13737) );
  AOI21_X1 U17233 ( .B1(n14015), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13737), .ZN(n13738) );
  NAND2_X1 U17234 ( .A1(n13739), .A2(n13738), .ZN(n13742) );
  NAND2_X1 U17235 ( .A1(n13742), .A2(n13741), .ZN(n14007) );
  OR2_X1 U17236 ( .A1(n16993), .A2(n13743), .ZN(n13744) );
  XNOR2_X2 U17237 ( .A(n14009), .B(n13746), .ZN(n20508) );
  MUX2_X1 U17238 ( .A(n14333), .B(P2_EBX_REG_2__SCAN_IN), .S(n16287), .Z(
        n13747) );
  AOI21_X1 U17239 ( .B1(n20508), .B2(n16311), .A(n13747), .ZN(n13748) );
  INV_X1 U17240 ( .A(n13748), .ZN(P2_U2885) );
  INV_X1 U17241 ( .A(n15372), .ZN(n15396) );
  AOI21_X1 U17242 ( .B1(n20770), .B2(n13749), .A(n15460), .ZN(n20792) );
  INV_X1 U17243 ( .A(n20792), .ZN(n13751) );
  NAND3_X1 U17244 ( .A1(n20744), .A2(n13749), .A3(n15366), .ZN(n13750) );
  OAI21_X1 U17245 ( .B1(n15396), .B2(n13751), .A(n13750), .ZN(n13755) );
  INV_X1 U17246 ( .A(n14284), .ZN(n13753) );
  AOI21_X1 U17247 ( .B1(n20756), .B2(n13753), .A(n13752), .ZN(n13754) );
  OAI211_X1 U17248 ( .C1(n20784), .C2(n13756), .A(n13755), .B(n13754), .ZN(
        P1_U3031) );
  INV_X1 U17249 ( .A(n13061), .ZN(n13757) );
  AOI21_X1 U17250 ( .B1(n13759), .B2(n13758), .A(n13757), .ZN(n16895) );
  INV_X1 U17251 ( .A(n16895), .ZN(n13761) );
  AOI22_X1 U17252 ( .A1(n16421), .A2(n16331), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19785), .ZN(n13760) );
  OAI21_X1 U17253 ( .B1(n13761), .B2(n16424), .A(n13760), .ZN(P2_U2907) );
  INV_X1 U17254 ( .A(n15926), .ZN(n13770) );
  NAND2_X1 U17255 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13762) );
  OAI211_X1 U17256 ( .C1(n13764), .C2(n16722), .A(n13763), .B(n13762), .ZN(
        n13769) );
  AOI211_X1 U17257 ( .C1(n13767), .C2(n13766), .A(n16707), .B(n13765), .ZN(
        n13768) );
  AOI211_X1 U17258 ( .C1(n13770), .C2(n16697), .A(n13769), .B(n13768), .ZN(
        n13771) );
  OAI21_X1 U17259 ( .B1(n13240), .B2(n16682), .A(n13771), .ZN(P2_U3012) );
  OR2_X1 U17260 ( .A1(n20796), .A2(n13774), .ZN(n13776) );
  NAND2_X1 U17261 ( .A1(n20796), .A2(DATAI_4_), .ZN(n13775) );
  NAND2_X1 U17262 ( .A1(n13776), .A2(n13775), .ZN(n14988) );
  NAND2_X1 U17263 ( .A1(n20713), .A2(n14988), .ZN(n13811) );
  AND2_X2 U17264 ( .A1(n13800), .A2(n13777), .ZN(n20723) );
  AOI22_X1 U17265 ( .A1(n20723), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U17266 ( .A1(n13811), .A2(n13778), .ZN(P1_U2956) );
  OR2_X1 U17267 ( .A1(n20796), .A2(n13779), .ZN(n13781) );
  NAND2_X1 U17268 ( .A1(n20796), .A2(DATAI_2_), .ZN(n13780) );
  NAND2_X1 U17269 ( .A1(n13781), .A2(n13780), .ZN(n14006) );
  NAND2_X1 U17270 ( .A1(n20713), .A2(n14006), .ZN(n13820) );
  AOI22_X1 U17271 ( .A1(n20723), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13782) );
  NAND2_X1 U17272 ( .A1(n13820), .A2(n13782), .ZN(P1_U2954) );
  OR2_X1 U17273 ( .A1(n20796), .A2(n13783), .ZN(n13785) );
  NAND2_X1 U17274 ( .A1(n20796), .A2(DATAI_7_), .ZN(n13784) );
  NAND2_X1 U17275 ( .A1(n13785), .A2(n13784), .ZN(n14973) );
  NAND2_X1 U17276 ( .A1(n20713), .A2(n14973), .ZN(n13809) );
  AOI22_X1 U17277 ( .A1(n20723), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13786) );
  NAND2_X1 U17278 ( .A1(n13809), .A2(n13786), .ZN(P1_U2959) );
  OR2_X1 U17279 ( .A1(n20796), .A2(n13787), .ZN(n13789) );
  NAND2_X1 U17280 ( .A1(n20796), .A2(DATAI_6_), .ZN(n13788) );
  NAND2_X1 U17281 ( .A1(n13789), .A2(n13788), .ZN(n14979) );
  NAND2_X1 U17282 ( .A1(n20713), .A2(n14979), .ZN(n13807) );
  AOI22_X1 U17283 ( .A1(n20723), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13790) );
  NAND2_X1 U17284 ( .A1(n13807), .A2(n13790), .ZN(P1_U2958) );
  OR2_X1 U17285 ( .A1(n20796), .A2(n17399), .ZN(n13792) );
  NAND2_X1 U17286 ( .A1(n20796), .A2(DATAI_3_), .ZN(n13791) );
  NAND2_X1 U17287 ( .A1(n13792), .A2(n13791), .ZN(n14048) );
  NAND2_X1 U17288 ( .A1(n20713), .A2(n14048), .ZN(n13818) );
  AOI22_X1 U17289 ( .A1(n20723), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U17290 ( .A1(n13818), .A2(n13793), .ZN(P1_U2955) );
  OR2_X1 U17291 ( .A1(n20796), .A2(n13794), .ZN(n13796) );
  NAND2_X1 U17292 ( .A1(n20796), .A2(DATAI_5_), .ZN(n13795) );
  NAND2_X1 U17293 ( .A1(n13796), .A2(n13795), .ZN(n14220) );
  NAND2_X1 U17294 ( .A1(n20713), .A2(n14220), .ZN(n13822) );
  AOI22_X1 U17295 ( .A1(n20723), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U17296 ( .A1(n13822), .A2(n13797), .ZN(P1_U2957) );
  INV_X1 U17297 ( .A(n20713), .ZN(n13802) );
  NOR2_X1 U17298 ( .A1(n20796), .A2(n13798), .ZN(n13799) );
  AOI21_X1 U17299 ( .B1(DATAI_15_), .B2(n20796), .A(n13799), .ZN(n15018) );
  INV_X1 U17300 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13801) );
  OAI222_X1 U17301 ( .A1(n13804), .A2(n20669), .B1(n13802), .B2(n15018), .C1(
        n13801), .C2(n13800), .ZN(P1_U2967) );
  NAND2_X1 U17302 ( .A1(n20713), .A2(n13803), .ZN(n13816) );
  AOI22_X1 U17303 ( .A1(n20723), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13805) );
  NAND2_X1 U17304 ( .A1(n13816), .A2(n13805), .ZN(P1_U2938) );
  AOI22_X1 U17305 ( .A1(n20723), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U17306 ( .A1(n13807), .A2(n13806), .ZN(P1_U2943) );
  AOI22_X1 U17307 ( .A1(n20723), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U17308 ( .A1(n13809), .A2(n13808), .ZN(P1_U2944) );
  AOI22_X1 U17309 ( .A1(n20723), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U17310 ( .A1(n13811), .A2(n13810), .ZN(P1_U2941) );
  NAND2_X1 U17311 ( .A1(n20713), .A2(n15010), .ZN(n13814) );
  AOI22_X1 U17312 ( .A1(n20723), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13812) );
  NAND2_X1 U17313 ( .A1(n13814), .A2(n13812), .ZN(P1_U2937) );
  AOI22_X1 U17314 ( .A1(n20723), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U17315 ( .A1(n13814), .A2(n13813), .ZN(P1_U2952) );
  AOI22_X1 U17316 ( .A1(n20723), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13815) );
  NAND2_X1 U17317 ( .A1(n13816), .A2(n13815), .ZN(P1_U2953) );
  AOI22_X1 U17318 ( .A1(n20723), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U17319 ( .A1(n13818), .A2(n13817), .ZN(P1_U2940) );
  AOI22_X1 U17320 ( .A1(n20723), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U17321 ( .A1(n13820), .A2(n13819), .ZN(P1_U2939) );
  AOI22_X1 U17322 ( .A1(n20723), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U17323 ( .A1(n13822), .A2(n13821), .ZN(P1_U2942) );
  NOR2_X1 U17324 ( .A1(n13823), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20785) );
  INV_X1 U17325 ( .A(n20785), .ZN(n13825) );
  NAND3_X1 U17326 ( .A1(n13825), .A2(n20738), .A3(n13824), .ZN(n13829) );
  AOI22_X1 U17327 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20731), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13826) );
  OAI21_X1 U17328 ( .B1(n20742), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13826), .ZN(n13827) );
  INV_X1 U17329 ( .A(n13827), .ZN(n13828) );
  OAI211_X1 U17330 ( .C1(n20797), .C2(n14255), .A(n13829), .B(n13828), .ZN(
        P1_U2998) );
  AND2_X1 U17331 ( .A1(n10214), .A2(n19102), .ZN(n13838) );
  AOI211_X1 U17332 ( .C1(n19681), .C2(n19106), .A(n13838), .B(n13830), .ZN(
        n13831) );
  NOR2_X1 U17333 ( .A1(n19677), .A2(n13831), .ZN(n17448) );
  NAND3_X1 U17334 ( .A1(n17448), .A2(n13832), .A3(n19516), .ZN(n13842) );
  OAI21_X1 U17335 ( .B1(n13833), .B2(n19117), .A(n19513), .ZN(n13841) );
  OR2_X1 U17336 ( .A1(n13835), .A2(n13834), .ZN(n13837) );
  NAND2_X1 U17337 ( .A1(n13837), .A2(n13836), .ZN(n19515) );
  NAND2_X1 U17338 ( .A1(n13838), .A2(n19127), .ZN(n13976) );
  INV_X1 U17339 ( .A(n13976), .ZN(n13839) );
  NAND2_X1 U17340 ( .A1(n19515), .A2(n13839), .ZN(n13840) );
  NAND3_X1 U17341 ( .A1(n13842), .A2(n13841), .A3(n13840), .ZN(n13843) );
  AOI22_X1 U17342 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17343 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13851) );
  INV_X1 U17344 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18015) );
  NAND2_X1 U17345 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13847) );
  NAND2_X1 U17346 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13846) );
  OAI211_X1 U17347 ( .C1(n9603), .C2(n18015), .A(n13847), .B(n13846), .ZN(
        n13848) );
  INV_X1 U17348 ( .A(n13848), .ZN(n13850) );
  INV_X1 U17349 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18014) );
  OR2_X1 U17350 ( .A1(n18227), .A2(n18014), .ZN(n13849) );
  NAND4_X1 U17351 ( .A1(n13852), .A2(n13851), .A3(n13850), .A4(n13849), .ZN(
        n13858) );
  AOI22_X1 U17352 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17353 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17354 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17355 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13853) );
  NAND4_X1 U17356 ( .A1(n13856), .A2(n13855), .A3(n13854), .A4(n13853), .ZN(
        n13857) );
  AOI22_X1 U17357 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13906), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13867) );
  INV_X1 U17358 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13862) );
  INV_X1 U17359 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13859) );
  OR2_X1 U17360 ( .A1(n18224), .A2(n13859), .ZN(n13861) );
  NAND2_X1 U17361 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13860) );
  OAI211_X1 U17362 ( .C1(n18227), .C2(n13862), .A(n13861), .B(n13860), .ZN(
        n13863) );
  INV_X1 U17363 ( .A(n13863), .ZN(n13866) );
  AOI22_X1 U17364 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14144), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13865) );
  NAND2_X1 U17365 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13864) );
  AOI22_X1 U17366 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17367 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17368 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U17369 ( .A1(n13869), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13870) );
  AND4_X1 U17370 ( .A1(n13873), .A2(n13872), .A3(n13871), .A4(n13870), .ZN(
        n13874) );
  NAND2_X2 U17371 ( .A1(n13875), .A2(n13874), .ZN(n14204) );
  INV_X1 U17372 ( .A(n14204), .ZN(n13905) );
  AOI22_X1 U17373 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17374 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17375 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17376 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13876) );
  NAND4_X1 U17377 ( .A1(n13879), .A2(n13878), .A3(n13877), .A4(n13876), .ZN(
        n13887) );
  AOI22_X1 U17378 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17379 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13884) );
  INV_X1 U17380 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17885) );
  INV_X1 U17381 ( .A(n13881), .ZN(n13883) );
  INV_X1 U17382 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17886) );
  OR2_X1 U17383 ( .A1(n18227), .A2(n17886), .ZN(n13882) );
  NAND4_X1 U17384 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13886) );
  AOI22_X1 U17385 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17386 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13895) );
  INV_X1 U17387 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13890) );
  NAND2_X1 U17388 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13889) );
  NAND2_X1 U17389 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13888) );
  OAI211_X1 U17390 ( .C1(n9603), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13891) );
  INV_X1 U17391 ( .A(n13891), .ZN(n13894) );
  INV_X1 U17392 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13892) );
  OR2_X1 U17393 ( .A1(n18227), .A2(n13892), .ZN(n13893) );
  NAND4_X1 U17394 ( .A1(n13896), .A2(n13895), .A3(n13894), .A4(n13893), .ZN(
        n13904) );
  AOI22_X1 U17395 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17396 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17397 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17398 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13899) );
  NAND4_X1 U17399 ( .A1(n13902), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13903) );
  NAND2_X1 U17400 ( .A1(n13905), .A2(n13939), .ZN(n13935) );
  AOI22_X1 U17401 ( .A1(n13906), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U17402 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13913) );
  INV_X1 U17403 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17899) );
  NAND2_X1 U17404 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13908) );
  NAND2_X1 U17405 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13907) );
  OAI211_X1 U17406 ( .C1(n9602), .C2(n17899), .A(n13908), .B(n13907), .ZN(
        n13909) );
  INV_X1 U17407 ( .A(n13909), .ZN(n13912) );
  INV_X1 U17408 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13910) );
  OR2_X1 U17409 ( .A1(n18227), .A2(n13910), .ZN(n13911) );
  NAND4_X1 U17410 ( .A1(n13914), .A2(n13913), .A3(n13912), .A4(n13911), .ZN(
        n13921) );
  AOI22_X1 U17411 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17412 ( .A1(n13915), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17413 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17414 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13916) );
  NAND4_X1 U17415 ( .A1(n13919), .A2(n13918), .A3(n13917), .A4(n13916), .ZN(
        n13920) );
  NAND2_X1 U17416 ( .A1(n13935), .A2(n13959), .ZN(n13945) );
  NOR2_X1 U17417 ( .A1(n18404), .A2(n13945), .ZN(n14169) );
  AOI22_X1 U17418 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17419 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13927) );
  INV_X1 U17420 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U17421 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13923) );
  NAND2_X1 U17422 ( .A1(n14144), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13922) );
  OAI211_X1 U17423 ( .C1(n9603), .C2(n17997), .A(n13923), .B(n13922), .ZN(
        n13924) );
  INV_X1 U17424 ( .A(n13924), .ZN(n13926) );
  INV_X1 U17425 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17996) );
  OR2_X1 U17426 ( .A1(n18227), .A2(n17996), .ZN(n13925) );
  NAND4_X1 U17427 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n13934) );
  AOI22_X1 U17428 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U17429 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U17430 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17431 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13929) );
  NAND4_X1 U17432 ( .A1(n13932), .A2(n13931), .A3(n13930), .A4(n13929), .ZN(
        n13933) );
  XOR2_X1 U17433 ( .A(n14169), .B(n14168), .Z(n14170) );
  XOR2_X1 U17434 ( .A(n21719), .B(n14170), .Z(n13947) );
  INV_X1 U17435 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21734) );
  OAI21_X1 U17436 ( .B1(n13935), .B2(n13959), .A(n13945), .ZN(n13944) );
  INV_X1 U17437 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19073) );
  INV_X1 U17438 ( .A(n13936), .ZN(n13938) );
  OAI21_X1 U17439 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13938), .A(
        n13937), .ZN(n18795) );
  INV_X1 U17440 ( .A(n14214), .ZN(n13984) );
  AOI21_X1 U17441 ( .B1(n13984), .B2(n18884), .A(n19053), .ZN(n13942) );
  INV_X1 U17442 ( .A(n13939), .ZN(n13940) );
  AOI21_X1 U17443 ( .B1(n18884), .B2(n19053), .A(n13940), .ZN(n13941) );
  OAI21_X1 U17444 ( .B1(n13942), .B2(n14198), .A(n13941), .ZN(n18796) );
  NOR2_X1 U17445 ( .A1(n18795), .A2(n18796), .ZN(n18794) );
  XOR2_X1 U17446 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13944), .Z(
        n18782) );
  XNOR2_X1 U17447 ( .A(n13945), .B(n18404), .ZN(n18773) );
  AOI21_X1 U17448 ( .B1(n13947), .B2(n13946), .A(n14171), .ZN(n18761) );
  INV_X1 U17449 ( .A(n18761), .ZN(n13983) );
  NAND2_X1 U17450 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19033) );
  INV_X1 U17451 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18774) );
  NOR3_X1 U17452 ( .A1(n21719), .A2(n21734), .A3(n18774), .ZN(n14166) );
  INV_X1 U17453 ( .A(n14166), .ZN(n13948) );
  NOR2_X1 U17454 ( .A1(n19033), .A2(n13948), .ZN(n14449) );
  AOI21_X1 U17455 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13952) );
  INV_X1 U17456 ( .A(n13952), .ZN(n19054) );
  NAND2_X1 U17457 ( .A1(n14166), .A2(n19054), .ZN(n14452) );
  NOR2_X1 U17458 ( .A1(n18994), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19064) );
  AOI21_X1 U17459 ( .B1(n9887), .B2(n14452), .A(n19064), .ZN(n13949) );
  OAI21_X1 U17460 ( .B1(n19062), .B2(n14449), .A(n13949), .ZN(n14182) );
  OAI21_X1 U17461 ( .B1(n19080), .B2(n14182), .A(n19075), .ZN(n13951) );
  INV_X1 U17462 ( .A(n13951), .ZN(n19023) );
  AOI21_X1 U17463 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18971), .A(
        n19081), .ZN(n19052) );
  OAI22_X1 U17464 ( .A1(n13952), .A2(n19061), .B1(n19033), .B2(n19052), .ZN(
        n19045) );
  NAND3_X1 U17465 ( .A1(n19070), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19045), .ZN(n19040) );
  NOR2_X1 U17466 ( .A1(n18774), .A2(n19040), .ZN(n19027) );
  AOI22_X1 U17467 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19023), .B1(
        n19027), .B2(n21719), .ZN(n13982) );
  XNOR2_X1 U17468 ( .A(n14198), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13986) );
  NAND2_X1 U17469 ( .A1(n13986), .A2(n17173), .ZN(n13985) );
  INV_X1 U17470 ( .A(n14198), .ZN(n13953) );
  NAND2_X1 U17471 ( .A1(n13953), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13954) );
  NAND2_X1 U17472 ( .A1(n13985), .A2(n13954), .ZN(n18798) );
  XNOR2_X1 U17473 ( .A(n13955), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18799) );
  NAND2_X1 U17474 ( .A1(n18798), .A2(n18799), .ZN(n18797) );
  INV_X1 U17475 ( .A(n13955), .ZN(n13956) );
  NAND2_X1 U17476 ( .A1(n13956), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13957) );
  NAND2_X1 U17477 ( .A1(n13958), .A2(n13959), .ZN(n13969) );
  INV_X1 U17478 ( .A(n13958), .ZN(n13960) );
  INV_X1 U17479 ( .A(n13959), .ZN(n18409) );
  NAND2_X1 U17480 ( .A1(n13960), .A2(n18409), .ZN(n13961) );
  NAND2_X1 U17481 ( .A1(n13969), .A2(n13961), .ZN(n13962) );
  XNOR2_X1 U17482 ( .A(n13964), .B(n13962), .ZN(n18784) );
  INV_X1 U17483 ( .A(n13962), .ZN(n13963) );
  NAND2_X1 U17484 ( .A1(n13964), .A2(n13963), .ZN(n13965) );
  XNOR2_X1 U17485 ( .A(n13969), .B(n18404), .ZN(n13966) );
  XNOR2_X1 U17486 ( .A(n13966), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18767) );
  INV_X1 U17487 ( .A(n13966), .ZN(n13967) );
  NAND2_X1 U17488 ( .A1(n13967), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13968) );
  INV_X1 U17489 ( .A(n13969), .ZN(n13971) );
  NAND2_X1 U17490 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  NAND2_X1 U17491 ( .A1(n13972), .A2(n18401), .ZN(n13973) );
  NAND2_X1 U17492 ( .A1(n14143), .A2(n13973), .ZN(n14121) );
  OAI21_X1 U17493 ( .B1(n13974), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n14125), .ZN(n13975) );
  INV_X1 U17494 ( .A(n13975), .ZN(n18759) );
  NOR2_X1 U17495 ( .A1(n13977), .A2(n13976), .ZN(n13978) );
  NAND2_X1 U17496 ( .A1(n13979), .A2(n13978), .ZN(n19514) );
  INV_X1 U17497 ( .A(n19514), .ZN(n17216) );
  INV_X1 U17498 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n13980) );
  NOR2_X1 U17499 ( .A1(n19075), .A2(n13980), .ZN(n18758) );
  AOI21_X1 U17500 ( .B1(n18759), .B2(n19074), .A(n18758), .ZN(n13981) );
  OAI211_X1 U17501 ( .C1(n19021), .C2(n13983), .A(n13982), .B(n13981), .ZN(
        P3_U2857) );
  NAND2_X1 U17502 ( .A1(n13984), .A2(n18884), .ZN(n17174) );
  XNOR2_X1 U17503 ( .A(n13986), .B(n17174), .ZN(n18811) );
  INV_X1 U17504 ( .A(n18811), .ZN(n13993) );
  OAI21_X1 U17505 ( .B1(n13986), .B2(n17173), .A(n13985), .ZN(n13987) );
  INV_X1 U17506 ( .A(n13987), .ZN(n18810) );
  INV_X1 U17507 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n13988) );
  NOR2_X1 U17508 ( .A1(n19075), .A2(n13988), .ZN(n18809) );
  AOI21_X1 U17509 ( .B1(n19074), .B2(n18810), .A(n18809), .ZN(n13992) );
  NAND2_X1 U17510 ( .A1(n18920), .A2(n19070), .ZN(n19035) );
  INV_X1 U17511 ( .A(n19035), .ZN(n14458) );
  OAI21_X1 U17512 ( .B1(n19081), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14458), .ZN(n13990) );
  NAND2_X1 U17513 ( .A1(n18994), .A2(n19061), .ZN(n18947) );
  NAND3_X1 U17514 ( .A1(n19070), .A2(n18884), .A3(n18947), .ZN(n19083) );
  AND2_X1 U17515 ( .A1(n19083), .A2(n19072), .ZN(n13989) );
  MUX2_X1 U17516 ( .A(n13990), .B(n13989), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13991) );
  OAI211_X1 U17517 ( .C1(n19021), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        P3_U2861) );
  INV_X1 U17518 ( .A(n15813), .ZN(n13995) );
  INV_X1 U17519 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19804) );
  INV_X1 U17520 ( .A(n16326), .ZN(n13994) );
  OAI222_X1 U17521 ( .A1(n13995), .A2(n16424), .B1(n19768), .B2(n19804), .C1(
        n19794), .C2(n13994), .ZN(P2_U2906) );
  INV_X1 U17522 ( .A(n13996), .ZN(n13997) );
  AOI21_X1 U17523 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n15295) );
  INV_X1 U17524 ( .A(n15295), .ZN(n14271) );
  NAND2_X1 U17525 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  NAND2_X1 U17526 ( .A1(n14000), .A2(n14003), .ZN(n20773) );
  INV_X1 U17527 ( .A(n20773), .ZN(n14004) );
  AOI22_X1 U17528 ( .A1(n20658), .A2(n14004), .B1(n14927), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14005) );
  OAI21_X1 U17529 ( .B1(n14271), .B2(n14935), .A(n14005), .ZN(P1_U2870) );
  INV_X1 U17530 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20690) );
  OAI222_X1 U17531 ( .A1(n15038), .A2(n14271), .B1(n15037), .B2(n20821), .C1(
        n13186), .C2(n20690), .ZN(P1_U2902) );
  INV_X1 U17532 ( .A(n14013), .ZN(n14012) );
  NAND2_X1 U17533 ( .A1(n14012), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20358) );
  NAND2_X1 U17534 ( .A1(n14013), .A2(n20505), .ZN(n14014) );
  AOI22_X1 U17535 ( .A1(n14015), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19846), .B2(n14014), .ZN(n14016) );
  NAND2_X1 U17536 ( .A1(n14018), .A2(n14019), .ZN(n14037) );
  MUX2_X1 U17537 ( .A(n11251), .B(n14022), .S(n16308), .Z(n14023) );
  OAI21_X1 U17538 ( .B1(n20169), .B2(n16301), .A(n14023), .ZN(P2_U2884) );
  OR2_X1 U17539 ( .A1(n13062), .A2(n14025), .ZN(n14026) );
  AND2_X1 U17540 ( .A1(n14024), .A2(n14026), .ZN(n16881) );
  INV_X1 U17541 ( .A(n16881), .ZN(n14031) );
  OR2_X1 U17542 ( .A1(n14325), .A2(n14027), .ZN(n14029) );
  NAND2_X1 U17543 ( .A1(n14325), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U17544 ( .A1(n14029), .A2(n14028), .ZN(n19829) );
  AOI22_X1 U17545 ( .A1(n16421), .A2(n19829), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19785), .ZN(n14030) );
  OAI21_X1 U17546 ( .B1(n14031), .B2(n16424), .A(n14030), .ZN(P2_U2905) );
  XOR2_X1 U17547 ( .A(n14032), .B(n14033), .Z(n15287) );
  INV_X1 U17548 ( .A(n15287), .ZN(n14264) );
  INV_X1 U17549 ( .A(n14189), .ZN(n14034) );
  AOI21_X1 U17550 ( .B1(n14000), .B2(n14035), .A(n14034), .ZN(n20755) );
  AOI22_X1 U17551 ( .A1(n20658), .A2(n20755), .B1(n14927), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14036) );
  OAI21_X1 U17552 ( .B1(n14264), .B2(n14935), .A(n14036), .ZN(P1_U2869) );
  OAI211_X1 U17553 ( .C1(n14039), .C2(n13342), .A(n14038), .B(n14037), .ZN(
        n14042) );
  INV_X1 U17554 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14040) );
  NOR2_X1 U17555 ( .A1(n9595), .A2(n14040), .ZN(n14041) );
  OR2_X1 U17556 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  NAND2_X1 U17557 ( .A1(n14042), .A2(n14041), .ZN(n14274) );
  NAND2_X1 U17558 ( .A1(n14043), .A2(n14274), .ZN(n19773) );
  NAND2_X1 U17559 ( .A1(n9646), .A2(n14044), .ZN(n14207) );
  OR2_X1 U17560 ( .A1(n9646), .A2(n14044), .ZN(n14045) );
  AND2_X1 U17561 ( .A1(n14207), .A2(n14045), .ZN(n16983) );
  INV_X1 U17562 ( .A(n16983), .ZN(n14046) );
  MUX2_X1 U17563 ( .A(n14046), .B(n15902), .S(n16287), .Z(n14047) );
  OAI21_X1 U17564 ( .B1(n19773), .B2(n16301), .A(n14047), .ZN(P2_U2883) );
  INV_X1 U17565 ( .A(n14048), .ZN(n20826) );
  INV_X1 U17566 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20687) );
  OAI222_X1 U17567 ( .A1(n15038), .A2(n14264), .B1(n15037), .B2(n20826), .C1(
        n13186), .C2(n20687), .ZN(P1_U2901) );
  NAND2_X1 U17568 ( .A1(n14024), .A2(n14050), .ZN(n14051) );
  NAND2_X1 U17569 ( .A1(n14049), .A2(n14051), .ZN(n16870) );
  OAI222_X1 U17570 ( .A1(n16870), .A2(n16424), .B1(n19768), .B2(n19800), .C1(
        n14052), .C2(n19794), .ZN(P2_U2904) );
  NOR2_X1 U17571 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21500), .ZN(n14065) );
  MUX2_X1 U17572 ( .A(n14053), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17284), .Z(n17289) );
  AOI22_X1 U17573 ( .A1(n14065), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17289), .B2(n21500), .ZN(n14059) );
  INV_X1 U17574 ( .A(n17284), .ZN(n14054) );
  MUX2_X1 U17575 ( .A(n14056), .B(n14055), .S(n14054), .Z(n17291) );
  INV_X1 U17576 ( .A(n17291), .ZN(n14057) );
  AOI22_X1 U17577 ( .A1(n14065), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21500), .B2(n14057), .ZN(n14058) );
  NOR2_X1 U17578 ( .A1(n14059), .A2(n14058), .ZN(n17298) );
  INV_X1 U17579 ( .A(n17298), .ZN(n14066) );
  AOI21_X1 U17580 ( .B1(n20640), .B2(n14061), .A(n17284), .ZN(n14062) );
  AOI211_X1 U17581 ( .C1(n17284), .C2(n14063), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n14062), .ZN(n14064) );
  AOI21_X1 U17582 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n14065), .A(
        n14064), .ZN(n17296) );
  OAI21_X1 U17583 ( .B1(n14066), .B2(n14060), .A(n17296), .ZN(n14069) );
  OAI21_X1 U17584 ( .B1(n14069), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14067), .ZN(
        n14068) );
  INV_X1 U17585 ( .A(n21587), .ZN(n14227) );
  NAND2_X1 U17586 ( .A1(n14068), .A2(n20975), .ZN(n20795) );
  NOR2_X1 U17587 ( .A1(n14069), .A2(n17321), .ZN(n17308) );
  AND2_X1 U17588 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21282), .ZN(n15558) );
  OAI22_X1 U17589 ( .A1(n14070), .A2(n15558), .B1(n9587), .B2(n21433), .ZN(
        n14071) );
  OAI21_X1 U17590 ( .B1(n17308), .B2(n14071), .A(n20795), .ZN(n14072) );
  OAI21_X1 U17591 ( .B1(n20795), .B2(n21327), .A(n14072), .ZN(P1_U3478) );
  INV_X1 U17592 ( .A(n16407), .ZN(n19855) );
  XNOR2_X1 U17593 ( .A(n20103), .B(n20510), .ZN(n14076) );
  NOR2_X1 U17594 ( .A1(n20494), .A2(n20513), .ZN(n14073) );
  AOI21_X1 U17595 ( .B1(n20494), .B2(n20513), .A(n14073), .ZN(n19789) );
  NAND2_X1 U17596 ( .A1(n19789), .A2(n19788), .ZN(n19787) );
  INV_X1 U17597 ( .A(n14073), .ZN(n14074) );
  NAND2_X1 U17598 ( .A1(n19787), .A2(n14074), .ZN(n14075) );
  NAND2_X1 U17599 ( .A1(n14076), .A2(n14075), .ZN(n16418) );
  OAI21_X1 U17600 ( .B1(n14076), .B2(n14075), .A(n16418), .ZN(n14077) );
  NAND2_X1 U17601 ( .A1(n14077), .A2(n19790), .ZN(n14079) );
  AOI22_X1 U17602 ( .A1(n19786), .A2(n20510), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19785), .ZN(n14078) );
  OAI211_X1 U17603 ( .C1(n19794), .C2(n19855), .A(n14079), .B(n14078), .ZN(
        P2_U2917) );
  OR2_X1 U17604 ( .A1(n13057), .A2(n14080), .ZN(n14081) );
  NAND2_X1 U17605 ( .A1(n14082), .A2(n14081), .ZN(n16897) );
  NAND2_X1 U17606 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14273) );
  INV_X1 U17607 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14083) );
  NOR2_X1 U17608 ( .A1(n14273), .A2(n14083), .ZN(n14084) );
  NAND3_X1 U17609 ( .A1(n16313), .A2(n16294), .A3(n14084), .ZN(n14087) );
  NAND2_X1 U17610 ( .A1(n14085), .A2(n16304), .ZN(n14086) );
  NOR2_X1 U17611 ( .A1(n14087), .A2(n14086), .ZN(n14091) );
  AND3_X1 U17612 ( .A1(n16120), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        n14091), .ZN(n14089) );
  AND4_X1 U17613 ( .A1(n16120), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .A4(n14091), .ZN(n14092) );
  NAND2_X1 U17614 ( .A1(n14018), .A2(n14092), .ZN(n14093) );
  OAI211_X1 U17615 ( .C1(n14095), .C2(n14096), .A(n15967), .B(n16311), .ZN(
        n14098) );
  NAND2_X1 U17616 ( .A1(n16287), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14097) );
  OAI211_X1 U17617 ( .C1(n16897), .C2(n16287), .A(n14098), .B(n14097), .ZN(
        P2_U2875) );
  NAND2_X1 U17618 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  AND2_X1 U17619 ( .A1(n14099), .A2(n14102), .ZN(n20736) );
  INV_X1 U17620 ( .A(n20736), .ZN(n14191) );
  INV_X1 U17621 ( .A(n14988), .ZN(n20831) );
  INV_X1 U17622 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20685) );
  OAI222_X1 U17623 ( .A1(n15038), .A2(n14191), .B1(n20831), .B2(n15037), .C1(
        n20685), .C2(n15036), .ZN(P1_U2900) );
  INV_X1 U17624 ( .A(n20169), .ZN(n20498) );
  INV_X1 U17625 ( .A(n14350), .ZN(n14354) );
  NAND2_X1 U17626 ( .A1(n17345), .A2(n14354), .ZN(n14118) );
  INV_X1 U17627 ( .A(n14372), .ZN(n14104) );
  AND2_X1 U17628 ( .A1(n14104), .A2(n14103), .ZN(n14340) );
  NOR2_X1 U17629 ( .A1(n14105), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14332) );
  XNOR2_X1 U17630 ( .A(n14332), .B(n14341), .ZN(n14115) );
  INV_X1 U17631 ( .A(n14107), .ZN(n14108) );
  OAI21_X1 U17632 ( .B1(n16201), .B2(n14341), .A(n14108), .ZN(n14109) );
  NAND2_X1 U17633 ( .A1(n14335), .A2(n14109), .ZN(n14114) );
  INV_X1 U17634 ( .A(n14110), .ZN(n14111) );
  OAI211_X1 U17635 ( .C1(n14112), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12676), .B(n14111), .ZN(n14113) );
  OAI211_X1 U17636 ( .C1(n14340), .C2(n14115), .A(n14114), .B(n14113), .ZN(
        n14116) );
  INV_X1 U17637 ( .A(n14116), .ZN(n14117) );
  NAND2_X1 U17638 ( .A1(n14118), .A2(n14117), .ZN(n14344) );
  AOI22_X1 U17639 ( .A1(n20498), .A2(n17016), .B1(n17050), .B2(n14344), .ZN(
        n14120) );
  NAND2_X1 U17640 ( .A1(n17010), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14119) );
  OAI21_X1 U17641 ( .B1(n14120), .B2(n17010), .A(n14119), .ZN(P2_U3596) );
  INV_X1 U17642 ( .A(n14121), .ZN(n14122) );
  NAND2_X1 U17643 ( .A1(n14123), .A2(n14122), .ZN(n14124) );
  INV_X1 U17644 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U17645 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14127) );
  NAND2_X1 U17646 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14126) );
  OAI211_X1 U17647 ( .C1(n18227), .C2(n14128), .A(n14127), .B(n14126), .ZN(
        n14129) );
  INV_X1 U17648 ( .A(n14129), .ZN(n14133) );
  AOI22_X1 U17649 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17650 ( .A1(n18220), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14144), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17651 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14130) );
  NAND4_X1 U17652 ( .A1(n14133), .A2(n14132), .A3(n14131), .A4(n14130), .ZN(
        n14140) );
  AOI22_X1 U17653 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14134), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17654 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17655 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13869), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17656 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14135) );
  NAND4_X1 U17657 ( .A1(n14138), .A2(n14137), .A3(n14136), .A4(n14135), .ZN(
        n14139) );
  XNOR2_X1 U17658 ( .A(n14143), .B(n18397), .ZN(n14141) );
  XNOR2_X1 U17659 ( .A(n14141), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18747) );
  INV_X1 U17660 ( .A(n14141), .ZN(n14142) );
  AOI22_X1 U17661 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17662 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14150) );
  INV_X1 U17663 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18094) );
  NAND2_X1 U17664 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n14146) );
  NAND2_X1 U17665 ( .A1(n10621), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14145) );
  OAI211_X1 U17666 ( .C1(n9602), .C2(n18094), .A(n14146), .B(n14145), .ZN(
        n14147) );
  INV_X1 U17667 ( .A(n14147), .ZN(n14149) );
  INV_X1 U17668 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17918) );
  OR2_X1 U17669 ( .A1(n18227), .A2(n17918), .ZN(n14148) );
  NAND4_X1 U17670 ( .A1(n14151), .A2(n14150), .A3(n14149), .A4(n14148), .ZN(
        n14157) );
  AOI22_X1 U17671 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17672 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17673 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17674 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17675 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  INV_X1 U17676 ( .A(n14158), .ZN(n14159) );
  NAND2_X1 U17677 ( .A1(n14159), .A2(n18394), .ZN(n14160) );
  NAND2_X1 U17678 ( .A1(n18663), .A2(n14160), .ZN(n14161) );
  NAND2_X1 U17679 ( .A1(n18740), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18739) );
  INV_X1 U17680 ( .A(n14161), .ZN(n14162) );
  NAND2_X1 U17681 ( .A1(n14163), .A2(n14162), .ZN(n14164) );
  NAND2_X2 U17682 ( .A1(n14165), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18664) );
  XNOR2_X1 U17683 ( .A(n17167), .B(n18644), .ZN(n17172) );
  INV_X1 U17684 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19015) );
  NAND2_X1 U17685 ( .A1(n14166), .A2(n19045), .ZN(n19014) );
  NOR3_X1 U17686 ( .A1(n19015), .A2(n19026), .A3(n19014), .ZN(n17249) );
  INV_X1 U17687 ( .A(n17249), .ZN(n14167) );
  OR2_X1 U17688 ( .A1(n19514), .A2(n17215), .ZN(n18987) );
  OAI22_X1 U17689 ( .A1(n14167), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18987), .B2(n17167), .ZN(n14187) );
  NAND2_X1 U17690 ( .A1(n14169), .A2(n14168), .ZN(n14173) );
  NOR2_X1 U17691 ( .A1(n18397), .A2(n14173), .ZN(n14177) );
  NAND2_X1 U17692 ( .A1(n14177), .A2(n17215), .ZN(n14446) );
  INV_X1 U17693 ( .A(n14446), .ZN(n14180) );
  AND2_X1 U17694 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14170), .ZN(
        n14172) );
  XNOR2_X1 U17695 ( .A(n14173), .B(n18397), .ZN(n14175) );
  NOR2_X1 U17696 ( .A1(n14174), .A2(n14175), .ZN(n14176) );
  XOR2_X1 U17697 ( .A(n14177), .B(n18394), .Z(n14178) );
  AOI21_X1 U17698 ( .B1(n14180), .B2(n14445), .A(n14179), .ZN(n14181) );
  AOI21_X1 U17699 ( .B1(n14181), .B2(n10023), .A(n14447), .ZN(n17168) );
  INV_X1 U17700 ( .A(n17168), .ZN(n14185) );
  AOI211_X1 U17701 ( .C1(n18920), .C2(n19026), .A(n19015), .B(n14182), .ZN(
        n19013) );
  OAI21_X1 U17702 ( .B1(n19013), .B2(n19035), .A(n19072), .ZN(n14183) );
  AOI22_X1 U17703 ( .A1(n14183), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13950), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n14184) );
  OAI21_X1 U17704 ( .B1(n14185), .B2(n19021), .A(n14184), .ZN(n14186) );
  AOI21_X1 U17705 ( .B1(n19070), .B2(n14187), .A(n14186), .ZN(n14188) );
  OAI21_X1 U17706 ( .B1(n17172), .B2(n18956), .A(n14188), .ZN(P3_U2854) );
  AOI21_X1 U17707 ( .B1(n14190), .B2(n14189), .A(n15541), .ZN(n20646) );
  INV_X1 U17708 ( .A(n20646), .ZN(n20747) );
  OAI222_X1 U17709 ( .A1(n20747), .A2(n14933), .B1(n20662), .B2(n11964), .C1(
        n14191), .C2(n14935), .ZN(P1_U2868) );
  NOR3_X1 U17710 ( .A1(n17259), .A2(n9889), .A3(n19102), .ZN(n14194) );
  OR2_X1 U17711 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  INV_X1 U17712 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18495) );
  INV_X1 U17713 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18472) );
  NOR2_X1 U17714 ( .A1(n18495), .A2(n18472), .ZN(n14202) );
  AOI211_X1 U17715 ( .C1(n18495), .C2(n18472), .A(n18319), .B(n14202), .ZN(
        n14197) );
  AOI21_X1 U17716 ( .B1(n18389), .B2(n14198), .A(n14197), .ZN(n14201) );
  NAND2_X1 U17717 ( .A1(n14199), .A2(n18357), .ZN(n18413) );
  AOI22_X1 U17718 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18378), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n10359), .ZN(n14200) );
  NAND2_X1 U17719 ( .A1(n14201), .A2(n14200), .ZN(P3_U2734) );
  NAND3_X1 U17720 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n18273) );
  OAI221_X1 U17721 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n14203), .C1(
        P3_EAX_REG_2__SCAN_IN), .C2(n14202), .A(n18408), .ZN(n14206) );
  AOI22_X1 U17722 ( .A1(n14204), .A2(n18389), .B1(BUF2_REG_2__SCAN_IN), .B2(
        n18378), .ZN(n14205) );
  OAI21_X1 U17723 ( .B1(n18407), .B2(n14206), .A(n14205), .ZN(P3_U2733) );
  XOR2_X1 U17724 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14274), .Z(n14213)
         );
  INV_X1 U17725 ( .A(n14207), .ZN(n14211) );
  INV_X1 U17726 ( .A(n14208), .ZN(n14210) );
  OAI21_X1 U17727 ( .B1(n14211), .B2(n14210), .A(n14209), .ZN(n17331) );
  MUX2_X1 U17728 ( .A(n11155), .B(n17331), .S(n16308), .Z(n14212) );
  OAI21_X1 U17729 ( .B1(n14213), .B2(n16301), .A(n14212), .ZN(P2_U2882) );
  AOI22_X1 U17730 ( .A1(n14214), .A2(n18389), .B1(BUF2_REG_0__SCAN_IN), .B2(
        n18378), .ZN(n14216) );
  NAND2_X1 U17731 ( .A1(n10359), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n14215) );
  OAI211_X1 U17732 ( .C1(n18319), .C2(P3_EAX_REG_0__SCAN_IN), .A(n14216), .B(
        n14215), .ZN(P3_U2735) );
  INV_X1 U17733 ( .A(n14217), .ZN(n14218) );
  AND2_X1 U17734 ( .A1(n14218), .A2(n14099), .ZN(n14219) );
  NOR2_X1 U17735 ( .A1(n14218), .A2(n14099), .ZN(n14930) );
  OR2_X1 U17736 ( .A1(n14219), .A2(n14930), .ZN(n15277) );
  INV_X1 U17737 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20683) );
  INV_X1 U17738 ( .A(n14220), .ZN(n20836) );
  OAI222_X1 U17739 ( .A1(n15277), .A2(n15038), .B1(n15036), .B2(n20683), .C1(
        n20836), .C2(n15037), .ZN(P1_U2899) );
  INV_X1 U17740 ( .A(n14221), .ZN(n14222) );
  NAND2_X1 U17741 ( .A1(n14222), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14224) );
  INV_X1 U17742 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14223) );
  NOR2_X1 U17743 ( .A1(n21282), .A2(n14227), .ZN(n17307) );
  INV_X1 U17744 ( .A(n17307), .ZN(n17304) );
  NAND2_X1 U17745 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21501), .ZN(n14229) );
  OAI21_X1 U17746 ( .B1(n14229), .B2(n14228), .A(n20786), .ZN(n14230) );
  INV_X1 U17747 ( .A(n14230), .ZN(n14231) );
  OAI21_X1 U17748 ( .B1(n17304), .B2(n21501), .A(n14231), .ZN(n14232) );
  INV_X1 U17749 ( .A(n14244), .ZN(n14233) );
  NAND2_X1 U17750 ( .A1(n14233), .A2(n9837), .ZN(n14234) );
  NAND2_X1 U17751 ( .A1(n20603), .A2(n14234), .ZN(n20652) );
  INV_X1 U17752 ( .A(n20652), .ZN(n14289) );
  INV_X1 U17753 ( .A(n14235), .ZN(n14236) );
  INV_X1 U17754 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14253) );
  INV_X1 U17755 ( .A(n14237), .ZN(n20787) );
  NAND2_X1 U17756 ( .A1(n21581), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14240) );
  AND2_X1 U17757 ( .A1(n21590), .A2(n21373), .ZN(n17302) );
  NOR2_X1 U17758 ( .A1(n14240), .A2(n17302), .ZN(n14238) );
  NOR2_X1 U17759 ( .A1(n14239), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14249) );
  INV_X1 U17760 ( .A(n14240), .ZN(n14241) );
  NOR2_X1 U17761 ( .A1(n14249), .A2(n14241), .ZN(n14242) );
  NAND2_X1 U17762 ( .A1(n14250), .A2(n14242), .ZN(n20627) );
  INV_X2 U17763 ( .A(n20627), .ZN(n14862) );
  NOR2_X1 U17764 ( .A1(n14244), .A2(n14243), .ZN(n20639) );
  INV_X1 U17765 ( .A(n20639), .ZN(n14259) );
  INV_X1 U17766 ( .A(n20594), .ZN(n14246) );
  AOI22_X1 U17767 ( .A1(n20611), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14246), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14247) );
  OAI21_X1 U17768 ( .B1(n14259), .B2(n14245), .A(n14247), .ZN(n14248) );
  AOI21_X1 U17769 ( .B1(n14862), .B2(P1_EBX_REG_1__SCAN_IN), .A(n14248), .ZN(
        n14251) );
  INV_X1 U17770 ( .A(n20593), .ZN(n14868) );
  INV_X1 U17771 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21571) );
  NAND2_X1 U17772 ( .A1(n14868), .A2(n21571), .ZN(n14256) );
  OAI211_X1 U17773 ( .C1(n20787), .C2(n20615), .A(n14251), .B(n14256), .ZN(
        n14252) );
  AOI21_X1 U17774 ( .B1(n14836), .B2(n14253), .A(n14252), .ZN(n14254) );
  OAI21_X1 U17775 ( .B1(n14289), .B2(n14255), .A(n14254), .ZN(P1_U2839) );
  NAND2_X1 U17776 ( .A1(n14256), .A2(n20594), .ZN(n14269) );
  INV_X1 U17777 ( .A(n21118), .ZN(n15559) );
  AOI22_X1 U17778 ( .A1(n14862), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20611), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U17779 ( .A1(n20647), .A2(n20755), .ZN(n14257) );
  OAI211_X1 U17780 ( .C1(n15559), .C2(n14259), .A(n14258), .B(n14257), .ZN(
        n14262) );
  NAND2_X1 U17781 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20638) );
  OAI21_X1 U17782 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20638), .ZN(n14260) );
  OAI22_X1 U17783 ( .A1(n20649), .A2(n15285), .B1(n14260), .B2(n20637), .ZN(
        n14261) );
  AOI211_X1 U17784 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n14269), .A(n14262), .B(
        n14261), .ZN(n14263) );
  OAI21_X1 U17785 ( .B1(n14264), .B2(n14289), .A(n14263), .ZN(P1_U2837) );
  INV_X1 U17786 ( .A(n21279), .ZN(n20805) );
  AOI22_X1 U17787 ( .A1(n20805), .A2(n20639), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20611), .ZN(n14266) );
  NAND2_X1 U17788 ( .A1(n14862), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14265) );
  OAI211_X1 U17789 ( .C1(n20615), .C2(n20773), .A(n14266), .B(n14265), .ZN(
        n14268) );
  OAI22_X1 U17790 ( .A1(n20649), .A2(n15290), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n20637), .ZN(n14267) );
  AOI211_X1 U17791 ( .C1(n14269), .C2(P1_REIP_REG_2__SCAN_IN), .A(n14268), .B(
        n14267), .ZN(n14270) );
  OAI21_X1 U17792 ( .B1(n14271), .B2(n14289), .A(n14270), .ZN(P1_U2838) );
  INV_X1 U17793 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14272) );
  NOR2_X1 U17794 ( .A1(n14274), .A2(n14272), .ZN(n14276) );
  INV_X1 U17795 ( .A(n16291), .ZN(n14275) );
  OAI211_X1 U17796 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14276), .A(
        n14275), .B(n16311), .ZN(n14282) );
  INV_X1 U17797 ( .A(n14291), .ZN(n14277) );
  AOI21_X1 U17798 ( .B1(n14278), .B2(n14209), .A(n14277), .ZN(n19762) );
  INV_X1 U17799 ( .A(n19762), .ZN(n14279) );
  MUX2_X1 U17800 ( .A(n14280), .B(n14279), .S(n16308), .Z(n14281) );
  NAND2_X1 U17801 ( .A1(n14282), .A2(n14281), .ZN(P2_U2881) );
  OAI21_X1 U17802 ( .B1(n14836), .B2(n20611), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U17803 ( .A1(n20593), .A2(n20594), .ZN(n20596) );
  AOI22_X1 U17804 ( .A1(n14862), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n20930), .B2(
        n20639), .ZN(n14283) );
  OAI21_X1 U17805 ( .B1(n20615), .B2(n14284), .A(n14283), .ZN(n14285) );
  AOI21_X1 U17806 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n20596), .A(n14285), .ZN(
        n14286) );
  OAI211_X1 U17807 ( .C1(n14289), .C2(n14288), .A(n14287), .B(n14286), .ZN(
        P1_U2840) );
  XNOR2_X1 U17808 ( .A(n16291), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14294) );
  AND2_X1 U17809 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  OR2_X1 U17810 ( .A1(n14292), .A2(n15856), .ZN(n16955) );
  MUX2_X1 U17811 ( .A(n16955), .B(n11255), .S(n16287), .Z(n14293) );
  OAI21_X1 U17812 ( .B1(n14294), .B2(n16301), .A(n14293), .ZN(P2_U2880) );
  AND2_X1 U17813 ( .A1(n13058), .A2(n14295), .ZN(n14297) );
  OR2_X1 U17814 ( .A1(n14297), .A2(n14296), .ZN(n16884) );
  NOR2_X1 U17815 ( .A1(n15967), .A2(n14298), .ZN(n14301) );
  NAND2_X1 U17816 ( .A1(n14301), .A2(n14317), .ZN(n14398) );
  OAI211_X1 U17817 ( .C1(n14301), .C2(n14317), .A(n14398), .B(n16311), .ZN(
        n14300) );
  NAND2_X1 U17818 ( .A1(n16287), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14299) );
  OAI211_X1 U17819 ( .C1(n16884), .C2(n16287), .A(n14300), .B(n14299), .ZN(
        P2_U2873) );
  NAND2_X1 U17820 ( .A1(n16584), .A2(n16308), .ZN(n14305) );
  INV_X1 U17821 ( .A(n15967), .ZN(n14303) );
  INV_X1 U17822 ( .A(n14301), .ZN(n14302) );
  OAI211_X1 U17823 ( .C1(n14303), .C2(n14318), .A(n14302), .B(n16311), .ZN(
        n14304) );
  OAI211_X1 U17824 ( .C1(n16308), .C2(n11258), .A(n14305), .B(n14304), .ZN(
        P2_U2874) );
  NOR2_X1 U17825 ( .A1(n14398), .A2(n14306), .ZN(n14399) );
  AOI22_X1 U17826 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17827 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U17828 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U17829 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14307) );
  NAND4_X1 U17830 ( .A1(n14310), .A2(n14309), .A3(n14308), .A4(n14307), .ZN(
        n14316) );
  AOI22_X1 U17831 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n14409), .ZN(n14314) );
  AOI22_X1 U17832 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U17833 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n16048), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17834 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14311) );
  NAND4_X1 U17835 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        n14315) );
  OR2_X1 U17836 ( .A1(n14316), .A2(n14315), .ZN(n14321) );
  NAND2_X1 U17837 ( .A1(n14401), .A2(n14317), .ZN(n15980) );
  AND2_X1 U17838 ( .A1(n14318), .A2(n14321), .ZN(n15979) );
  INV_X1 U17839 ( .A(n15979), .ZN(n14319) );
  NOR3_X1 U17840 ( .A1(n15967), .A2(n15980), .A3(n14319), .ZN(n14416) );
  INV_X1 U17841 ( .A(n14416), .ZN(n14320) );
  OAI21_X1 U17842 ( .B1(n14399), .B2(n14321), .A(n14320), .ZN(n16290) );
  AOI21_X1 U17843 ( .B1(n14324), .B2(n14049), .A(n14323), .ZN(n16864) );
  INV_X1 U17844 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U17845 ( .A1(n16408), .A2(n17019), .B1(n19785), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14328) );
  NAND2_X1 U17846 ( .A1(n16395), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14327) );
  OAI211_X1 U17847 ( .C1(n16392), .C2(n14329), .A(n14328), .B(n14327), .ZN(
        n14330) );
  AOI21_X1 U17848 ( .B1(n16864), .B2(n19786), .A(n14330), .ZN(n14331) );
  OAI21_X1 U17849 ( .B1(n16398), .B2(n16290), .A(n14331), .ZN(P2_U2903) );
  NOR2_X1 U17850 ( .A1(n14332), .A2(n16201), .ZN(n14339) );
  NAND2_X1 U17851 ( .A1(n14333), .A2(n14354), .ZN(n14338) );
  XNOR2_X1 U17852 ( .A(n14334), .B(n17004), .ZN(n14336) );
  AOI22_X1 U17853 ( .A1(n12676), .A2(n14336), .B1(n14335), .B2(n14339), .ZN(
        n14337) );
  OAI211_X1 U17854 ( .C1(n14340), .C2(n14339), .A(n14338), .B(n14337), .ZN(
        n17008) );
  MUX2_X1 U17855 ( .A(n17008), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14377), .Z(n14360) );
  INV_X1 U17856 ( .A(n14360), .ZN(n14381) );
  OR2_X1 U17857 ( .A1(n14344), .A2(n14377), .ZN(n14343) );
  NAND2_X1 U17858 ( .A1(n14377), .A2(n14341), .ZN(n14342) );
  NAND2_X1 U17859 ( .A1(n14343), .A2(n14342), .ZN(n14380) );
  INV_X1 U17860 ( .A(n14344), .ZN(n14358) );
  INV_X1 U17861 ( .A(n12681), .ZN(n14346) );
  NAND2_X1 U17862 ( .A1(n14346), .A2(n14345), .ZN(n14352) );
  AOI22_X1 U17863 ( .A1(n12676), .A2(n14348), .B1(n14352), .B2(n14347), .ZN(
        n14349) );
  OAI21_X1 U17864 ( .B1(n15946), .B2(n14350), .A(n14349), .ZN(n17000) );
  MUX2_X1 U17865 ( .A(n12676), .B(n14352), .S(n14351), .Z(n14353) );
  AOI21_X1 U17866 ( .B1(n15962), .B2(n14354), .A(n14353), .ZN(n16991) );
  AOI21_X1 U17867 ( .B1(n16991), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14356) );
  AOI21_X1 U17868 ( .B1(n16991), .B2(n20199), .A(n14377), .ZN(n14355) );
  OAI21_X1 U17869 ( .B1(n17000), .B2(n14356), .A(n14355), .ZN(n14357) );
  AOI21_X1 U17870 ( .B1(n14358), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n14357), .ZN(n14359) );
  AOI222_X1 U17871 ( .A1(n14360), .A2(n14359), .B1(n14360), .B2(n19950), .C1(
        n14359), .C2(n20512), .ZN(n14361) );
  OAI21_X1 U17872 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14380), .A(
        n14361), .ZN(n14362) );
  NAND2_X1 U17873 ( .A1(n14362), .A2(n17317), .ZN(n14379) );
  INV_X1 U17874 ( .A(n14363), .ZN(n14369) );
  NOR4_X1 U17875 ( .A1(n14364), .A2(n14366), .A3(n14365), .A4(n14374), .ZN(
        n19707) );
  OAI21_X1 U17876 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19707), .ZN(n14368) );
  OAI211_X1 U17877 ( .C1(n20550), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        n14376) );
  MUX2_X1 U17878 ( .A(n14372), .B(n14371), .S(n14370), .Z(n14373) );
  AOI21_X1 U17879 ( .B1(n14374), .B2(n12680), .A(n14373), .ZN(n20540) );
  INV_X1 U17880 ( .A(n20540), .ZN(n14375) );
  AOI211_X1 U17881 ( .C1(n14377), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14376), .B(n14375), .ZN(n14378) );
  OAI211_X1 U17882 ( .C1(n14381), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        n14392) );
  OAI21_X1 U17883 ( .B1(n14392), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14384) );
  NOR2_X1 U17884 ( .A1(n14382), .A2(n20552), .ZN(n14383) );
  OAI211_X1 U17885 ( .C1(n14386), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n17054) );
  OAI21_X1 U17886 ( .B1(n17016), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20551), 
        .ZN(n14388) );
  OAI21_X1 U17887 ( .B1(n17054), .B2(n20547), .A(n14388), .ZN(n14394) );
  INV_X1 U17888 ( .A(n14389), .ZN(n14391) );
  OAI22_X1 U17889 ( .A1(n20538), .A2(n17316), .B1(n17052), .B2(n20547), .ZN(
        n14390) );
  AOI211_X1 U17890 ( .C1(n14392), .C2(n17055), .A(n14391), .B(n14390), .ZN(
        n14393) );
  OAI211_X1 U17891 ( .C1(n17054), .C2(n20559), .A(n14394), .B(n14393), .ZN(
        P2_U3176) );
  OR2_X1 U17892 ( .A1(n14296), .A2(n14396), .ZN(n14397) );
  NAND2_X1 U17893 ( .A1(n14395), .A2(n14397), .ZN(n16868) );
  INV_X1 U17894 ( .A(n14398), .ZN(n14402) );
  INV_X1 U17895 ( .A(n14399), .ZN(n14400) );
  OAI211_X1 U17896 ( .C1(n14402), .C2(n14401), .A(n14400), .B(n16311), .ZN(
        n14404) );
  NAND2_X1 U17897 ( .A1(n16287), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14403) );
  OAI211_X1 U17898 ( .C1(n16868), .C2(n16287), .A(n14404), .B(n14403), .ZN(
        P2_U2872) );
  AOI22_X1 U17899 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17900 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17901 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17902 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14405) );
  NAND4_X1 U17903 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14415) );
  AOI22_X1 U17904 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n14409), .ZN(n14413) );
  AOI22_X1 U17905 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17906 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16048), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U17907 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14410) );
  NAND4_X1 U17908 ( .A1(n14413), .A2(n14412), .A3(n14411), .A4(n14410), .ZN(
        n14414) );
  OR2_X1 U17909 ( .A1(n14415), .A2(n14414), .ZN(n15978) );
  NAND2_X1 U17910 ( .A1(n14416), .A2(n15978), .ZN(n16282) );
  OAI21_X1 U17911 ( .B1(n14416), .B2(n15978), .A(n16282), .ZN(n16284) );
  INV_X1 U17912 ( .A(n14417), .ZN(n14420) );
  INV_X1 U17913 ( .A(n14323), .ZN(n14419) );
  AOI21_X1 U17914 ( .B1(n14420), .B2(n14419), .A(n14418), .ZN(n16853) );
  NAND2_X1 U17915 ( .A1(n16853), .A2(n19786), .ZN(n14425) );
  INV_X1 U17916 ( .A(n16408), .ZN(n16390) );
  OAI22_X1 U17917 ( .A1(n16390), .A2(n19852), .B1(n14421), .B2(n19768), .ZN(
        n14423) );
  NOR2_X1 U17918 ( .A1(n16392), .A2(n21618), .ZN(n14422) );
  AOI211_X1 U17919 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n16395), .A(n14423), .B(
        n14422), .ZN(n14424) );
  OAI211_X1 U17920 ( .C1(n16284), .C2(n16398), .A(n14425), .B(n14424), .ZN(
        P2_U2902) );
  NAND2_X1 U17921 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18668) );
  INV_X1 U17922 ( .A(n18668), .ZN(n18673) );
  NOR2_X1 U17923 ( .A1(n19010), .A2(n17144), .ZN(n17129) );
  NAND2_X1 U17924 ( .A1(n17129), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18717) );
  INV_X1 U17925 ( .A(n17065), .ZN(n17251) );
  INV_X1 U17926 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18675) );
  NOR2_X1 U17927 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18671) );
  NOR3_X1 U17928 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18665) );
  NAND3_X1 U17929 ( .A1(n18675), .A2(n18671), .A3(n18665), .ZN(n14426) );
  AOI21_X2 U17930 ( .B1(n18645), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14429), .ZN(n17247) );
  INV_X1 U17931 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U17932 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18628) );
  NAND2_X1 U17933 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18882) );
  INV_X1 U17934 ( .A(n18882), .ZN(n18866) );
  AND3_X1 U17935 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18866), .ZN(n14455) );
  INV_X1 U17936 ( .A(n18628), .ZN(n14451) );
  AND2_X1 U17937 ( .A1(n18828), .A2(n14451), .ZN(n17066) );
  NAND2_X1 U17938 ( .A1(n17066), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18539) );
  NAND2_X1 U17939 ( .A1(n18663), .A2(n18862), .ZN(n18625) );
  NOR2_X1 U17940 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18625), .ZN(
        n14431) );
  INV_X1 U17941 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U17942 ( .A1(n14431), .A2(n18864), .ZN(n18585) );
  NOR2_X1 U17943 ( .A1(n18585), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18569) );
  INV_X1 U17944 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18872) );
  INV_X1 U17945 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18844) );
  NAND3_X1 U17946 ( .A1(n18569), .A2(n18872), .A3(n18844), .ZN(n14432) );
  OAI21_X1 U17947 ( .B1(n18645), .B2(n18539), .A(n14432), .ZN(n14433) );
  INV_X1 U17948 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14434) );
  NAND2_X1 U17949 ( .A1(n14435), .A2(n18663), .ZN(n18541) );
  OAI211_X1 U17950 ( .C1(n18542), .C2(n14436), .A(n18541), .B(n10544), .ZN(
        n14437) );
  INV_X1 U17951 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18818) );
  INV_X1 U17952 ( .A(n18542), .ZN(n14438) );
  OAI21_X1 U17953 ( .B1(n14438), .B2(n14436), .A(n18644), .ZN(n14440) );
  AND2_X1 U17954 ( .A1(n14440), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14439) );
  NAND2_X1 U17955 ( .A1(n17114), .A2(n18644), .ZN(n17214) );
  AND2_X1 U17956 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17185) );
  NAND2_X1 U17957 ( .A1(n17185), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14466) );
  NOR2_X2 U17958 ( .A1(n17214), .A2(n14466), .ZN(n17060) );
  NAND2_X1 U17959 ( .A1(n18525), .A2(n14440), .ZN(n14441) );
  INV_X1 U17960 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17240) );
  NOR2_X1 U17961 ( .A1(n18644), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14443) );
  INV_X1 U17962 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17188) );
  NOR2_X1 U17963 ( .A1(n18844), .A2(n14434), .ZN(n18827) );
  NAND3_X1 U17964 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n18827), .ZN(n17241) );
  INV_X1 U17965 ( .A(n17241), .ZN(n17233) );
  NAND2_X1 U17966 ( .A1(n17066), .A2(n17233), .ZN(n14459) );
  NOR2_X1 U17967 ( .A1(n18927), .A2(n14459), .ZN(n17104) );
  INV_X1 U17968 ( .A(n17104), .ZN(n17239) );
  NOR2_X1 U17969 ( .A1(n17239), .A2(n14466), .ZN(n17182) );
  NAND2_X1 U17970 ( .A1(n17182), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14448) );
  XNOR2_X1 U17971 ( .A(n14448), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14489) );
  INV_X1 U17972 ( .A(n14449), .ZN(n14450) );
  NAND3_X1 U17973 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14453) );
  NOR2_X1 U17974 ( .A1(n14450), .A2(n14453), .ZN(n18981) );
  NAND2_X1 U17975 ( .A1(n17065), .A2(n18981), .ZN(n18883) );
  OR2_X1 U17976 ( .A1(n14459), .A2(n18883), .ZN(n14465) );
  INV_X1 U17977 ( .A(n18828), .ZN(n14454) );
  AND2_X1 U17978 ( .A1(n14451), .A2(n17065), .ZN(n17209) );
  NOR2_X1 U17979 ( .A1(n14453), .A2(n14452), .ZN(n18915) );
  NAND2_X1 U17980 ( .A1(n17209), .A2(n18915), .ZN(n14462) );
  AND2_X1 U17981 ( .A1(n14462), .A2(n9887), .ZN(n18861) );
  AOI21_X1 U17982 ( .B1(n9887), .B2(n14454), .A(n18861), .ZN(n18846) );
  OAI21_X1 U17983 ( .B1(n17233), .B2(n19061), .A(n18846), .ZN(n17235) );
  INV_X1 U17984 ( .A(n14455), .ZN(n18869) );
  NAND2_X1 U17985 ( .A1(n18981), .A2(n17209), .ZN(n17208) );
  NOR2_X1 U17986 ( .A1(n18869), .A2(n17208), .ZN(n17232) );
  NAND2_X1 U17987 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17232), .ZN(
        n18857) );
  NOR2_X1 U17988 ( .A1(n18872), .A2(n18857), .ZN(n14463) );
  NOR2_X1 U17989 ( .A1(n17241), .A2(n17240), .ZN(n17211) );
  AOI21_X1 U17990 ( .B1(n14463), .B2(n17211), .A(n18994), .ZN(n14456) );
  AOI211_X1 U17991 ( .C1(n19081), .C2(n14465), .A(n17235), .B(n14456), .ZN(
        n17197) );
  NAND2_X1 U17992 ( .A1(n14458), .A2(n14466), .ZN(n14457) );
  OAI211_X1 U17993 ( .C1(n17197), .C2(n19080), .A(n19072), .B(n14457), .ZN(
        n17183) );
  AOI21_X1 U17994 ( .B1(n14458), .B2(n17188), .A(n17183), .ZN(n14471) );
  INV_X1 U17995 ( .A(n18645), .ZN(n18929) );
  INV_X1 U17996 ( .A(n14459), .ZN(n14460) );
  INV_X1 U17997 ( .A(n14466), .ZN(n17189) );
  NAND2_X1 U17998 ( .A1(n17237), .A2(n17189), .ZN(n17180) );
  OR2_X1 U17999 ( .A1(n17180), .A2(n17188), .ZN(n14461) );
  XNOR2_X1 U18000 ( .A(n14461), .B(n14470), .ZN(n14487) );
  NOR2_X1 U18001 ( .A1(n19061), .A2(n14462), .ZN(n17206) );
  AOI22_X1 U18002 ( .A1(n17206), .A2(n18828), .B1(n14463), .B2(n18971), .ZN(
        n14464) );
  OAI22_X1 U18003 ( .A1(n18943), .A2(n14465), .B1(n14464), .B2(n17241), .ZN(
        n17184) );
  NAND3_X1 U18004 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n14470), .A3(
        n17184), .ZN(n14467) );
  OAI22_X1 U18005 ( .A1(n14487), .A2(n18987), .B1(n14467), .B2(n14466), .ZN(
        n14468) );
  NAND2_X1 U18006 ( .A1(n14468), .A2(n19070), .ZN(n14469) );
  NAND2_X1 U18007 ( .A1(n13950), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n14480) );
  OAI211_X1 U18008 ( .C1(n14471), .C2(n14470), .A(n14469), .B(n14480), .ZN(
        n14472) );
  AOI21_X1 U18009 ( .B1(n14489), .B2(n19079), .A(n14472), .ZN(n14473) );
  OAI21_X1 U18010 ( .B1(n14491), .B2(n18956), .A(n14473), .ZN(P3_U2831) );
  INV_X1 U18011 ( .A(n19515), .ZN(n14474) );
  NAND2_X1 U18012 ( .A1(n19692), .A2(n19660), .ZN(n17446) );
  NAND2_X1 U18013 ( .A1(n17256), .A2(n17446), .ZN(n19087) );
  NAND2_X1 U18014 ( .A1(n19087), .A2(n19657), .ZN(n14476) );
  NAND2_X1 U18015 ( .A1(n19657), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19570) );
  INV_X1 U18016 ( .A(n19570), .ZN(n18704) );
  INV_X1 U18017 ( .A(n18573), .ZN(n18598) );
  NOR2_X1 U18018 ( .A1(n18598), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17080) );
  NAND3_X1 U18019 ( .A1(n14477), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17079) );
  NOR2_X1 U18020 ( .A1(n17478), .A2(n17079), .ZN(n14482) );
  INV_X1 U18021 ( .A(n14482), .ZN(n14478) );
  AOI22_X1 U18022 ( .A1(n17078), .A2(n14478), .B1(n18704), .B2(n17081), .ZN(
        n14479) );
  NAND2_X1 U18023 ( .A1(n18807), .A2(n14479), .ZN(n17085) );
  NOR2_X1 U18024 ( .A1(n17080), .A2(n17085), .ZN(n17068) );
  OAI21_X1 U18025 ( .B1(n17068), .B2(n14481), .A(n14480), .ZN(n14485) );
  AOI21_X2 U18026 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18573), .A(
        n17078), .ZN(n18649) );
  INV_X1 U18027 ( .A(n18649), .ZN(n18699) );
  NAND2_X1 U18028 ( .A1(n14482), .A2(n18699), .ZN(n17063) );
  XNOR2_X1 U18029 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14483) );
  NOR2_X1 U18030 ( .A1(n17063), .A2(n14483), .ZN(n14484) );
  AOI211_X1 U18031 ( .C1(n18730), .C2(n17748), .A(n14485), .B(n14484), .ZN(
        n14486) );
  OAI21_X1 U18032 ( .B1(n18696), .B2(n14487), .A(n14486), .ZN(n14488) );
  AOI21_X1 U18033 ( .B1(n18812), .B2(n14489), .A(n14488), .ZN(n14490) );
  OAI21_X1 U18034 ( .B1(n14491), .B2(n18732), .A(n14490), .ZN(P3_U2799) );
  NAND2_X1 U18035 ( .A1(n14492), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14494) );
  NAND2_X1 U18036 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  XNOR2_X1 U18037 ( .A(n14495), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14544) );
  NAND2_X1 U18038 ( .A1(n14576), .A2(n14496), .ZN(n14501) );
  AOI22_X1 U18039 ( .A1(n14498), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14497), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14499) );
  INV_X1 U18040 ( .A(n14499), .ZN(n14500) );
  NAND2_X1 U18041 ( .A1(n20731), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U18042 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14502) );
  OAI211_X1 U18043 ( .C1(n14503), .C2(n20742), .A(n14538), .B(n14502), .ZN(
        n14504) );
  OAI21_X1 U18044 ( .B1(n14544), .B2(n20574), .A(n14505), .ZN(P1_U2968) );
  OR2_X1 U18045 ( .A1(n14588), .A2(n14506), .ZN(n14507) );
  NAND2_X1 U18046 ( .A1(n14592), .A2(n14508), .ZN(n14509) );
  AOI22_X1 U18047 ( .A1(n10551), .A2(n20658), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14927), .ZN(n14511) );
  OAI21_X1 U18048 ( .B1(n15055), .B2(n14935), .A(n14511), .ZN(P1_U2844) );
  INV_X1 U18049 ( .A(n15057), .ZN(n14523) );
  AOI22_X1 U18050 ( .A1(n14862), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20611), .ZN(n14522) );
  INV_X1 U18051 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15061) );
  NAND3_X1 U18052 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20631) );
  NOR2_X1 U18053 ( .A1(n21571), .A2(n20631), .ZN(n20592) );
  NAND4_X1 U18054 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20592), .A3(
        P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14873) );
  INV_X1 U18055 ( .A(n14873), .ZN(n14512) );
  NAND2_X1 U18056 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14512), .ZN(n14863) );
  NAND2_X1 U18057 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14513) );
  NOR2_X1 U18058 ( .A1(n14863), .A2(n14513), .ZN(n14815) );
  INV_X1 U18059 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21544) );
  NAND2_X1 U18060 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14756) );
  NAND2_X1 U18061 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14736) );
  NOR3_X1 U18062 ( .A1(n21544), .A2(n14756), .A3(n14736), .ZN(n14716) );
  NAND3_X1 U18063 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n14716), .ZN(n14515) );
  NAND2_X1 U18064 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14514) );
  NOR2_X1 U18065 ( .A1(n14515), .A2(n14514), .ZN(n14516) );
  NAND2_X1 U18066 ( .A1(n14815), .A2(n14516), .ZN(n14664) );
  NAND2_X1 U18067 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14650) );
  INV_X1 U18068 ( .A(n14650), .ZN(n14669) );
  NAND3_X1 U18069 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(n14669), .ZN(n14517) );
  OR2_X1 U18070 ( .A1(n14664), .A2(n14517), .ZN(n14627) );
  NAND2_X1 U18071 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14518) );
  NOR2_X1 U18072 ( .A1(n14627), .A2(n14518), .ZN(n14610) );
  NAND2_X1 U18073 ( .A1(n14610), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14595) );
  NOR3_X1 U18074 ( .A1(n20593), .A2(n15061), .A3(n14595), .ZN(n14520) );
  INV_X1 U18075 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21605) );
  OR3_X1 U18076 ( .A1(n14595), .A2(n15061), .A3(n21605), .ZN(n14559) );
  INV_X1 U18077 ( .A(n14559), .ZN(n14579) );
  OR2_X1 U18078 ( .A1(n20593), .A2(n14579), .ZN(n14519) );
  NAND2_X1 U18079 ( .A1(n14519), .A2(n20594), .ZN(n14585) );
  OAI21_X1 U18080 ( .B1(n14520), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14585), 
        .ZN(n14521) );
  OAI211_X1 U18081 ( .C1(n20649), .C2(n14523), .A(n14522), .B(n14521), .ZN(
        n14524) );
  AOI21_X1 U18082 ( .B1(n10551), .B2(n20647), .A(n14524), .ZN(n14525) );
  OAI21_X1 U18083 ( .B1(n15055), .B2(n20603), .A(n14525), .ZN(P1_U2812) );
  NAND2_X1 U18084 ( .A1(n14527), .A2(n14526), .ZN(n14528) );
  NAND2_X1 U18085 ( .A1(n14529), .A2(n14528), .ZN(n14534) );
  AOI22_X1 U18086 ( .A1(n14531), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14530), .ZN(n14532) );
  INV_X1 U18087 ( .A(n14532), .ZN(n14533) );
  XNOR2_X2 U18088 ( .A(n14534), .B(n14533), .ZN(n14888) );
  NAND2_X1 U18089 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14541) );
  NAND3_X1 U18090 ( .A1(n14537), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14536), .ZN(n14539) );
  OAI211_X1 U18091 ( .C1(n14541), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        n14542) );
  OAI21_X1 U18092 ( .B1(n14544), .B2(n20784), .A(n14543), .ZN(P1_U3000) );
  INV_X1 U18093 ( .A(DATAI_31_), .ZN(n14549) );
  AND2_X1 U18094 ( .A1(n15036), .A2(n14545), .ZN(n14546) );
  NAND2_X1 U18095 ( .A1(n14557), .A2(n14546), .ZN(n14548) );
  AOI22_X1 U18096 ( .A1(n15016), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15009), .ZN(n14547) );
  OAI211_X1 U18097 ( .C1(n15014), .C2(n14549), .A(n14548), .B(n14547), .ZN(
        P1_U2873) );
  AOI22_X1 U18098 ( .A1(n16395), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19785), .ZN(n14551) );
  NAND2_X1 U18099 ( .A1(n16409), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14550) );
  OAI211_X1 U18100 ( .C1(n14552), .C2(n19770), .A(n14551), .B(n14550), .ZN(
        P2_U2888) );
  NAND2_X1 U18101 ( .A1(n16287), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14553) );
  OAI21_X1 U18102 ( .B1(n13162), .B2(n16287), .A(n14553), .ZN(P2_U2856) );
  OR2_X1 U18103 ( .A1(n14713), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14556) );
  INV_X1 U18104 ( .A(n14554), .ZN(n14555) );
  MUX2_X1 U18105 ( .A(n14556), .B(n14555), .S(n21588), .Z(P1_U3487) );
  INV_X1 U18106 ( .A(n14557), .ZN(n14565) );
  AOI21_X1 U18107 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(P1_REIP_REG_30__SCAN_IN), 
        .A(n20593), .ZN(n14558) );
  NOR2_X1 U18108 ( .A1(n14558), .A2(n14585), .ZN(n14568) );
  INV_X1 U18109 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U18110 ( .A1(n14862), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20611), .ZN(n14561) );
  NOR3_X1 U18111 ( .A1(n20593), .A2(n14578), .A3(n14559), .ZN(n14570) );
  NAND3_X1 U18112 ( .A1(n14570), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14562), 
        .ZN(n14560) );
  OAI211_X1 U18113 ( .C1(n14568), .C2(n14562), .A(n14561), .B(n14560), .ZN(
        n14563) );
  AOI21_X1 U18114 ( .B1(n14888), .B2(n20647), .A(n14563), .ZN(n14564) );
  OAI21_X1 U18115 ( .B1(n14565), .B2(n20603), .A(n14564), .ZN(P1_U2809) );
  INV_X1 U18116 ( .A(n14566), .ZN(n14893) );
  INV_X1 U18117 ( .A(n14567), .ZN(n14573) );
  INV_X1 U18118 ( .A(n14568), .ZN(n14569) );
  OAI21_X1 U18119 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14570), .A(n14569), 
        .ZN(n14572) );
  AOI22_X1 U18120 ( .A1(n14862), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20611), .ZN(n14571) );
  OAI211_X1 U18121 ( .C1(n14573), .C2(n20649), .A(n14572), .B(n14571), .ZN(
        n14574) );
  AOI21_X1 U18122 ( .B1(n14891), .B2(n20647), .A(n14574), .ZN(n14575) );
  OAI21_X1 U18123 ( .B1(n14893), .B2(n20603), .A(n14575), .ZN(P1_U2810) );
  AOI21_X1 U18124 ( .B1(n14577), .B2(n9660), .A(n14576), .ZN(n15043) );
  INV_X1 U18125 ( .A(n15043), .ZN(n14896) );
  NAND2_X1 U18126 ( .A1(n14579), .A2(n14578), .ZN(n14583) );
  INV_X1 U18127 ( .A(n15041), .ZN(n14580) );
  NAND2_X1 U18128 ( .A1(n14836), .A2(n14580), .ZN(n14582) );
  AOI22_X1 U18129 ( .A1(n14862), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20611), .ZN(n14581) );
  OAI211_X1 U18130 ( .C1(n20593), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14584) );
  AOI21_X1 U18131 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14585), .A(n14584), 
        .ZN(n14587) );
  NAND2_X1 U18132 ( .A1(n14894), .A2(n20647), .ZN(n14586) );
  OAI211_X1 U18133 ( .C1(n14896), .C2(n20603), .A(n14587), .B(n14586), .ZN(
        P1_U2811) );
  AOI21_X1 U18134 ( .B1(n14589), .B2(n14603), .A(n14588), .ZN(n15065) );
  INV_X1 U18135 ( .A(n15065), .ZN(n14899) );
  NAND2_X1 U18136 ( .A1(n14608), .A2(n14590), .ZN(n14591) );
  NAND2_X1 U18137 ( .A1(n14592), .A2(n14591), .ZN(n14897) );
  INV_X1 U18138 ( .A(n14897), .ZN(n15310) );
  OR2_X1 U18139 ( .A1(n20649), .A2(n15063), .ZN(n14599) );
  AOI22_X1 U18140 ( .A1(n14862), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20611), .ZN(n14598) );
  INV_X1 U18141 ( .A(n14595), .ZN(n14593) );
  OR2_X1 U18142 ( .A1(n20593), .A2(n14593), .ZN(n14594) );
  NAND2_X1 U18143 ( .A1(n14594), .A2(n20594), .ZN(n14612) );
  NAND2_X1 U18144 ( .A1(n14612), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14597) );
  OR3_X1 U18145 ( .A1(n20593), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14595), .ZN(
        n14596) );
  NAND4_X1 U18146 ( .A1(n14599), .A2(n14598), .A3(n14597), .A4(n14596), .ZN(
        n14600) );
  AOI21_X1 U18147 ( .B1(n15310), .B2(n20647), .A(n14600), .ZN(n14601) );
  OAI21_X1 U18148 ( .B1(n14899), .B2(n20603), .A(n14601), .ZN(P1_U2813) );
  OAI21_X1 U18149 ( .B1(n14602), .B2(n14604), .A(n14603), .ZN(n14956) );
  OR2_X1 U18150 ( .A1(n14605), .A2(n14606), .ZN(n14607) );
  AND2_X1 U18151 ( .A1(n14608), .A2(n14607), .ZN(n15317) );
  INV_X1 U18152 ( .A(n14609), .ZN(n15074) );
  AOI22_X1 U18153 ( .A1(n14862), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20611), .ZN(n14615) );
  INV_X1 U18154 ( .A(n14610), .ZN(n14611) );
  NOR2_X1 U18155 ( .A1(n20593), .A2(n14611), .ZN(n14613) );
  OAI21_X1 U18156 ( .B1(n14613), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14612), 
        .ZN(n14614) );
  OAI211_X1 U18157 ( .C1(n20649), .C2(n15074), .A(n14615), .B(n14614), .ZN(
        n14616) );
  AOI21_X1 U18158 ( .B1(n15317), .B2(n20647), .A(n14616), .ZN(n14617) );
  OAI21_X1 U18159 ( .B1(n14956), .B2(n20603), .A(n14617), .ZN(P1_U2814) );
  AOI21_X1 U18160 ( .B1(n14619), .B2(n14618), .A(n14602), .ZN(n15085) );
  INV_X1 U18161 ( .A(n15085), .ZN(n14967) );
  NOR2_X1 U18162 ( .A1(n14641), .A2(n14620), .ZN(n14621) );
  OR2_X1 U18163 ( .A1(n14605), .A2(n14621), .ZN(n14901) );
  INV_X1 U18164 ( .A(n14901), .ZN(n15326) );
  OAI21_X1 U18165 ( .B1(n14627), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14622) );
  OAI21_X1 U18166 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(P1_REIP_REG_24__SCAN_IN), 
        .A(n14622), .ZN(n14625) );
  NAND2_X1 U18167 ( .A1(n14862), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14624) );
  NAND2_X1 U18168 ( .A1(n20611), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14623) );
  OAI211_X1 U18169 ( .C1(n14625), .C2(n20593), .A(n14624), .B(n14623), .ZN(
        n14626) );
  INV_X1 U18170 ( .A(n14626), .ZN(n14630) );
  INV_X1 U18171 ( .A(n14627), .ZN(n14636) );
  OR2_X1 U18172 ( .A1(n20593), .A2(n14636), .ZN(n14628) );
  NAND2_X1 U18173 ( .A1(n14628), .A2(n20594), .ZN(n14651) );
  NAND2_X1 U18174 ( .A1(n14651), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14629) );
  OAI211_X1 U18175 ( .C1(n20649), .C2(n15083), .A(n14630), .B(n14629), .ZN(
        n14631) );
  AOI21_X1 U18176 ( .B1(n15326), .B2(n20647), .A(n14631), .ZN(n14632) );
  OAI21_X1 U18177 ( .B1(n14967), .B2(n20603), .A(n14632), .ZN(P1_U2815) );
  OAI21_X1 U18178 ( .B1(n14633), .B2(n14634), .A(n14618), .ZN(n15092) );
  INV_X1 U18179 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U18180 ( .A1(n14636), .A2(n14635), .ZN(n14639) );
  NAND2_X1 U18181 ( .A1(n14836), .A2(n15095), .ZN(n14638) );
  AOI22_X1 U18182 ( .A1(n14862), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20611), .ZN(n14637) );
  OAI211_X1 U18183 ( .C1(n20593), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14640) );
  AOI21_X1 U18184 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14651), .A(n14640), 
        .ZN(n14644) );
  AOI21_X1 U18185 ( .B1(n14642), .B2(n14647), .A(n14641), .ZN(n15338) );
  NAND2_X1 U18186 ( .A1(n15338), .A2(n20647), .ZN(n14643) );
  OAI211_X1 U18187 ( .C1(n15092), .C2(n20603), .A(n14644), .B(n14643), .ZN(
        P1_U2816) );
  AOI21_X1 U18188 ( .B1(n14646), .B2(n14645), .A(n14633), .ZN(n15102) );
  INV_X1 U18189 ( .A(n15102), .ZN(n14904) );
  INV_X1 U18190 ( .A(n14647), .ZN(n14648) );
  AOI21_X1 U18191 ( .B1(n14649), .B2(n14662), .A(n14648), .ZN(n15346) );
  OR2_X1 U18192 ( .A1(n20593), .A2(n14664), .ZN(n14668) );
  INV_X1 U18193 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15110) );
  NOR3_X1 U18194 ( .A1(n14668), .A2(n14650), .A3(n15110), .ZN(n14652) );
  OAI21_X1 U18195 ( .B1(n14652), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14651), 
        .ZN(n14654) );
  AOI22_X1 U18196 ( .A1(n14862), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20611), .ZN(n14653) );
  OAI211_X1 U18197 ( .C1(n20649), .C2(n15100), .A(n14654), .B(n14653), .ZN(
        n14655) );
  AOI21_X1 U18198 ( .B1(n15346), .B2(n20647), .A(n14655), .ZN(n14656) );
  OAI21_X1 U18199 ( .B1(n14904), .B2(n20603), .A(n14656), .ZN(P1_U2817) );
  OAI21_X1 U18200 ( .B1(n14657), .B2(n14658), .A(n14645), .ZN(n14978) );
  OR2_X1 U18201 ( .A1(n14659), .A2(n14660), .ZN(n14661) );
  NAND2_X1 U18202 ( .A1(n14662), .A2(n14661), .ZN(n15356) );
  INV_X1 U18203 ( .A(n15356), .ZN(n14675) );
  INV_X1 U18204 ( .A(n14663), .ZN(n15112) );
  OR2_X1 U18205 ( .A1(n20649), .A2(n15112), .ZN(n14673) );
  AOI22_X1 U18206 ( .A1(n14862), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20611), .ZN(n14672) );
  INV_X1 U18207 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U18208 ( .A1(n14664), .A2(n15127), .ZN(n14665) );
  OR2_X1 U18209 ( .A1(n20593), .A2(n14665), .ZN(n14666) );
  NAND2_X1 U18210 ( .A1(n14666), .A2(n20594), .ZN(n14693) );
  NOR2_X1 U18211 ( .A1(n20593), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14667) );
  OAI21_X1 U18212 ( .B1(n14693), .B2(n14667), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14671) );
  INV_X1 U18213 ( .A(n14668), .ZN(n14694) );
  NAND3_X1 U18214 ( .A1(n14694), .A2(n15110), .A3(n14669), .ZN(n14670) );
  NAND4_X1 U18215 ( .A1(n14673), .A2(n14672), .A3(n14671), .A4(n14670), .ZN(
        n14674) );
  AOI21_X1 U18216 ( .B1(n14675), .B2(n20647), .A(n14674), .ZN(n14676) );
  OAI21_X1 U18217 ( .B1(n14978), .B2(n20603), .A(n14676), .ZN(P1_U2818) );
  AOI21_X1 U18218 ( .B1(n14678), .B2(n14677), .A(n14657), .ZN(n14679) );
  INV_X1 U18219 ( .A(n14679), .ZN(n15124) );
  NOR2_X1 U18220 ( .A1(n14680), .A2(n14681), .ZN(n14682) );
  OR2_X1 U18221 ( .A1(n14659), .A2(n14682), .ZN(n15364) );
  INV_X1 U18222 ( .A(n15364), .ZN(n14688) );
  INV_X1 U18223 ( .A(n15120), .ZN(n14683) );
  AOI22_X1 U18224 ( .A1(n14836), .A2(n14683), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n14693), .ZN(n14686) );
  AOI22_X1 U18225 ( .A1(n14862), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20611), .ZN(n14685) );
  INV_X1 U18226 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15119) );
  NAND3_X1 U18227 ( .A1(n14694), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n15119), 
        .ZN(n14684) );
  NAND3_X1 U18228 ( .A1(n14686), .A2(n14685), .A3(n14684), .ZN(n14687) );
  AOI21_X1 U18229 ( .B1(n14688), .B2(n20647), .A(n14687), .ZN(n14689) );
  OAI21_X1 U18230 ( .B1(n15124), .B2(n20603), .A(n14689), .ZN(P1_U2819) );
  OAI21_X1 U18231 ( .B1(n14690), .B2(n14691), .A(n14677), .ZN(n15132) );
  AOI21_X1 U18232 ( .B1(n14692), .B2(n14703), .A(n14680), .ZN(n14907) );
  INV_X1 U18233 ( .A(n15129), .ZN(n14697) );
  AOI22_X1 U18234 ( .A1(n14862), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20611), .ZN(n14696) );
  OAI21_X1 U18235 ( .B1(n14694), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14693), 
        .ZN(n14695) );
  OAI211_X1 U18236 ( .C1(n20649), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14698) );
  AOI21_X1 U18237 ( .B1(n14907), .B2(n20647), .A(n14698), .ZN(n14699) );
  OAI21_X1 U18238 ( .B1(n15132), .B2(n20603), .A(n14699), .ZN(P1_U2820) );
  NOR2_X1 U18239 ( .A1(n14700), .A2(n14701), .ZN(n14702) );
  OR2_X1 U18240 ( .A1(n14690), .A2(n14702), .ZN(n14993) );
  INV_X1 U18241 ( .A(n14703), .ZN(n14704) );
  AOI21_X1 U18242 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n15390) );
  INV_X1 U18243 ( .A(n14815), .ZN(n14707) );
  OR2_X1 U18244 ( .A1(n20593), .A2(n14707), .ZN(n14829) );
  NAND2_X1 U18245 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14708) );
  NOR2_X1 U18246 ( .A1(n14829), .A2(n14708), .ZN(n14800) );
  INV_X1 U18247 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15143) );
  NAND3_X1 U18248 ( .A1(n14800), .A2(n14716), .A3(n15143), .ZN(n14727) );
  AND2_X1 U18249 ( .A1(n20594), .A2(n14815), .ZN(n14832) );
  INV_X1 U18250 ( .A(n14708), .ZN(n14709) );
  NAND2_X1 U18251 ( .A1(n14832), .A2(n14709), .ZN(n14710) );
  NAND2_X1 U18252 ( .A1(n20596), .A2(n14710), .ZN(n14797) );
  INV_X1 U18253 ( .A(n14716), .ZN(n14711) );
  NAND2_X1 U18254 ( .A1(n20596), .A2(n14711), .ZN(n14712) );
  AND2_X1 U18255 ( .A1(n14797), .A2(n14712), .ZN(n14737) );
  INV_X1 U18256 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21547) );
  AOI21_X1 U18257 ( .B1(n14727), .B2(n14737), .A(n21547), .ZN(n14720) );
  NOR2_X1 U18258 ( .A1(n20655), .A2(n14714), .ZN(n14715) );
  AOI211_X1 U18259 ( .C1(n14862), .C2(P1_EBX_REG_19__SCAN_IN), .A(n20629), .B(
        n14715), .ZN(n14718) );
  NAND4_X1 U18260 ( .A1(n14800), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n14716), 
        .A4(n21547), .ZN(n14717) );
  OAI211_X1 U18261 ( .C1(n20649), .C2(n15136), .A(n14718), .B(n14717), .ZN(
        n14719) );
  AOI211_X1 U18262 ( .C1(n15390), .C2(n20647), .A(n14720), .B(n14719), .ZN(
        n14721) );
  OAI21_X1 U18263 ( .B1(n14993), .B2(n20603), .A(n14721), .ZN(P1_U2821) );
  AOI21_X1 U18264 ( .B1(n14723), .B2(n14722), .A(n14700), .ZN(n15142) );
  INV_X1 U18265 ( .A(n15142), .ZN(n14911) );
  XOR2_X1 U18266 ( .A(n14724), .B(n14735), .Z(n15411) );
  NAND2_X1 U18267 ( .A1(n14862), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14725) );
  OAI211_X1 U18268 ( .C1(n20655), .C2(n15144), .A(n14725), .B(n20641), .ZN(
        n14726) );
  AOI21_X1 U18269 ( .B1(n14836), .B2(n15146), .A(n14726), .ZN(n14728) );
  OAI211_X1 U18270 ( .C1(n14737), .C2(n15143), .A(n14728), .B(n14727), .ZN(
        n14729) );
  AOI21_X1 U18271 ( .B1(n15411), .B2(n20647), .A(n14729), .ZN(n14730) );
  OAI21_X1 U18272 ( .B1(n14911), .B2(n20603), .A(n14730), .ZN(P1_U2822) );
  AOI21_X1 U18273 ( .B1(n14732), .B2(n14731), .A(n10531), .ZN(n15160) );
  INV_X1 U18274 ( .A(n15160), .ZN(n15008) );
  AND2_X1 U18275 ( .A1(n14749), .A2(n14733), .ZN(n14734) );
  NOR2_X1 U18276 ( .A1(n14735), .A2(n14734), .ZN(n15416) );
  NAND3_X1 U18277 ( .A1(n14800), .A2(P1_REIP_REG_13__SCAN_IN), .A3(
        P1_REIP_REG_14__SCAN_IN), .ZN(n14755) );
  NOR2_X1 U18278 ( .A1(n14755), .A2(n14736), .ZN(n14739) );
  INV_X1 U18279 ( .A(n14737), .ZN(n14738) );
  OAI21_X1 U18280 ( .B1(n14739), .B2(P1_REIP_REG_17__SCAN_IN), .A(n14738), 
        .ZN(n14743) );
  OAI21_X1 U18281 ( .B1(n20655), .B2(n14740), .A(n20641), .ZN(n14741) );
  AOI21_X1 U18282 ( .B1(n14862), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14741), .ZN(
        n14742) );
  OAI211_X1 U18283 ( .C1(n20649), .C2(n15158), .A(n14743), .B(n14742), .ZN(
        n14744) );
  AOI21_X1 U18284 ( .B1(n15416), .B2(n20647), .A(n14744), .ZN(n14745) );
  OAI21_X1 U18285 ( .B1(n15008), .B2(n20603), .A(n14745), .ZN(P1_U2823) );
  OAI21_X1 U18286 ( .B1(n14746), .B2(n14747), .A(n14731), .ZN(n15173) );
  INV_X1 U18287 ( .A(n14749), .ZN(n14750) );
  AOI21_X1 U18288 ( .B1(n14751), .B2(n14748), .A(n14750), .ZN(n15427) );
  NAND2_X1 U18289 ( .A1(n14862), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14752) );
  OAI211_X1 U18290 ( .C1(n20655), .C2(n15168), .A(n14752), .B(n20641), .ZN(
        n14754) );
  INV_X1 U18291 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21540) );
  NOR3_X1 U18292 ( .A1(n14755), .A2(P1_REIP_REG_16__SCAN_IN), .A3(n21540), 
        .ZN(n14753) );
  AOI211_X1 U18293 ( .C1(n14836), .C2(n15171), .A(n14754), .B(n14753), .ZN(
        n14759) );
  NOR2_X1 U18294 ( .A1(n14755), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14771) );
  NAND2_X1 U18295 ( .A1(n20596), .A2(n14756), .ZN(n14757) );
  NAND2_X1 U18296 ( .A1(n14797), .A2(n14757), .ZN(n14787) );
  OAI21_X1 U18297 ( .B1(n14771), .B2(n14787), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14758) );
  NAND2_X1 U18298 ( .A1(n14759), .A2(n14758), .ZN(n14760) );
  AOI21_X1 U18299 ( .B1(n20647), .B2(n15427), .A(n14760), .ZN(n14761) );
  OAI21_X1 U18300 ( .B1(n15173), .B2(n20603), .A(n14761), .ZN(P1_U2824) );
  NAND2_X1 U18301 ( .A1(n14762), .A2(n14763), .ZN(n14764) );
  NAND2_X1 U18302 ( .A1(n14748), .A2(n14764), .ZN(n15433) );
  INV_X1 U18303 ( .A(n14765), .ZN(n14790) );
  INV_X1 U18304 ( .A(n14793), .ZN(n14824) );
  AND2_X1 U18305 ( .A1(n14765), .A2(n14789), .ZN(n14792) );
  INV_X1 U18306 ( .A(n14792), .ZN(n14766) );
  OAI21_X1 U18307 ( .B1(n14790), .B2(n14824), .A(n14766), .ZN(n14767) );
  NAND3_X1 U18308 ( .A1(n14767), .A2(n14796), .A3(n14794), .ZN(n14795) );
  OR2_X1 U18309 ( .A1(n14795), .A2(n14777), .ZN(n14775) );
  AOI21_X1 U18310 ( .B1(n14775), .B2(n14768), .A(n14746), .ZN(n15183) );
  NAND2_X1 U18311 ( .A1(n15183), .A2(n20620), .ZN(n14774) );
  AOI21_X1 U18312 ( .B1(n20611), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20629), .ZN(n14770) );
  NAND2_X1 U18313 ( .A1(n14862), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14769) );
  OAI211_X1 U18314 ( .C1(n20649), .C2(n15181), .A(n14770), .B(n14769), .ZN(
        n14772) );
  AOI211_X1 U18315 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n14787), .A(n14772), 
        .B(n14771), .ZN(n14773) );
  OAI211_X1 U18316 ( .C1(n15433), .C2(n20615), .A(n14774), .B(n14773), .ZN(
        P1_U2825) );
  INV_X1 U18317 ( .A(n14775), .ZN(n14776) );
  AOI21_X1 U18318 ( .B1(n14777), .B2(n14795), .A(n14776), .ZN(n15196) );
  INV_X1 U18319 ( .A(n15196), .ZN(n15021) );
  INV_X1 U18320 ( .A(n14800), .ZN(n14779) );
  INV_X1 U18321 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21537) );
  INV_X1 U18322 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14778) );
  OAI21_X1 U18323 ( .B1(n14779), .B2(n21537), .A(n14778), .ZN(n14786) );
  AOI21_X1 U18324 ( .B1(n20611), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20629), .ZN(n14781) );
  NAND2_X1 U18325 ( .A1(n14862), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14780) );
  OAI211_X1 U18326 ( .C1(n20649), .C2(n15194), .A(n14781), .B(n14780), .ZN(
        n14785) );
  OAI21_X1 U18327 ( .B1(n14782), .B2(n14783), .A(n14762), .ZN(n15441) );
  NOR2_X1 U18328 ( .A1(n15441), .A2(n20615), .ZN(n14784) );
  AOI211_X1 U18329 ( .C1(n14787), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        n14788) );
  OAI21_X1 U18330 ( .B1(n15021), .B2(n20603), .A(n14788), .ZN(P1_U2826) );
  INV_X1 U18331 ( .A(n14789), .ZN(n14791) );
  AOI21_X1 U18332 ( .B1(n14791), .B2(n14790), .A(n14792), .ZN(n14825) );
  AOI21_X1 U18333 ( .B1(n14825), .B2(n14793), .A(n14792), .ZN(n14814) );
  INV_X1 U18334 ( .A(n14794), .ZN(n14813) );
  NOR2_X1 U18335 ( .A1(n14814), .A2(n14813), .ZN(n14812) );
  OAI21_X1 U18336 ( .B1(n14812), .B2(n14796), .A(n14795), .ZN(n15209) );
  INV_X1 U18337 ( .A(n14797), .ZN(n14821) );
  NAND2_X1 U18338 ( .A1(n20611), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14798) );
  NAND2_X1 U18339 ( .A1(n20641), .A2(n14798), .ZN(n14799) );
  AOI21_X1 U18340 ( .B1(n14862), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14799), .ZN(
        n14802) );
  NAND2_X1 U18341 ( .A1(n14800), .A2(n21537), .ZN(n14801) );
  OAI211_X1 U18342 ( .C1(n20649), .C2(n15204), .A(n14802), .B(n14801), .ZN(
        n14809) );
  INV_X1 U18343 ( .A(n14804), .ZN(n14811) );
  INV_X1 U18344 ( .A(n14805), .ZN(n14806) );
  AOI21_X1 U18345 ( .B1(n14803), .B2(n14811), .A(n14806), .ZN(n14807) );
  OR2_X1 U18346 ( .A1(n14782), .A2(n14807), .ZN(n15455) );
  NOR2_X1 U18347 ( .A1(n15455), .A2(n20615), .ZN(n14808) );
  AOI211_X1 U18348 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n14821), .A(n14809), 
        .B(n14808), .ZN(n14810) );
  OAI21_X1 U18349 ( .B1(n15209), .B2(n20603), .A(n14810), .ZN(P1_U2827) );
  XNOR2_X1 U18350 ( .A(n14803), .B(n14811), .ZN(n15466) );
  AOI21_X1 U18351 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n15218) );
  NAND2_X1 U18352 ( .A1(n15218), .A2(n20620), .ZN(n14823) );
  NAND2_X1 U18353 ( .A1(n14815), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n14816) );
  INV_X1 U18354 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15214) );
  OAI21_X1 U18355 ( .B1(n20593), .B2(n14816), .A(n15214), .ZN(n14820) );
  AOI21_X1 U18356 ( .B1(n20611), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20629), .ZN(n14818) );
  NAND2_X1 U18357 ( .A1(n14862), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14817) );
  OAI211_X1 U18358 ( .C1(n20649), .C2(n15216), .A(n14818), .B(n14817), .ZN(
        n14819) );
  AOI21_X1 U18359 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14822) );
  OAI211_X1 U18360 ( .C1(n15466), .C2(n20615), .A(n14823), .B(n14822), .ZN(
        P1_U2828) );
  XNOR2_X1 U18361 ( .A(n14825), .B(n14824), .ZN(n15226) );
  INV_X1 U18362 ( .A(n15224), .ZN(n14837) );
  OAI21_X1 U18363 ( .B1(n20655), .B2(n14826), .A(n20641), .ZN(n14827) );
  AOI21_X1 U18364 ( .B1(n14862), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14827), .ZN(
        n14828) );
  OAI21_X1 U18365 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n14829), .A(n14828), 
        .ZN(n14835) );
  AND2_X1 U18366 ( .A1(n14844), .A2(n14830), .ZN(n14831) );
  OR2_X1 U18367 ( .A1(n14831), .A2(n14803), .ZN(n15476) );
  INV_X1 U18368 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21534) );
  INV_X1 U18369 ( .A(n14832), .ZN(n14833) );
  NAND2_X1 U18370 ( .A1(n20596), .A2(n14833), .ZN(n14853) );
  OAI22_X1 U18371 ( .A1(n15476), .A2(n20615), .B1(n21534), .B2(n14853), .ZN(
        n14834) );
  AOI211_X1 U18372 ( .C1(n14837), .C2(n14836), .A(n14835), .B(n14834), .ZN(
        n14838) );
  OAI21_X1 U18373 ( .B1(n15029), .B2(n20603), .A(n14838), .ZN(P1_U2829) );
  INV_X1 U18374 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15241) );
  NOR2_X1 U18375 ( .A1(n14863), .A2(n15241), .ZN(n14839) );
  AOI21_X1 U18376 ( .B1(n14868), .B2(n14839), .A(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14854) );
  AND2_X1 U18377 ( .A1(n14840), .A2(n14841), .ZN(n14842) );
  NOR2_X1 U18378 ( .A1(n14765), .A2(n14842), .ZN(n15237) );
  NAND2_X1 U18379 ( .A1(n15237), .A2(n20620), .ZN(n14852) );
  INV_X1 U18380 ( .A(n14844), .ZN(n14845) );
  AOI21_X1 U18381 ( .B1(n14846), .B2(n14843), .A(n14845), .ZN(n15490) );
  NAND2_X1 U18382 ( .A1(n14862), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14847) );
  OAI211_X1 U18383 ( .C1(n20655), .C2(n14848), .A(n14847), .B(n20641), .ZN(
        n14850) );
  NOR2_X1 U18384 ( .A1(n20649), .A2(n15235), .ZN(n14849) );
  AOI211_X1 U18385 ( .C1(n15490), .C2(n20647), .A(n14850), .B(n14849), .ZN(
        n14851) );
  OAI211_X1 U18386 ( .C1(n14854), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        P1_U2830) );
  INV_X1 U18387 ( .A(n14840), .ZN(n14856) );
  AOI21_X1 U18388 ( .B1(n14857), .B2(n14855), .A(n14856), .ZN(n15245) );
  INV_X1 U18389 ( .A(n15245), .ZN(n15033) );
  INV_X1 U18390 ( .A(n14863), .ZN(n14858) );
  OR2_X1 U18391 ( .A1(n20593), .A2(n14858), .ZN(n14859) );
  NAND2_X1 U18392 ( .A1(n14859), .A2(n20594), .ZN(n14882) );
  NAND2_X1 U18393 ( .A1(n20611), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14860) );
  NAND2_X1 U18394 ( .A1(n20641), .A2(n14860), .ZN(n14861) );
  AOI21_X1 U18395 ( .B1(n14862), .B2(P1_EBX_REG_9__SCAN_IN), .A(n14861), .ZN(
        n14870) );
  NOR2_X1 U18396 ( .A1(n14863), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14867) );
  OR2_X1 U18397 ( .A1(n14864), .A2(n14865), .ZN(n14866) );
  AND2_X1 U18398 ( .A1(n14843), .A2(n14866), .ZN(n15499) );
  AOI22_X1 U18399 ( .A1(n14868), .A2(n14867), .B1(n15499), .B2(n20647), .ZN(
        n14869) );
  OAI211_X1 U18400 ( .C1(n20649), .C2(n15243), .A(n14870), .B(n14869), .ZN(
        n14871) );
  AOI21_X1 U18401 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n14882), .A(n14871), .ZN(
        n14872) );
  OAI21_X1 U18402 ( .B1(n15033), .B2(n20603), .A(n14872), .ZN(P1_U2831) );
  NOR3_X1 U18403 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20593), .A3(n14873), .ZN(
        n14874) );
  AOI211_X1 U18404 ( .C1(n20611), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20629), .B(n14874), .ZN(n14887) );
  NAND2_X1 U18405 ( .A1(n14930), .A2(n14875), .ZN(n14929) );
  INV_X1 U18406 ( .A(n14876), .ZN(n14922) );
  INV_X1 U18407 ( .A(n14877), .ZN(n14878) );
  AOI21_X1 U18408 ( .B1(n14924), .B2(n14878), .A(n12214), .ZN(n15254) );
  NOR2_X1 U18409 ( .A1(n14879), .A2(n14880), .ZN(n14881) );
  OR2_X1 U18410 ( .A1(n14864), .A2(n14881), .ZN(n14921) );
  INV_X1 U18411 ( .A(n14921), .ZN(n15509) );
  AOI22_X1 U18412 ( .A1(n20647), .A2(n15509), .B1(n14862), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14884) );
  NAND2_X1 U18413 ( .A1(n14882), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n14883) );
  OAI211_X1 U18414 ( .C1(n20649), .C2(n15252), .A(n14884), .B(n14883), .ZN(
        n14885) );
  AOI21_X1 U18415 ( .B1(n15254), .B2(n20620), .A(n14885), .ZN(n14886) );
  NAND2_X1 U18416 ( .A1(n14887), .A2(n14886), .ZN(P1_U2832) );
  INV_X1 U18417 ( .A(n14888), .ZN(n14890) );
  INV_X1 U18418 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14889) );
  OAI22_X1 U18419 ( .A1(n14890), .A2(n14933), .B1(n20662), .B2(n14889), .ZN(
        P1_U2841) );
  AOI22_X1 U18420 ( .A1(n14891), .A2(n20658), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14927), .ZN(n14892) );
  OAI21_X1 U18421 ( .B1(n14893), .B2(n14935), .A(n14892), .ZN(P1_U2842) );
  AOI22_X1 U18422 ( .A1(n14894), .A2(n20658), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14927), .ZN(n14895) );
  OAI21_X1 U18423 ( .B1(n14896), .B2(n14935), .A(n14895), .ZN(P1_U2843) );
  INV_X1 U18424 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14898) );
  OAI222_X1 U18425 ( .A1(n14935), .A2(n14899), .B1(n14898), .B2(n20662), .C1(
        n14897), .C2(n14933), .ZN(P1_U2845) );
  AOI22_X1 U18426 ( .A1(n15317), .A2(n20658), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14927), .ZN(n14900) );
  OAI21_X1 U18427 ( .B1(n14956), .B2(n14935), .A(n14900), .ZN(P1_U2846) );
  INV_X1 U18428 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21648) );
  OAI222_X1 U18429 ( .A1(n14935), .A2(n14967), .B1(n21648), .B2(n20662), .C1(
        n14901), .C2(n14933), .ZN(P1_U2847) );
  INV_X1 U18430 ( .A(n15338), .ZN(n14902) );
  OAI222_X1 U18431 ( .A1(n14935), .A2(n15092), .B1(n21704), .B2(n20662), .C1(
        n14902), .C2(n14933), .ZN(P1_U2848) );
  AOI22_X1 U18432 ( .A1(n15346), .A2(n20658), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14927), .ZN(n14903) );
  OAI21_X1 U18433 ( .B1(n14904), .B2(n14935), .A(n14903), .ZN(P1_U2849) );
  OAI222_X1 U18434 ( .A1(n14978), .A2(n14935), .B1(n14905), .B2(n20662), .C1(
        n15356), .C2(n14933), .ZN(P1_U2850) );
  INV_X1 U18435 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14906) );
  OAI222_X1 U18436 ( .A1(n14935), .A2(n15124), .B1(n14906), .B2(n20662), .C1(
        n15364), .C2(n14933), .ZN(P1_U2851) );
  INV_X1 U18437 ( .A(n14907), .ZN(n15383) );
  OAI222_X1 U18438 ( .A1(n15132), .A2(n14935), .B1(n14908), .B2(n20662), .C1(
        n15383), .C2(n14933), .ZN(P1_U2852) );
  AOI22_X1 U18439 ( .A1(n15390), .A2(n20658), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14927), .ZN(n14909) );
  OAI21_X1 U18440 ( .B1(n14993), .B2(n14935), .A(n14909), .ZN(P1_U2853) );
  AOI22_X1 U18441 ( .A1(n15411), .A2(n20658), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14927), .ZN(n14910) );
  OAI21_X1 U18442 ( .B1(n14911), .B2(n14935), .A(n14910), .ZN(P1_U2854) );
  AOI22_X1 U18443 ( .A1(n15416), .A2(n20658), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14927), .ZN(n14912) );
  OAI21_X1 U18444 ( .B1(n15008), .B2(n14935), .A(n14912), .ZN(P1_U2855) );
  AOI22_X1 U18445 ( .A1(n15427), .A2(n20658), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14927), .ZN(n14913) );
  OAI21_X1 U18446 ( .B1(n15173), .B2(n14935), .A(n14913), .ZN(P1_U2856) );
  INV_X1 U18447 ( .A(n15183), .ZN(n15019) );
  INV_X1 U18448 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14914) );
  OAI222_X1 U18449 ( .A1(n15019), .A2(n14935), .B1(n14914), .B2(n20662), .C1(
        n15433), .C2(n14933), .ZN(P1_U2857) );
  OAI222_X1 U18450 ( .A1(n15021), .A2(n14935), .B1(n14915), .B2(n20662), .C1(
        n15441), .C2(n14933), .ZN(P1_U2858) );
  INV_X1 U18451 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14916) );
  OAI222_X1 U18452 ( .A1(n15209), .A2(n14935), .B1(n14916), .B2(n20662), .C1(
        n15455), .C2(n14933), .ZN(P1_U2859) );
  INV_X1 U18453 ( .A(n15218), .ZN(n15026) );
  OAI222_X1 U18454 ( .A1(n15026), .A2(n14935), .B1(n14917), .B2(n20662), .C1(
        n14933), .C2(n15466), .ZN(P1_U2860) );
  INV_X1 U18455 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14918) );
  OAI222_X1 U18456 ( .A1(n15029), .A2(n14935), .B1(n14918), .B2(n20662), .C1(
        n15476), .C2(n14933), .ZN(P1_U2861) );
  INV_X1 U18457 ( .A(n15237), .ZN(n15032) );
  AOI22_X1 U18458 ( .A1(n15490), .A2(n20658), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14927), .ZN(n14919) );
  OAI21_X1 U18459 ( .B1(n15032), .B2(n14935), .A(n14919), .ZN(P1_U2862) );
  AOI22_X1 U18460 ( .A1(n15499), .A2(n20658), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14927), .ZN(n14920) );
  OAI21_X1 U18461 ( .B1(n15033), .B2(n14935), .A(n14920), .ZN(P1_U2863) );
  INV_X1 U18462 ( .A(n15254), .ZN(n15035) );
  OAI222_X1 U18463 ( .A1(n15035), .A2(n14935), .B1(n20662), .B2(n11980), .C1(
        n14921), .C2(n14933), .ZN(P1_U2864) );
  NAND2_X1 U18464 ( .A1(n14929), .A2(n14922), .ZN(n14923) );
  NAND2_X1 U18465 ( .A1(n14924), .A2(n14923), .ZN(n20604) );
  AOI21_X1 U18466 ( .B1(n14926), .B2(n14925), .A(n14879), .ZN(n20597) );
  AOI22_X1 U18467 ( .A1(n20597), .A2(n20658), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14927), .ZN(n14928) );
  OAI21_X1 U18468 ( .B1(n20604), .B2(n14935), .A(n14928), .ZN(P1_U2865) );
  OAI21_X1 U18469 ( .B1(n14930), .B2(n14875), .A(n14929), .ZN(n20610) );
  XNOR2_X1 U18470 ( .A(n14931), .B(n14932), .ZN(n20614) );
  OAI222_X1 U18471 ( .A1(n20610), .A2(n14935), .B1(n14934), .B2(n20662), .C1(
        n14933), .C2(n20614), .ZN(P1_U2866) );
  INV_X1 U18472 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14942) );
  NAND2_X1 U18473 ( .A1(n15043), .A2(n14997), .ZN(n14941) );
  OR2_X1 U18474 ( .A1(n20796), .A2(n14936), .ZN(n14938) );
  NAND2_X1 U18475 ( .A1(n20796), .A2(DATAI_13_), .ZN(n14937) );
  NAND2_X1 U18476 ( .A1(n14938), .A2(n14937), .ZN(n20709) );
  INV_X1 U18477 ( .A(n20709), .ZN(n15023) );
  OAI22_X1 U18478 ( .A1(n15003), .A2(n15023), .B1(n15036), .B2(n13450), .ZN(
        n14939) );
  AOI21_X1 U18479 ( .B1(n15005), .B2(DATAI_29_), .A(n14939), .ZN(n14940) );
  OAI211_X1 U18480 ( .C1(n15001), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        P1_U2875) );
  INV_X1 U18481 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16334) );
  INV_X1 U18482 ( .A(n15055), .ZN(n14943) );
  NAND2_X1 U18483 ( .A1(n14943), .A2(n14997), .ZN(n14948) );
  OR2_X1 U18484 ( .A1(n20796), .A2(n21639), .ZN(n14945) );
  NAND2_X1 U18485 ( .A1(n20796), .A2(DATAI_12_), .ZN(n14944) );
  NAND2_X1 U18486 ( .A1(n14945), .A2(n14944), .ZN(n20707) );
  INV_X1 U18487 ( .A(n20707), .ZN(n15025) );
  OAI22_X1 U18488 ( .A1(n15003), .A2(n15025), .B1(n15036), .B2(n13448), .ZN(
        n14946) );
  AOI21_X1 U18489 ( .B1(n15005), .B2(DATAI_28_), .A(n14946), .ZN(n14947) );
  OAI211_X1 U18490 ( .C1(n15001), .C2(n16334), .A(n14948), .B(n14947), .ZN(
        P1_U2876) );
  INV_X1 U18491 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14955) );
  NAND2_X1 U18492 ( .A1(n15065), .A2(n14997), .ZN(n14954) );
  OR2_X1 U18493 ( .A1(n20796), .A2(n14949), .ZN(n14951) );
  NAND2_X1 U18494 ( .A1(n20796), .A2(DATAI_11_), .ZN(n14950) );
  NAND2_X1 U18495 ( .A1(n14951), .A2(n14950), .ZN(n20705) );
  INV_X1 U18496 ( .A(n20705), .ZN(n15028) );
  OAI22_X1 U18497 ( .A1(n15003), .A2(n15028), .B1(n15036), .B2(n13452), .ZN(
        n14952) );
  AOI21_X1 U18498 ( .B1(n15005), .B2(DATAI_27_), .A(n14952), .ZN(n14953) );
  OAI211_X1 U18499 ( .C1(n15001), .C2(n14955), .A(n14954), .B(n14953), .ZN(
        P1_U2877) );
  INV_X1 U18500 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16350) );
  INV_X1 U18501 ( .A(n14956), .ZN(n15076) );
  NAND2_X1 U18502 ( .A1(n15076), .A2(n14997), .ZN(n14961) );
  OR2_X1 U18503 ( .A1(n20796), .A2(n17389), .ZN(n14958) );
  NAND2_X1 U18504 ( .A1(n20796), .A2(DATAI_10_), .ZN(n14957) );
  NAND2_X1 U18505 ( .A1(n14958), .A2(n14957), .ZN(n20703) );
  INV_X1 U18506 ( .A(n20703), .ZN(n15031) );
  OAI22_X1 U18507 ( .A1(n15003), .A2(n15031), .B1(n15036), .B2(n13435), .ZN(
        n14959) );
  AOI21_X1 U18508 ( .B1(n15005), .B2(DATAI_26_), .A(n14959), .ZN(n14960) );
  OAI211_X1 U18509 ( .C1(n15001), .C2(n16350), .A(n14961), .B(n14960), .ZN(
        P1_U2878) );
  NOR2_X1 U18510 ( .A1(n20796), .A2(n17391), .ZN(n14962) );
  AOI21_X1 U18511 ( .B1(DATAI_9_), .B2(n20796), .A(n14962), .ZN(n20700) );
  INV_X1 U18512 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14963) );
  OAI22_X1 U18513 ( .A1(n15003), .A2(n20700), .B1(n15036), .B2(n14963), .ZN(
        n14964) );
  AOI21_X1 U18514 ( .B1(n15005), .B2(DATAI_25_), .A(n14964), .ZN(n14966) );
  NAND2_X1 U18515 ( .A1(n15016), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14965) );
  OAI211_X1 U18516 ( .C1(n14967), .C2(n15038), .A(n14966), .B(n14965), .ZN(
        P1_U2879) );
  NOR2_X1 U18517 ( .A1(n20796), .A2(n17393), .ZN(n14968) );
  AOI21_X1 U18518 ( .B1(DATAI_8_), .B2(n20796), .A(n14968), .ZN(n20697) );
  INV_X1 U18519 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14969) );
  OAI22_X1 U18520 ( .A1(n15003), .A2(n20697), .B1(n15036), .B2(n14969), .ZN(
        n14970) );
  AOI21_X1 U18521 ( .B1(n15005), .B2(DATAI_24_), .A(n14970), .ZN(n14972) );
  NAND2_X1 U18522 ( .A1(n15016), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14971) );
  OAI211_X1 U18523 ( .C1(n15092), .C2(n15038), .A(n14972), .B(n14971), .ZN(
        P1_U2880) );
  INV_X1 U18524 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16372) );
  NAND2_X1 U18525 ( .A1(n15102), .A2(n14997), .ZN(n14977) );
  OAI22_X1 U18526 ( .A1(n15003), .A2(n20849), .B1(n15036), .B2(n14974), .ZN(
        n14975) );
  AOI21_X1 U18527 ( .B1(n15005), .B2(DATAI_23_), .A(n14975), .ZN(n14976) );
  OAI211_X1 U18528 ( .C1(n15001), .C2(n16372), .A(n14977), .B(n14976), .ZN(
        P1_U2881) );
  INV_X1 U18529 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14983) );
  INV_X1 U18530 ( .A(n14978), .ZN(n15114) );
  NAND2_X1 U18531 ( .A1(n15114), .A2(n14997), .ZN(n14982) );
  INV_X1 U18532 ( .A(n14979), .ZN(n20841) );
  OAI22_X1 U18533 ( .A1(n15003), .A2(n20841), .B1(n15036), .B2(n13446), .ZN(
        n14980) );
  AOI21_X1 U18534 ( .B1(n15005), .B2(DATAI_22_), .A(n14980), .ZN(n14981) );
  OAI211_X1 U18535 ( .C1(n15001), .C2(n14983), .A(n14982), .B(n14981), .ZN(
        P1_U2882) );
  OAI22_X1 U18536 ( .A1(n15003), .A2(n20836), .B1(n15036), .B2(n14984), .ZN(
        n14985) );
  AOI21_X1 U18537 ( .B1(n15005), .B2(DATAI_21_), .A(n14985), .ZN(n14987) );
  NAND2_X1 U18538 ( .A1(n15016), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14986) );
  OAI211_X1 U18539 ( .C1(n15124), .C2(n15038), .A(n14987), .B(n14986), .ZN(
        P1_U2883) );
  INV_X1 U18540 ( .A(DATAI_20_), .ZN(n14990) );
  INV_X1 U18541 ( .A(n15003), .ZN(n15011) );
  AOI22_X1 U18542 ( .A1(n15011), .A2(n14988), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15009), .ZN(n14989) );
  OAI21_X1 U18543 ( .B1(n15014), .B2(n14990), .A(n14989), .ZN(n14991) );
  AOI21_X1 U18544 ( .B1(n15016), .B2(BUF1_REG_20__SCAN_IN), .A(n14991), .ZN(
        n14992) );
  OAI21_X1 U18545 ( .B1(n15132), .B2(n15038), .A(n14992), .ZN(P1_U2884) );
  INV_X1 U18546 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16403) );
  INV_X1 U18547 ( .A(n14993), .ZN(n15138) );
  NAND2_X1 U18548 ( .A1(n15138), .A2(n14997), .ZN(n14996) );
  OAI22_X1 U18549 ( .A1(n15003), .A2(n20826), .B1(n15036), .B2(n13440), .ZN(
        n14994) );
  AOI21_X1 U18550 ( .B1(n15005), .B2(DATAI_19_), .A(n14994), .ZN(n14995) );
  OAI211_X1 U18551 ( .C1(n15001), .C2(n16403), .A(n14996), .B(n14995), .ZN(
        P1_U2885) );
  INV_X1 U18552 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16412) );
  NAND2_X1 U18553 ( .A1(n15142), .A2(n14997), .ZN(n15000) );
  OAI22_X1 U18554 ( .A1(n15003), .A2(n20821), .B1(n15036), .B2(n13438), .ZN(
        n14998) );
  AOI21_X1 U18555 ( .B1(n15005), .B2(DATAI_18_), .A(n14998), .ZN(n14999) );
  OAI211_X1 U18556 ( .C1(n15001), .C2(n16412), .A(n15000), .B(n14999), .ZN(
        P1_U2886) );
  OAI22_X1 U18557 ( .A1(n15003), .A2(n20816), .B1(n15036), .B2(n15002), .ZN(
        n15004) );
  AOI21_X1 U18558 ( .B1(n15005), .B2(DATAI_17_), .A(n15004), .ZN(n15007) );
  NAND2_X1 U18559 ( .A1(n15016), .A2(BUF1_REG_17__SCAN_IN), .ZN(n15006) );
  OAI211_X1 U18560 ( .C1(n15008), .C2(n15038), .A(n15007), .B(n15006), .ZN(
        P1_U2887) );
  INV_X1 U18561 ( .A(DATAI_16_), .ZN(n15013) );
  AOI22_X1 U18562 ( .A1(n15011), .A2(n15010), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15009), .ZN(n15012) );
  OAI21_X1 U18563 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15015) );
  AOI21_X1 U18564 ( .B1(n15016), .B2(BUF1_REG_16__SCAN_IN), .A(n15015), .ZN(
        n15017) );
  OAI21_X1 U18565 ( .B1(n15173), .B2(n15038), .A(n15017), .ZN(P1_U2888) );
  OAI222_X1 U18566 ( .A1(n15038), .A2(n15019), .B1(n15037), .B2(n15018), .C1(
        n20669), .C2(n15036), .ZN(P1_U2889) );
  INV_X1 U18567 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15020) );
  OAI222_X1 U18568 ( .A1(n15021), .A2(n15038), .B1(n20711), .B2(n15037), .C1(
        n15020), .C2(n15036), .ZN(P1_U2890) );
  INV_X1 U18569 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15022) );
  OAI222_X1 U18570 ( .A1(n15038), .A2(n15209), .B1(n15023), .B2(n15037), .C1(
        n15022), .C2(n15036), .ZN(P1_U2891) );
  INV_X1 U18571 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15024) );
  OAI222_X1 U18572 ( .A1(n15026), .A2(n15038), .B1(n15025), .B2(n15037), .C1(
        n15024), .C2(n15036), .ZN(P1_U2892) );
  INV_X1 U18573 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15027) );
  OAI222_X1 U18574 ( .A1(n15038), .A2(n15029), .B1(n15028), .B2(n15037), .C1(
        n15027), .C2(n15036), .ZN(P1_U2893) );
  INV_X1 U18575 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15030) );
  OAI222_X1 U18576 ( .A1(n15038), .A2(n15032), .B1(n15031), .B2(n15037), .C1(
        n15030), .C2(n15036), .ZN(P1_U2894) );
  OAI222_X1 U18577 ( .A1(n15038), .A2(n15033), .B1(n20700), .B2(n15037), .C1(
        n20676), .C2(n15036), .ZN(P1_U2895) );
  INV_X1 U18578 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15034) );
  OAI222_X1 U18579 ( .A1(n15035), .A2(n15038), .B1(n20697), .B2(n15037), .C1(
        n15034), .C2(n15036), .ZN(P1_U2896) );
  INV_X1 U18580 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U18581 ( .A1(n15038), .A2(n20604), .B1(n20849), .B2(n15037), .C1(
        n15036), .C2(n20679), .ZN(P1_U2897) );
  INV_X1 U18582 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20681) );
  OAI222_X1 U18583 ( .A1(n20610), .A2(n15038), .B1(n20841), .B2(n15037), .C1(
        n20681), .C2(n15036), .ZN(P1_U2898) );
  AOI21_X1 U18584 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15039), .ZN(n15040) );
  OAI21_X1 U18585 ( .B1(n15041), .B2(n20742), .A(n15040), .ZN(n15042) );
  AOI21_X1 U18586 ( .B1(n15043), .B2(n20737), .A(n15042), .ZN(n15044) );
  OAI21_X1 U18587 ( .B1(n15045), .B2(n20574), .A(n15044), .ZN(P1_U2970) );
  OAI21_X1 U18588 ( .B1(n15220), .B2(n10455), .A(n15098), .ZN(n15051) );
  NAND4_X1 U18589 ( .A1(n11850), .A2(n15320), .A3(n15330), .A4(n15070), .ZN(
        n15047) );
  NAND2_X1 U18590 ( .A1(n15051), .A2(n15047), .ZN(n15050) );
  INV_X1 U18591 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15048) );
  MUX2_X1 U18592 ( .A(n15048), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15239), .Z(n15049) );
  OAI211_X1 U18593 ( .C1(n15051), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15050), .B(n15049), .ZN(n15053) );
  XNOR2_X1 U18594 ( .A(n15053), .B(n15052), .ZN(n15304) );
  NAND2_X1 U18595 ( .A1(n20731), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15297) );
  OAI21_X1 U18596 ( .B1(n15169), .B2(n15054), .A(n15297), .ZN(n15056) );
  NOR2_X1 U18597 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  NOR2_X1 U18598 ( .A1(n20786), .A2(n15061), .ZN(n15305) );
  AOI21_X1 U18599 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15305), .ZN(n15062) );
  OAI21_X1 U18600 ( .B1(n20742), .B2(n15063), .A(n15062), .ZN(n15064) );
  AOI21_X1 U18601 ( .B1(n15065), .B2(n20737), .A(n15064), .ZN(n15066) );
  INV_X1 U18602 ( .A(n15098), .ZN(n15087) );
  OAI21_X1 U18603 ( .B1(n15087), .B2(n15067), .A(n15239), .ZN(n15068) );
  NAND2_X1 U18604 ( .A1(n15069), .A2(n15068), .ZN(n15071) );
  XNOR2_X1 U18605 ( .A(n15071), .B(n15070), .ZN(n15319) );
  INV_X1 U18606 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U18607 ( .A1(n20786), .A2(n15072), .ZN(n15316) );
  AOI21_X1 U18608 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15316), .ZN(n15073) );
  OAI21_X1 U18609 ( .B1(n20742), .B2(n15074), .A(n15073), .ZN(n15075) );
  AOI21_X1 U18610 ( .B1(n15076), .B2(n20737), .A(n15075), .ZN(n15077) );
  OAI21_X1 U18611 ( .B1(n20574), .B2(n15319), .A(n15077), .ZN(P1_U2973) );
  INV_X1 U18612 ( .A(n15078), .ZN(n15079) );
  NAND2_X1 U18613 ( .A1(n15079), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15089) );
  XNOR2_X1 U18614 ( .A(n15080), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15329) );
  INV_X1 U18615 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U18616 ( .A1(n20786), .A2(n15081), .ZN(n15323) );
  AOI21_X1 U18617 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15323), .ZN(n15082) );
  OAI21_X1 U18618 ( .B1(n20742), .B2(n15083), .A(n15082), .ZN(n15084) );
  AOI21_X1 U18619 ( .B1(n15085), .B2(n20737), .A(n15084), .ZN(n15086) );
  OAI21_X1 U18620 ( .B1(n20574), .B2(n15329), .A(n15086), .ZN(P1_U2974) );
  NAND2_X1 U18621 ( .A1(n15089), .A2(n15087), .ZN(n15088) );
  MUX2_X1 U18622 ( .A(n15089), .B(n15088), .S(n15220), .Z(n15090) );
  XNOR2_X1 U18623 ( .A(n15090), .B(n15330), .ZN(n15340) );
  NAND2_X1 U18624 ( .A1(n20731), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15335) );
  OAI21_X1 U18625 ( .B1(n15169), .B2(n15091), .A(n15335), .ZN(n15094) );
  NOR2_X1 U18626 ( .A1(n15092), .A2(n20797), .ZN(n15093) );
  AOI211_X1 U18627 ( .C1(n15172), .C2(n15095), .A(n15094), .B(n15093), .ZN(
        n15096) );
  OAI21_X1 U18628 ( .B1(n20574), .B2(n15340), .A(n15096), .ZN(P1_U2975) );
  XNOR2_X1 U18629 ( .A(n15239), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15097) );
  XNOR2_X1 U18630 ( .A(n15098), .B(n15097), .ZN(n15348) );
  INV_X1 U18631 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21722) );
  NOR2_X1 U18632 ( .A1(n20786), .A2(n21722), .ZN(n15341) );
  AOI21_X1 U18633 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15341), .ZN(n15099) );
  OAI21_X1 U18634 ( .B1(n20742), .B2(n15100), .A(n15099), .ZN(n15101) );
  AOI21_X1 U18635 ( .B1(n15102), .B2(n20737), .A(n15101), .ZN(n15103) );
  OAI21_X1 U18636 ( .B1(n15348), .B2(n20574), .A(n15103), .ZN(P1_U2976) );
  INV_X1 U18637 ( .A(n15117), .ZN(n15106) );
  OAI21_X1 U18638 ( .B1(n15106), .B2(n15105), .A(n15239), .ZN(n15108) );
  NAND2_X1 U18639 ( .A1(n15108), .A2(n15107), .ZN(n15109) );
  XNOR2_X1 U18640 ( .A(n15109), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15349) );
  INV_X1 U18641 ( .A(n15349), .ZN(n15116) );
  NOR2_X1 U18642 ( .A1(n20786), .A2(n15110), .ZN(n15353) );
  AOI21_X1 U18643 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15353), .ZN(n15111) );
  OAI21_X1 U18644 ( .B1(n20742), .B2(n15112), .A(n15111), .ZN(n15113) );
  AOI21_X1 U18645 ( .B1(n15114), .B2(n20737), .A(n15113), .ZN(n15115) );
  OAI21_X1 U18646 ( .B1(n15116), .B2(n20574), .A(n15115), .ZN(P1_U2977) );
  XOR2_X1 U18647 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15118), .Z(
        n15357) );
  NAND2_X1 U18648 ( .A1(n15357), .A2(n20738), .ZN(n15123) );
  NOR2_X1 U18649 ( .A1(n20786), .A2(n15119), .ZN(n15360) );
  NOR2_X1 U18650 ( .A1(n20742), .A2(n15120), .ZN(n15121) );
  AOI211_X1 U18651 ( .C1(n20732), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15360), .B(n15121), .ZN(n15122) );
  OAI211_X1 U18652 ( .C1(n20797), .C2(n15124), .A(n15123), .B(n15122), .ZN(
        P1_U2978) );
  OAI21_X1 U18653 ( .B1(n15126), .B2(n11844), .A(n15125), .ZN(n15365) );
  NAND2_X1 U18654 ( .A1(n15365), .A2(n20738), .ZN(n15131) );
  NOR2_X1 U18655 ( .A1(n20786), .A2(n15127), .ZN(n15379) );
  NOR2_X1 U18656 ( .A1(n15169), .A2(n21627), .ZN(n15128) );
  AOI211_X1 U18657 ( .C1(n15172), .C2(n15129), .A(n15379), .B(n15128), .ZN(
        n15130) );
  OAI211_X1 U18658 ( .C1(n20797), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        P1_U2979) );
  NAND2_X1 U18659 ( .A1(n15104), .A2(n11843), .ZN(n15133) );
  MUX2_X1 U18660 ( .A(n15104), .B(n15133), .S(n15220), .Z(n15134) );
  XNOR2_X1 U18661 ( .A(n15134), .B(n11842), .ZN(n15393) );
  NOR2_X1 U18662 ( .A1(n20786), .A2(n21547), .ZN(n15387) );
  AOI21_X1 U18663 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15387), .ZN(n15135) );
  OAI21_X1 U18664 ( .B1(n20742), .B2(n15136), .A(n15135), .ZN(n15137) );
  AOI21_X1 U18665 ( .B1(n15138), .B2(n20737), .A(n15137), .ZN(n15139) );
  OAI21_X1 U18666 ( .B1(n15393), .B2(n20574), .A(n15139), .ZN(P1_U2980) );
  OAI21_X1 U18667 ( .B1(n15141), .B2(n15140), .A(n15104), .ZN(n15414) );
  NAND2_X1 U18668 ( .A1(n15142), .A2(n20737), .ZN(n15148) );
  NOR2_X1 U18669 ( .A1(n20786), .A2(n15143), .ZN(n15410) );
  NOR2_X1 U18670 ( .A1(n15169), .A2(n15144), .ZN(n15145) );
  AOI211_X1 U18671 ( .C1(n15172), .C2(n15146), .A(n15410), .B(n15145), .ZN(
        n15147) );
  OAI211_X1 U18672 ( .C1(n15414), .C2(n20574), .A(n15148), .B(n15147), .ZN(
        P1_U2981) );
  INV_X1 U18673 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15503) );
  INV_X1 U18674 ( .A(n15150), .ZN(n15151) );
  NOR2_X1 U18675 ( .A1(n15220), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15190) );
  INV_X1 U18676 ( .A(n15153), .ZN(n15186) );
  XNOR2_X1 U18677 ( .A(n15156), .B(n21716), .ZN(n15421) );
  NOR2_X1 U18678 ( .A1(n20786), .A2(n21544), .ZN(n15415) );
  AOI21_X1 U18679 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15415), .ZN(n15157) );
  OAI21_X1 U18680 ( .B1(n20742), .B2(n15158), .A(n15157), .ZN(n15159) );
  AOI21_X1 U18681 ( .B1(n15160), .B2(n20737), .A(n15159), .ZN(n15161) );
  OAI21_X1 U18682 ( .B1(n15421), .B2(n20574), .A(n15161), .ZN(P1_U2982) );
  INV_X1 U18683 ( .A(n15162), .ZN(n15163) );
  NOR2_X1 U18684 ( .A1(n15163), .A2(n15424), .ZN(n15166) );
  OAI21_X1 U18685 ( .B1(n15166), .B2(n15165), .A(n15164), .ZN(n15430) );
  INV_X1 U18686 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15167) );
  NOR2_X1 U18687 ( .A1(n20786), .A2(n15167), .ZN(n15425) );
  NOR2_X1 U18688 ( .A1(n15169), .A2(n15168), .ZN(n15170) );
  AOI211_X1 U18689 ( .C1(n15172), .C2(n15171), .A(n15425), .B(n15170), .ZN(
        n15176) );
  INV_X1 U18690 ( .A(n15173), .ZN(n15174) );
  NAND2_X1 U18691 ( .A1(n15174), .A2(n20737), .ZN(n15175) );
  OAI211_X1 U18692 ( .C1(n15430), .C2(n20574), .A(n15176), .B(n15175), .ZN(
        P1_U2983) );
  XNOR2_X1 U18693 ( .A(n15239), .B(n15177), .ZN(n15178) );
  XNOR2_X1 U18694 ( .A(n15179), .B(n15178), .ZN(n15438) );
  OR2_X1 U18695 ( .A1(n20786), .A2(n21540), .ZN(n15432) );
  NAND2_X1 U18696 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15180) );
  OAI211_X1 U18697 ( .C1(n20742), .C2(n15181), .A(n15432), .B(n15180), .ZN(
        n15182) );
  AOI21_X1 U18698 ( .B1(n15183), .B2(n20737), .A(n15182), .ZN(n15184) );
  OAI21_X1 U18699 ( .B1(n15438), .B2(n20574), .A(n15184), .ZN(P1_U2984) );
  OAI21_X1 U18700 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15192) );
  INV_X1 U18701 ( .A(n15188), .ZN(n15189) );
  NOR2_X1 U18702 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  XNOR2_X1 U18703 ( .A(n15192), .B(n15191), .ZN(n15448) );
  NAND2_X1 U18704 ( .A1(n20731), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U18705 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15193) );
  OAI211_X1 U18706 ( .C1(n20742), .C2(n15194), .A(n15440), .B(n15193), .ZN(
        n15195) );
  AOI21_X1 U18707 ( .B1(n15196), .B2(n20737), .A(n15195), .ZN(n15197) );
  OAI21_X1 U18708 ( .B1(n15448), .B2(n20574), .A(n15197), .ZN(P1_U2985) );
  INV_X1 U18709 ( .A(n15198), .ZN(n15199) );
  AOI22_X1 U18710 ( .A1(n15229), .A2(n15200), .B1(n15220), .B2(n15199), .ZN(
        n15212) );
  INV_X1 U18711 ( .A(n15202), .ZN(n15201) );
  AOI21_X1 U18712 ( .B1(n15220), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15201), .ZN(n15211) );
  NAND2_X1 U18713 ( .A1(n15212), .A2(n15211), .ZN(n15210) );
  NAND2_X1 U18714 ( .A1(n15210), .A2(n15202), .ZN(n15203) );
  NAND2_X1 U18715 ( .A1(n15458), .A2(n20738), .ZN(n15208) );
  OR2_X1 U18716 ( .A1(n20786), .A2(n21537), .ZN(n15449) );
  INV_X1 U18717 ( .A(n15449), .ZN(n15206) );
  NOR2_X1 U18718 ( .A1(n20742), .A2(n15204), .ZN(n15205) );
  AOI211_X1 U18719 ( .C1(n20732), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15206), .B(n15205), .ZN(n15207) );
  OAI211_X1 U18720 ( .C1(n20797), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        P1_U2986) );
  OAI21_X1 U18721 ( .B1(n15212), .B2(n15211), .A(n15210), .ZN(n15213) );
  INV_X1 U18722 ( .A(n15213), .ZN(n15474) );
  NOR2_X1 U18723 ( .A1(n20786), .A2(n15214), .ZN(n15468) );
  AOI21_X1 U18724 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15468), .ZN(n15215) );
  OAI21_X1 U18725 ( .B1(n20742), .B2(n15216), .A(n15215), .ZN(n15217) );
  AOI21_X1 U18726 ( .B1(n15218), .B2(n20737), .A(n15217), .ZN(n15219) );
  OAI21_X1 U18727 ( .B1(n15474), .B2(n20574), .A(n15219), .ZN(P1_U2987) );
  NOR2_X1 U18728 ( .A1(n15220), .A2(n15493), .ZN(n15221) );
  NOR3_X1 U18729 ( .A1(n10278), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15239), .ZN(n15232) );
  AOI21_X1 U18730 ( .B1(n15229), .B2(n15221), .A(n15232), .ZN(n15222) );
  XOR2_X1 U18731 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15222), .Z(
        n15483) );
  OR2_X1 U18732 ( .A1(n20786), .A2(n21534), .ZN(n15475) );
  NAND2_X1 U18733 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15223) );
  OAI211_X1 U18734 ( .C1(n20742), .C2(n15224), .A(n15475), .B(n15223), .ZN(
        n15225) );
  AOI21_X1 U18735 ( .B1(n15226), .B2(n20737), .A(n15225), .ZN(n15227) );
  OAI21_X1 U18736 ( .B1(n15483), .B2(n20574), .A(n15227), .ZN(P1_U2988) );
  NOR2_X1 U18737 ( .A1(n15228), .A2(n15493), .ZN(n15231) );
  XNOR2_X1 U18738 ( .A(n15229), .B(n15493), .ZN(n15230) );
  MUX2_X1 U18739 ( .A(n15231), .B(n15230), .S(n15239), .Z(n15233) );
  NOR2_X1 U18740 ( .A1(n15233), .A2(n15232), .ZN(n15497) );
  NAND2_X1 U18741 ( .A1(n20731), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15492) );
  NAND2_X1 U18742 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15234) );
  OAI211_X1 U18743 ( .C1(n20742), .C2(n15235), .A(n15492), .B(n15234), .ZN(
        n15236) );
  AOI21_X1 U18744 ( .B1(n15237), .B2(n20737), .A(n15236), .ZN(n15238) );
  OAI21_X1 U18745 ( .B1(n15497), .B2(n20574), .A(n15238), .ZN(P1_U2989) );
  XNOR2_X1 U18746 ( .A(n15239), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15240) );
  XNOR2_X1 U18747 ( .A(n15149), .B(n15240), .ZN(n15506) );
  NOR2_X1 U18748 ( .A1(n20786), .A2(n15241), .ZN(n15498) );
  AOI21_X1 U18749 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15498), .ZN(n15242) );
  OAI21_X1 U18750 ( .B1(n20742), .B2(n15243), .A(n15242), .ZN(n15244) );
  AOI21_X1 U18751 ( .B1(n15245), .B2(n20737), .A(n15244), .ZN(n15246) );
  OAI21_X1 U18752 ( .B1(n15506), .B2(n20574), .A(n15246), .ZN(P1_U2990) );
  XNOR2_X1 U18753 ( .A(n15247), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15248) );
  XNOR2_X1 U18754 ( .A(n15249), .B(n15248), .ZN(n15523) );
  INV_X1 U18755 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15250) );
  NOR2_X1 U18756 ( .A1(n20786), .A2(n15250), .ZN(n15508) );
  AOI21_X1 U18757 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15508), .ZN(n15251) );
  OAI21_X1 U18758 ( .B1(n20742), .B2(n15252), .A(n15251), .ZN(n15253) );
  AOI21_X1 U18759 ( .B1(n15254), .B2(n20737), .A(n15253), .ZN(n15255) );
  OAI21_X1 U18760 ( .B1(n15523), .B2(n20574), .A(n15255), .ZN(P1_U2991) );
  NAND2_X1 U18761 ( .A1(n15257), .A2(n15256), .ZN(n15259) );
  XOR2_X1 U18762 ( .A(n15259), .B(n15258), .Z(n15529) );
  INV_X1 U18763 ( .A(n20604), .ZN(n15262) );
  INV_X1 U18764 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20609) );
  NOR2_X1 U18765 ( .A1(n20786), .A2(n20609), .ZN(n15525) );
  AOI21_X1 U18766 ( .B1(n20732), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n15525), .ZN(n15260) );
  OAI21_X1 U18767 ( .B1(n20742), .B2(n20602), .A(n15260), .ZN(n15261) );
  AOI21_X1 U18768 ( .B1(n15262), .B2(n20737), .A(n15261), .ZN(n15263) );
  OAI21_X1 U18769 ( .B1(n15529), .B2(n20574), .A(n15263), .ZN(P1_U2992) );
  XNOR2_X1 U18770 ( .A(n15264), .B(n15534), .ZN(n15265) );
  XNOR2_X1 U18771 ( .A(n15266), .B(n15265), .ZN(n15538) );
  NAND2_X1 U18772 ( .A1(n15538), .A2(n20738), .ZN(n15270) );
  INV_X1 U18773 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n15267) );
  NOR2_X1 U18774 ( .A1(n20786), .A2(n15267), .ZN(n15531) );
  NOR2_X1 U18775 ( .A1(n20742), .A2(n20623), .ZN(n15268) );
  AOI211_X1 U18776 ( .C1(n20732), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15531), .B(n15268), .ZN(n15269) );
  OAI211_X1 U18777 ( .C1(n20797), .C2(n20610), .A(n15270), .B(n15269), .ZN(
        P1_U2993) );
  XNOR2_X1 U18778 ( .A(n15271), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20735) );
  INV_X1 U18779 ( .A(n15272), .ZN(n20734) );
  NOR2_X1 U18780 ( .A1(n20735), .A2(n20734), .ZN(n20733) );
  AOI21_X1 U18781 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15271), .A(
        n20733), .ZN(n15276) );
  XNOR2_X1 U18782 ( .A(n15274), .B(n15273), .ZN(n15275) );
  XNOR2_X1 U18783 ( .A(n15276), .B(n15275), .ZN(n15548) );
  INV_X1 U18784 ( .A(n15277), .ZN(n20660) );
  NAND2_X1 U18785 ( .A1(n20731), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15542) );
  NAND2_X1 U18786 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15278) );
  OAI211_X1 U18787 ( .C1(n20742), .C2(n20636), .A(n15542), .B(n15278), .ZN(
        n15279) );
  AOI21_X1 U18788 ( .B1(n20660), .B2(n20737), .A(n15279), .ZN(n15280) );
  OAI21_X1 U18789 ( .B1(n15548), .B2(n20574), .A(n15280), .ZN(P1_U2994) );
  OAI21_X1 U18790 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n20757) );
  NAND2_X1 U18791 ( .A1(n20731), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20753) );
  NAND2_X1 U18792 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15284) );
  OAI211_X1 U18793 ( .C1(n20742), .C2(n15285), .A(n20753), .B(n15284), .ZN(
        n15286) );
  AOI21_X1 U18794 ( .B1(n15287), .B2(n20737), .A(n15286), .ZN(n15288) );
  OAI21_X1 U18795 ( .B1(n20757), .B2(n20574), .A(n15288), .ZN(P1_U2996) );
  AOI22_X1 U18796 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20731), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15289) );
  OAI21_X1 U18797 ( .B1(n20742), .B2(n15290), .A(n15289), .ZN(n15294) );
  INV_X1 U18798 ( .A(n20776), .ZN(n15292) );
  NOR3_X1 U18799 ( .A1(n20771), .A2(n15292), .A3(n20574), .ZN(n15293) );
  AOI211_X1 U18800 ( .C1(n20737), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        n15296) );
  INV_X1 U18801 ( .A(n15296), .ZN(P1_U2997) );
  INV_X1 U18802 ( .A(n15297), .ZN(n15301) );
  NOR3_X1 U18803 ( .A1(n15308), .A2(n15299), .A3(n15298), .ZN(n15300) );
  AOI211_X1 U18804 ( .C1(n15306), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15301), .B(n15300), .ZN(n15303) );
  NAND2_X1 U18805 ( .A1(n10551), .A2(n20756), .ZN(n15302) );
  OAI211_X1 U18806 ( .C1(n15304), .C2(n20784), .A(n15303), .B(n15302), .ZN(
        P1_U3003) );
  AOI21_X1 U18807 ( .B1(n15306), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15305), .ZN(n15307) );
  OAI21_X1 U18808 ( .B1(n15308), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15307), .ZN(n15309) );
  AOI21_X1 U18809 ( .B1(n15310), .B2(n20756), .A(n15309), .ZN(n15311) );
  OAI21_X1 U18810 ( .B1(n15312), .B2(n20784), .A(n15311), .ZN(P1_U3004) );
  INV_X1 U18811 ( .A(n15344), .ZN(n15331) );
  AOI21_X1 U18812 ( .B1(n15331), .B2(n10455), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15314) );
  NOR2_X1 U18813 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  AOI211_X1 U18814 ( .C1(n15317), .C2(n20756), .A(n15316), .B(n15315), .ZN(
        n15318) );
  OAI21_X1 U18815 ( .B1(n15319), .B2(n20784), .A(n15318), .ZN(P1_U3005) );
  NAND2_X1 U18816 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15321) );
  OAI21_X1 U18817 ( .B1(n15344), .B2(n15321), .A(n15320), .ZN(n15325) );
  NAND2_X1 U18818 ( .A1(n15332), .A2(n15322), .ZN(n15324) );
  AOI21_X1 U18819 ( .B1(n15325), .B2(n15324), .A(n15323), .ZN(n15328) );
  NAND2_X1 U18820 ( .A1(n15326), .A2(n20756), .ZN(n15327) );
  OAI211_X1 U18821 ( .C1(n15329), .C2(n20784), .A(n15328), .B(n15327), .ZN(
        P1_U3006) );
  NAND3_X1 U18822 ( .A1(n15331), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15330), .ZN(n15336) );
  INV_X1 U18823 ( .A(n15332), .ZN(n15342) );
  AOI21_X1 U18824 ( .B1(n20766), .B2(n20744), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15333) );
  OAI21_X1 U18825 ( .B1(n15342), .B2(n15333), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15334) );
  NAND3_X1 U18826 ( .A1(n15336), .A2(n15335), .A3(n15334), .ZN(n15337) );
  AOI21_X1 U18827 ( .B1(n15338), .B2(n20756), .A(n15337), .ZN(n15339) );
  OAI21_X1 U18828 ( .B1(n15340), .B2(n20784), .A(n15339), .ZN(P1_U3007) );
  AOI21_X1 U18829 ( .B1(n15342), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15341), .ZN(n15343) );
  OAI21_X1 U18830 ( .B1(n15344), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15343), .ZN(n15345) );
  AOI21_X1 U18831 ( .B1(n15346), .B2(n20756), .A(n15345), .ZN(n15347) );
  OAI21_X1 U18832 ( .B1(n15348), .B2(n20784), .A(n15347), .ZN(P1_U3008) );
  NAND2_X1 U18833 ( .A1(n15349), .A2(n20760), .ZN(n15355) );
  INV_X1 U18834 ( .A(n15350), .ZN(n15361) );
  XNOR2_X1 U18835 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U18836 ( .A1(n15358), .A2(n15351), .ZN(n15352) );
  AOI211_X1 U18837 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15361), .A(
        n15353), .B(n15352), .ZN(n15354) );
  OAI211_X1 U18838 ( .C1(n20788), .C2(n15356), .A(n15355), .B(n15354), .ZN(
        P1_U3009) );
  NAND2_X1 U18839 ( .A1(n15357), .A2(n20760), .ZN(n15363) );
  NOR2_X1 U18840 ( .A1(n15358), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15359) );
  AOI211_X1 U18841 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15361), .A(
        n15360), .B(n15359), .ZN(n15362) );
  OAI211_X1 U18842 ( .C1(n20788), .C2(n15364), .A(n15363), .B(n15362), .ZN(
        P1_U3010) );
  NAND2_X1 U18843 ( .A1(n15365), .A2(n20760), .ZN(n15382) );
  INV_X1 U18844 ( .A(n15366), .ZN(n15399) );
  NAND2_X1 U18845 ( .A1(n15394), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15398) );
  INV_X1 U18846 ( .A(n15398), .ZN(n15367) );
  NAND2_X1 U18847 ( .A1(n15399), .A2(n15367), .ZN(n15369) );
  NAND2_X1 U18848 ( .A1(n15369), .A2(n15368), .ZN(n15404) );
  INV_X1 U18849 ( .A(n15404), .ZN(n15376) );
  NAND2_X1 U18850 ( .A1(n15370), .A2(n11842), .ZN(n15384) );
  INV_X1 U18851 ( .A(n15371), .ZN(n15373) );
  OAI22_X1 U18852 ( .A1(n20744), .A2(n15373), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15372), .ZN(n15374) );
  AOI211_X1 U18853 ( .C1(n15375), .C2(n15510), .A(n15460), .B(n15374), .ZN(
        n15385) );
  OAI21_X1 U18854 ( .B1(n15376), .B2(n15384), .A(n15385), .ZN(n15380) );
  NOR2_X1 U18855 ( .A1(n15377), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15378) );
  AOI211_X1 U18856 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15380), .A(
        n15379), .B(n15378), .ZN(n15381) );
  OAI211_X1 U18857 ( .C1(n20788), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        P1_U3011) );
  INV_X1 U18858 ( .A(n15384), .ZN(n15389) );
  NOR2_X1 U18859 ( .A1(n15385), .A2(n11842), .ZN(n15386) );
  AOI211_X1 U18860 ( .C1(n15389), .C2(n15388), .A(n15387), .B(n15386), .ZN(
        n15392) );
  NAND2_X1 U18861 ( .A1(n15390), .A2(n20756), .ZN(n15391) );
  OAI211_X1 U18862 ( .C1(n15393), .C2(n20784), .A(n15392), .B(n15391), .ZN(
        P1_U3012) );
  NAND2_X1 U18863 ( .A1(n15394), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15395) );
  NAND2_X1 U18864 ( .A1(n15396), .A2(n15395), .ZN(n15451) );
  INV_X1 U18865 ( .A(n15397), .ZN(n15403) );
  NAND2_X1 U18866 ( .A1(n15399), .A2(n15398), .ZN(n15402) );
  INV_X1 U18867 ( .A(n15445), .ZN(n15400) );
  NAND2_X1 U18868 ( .A1(n20770), .A2(n15400), .ZN(n15401) );
  AND4_X1 U18869 ( .A1(n15451), .A2(n15403), .A3(n15402), .A4(n15401), .ZN(
        n15454) );
  NAND2_X1 U18870 ( .A1(n15404), .A2(n15453), .ZN(n15450) );
  AND2_X1 U18871 ( .A1(n15454), .A2(n15450), .ZN(n15439) );
  NAND2_X1 U18872 ( .A1(n20782), .A2(n15444), .ZN(n15405) );
  NAND2_X1 U18873 ( .A1(n15439), .A2(n15405), .ZN(n15436) );
  AND2_X1 U18874 ( .A1(n20782), .A2(n15406), .ZN(n15407) );
  OR2_X1 U18875 ( .A1(n15436), .A2(n15407), .ZN(n15418) );
  AND2_X1 U18876 ( .A1(n15408), .A2(n11843), .ZN(n15409) );
  AOI211_X1 U18877 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15418), .A(
        n15410), .B(n15409), .ZN(n15413) );
  NAND2_X1 U18878 ( .A1(n15411), .A2(n20756), .ZN(n15412) );
  OAI211_X1 U18879 ( .C1(n15414), .C2(n20784), .A(n15413), .B(n15412), .ZN(
        P1_U3013) );
  AOI21_X1 U18880 ( .B1(n15416), .B2(n20756), .A(n15415), .ZN(n15420) );
  NAND2_X1 U18881 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15422) );
  OAI21_X1 U18882 ( .B1(n15431), .B2(n15422), .A(n21716), .ZN(n15417) );
  NAND2_X1 U18883 ( .A1(n15418), .A2(n15417), .ZN(n15419) );
  OAI211_X1 U18884 ( .C1(n15421), .C2(n20784), .A(n15420), .B(n15419), .ZN(
        P1_U3014) );
  INV_X1 U18885 ( .A(n15422), .ZN(n15423) );
  NOR3_X1 U18886 ( .A1(n15431), .A2(n15424), .A3(n15423), .ZN(n15426) );
  NOR2_X1 U18887 ( .A1(n15426), .A2(n15425), .ZN(n15429) );
  AOI22_X1 U18888 ( .A1(n15427), .A2(n20756), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15436), .ZN(n15428) );
  OAI211_X1 U18889 ( .C1(n15430), .C2(n20784), .A(n15429), .B(n15428), .ZN(
        P1_U3015) );
  NOR2_X1 U18890 ( .A1(n15431), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15435) );
  OAI21_X1 U18891 ( .B1(n15433), .B2(n20788), .A(n15432), .ZN(n15434) );
  AOI211_X1 U18892 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15436), .A(
        n15435), .B(n15434), .ZN(n15437) );
  OAI21_X1 U18893 ( .B1(n15438), .B2(n20784), .A(n15437), .ZN(P1_U3016) );
  INV_X1 U18894 ( .A(n15439), .ZN(n15443) );
  OAI21_X1 U18895 ( .B1(n15441), .B2(n20788), .A(n15440), .ZN(n15442) );
  AOI21_X1 U18896 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15443), .A(
        n15442), .ZN(n15447) );
  NAND2_X1 U18897 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15486) );
  NAND2_X1 U18898 ( .A1(n15516), .A2(n20744), .ZN(n15543) );
  NAND4_X1 U18899 ( .A1(n15543), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15445), .A4(n15444), .ZN(n15446) );
  OAI211_X1 U18900 ( .C1(n15448), .C2(n20784), .A(n15447), .B(n15446), .ZN(
        P1_U3017) );
  OAI211_X1 U18901 ( .C1(n15452), .C2(n15451), .A(n15450), .B(n15449), .ZN(
        n15457) );
  OAI22_X1 U18902 ( .A1(n15455), .A2(n20788), .B1(n15454), .B2(n15453), .ZN(
        n15456) );
  AOI211_X1 U18903 ( .C1(n15458), .C2(n20760), .A(n15457), .B(n15456), .ZN(
        n15459) );
  INV_X1 U18904 ( .A(n15459), .ZN(P1_U3018) );
  INV_X1 U18905 ( .A(n15460), .ZN(n15488) );
  INV_X1 U18906 ( .A(n15461), .ZN(n15464) );
  INV_X1 U18907 ( .A(n15462), .ZN(n15463) );
  AOI22_X1 U18908 ( .A1(n15510), .A2(n15464), .B1(n20770), .B2(n15463), .ZN(
        n15465) );
  NAND2_X1 U18909 ( .A1(n15488), .A2(n15465), .ZN(n15481) );
  NOR2_X1 U18910 ( .A1(n15466), .A2(n20788), .ZN(n15467) );
  AOI211_X1 U18911 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15481), .A(
        n15468), .B(n15467), .ZN(n15473) );
  NOR2_X1 U18912 ( .A1(n20766), .A2(n15469), .ZN(n15471) );
  NAND2_X1 U18913 ( .A1(n15543), .A2(n15511), .ZN(n15530) );
  OAI21_X1 U18914 ( .B1(n15530), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15470) );
  OAI211_X1 U18915 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15471), .A(
        n15470), .B(n15477), .ZN(n15472) );
  OAI211_X1 U18916 ( .C1(n15474), .C2(n20784), .A(n15473), .B(n15472), .ZN(
        P1_U3019) );
  OAI21_X1 U18917 ( .B1(n15476), .B2(n20788), .A(n15475), .ZN(n15480) );
  INV_X1 U18918 ( .A(n15477), .ZN(n15478) );
  NOR3_X1 U18919 ( .A1(n15530), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15478), .ZN(n15479) );
  AOI211_X1 U18920 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15481), .A(
        n15480), .B(n15479), .ZN(n15482) );
  OAI21_X1 U18921 ( .B1(n15483), .B2(n20784), .A(n15482), .ZN(P1_U3020) );
  XNOR2_X1 U18922 ( .A(n15493), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15495) );
  INV_X1 U18923 ( .A(n15485), .ZN(n15484) );
  NOR2_X1 U18924 ( .A1(n15530), .A2(n15484), .ZN(n15504) );
  NAND2_X1 U18925 ( .A1(n15511), .A2(n15485), .ZN(n15489) );
  NAND2_X1 U18926 ( .A1(n15510), .A2(n15486), .ZN(n15487) );
  NAND2_X1 U18927 ( .A1(n15488), .A2(n15487), .ZN(n20768) );
  AOI21_X1 U18928 ( .B1(n20782), .B2(n15489), .A(n20768), .ZN(n15501) );
  NAND2_X1 U18929 ( .A1(n15490), .A2(n20756), .ZN(n15491) );
  OAI211_X1 U18930 ( .C1(n15501), .C2(n15493), .A(n15492), .B(n15491), .ZN(
        n15494) );
  AOI21_X1 U18931 ( .B1(n15495), .B2(n15504), .A(n15494), .ZN(n15496) );
  OAI21_X1 U18932 ( .B1(n15497), .B2(n20784), .A(n15496), .ZN(P1_U3021) );
  AOI21_X1 U18933 ( .B1(n15499), .B2(n20756), .A(n15498), .ZN(n15500) );
  OAI21_X1 U18934 ( .B1(n15501), .B2(n15503), .A(n15500), .ZN(n15502) );
  AOI21_X1 U18935 ( .B1(n15504), .B2(n15503), .A(n15502), .ZN(n15505) );
  OAI21_X1 U18936 ( .B1(n15506), .B2(n20784), .A(n15505), .ZN(P1_U3022) );
  NOR4_X1 U18937 ( .A1(n15530), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n15534), .A4(n15519), .ZN(n15507) );
  AOI211_X1 U18938 ( .C1(n20756), .C2(n15509), .A(n15508), .B(n15507), .ZN(
        n15522) );
  NAND2_X1 U18939 ( .A1(n15510), .A2(n20745), .ZN(n15514) );
  INV_X1 U18940 ( .A(n15511), .ZN(n15512) );
  NAND2_X1 U18941 ( .A1(n20770), .A2(n15512), .ZN(n15513) );
  NAND2_X1 U18942 ( .A1(n15514), .A2(n15513), .ZN(n15515) );
  OR2_X1 U18943 ( .A1(n20768), .A2(n15515), .ZN(n15546) );
  NOR2_X1 U18944 ( .A1(n15516), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15517) );
  NOR2_X1 U18945 ( .A1(n15546), .A2(n15517), .ZN(n15535) );
  OAI21_X1 U18946 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15518), .A(
        n15535), .ZN(n15526) );
  NAND2_X1 U18947 ( .A1(n15519), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15520) );
  NOR2_X1 U18948 ( .A1(n15530), .A2(n15520), .ZN(n15524) );
  OAI21_X1 U18949 ( .B1(n15526), .B2(n15524), .A(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15521) );
  OAI211_X1 U18950 ( .C1(n15523), .C2(n20784), .A(n15522), .B(n15521), .ZN(
        P1_U3023) );
  AOI211_X1 U18951 ( .C1(n20756), .C2(n20597), .A(n15525), .B(n15524), .ZN(
        n15528) );
  NAND2_X1 U18952 ( .A1(n15526), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15527) );
  OAI211_X1 U18953 ( .C1(n15529), .C2(n20784), .A(n15528), .B(n15527), .ZN(
        P1_U3024) );
  NOR2_X1 U18954 ( .A1(n15530), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15537) );
  INV_X1 U18955 ( .A(n20614), .ZN(n15532) );
  AOI21_X1 U18956 ( .B1(n20756), .B2(n15532), .A(n15531), .ZN(n15533) );
  OAI21_X1 U18957 ( .B1(n15535), .B2(n15534), .A(n15533), .ZN(n15536) );
  AOI211_X1 U18958 ( .C1(n15538), .C2(n20760), .A(n15537), .B(n15536), .ZN(
        n15539) );
  INV_X1 U18959 ( .A(n15539), .ZN(P1_U3025) );
  OAI21_X1 U18960 ( .B1(n15541), .B2(n15540), .A(n14931), .ZN(n20624) );
  OAI21_X1 U18961 ( .B1(n20788), .B2(n20624), .A(n15542), .ZN(n15545) );
  NAND2_X1 U18962 ( .A1(n15543), .A2(n20743), .ZN(n20758) );
  NOR3_X1 U18963 ( .A1(n20758), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n20745), .ZN(n15544) );
  AOI211_X1 U18964 ( .C1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15546), .A(
        n15545), .B(n15544), .ZN(n15547) );
  OAI21_X1 U18965 ( .B1(n15548), .B2(n20784), .A(n15547), .ZN(P1_U3026) );
  NAND2_X1 U18966 ( .A1(n15549), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15552) );
  NAND2_X1 U18967 ( .A1(n15552), .A2(n9585), .ZN(n21432) );
  NOR2_X1 U18968 ( .A1(n15549), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15550) );
  OAI22_X1 U18969 ( .A1(n21432), .A2(n15550), .B1(n14245), .B2(n15558), .ZN(
        n15551) );
  MUX2_X1 U18970 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15551), .S(
        n20795), .Z(P1_U3477) );
  INV_X1 U18971 ( .A(n15552), .ZN(n15557) );
  NAND2_X1 U18972 ( .A1(n15557), .A2(n9585), .ZN(n21241) );
  MUX2_X1 U18973 ( .A(n21241), .B(n21432), .S(n20799), .Z(n15553) );
  OAI21_X1 U18974 ( .B1(n21279), .B2(n15558), .A(n15553), .ZN(n15554) );
  MUX2_X1 U18975 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15554), .S(
        n20795), .Z(P1_U3476) );
  NOR2_X1 U18976 ( .A1(n15549), .A2(n21373), .ZN(n15556) );
  AOI22_X1 U18977 ( .A1(n15557), .A2(n21088), .B1(n21372), .B2(n15556), .ZN(
        n21013) );
  NOR2_X1 U18978 ( .A1(n21013), .A2(n21233), .ZN(n15561) );
  OAI22_X1 U18979 ( .A1(n15561), .A2(n15560), .B1(n15559), .B2(n15558), .ZN(
        n15562) );
  MUX2_X1 U18980 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15562), .S(
        n20795), .Z(P1_U3475) );
  INV_X1 U18981 ( .A(n14060), .ZN(n15565) );
  INV_X1 U18982 ( .A(n15563), .ZN(n15564) );
  NAND2_X1 U18983 ( .A1(n15565), .A2(n15564), .ZN(n15571) );
  OAI21_X1 U18984 ( .B1(n15567), .B2(n15571), .A(n15566), .ZN(n15568) );
  AOI21_X1 U18985 ( .B1(n21375), .B2(n15569), .A(n15568), .ZN(n17283) );
  INV_X1 U18986 ( .A(n15570), .ZN(n15577) );
  INV_X1 U18987 ( .A(n15571), .ZN(n15574) );
  AOI22_X1 U18988 ( .A1(n15575), .A2(n15574), .B1(n15573), .B2(n15572), .ZN(
        n15576) );
  OAI21_X1 U18989 ( .B1(n17283), .B2(n15577), .A(n15576), .ZN(n15579) );
  MUX2_X1 U18990 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15579), .S(
        n15578), .Z(P1_U3473) );
  INV_X1 U18991 ( .A(HOLD), .ZN(n21512) );
  OAI211_X1 U18992 ( .C1(n21520), .C2(n21512), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15581) );
  NAND3_X1 U18993 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n21520), .ZN(
        n15580) );
  NAND2_X1 U18994 ( .A1(n17309), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21510) );
  NAND4_X1 U18995 ( .A1(n15582), .A2(n15581), .A3(n15580), .A4(n21510), .ZN(
        P1_U3195) );
  INV_X1 U18996 ( .A(n15583), .ZN(n15584) );
  INV_X1 U18997 ( .A(n16723), .ZN(n16219) );
  INV_X1 U18998 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18999 ( .A1(n19737), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19746), .ZN(n15588) );
  OAI21_X1 U19000 ( .B1(n15589), .B2(n19767), .A(n15588), .ZN(n15593) );
  NOR2_X1 U19001 ( .A1(n16731), .A2(n15954), .ZN(n15592) );
  INV_X1 U19002 ( .A(n16435), .ZN(n15596) );
  AOI21_X1 U19003 ( .B1(n15595), .B2(n15596), .A(n19734), .ZN(n15597) );
  OAI21_X1 U19004 ( .B1(n15597), .B2(n15952), .A(n13091), .ZN(n15598) );
  OAI211_X1 U19005 ( .C1(n16219), .C2(n15945), .A(n15599), .B(n15598), .ZN(
        P2_U2826) );
  OAI21_X1 U19006 ( .B1(n9675), .B2(n15601), .A(n15600), .ZN(n16739) );
  NOR2_X1 U19007 ( .A1(n15602), .A2(n15603), .ZN(n15604) );
  OR2_X1 U19008 ( .A1(n15590), .A2(n15604), .ZN(n16738) );
  INV_X1 U19009 ( .A(n16738), .ZN(n16336) );
  OAI22_X1 U19010 ( .A1(n19748), .A2(n16444), .B1(n15955), .B2(n15605), .ZN(
        n15606) );
  AOI21_X1 U19011 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15606), .ZN(n15607) );
  OAI21_X1 U19012 ( .B1(n15608), .B2(n15941), .A(n15607), .ZN(n15609) );
  AOI21_X1 U19013 ( .B1(n16336), .B2(n19760), .A(n15609), .ZN(n15614) );
  INV_X1 U19014 ( .A(n16445), .ZN(n15611) );
  AOI21_X1 U19015 ( .B1(n15610), .B2(n15611), .A(n19734), .ZN(n15612) );
  OAI21_X1 U19016 ( .B1(n15612), .B2(n15952), .A(n15595), .ZN(n15613) );
  OAI211_X1 U19017 ( .C1(n16739), .C2(n15945), .A(n15614), .B(n15613), .ZN(
        P2_U2827) );
  NOR2_X1 U19018 ( .A1(n9622), .A2(n15615), .ZN(n15616) );
  AND2_X1 U19019 ( .A1(n15617), .A2(n15618), .ZN(n15619) );
  NOR2_X1 U19020 ( .A1(n15602), .A2(n15619), .ZN(n16747) );
  INV_X1 U19021 ( .A(n16454), .ZN(n15621) );
  AOI21_X1 U19022 ( .B1(n15620), .B2(n15621), .A(n19734), .ZN(n15622) );
  OAI21_X1 U19023 ( .B1(n15622), .B2(n15952), .A(n15610), .ZN(n15626) );
  INV_X1 U19024 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20476) );
  OAI22_X1 U19025 ( .A1(n19748), .A2(n20476), .B1(n15955), .B2(n15623), .ZN(
        n15624) );
  AOI21_X1 U19026 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15624), .ZN(n15625) );
  OAI211_X1 U19027 ( .C1(n15941), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        n15628) );
  AOI21_X1 U19028 ( .B1(n16747), .B2(n19760), .A(n15628), .ZN(n15629) );
  OAI21_X1 U19029 ( .B1(n16748), .B2(n15945), .A(n15629), .ZN(P2_U2828) );
  NOR2_X1 U19030 ( .A1(n9617), .A2(n15630), .ZN(n15631) );
  NAND2_X1 U19031 ( .A1(n15633), .A2(n15632), .ZN(n15634) );
  NAND2_X1 U19032 ( .A1(n15617), .A2(n15634), .ZN(n16762) );
  INV_X1 U19033 ( .A(n16762), .ZN(n16352) );
  INV_X1 U19034 ( .A(n16465), .ZN(n15636) );
  AOI21_X1 U19035 ( .B1(n15635), .B2(n15636), .A(n19734), .ZN(n15637) );
  OAI21_X1 U19036 ( .B1(n15637), .B2(n15952), .A(n15620), .ZN(n15640) );
  INV_X1 U19037 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20473) );
  OAI22_X1 U19038 ( .A1(n19748), .A2(n20473), .B1(n15955), .B2(n16240), .ZN(
        n15638) );
  AOI21_X1 U19039 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15638), .ZN(n15639) );
  OAI211_X1 U19040 ( .C1(n15941), .C2(n15641), .A(n15640), .B(n15639), .ZN(
        n15642) );
  AOI21_X1 U19041 ( .B1(n16352), .B2(n19760), .A(n15642), .ZN(n15643) );
  OAI21_X1 U19042 ( .B1(n16752), .B2(n15945), .A(n15643), .ZN(P2_U2829) );
  XNOR2_X1 U19043 ( .A(n15644), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n15652) );
  INV_X1 U19044 ( .A(n15646), .ZN(n15647) );
  AOI21_X1 U19045 ( .B1(n15645), .B2(n15647), .A(n19734), .ZN(n15648) );
  OAI21_X1 U19046 ( .B1(n15648), .B2(n15952), .A(n15635), .ZN(n15651) );
  OAI22_X1 U19047 ( .A1(n19748), .A2(n20471), .B1(n15955), .B2(n21691), .ZN(
        n15649) );
  AOI21_X1 U19048 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15649), .ZN(n15650) );
  OAI211_X1 U19049 ( .C1(n15652), .C2(n15941), .A(n15651), .B(n15650), .ZN(
        n15653) );
  AOI21_X1 U19050 ( .B1(n16244), .B2(n19761), .A(n15653), .ZN(n15654) );
  OAI21_X1 U19051 ( .B1(n16358), .B2(n15954), .A(n15654), .ZN(P2_U2830) );
  INV_X1 U19052 ( .A(n13142), .ZN(n15656) );
  AOI21_X1 U19053 ( .B1(n15657), .B2(n15655), .A(n15656), .ZN(n16777) );
  AND2_X1 U19054 ( .A1(n15658), .A2(n15659), .ZN(n15660) );
  OR2_X1 U19055 ( .A1(n15660), .A2(n13144), .ZN(n16775) );
  NAND2_X1 U19056 ( .A1(n19746), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U19057 ( .A1(n19737), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15661) );
  OAI211_X1 U19058 ( .C1(n19767), .C2(n15663), .A(n15662), .B(n15661), .ZN(
        n15664) );
  AOI21_X1 U19059 ( .B1(n15665), .B2(n19750), .A(n15664), .ZN(n15670) );
  INV_X1 U19060 ( .A(n16480), .ZN(n15667) );
  AOI21_X1 U19061 ( .B1(n15666), .B2(n15667), .A(n19734), .ZN(n15668) );
  OAI21_X1 U19062 ( .B1(n15668), .B2(n15952), .A(n15645), .ZN(n15669) );
  OAI211_X1 U19063 ( .C1(n16775), .C2(n15954), .A(n15670), .B(n15669), .ZN(
        n15671) );
  AOI21_X1 U19064 ( .B1(n16777), .B2(n19761), .A(n15671), .ZN(n15672) );
  INV_X1 U19065 ( .A(n15672), .ZN(P2_U2831) );
  OAI21_X1 U19066 ( .B1(n13015), .B2(n9755), .A(n15658), .ZN(n16787) );
  OAI21_X1 U19067 ( .B1(n15674), .B2(n15675), .A(n15655), .ZN(n16259) );
  INV_X1 U19068 ( .A(n16259), .ZN(n16789) );
  NAND2_X1 U19069 ( .A1(n16789), .A2(n19761), .ZN(n15686) );
  AOI22_X1 U19070 ( .A1(n19737), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19746), .ZN(n15676) );
  OAI21_X1 U19071 ( .B1(n15677), .B2(n19767), .A(n15676), .ZN(n15683) );
  INV_X1 U19072 ( .A(n15678), .ZN(n15679) );
  OAI21_X1 U19073 ( .B1(n15679), .B2(n16486), .A(n19757), .ZN(n15681) );
  INV_X1 U19074 ( .A(n15666), .ZN(n15680) );
  AOI21_X1 U19075 ( .B1(n10546), .B2(n15681), .A(n15680), .ZN(n15682) );
  AOI211_X1 U19076 ( .C1(n19750), .C2(n15684), .A(n15683), .B(n15682), .ZN(
        n15685) );
  OAI211_X1 U19077 ( .C1(n15954), .C2(n16787), .A(n15686), .B(n15685), .ZN(
        P2_U2832) );
  INV_X1 U19078 ( .A(n15687), .ZN(n15690) );
  INV_X1 U19079 ( .A(n15688), .ZN(n15689) );
  AOI21_X1 U19080 ( .B1(n15690), .B2(n15689), .A(n15674), .ZN(n16805) );
  OR2_X1 U19081 ( .A1(n15691), .A2(n15692), .ZN(n15693) );
  NAND2_X1 U19082 ( .A1(n15673), .A2(n15693), .ZN(n16803) );
  NOR2_X1 U19083 ( .A1(n16803), .A2(n15954), .ZN(n15703) );
  INV_X1 U19084 ( .A(n16498), .ZN(n15695) );
  AOI21_X1 U19085 ( .B1(n15694), .B2(n15695), .A(n19734), .ZN(n15696) );
  OAI21_X1 U19086 ( .B1(n15696), .B2(n15952), .A(n15678), .ZN(n15700) );
  OAI22_X1 U19087 ( .A1(n19748), .A2(n20466), .B1(n15955), .B2(n15697), .ZN(
        n15698) );
  AOI21_X1 U19088 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15698), .ZN(n15699) );
  OAI211_X1 U19089 ( .C1(n15941), .C2(n15701), .A(n15700), .B(n15699), .ZN(
        n15702) );
  AOI211_X1 U19090 ( .C1(n16805), .C2(n19761), .A(n15703), .B(n15702), .ZN(
        n15704) );
  INV_X1 U19091 ( .A(n15704), .ZN(P2_U2833) );
  AOI21_X1 U19092 ( .B1(n15705), .B2(n9615), .A(n15688), .ZN(n16818) );
  INV_X1 U19093 ( .A(n16818), .ZN(n16269) );
  INV_X1 U19094 ( .A(n15691), .ZN(n15708) );
  NAND2_X1 U19095 ( .A1(n13011), .A2(n15706), .ZN(n15707) );
  NAND2_X1 U19096 ( .A1(n15708), .A2(n15707), .ZN(n16815) );
  INV_X1 U19097 ( .A(n16815), .ZN(n15718) );
  INV_X1 U19098 ( .A(n16510), .ZN(n15710) );
  AOI21_X1 U19099 ( .B1(n15709), .B2(n15710), .A(n19734), .ZN(n15711) );
  OAI21_X1 U19100 ( .B1(n15711), .B2(n15952), .A(n15694), .ZN(n15715) );
  OAI22_X1 U19101 ( .A1(n19748), .A2(n20464), .B1(n15955), .B2(n15712), .ZN(
        n15713) );
  AOI21_X1 U19102 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15713), .ZN(n15714) );
  OAI211_X1 U19103 ( .C1(n15941), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        n15717) );
  AOI21_X1 U19104 ( .B1(n15718), .B2(n19760), .A(n15717), .ZN(n15719) );
  OAI21_X1 U19105 ( .B1(n16269), .B2(n15945), .A(n15719), .ZN(P2_U2834) );
  NAND2_X1 U19106 ( .A1(n15720), .A2(n15721), .ZN(n15722) );
  NAND2_X1 U19107 ( .A1(n15723), .A2(n15722), .ZN(n16823) );
  OR2_X1 U19108 ( .A1(n15739), .A2(n15724), .ZN(n15725) );
  NAND2_X1 U19109 ( .A1(n16829), .A2(n19761), .ZN(n15737) );
  AOI21_X1 U19110 ( .B1(n15726), .B2(n10398), .A(n19734), .ZN(n15728) );
  OAI21_X1 U19111 ( .B1(n15952), .B2(n15728), .A(n15727), .ZN(n15732) );
  OAI21_X1 U19112 ( .B1(n15955), .B2(n15729), .A(n17339), .ZN(n15730) );
  AOI21_X1 U19113 ( .B1(n19737), .B2(P2_REIP_REG_19__SCAN_IN), .A(n15730), 
        .ZN(n15731) );
  OAI211_X1 U19114 ( .C1(n19767), .C2(n15733), .A(n15732), .B(n15731), .ZN(
        n15734) );
  AOI21_X1 U19115 ( .B1(n19750), .B2(n15735), .A(n15734), .ZN(n15736) );
  OAI211_X1 U19116 ( .C1(n15954), .C2(n16823), .A(n15737), .B(n15736), .ZN(
        P2_U2836) );
  AND2_X1 U19117 ( .A1(n15756), .A2(n15738), .ZN(n15740) );
  OR2_X1 U19118 ( .A1(n15740), .A2(n15739), .ZN(n16839) );
  OR2_X1 U19119 ( .A1(n14418), .A2(n15741), .ZN(n15742) );
  AND2_X1 U19120 ( .A1(n15720), .A2(n15742), .ZN(n16836) );
  NAND2_X1 U19121 ( .A1(n15912), .A2(n15743), .ZN(n15746) );
  INV_X1 U19122 ( .A(n15743), .ZN(n15744) );
  AOI21_X1 U19123 ( .B1(n19757), .B2(n15744), .A(n15952), .ZN(n15745) );
  MUX2_X1 U19124 ( .A(n15746), .B(n15745), .S(n16534), .Z(n15750) );
  AOI21_X1 U19125 ( .B1(n19746), .B2(P2_EBX_REG_18__SCAN_IN), .A(n19745), .ZN(
        n15747) );
  OAI21_X1 U19126 ( .B1(n12853), .B2(n19748), .A(n15747), .ZN(n15748) );
  AOI21_X1 U19127 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15951), .A(
        n15748), .ZN(n15749) );
  OAI211_X1 U19128 ( .C1(n15751), .C2(n15941), .A(n15750), .B(n15749), .ZN(
        n15752) );
  AOI21_X1 U19129 ( .B1(n16836), .B2(n19760), .A(n15752), .ZN(n15753) );
  OAI21_X1 U19130 ( .B1(n16839), .B2(n15945), .A(n15753), .ZN(P2_U2837) );
  INV_X1 U19131 ( .A(n15756), .ZN(n15757) );
  AOI21_X1 U19132 ( .B1(n15758), .B2(n15755), .A(n15757), .ZN(n16540) );
  INV_X1 U19133 ( .A(n16540), .ZN(n16855) );
  AOI21_X1 U19134 ( .B1(n19757), .B2(n15759), .A(n15952), .ZN(n15762) );
  INV_X1 U19135 ( .A(n15759), .ZN(n15760) );
  NAND2_X1 U19136 ( .A1(n15912), .A2(n15760), .ZN(n15761) );
  MUX2_X1 U19137 ( .A(n15762), .B(n15761), .S(n16543), .Z(n15766) );
  AOI21_X1 U19138 ( .B1(n19746), .B2(P2_EBX_REG_17__SCAN_IN), .A(n19745), .ZN(
        n15763) );
  OAI21_X1 U19139 ( .B1(n20459), .B2(n19748), .A(n15763), .ZN(n15764) );
  AOI21_X1 U19140 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n15951), .A(
        n15764), .ZN(n15765) );
  OAI211_X1 U19141 ( .C1(n15941), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        n15768) );
  AOI21_X1 U19142 ( .B1(n16853), .B2(n19760), .A(n15768), .ZN(n15769) );
  OAI21_X1 U19143 ( .B1(n16855), .B2(n15945), .A(n15769), .ZN(P2_U2838) );
  AOI21_X1 U19144 ( .B1(n15770), .B2(n14395), .A(n15754), .ZN(n16549) );
  INV_X1 U19145 ( .A(n16549), .ZN(n16866) );
  AOI21_X1 U19146 ( .B1(n19757), .B2(n15771), .A(n15952), .ZN(n15773) );
  INV_X1 U19147 ( .A(n15771), .ZN(n15772) );
  NAND2_X1 U19148 ( .A1(n15912), .A2(n15772), .ZN(n15785) );
  MUX2_X1 U19149 ( .A(n15773), .B(n15785), .S(n16552), .Z(n15777) );
  NAND2_X1 U19150 ( .A1(n19746), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15774) );
  OAI211_X1 U19151 ( .C1(n19748), .C2(n20457), .A(n17339), .B(n15774), .ZN(
        n15775) );
  AOI21_X1 U19152 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15951), .A(
        n15775), .ZN(n15776) );
  OAI211_X1 U19153 ( .C1(n15941), .C2(n15778), .A(n15777), .B(n15776), .ZN(
        n15779) );
  AOI21_X1 U19154 ( .B1(n16864), .B2(n19760), .A(n15779), .ZN(n15780) );
  OAI21_X1 U19155 ( .B1(n16866), .B2(n15945), .A(n15780), .ZN(P2_U2839) );
  INV_X1 U19156 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20455) );
  AOI21_X1 U19157 ( .B1(n19746), .B2(P2_EBX_REG_15__SCAN_IN), .A(n19745), .ZN(
        n15781) );
  OAI21_X1 U19158 ( .B1(n20455), .B2(n19748), .A(n15781), .ZN(n15782) );
  AOI21_X1 U19159 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n15951), .A(
        n15782), .ZN(n15783) );
  OAI21_X1 U19160 ( .B1(n15784), .B2(n15941), .A(n15783), .ZN(n15788) );
  AOI21_X1 U19161 ( .B1(n10543), .B2(n15786), .A(n15785), .ZN(n15787) );
  AOI211_X1 U19162 ( .C1(n15952), .C2(n10543), .A(n15788), .B(n15787), .ZN(
        n15791) );
  INV_X1 U19163 ( .A(n16868), .ZN(n15789) );
  NAND2_X1 U19164 ( .A1(n15789), .A2(n19761), .ZN(n15790) );
  OAI211_X1 U19165 ( .C1(n15954), .C2(n16870), .A(n15791), .B(n15790), .ZN(
        P2_U2840) );
  NAND2_X1 U19166 ( .A1(n15792), .A2(n19750), .ZN(n15796) );
  OAI21_X1 U19167 ( .B1(n15955), .B2(n15793), .A(n17339), .ZN(n15794) );
  AOI21_X1 U19168 ( .B1(n19737), .B2(P2_REIP_REG_14__SCAN_IN), .A(n15794), 
        .ZN(n15795) );
  OAI211_X1 U19169 ( .C1(n19767), .C2(n16573), .A(n15796), .B(n15795), .ZN(
        n15802) );
  INV_X1 U19170 ( .A(n15798), .ZN(n15797) );
  NOR2_X1 U19171 ( .A1(n15965), .A2(n15797), .ZN(n15800) );
  OAI21_X1 U19172 ( .B1(n19734), .B2(n15798), .A(n10546), .ZN(n15799) );
  MUX2_X1 U19173 ( .A(n15800), .B(n15799), .S(n16575), .Z(n15801) );
  AOI211_X1 U19174 ( .C1(n19760), .C2(n16881), .A(n15802), .B(n15801), .ZN(
        n15803) );
  OAI21_X1 U19175 ( .B1(n16884), .B2(n15945), .A(n15803), .ZN(P2_U2841) );
  AOI21_X1 U19176 ( .B1(n19757), .B2(n15804), .A(n15952), .ZN(n15807) );
  INV_X1 U19177 ( .A(n15804), .ZN(n15805) );
  NAND2_X1 U19178 ( .A1(n15912), .A2(n15805), .ZN(n15806) );
  MUX2_X1 U19179 ( .A(n15807), .B(n15806), .S(n16582), .Z(n15815) );
  NAND2_X1 U19180 ( .A1(n19737), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15808) );
  OAI211_X1 U19181 ( .C1(n15955), .C2(n11258), .A(n15808), .B(n17339), .ZN(
        n15809) );
  AOI21_X1 U19182 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n15951), .A(
        n15809), .ZN(n15810) );
  OAI21_X1 U19183 ( .B1(n15811), .B2(n15941), .A(n15810), .ZN(n15812) );
  AOI21_X1 U19184 ( .B1(n15813), .B2(n19760), .A(n15812), .ZN(n15814) );
  OAI211_X1 U19185 ( .C1(n15945), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        P2_U2842) );
  AOI21_X1 U19186 ( .B1(n19757), .B2(n15817), .A(n15952), .ZN(n15819) );
  MUX2_X1 U19187 ( .A(n15819), .B(n15818), .S(n16592), .Z(n15826) );
  INV_X1 U19188 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20449) );
  AOI21_X1 U19189 ( .B1(n19746), .B2(P2_EBX_REG_12__SCAN_IN), .A(n19745), .ZN(
        n15820) );
  OAI21_X1 U19190 ( .B1(n20449), .B2(n19748), .A(n15820), .ZN(n15821) );
  AOI21_X1 U19191 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15951), .A(
        n15821), .ZN(n15822) );
  OAI21_X1 U19192 ( .B1(n15823), .B2(n15941), .A(n15822), .ZN(n15824) );
  AOI21_X1 U19193 ( .B1(n16895), .B2(n19760), .A(n15824), .ZN(n15825) );
  OAI211_X1 U19194 ( .C1(n15945), .C2(n16897), .A(n15826), .B(n15825), .ZN(
        P2_U2843) );
  NAND2_X1 U19195 ( .A1(n15912), .A2(n15827), .ZN(n15830) );
  INV_X1 U19196 ( .A(n15827), .ZN(n15828) );
  AOI21_X1 U19197 ( .B1(n19757), .B2(n15828), .A(n15952), .ZN(n15829) );
  MUX2_X1 U19198 ( .A(n15830), .B(n15829), .S(n16621), .Z(n15840) );
  AND2_X1 U19199 ( .A1(n15831), .A2(n15832), .ZN(n15833) );
  OR2_X1 U19200 ( .A1(n15833), .A2(n13278), .ZN(n16623) );
  INV_X1 U19201 ( .A(n16623), .ZN(n16921) );
  AOI21_X1 U19202 ( .B1(n19746), .B2(P2_EBX_REG_10__SCAN_IN), .A(n19745), .ZN(
        n15834) );
  OAI21_X1 U19203 ( .B1(n20446), .B2(n19748), .A(n15834), .ZN(n15835) );
  AOI21_X1 U19204 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15951), .A(
        n15835), .ZN(n15836) );
  OAI21_X1 U19205 ( .B1(n15837), .B2(n15941), .A(n15836), .ZN(n15838) );
  AOI21_X1 U19206 ( .B1(n16921), .B2(n19761), .A(n15838), .ZN(n15839) );
  OAI211_X1 U19207 ( .C1(n16924), .C2(n15954), .A(n15840), .B(n15839), .ZN(
        P2_U2845) );
  INV_X1 U19208 ( .A(n19753), .ZN(n16996) );
  NOR2_X1 U19209 ( .A1(n16996), .A2(n15841), .ZN(n15842) );
  XOR2_X1 U19210 ( .A(n16634), .B(n15842), .Z(n15854) );
  INV_X1 U19211 ( .A(n15843), .ZN(n16932) );
  NAND2_X1 U19212 ( .A1(n19737), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n15844) );
  OAI211_X1 U19213 ( .C1(n15955), .C2(n10497), .A(n15844), .B(n17339), .ZN(
        n15845) );
  AOI21_X1 U19214 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n15951), .A(
        n15845), .ZN(n15846) );
  OAI21_X1 U19215 ( .B1(n15847), .B2(n15941), .A(n15846), .ZN(n15852) );
  NAND2_X1 U19216 ( .A1(n15848), .A2(n15849), .ZN(n15850) );
  NAND2_X1 U19217 ( .A1(n15831), .A2(n15850), .ZN(n16935) );
  NOR2_X1 U19218 ( .A1(n16935), .A2(n15945), .ZN(n15851) );
  AOI211_X1 U19219 ( .C1(n19760), .C2(n16932), .A(n15852), .B(n15851), .ZN(
        n15853) );
  OAI21_X1 U19220 ( .B1(n15854), .B2(n19734), .A(n15853), .ZN(P2_U2846) );
  OR2_X1 U19221 ( .A1(n15856), .A2(n15855), .ZN(n15857) );
  INV_X1 U19222 ( .A(n16650), .ZN(n16949) );
  NAND2_X1 U19223 ( .A1(n15912), .A2(n15858), .ZN(n15862) );
  INV_X1 U19224 ( .A(n15858), .ZN(n15859) );
  AOI21_X1 U19225 ( .B1(n19757), .B2(n15859), .A(n15952), .ZN(n15861) );
  MUX2_X1 U19226 ( .A(n15862), .B(n15861), .S(n15860), .Z(n15871) );
  INV_X1 U19227 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15868) );
  NAND2_X1 U19228 ( .A1(n15863), .A2(n19750), .ZN(n15867) );
  OAI21_X1 U19229 ( .B1(n15955), .B2(n15864), .A(n17339), .ZN(n15865) );
  AOI21_X1 U19230 ( .B1(n19737), .B2(P2_REIP_REG_8__SCAN_IN), .A(n15865), .ZN(
        n15866) );
  OAI211_X1 U19231 ( .C1(n19767), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        n15869) );
  AOI21_X1 U19232 ( .B1(n16946), .B2(n19760), .A(n15869), .ZN(n15870) );
  OAI211_X1 U19233 ( .C1(n16949), .C2(n15945), .A(n15871), .B(n15870), .ZN(
        P2_U2847) );
  NAND2_X1 U19234 ( .A1(n15912), .A2(n19756), .ZN(n15874) );
  INV_X1 U19235 ( .A(n19756), .ZN(n15872) );
  AOI21_X1 U19236 ( .B1(n19757), .B2(n15872), .A(n15952), .ZN(n15873) );
  MUX2_X1 U19237 ( .A(n15874), .B(n15873), .S(n16662), .Z(n15881) );
  OAI21_X1 U19238 ( .B1(n15955), .B2(n11255), .A(n17339), .ZN(n15875) );
  AOI21_X1 U19239 ( .B1(n19737), .B2(P2_REIP_REG_7__SCAN_IN), .A(n15875), .ZN(
        n15876) );
  OAI21_X1 U19240 ( .B1(n16660), .B2(n19767), .A(n15876), .ZN(n15878) );
  NOR2_X1 U19241 ( .A1(n16957), .A2(n15954), .ZN(n15877) );
  AOI211_X1 U19242 ( .C1(n19750), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        n15880) );
  OAI211_X1 U19243 ( .C1(n16955), .C2(n15945), .A(n15881), .B(n15880), .ZN(
        P2_U2848) );
  NOR2_X1 U19244 ( .A1(n16996), .A2(n15882), .ZN(n15883) );
  XOR2_X1 U19245 ( .A(n16684), .B(n15883), .Z(n15894) );
  INV_X1 U19246 ( .A(n15885), .ZN(n15886) );
  XNOR2_X1 U19247 ( .A(n15884), .B(n15886), .ZN(n17328) );
  NAND2_X1 U19248 ( .A1(n19737), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n15887) );
  OAI211_X1 U19249 ( .C1(n15955), .C2(n11155), .A(n15887), .B(n17339), .ZN(
        n15888) );
  AOI21_X1 U19250 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n15951), .A(
        n15888), .ZN(n15889) );
  OAI21_X1 U19251 ( .B1(n15890), .B2(n15941), .A(n15889), .ZN(n15892) );
  NOR2_X1 U19252 ( .A1(n17331), .A2(n15945), .ZN(n15891) );
  AOI211_X1 U19253 ( .C1(n19760), .C2(n17328), .A(n15892), .B(n15891), .ZN(
        n15893) );
  OAI21_X1 U19254 ( .B1(n15894), .B2(n19734), .A(n15893), .ZN(P2_U2850) );
  NAND2_X1 U19255 ( .A1(n15912), .A2(n15895), .ZN(n15898) );
  INV_X1 U19256 ( .A(n15895), .ZN(n15896) );
  AOI21_X1 U19257 ( .B1(n19757), .B2(n15896), .A(n15952), .ZN(n15897) );
  MUX2_X1 U19258 ( .A(n15898), .B(n15897), .S(n16696), .Z(n15909) );
  NAND2_X1 U19259 ( .A1(n15899), .A2(n15900), .ZN(n15901) );
  NAND2_X1 U19260 ( .A1(n15884), .A2(n15901), .ZN(n19771) );
  NOR2_X1 U19261 ( .A1(n19771), .A2(n15954), .ZN(n15907) );
  OAI21_X1 U19262 ( .B1(n15955), .B2(n15902), .A(n17339), .ZN(n15904) );
  NOR2_X1 U19263 ( .A1(n19767), .A2(n16699), .ZN(n15903) );
  AOI211_X1 U19264 ( .C1(n19737), .C2(P2_REIP_REG_4__SCAN_IN), .A(n15904), .B(
        n15903), .ZN(n15905) );
  OAI21_X1 U19265 ( .B1(n16693), .B2(n15941), .A(n15905), .ZN(n15906) );
  AOI211_X1 U19266 ( .C1(n16983), .C2(n19761), .A(n15907), .B(n15906), .ZN(
        n15908) );
  OAI211_X1 U19267 ( .C1(n19773), .C2(n15959), .A(n15909), .B(n15908), .ZN(
        P2_U2851) );
  AOI21_X1 U19268 ( .B1(n19757), .B2(n15910), .A(n15952), .ZN(n15914) );
  INV_X1 U19269 ( .A(n15910), .ZN(n15911) );
  NAND2_X1 U19270 ( .A1(n15912), .A2(n15911), .ZN(n15913) );
  MUX2_X1 U19271 ( .A(n15914), .B(n15913), .S(n16716), .Z(n15923) );
  NAND2_X1 U19272 ( .A1(n15916), .A2(n15915), .ZN(n15917) );
  NAND2_X1 U19273 ( .A1(n15899), .A2(n15917), .ZN(n20502) );
  OAI22_X1 U19274 ( .A1(n19748), .A2(n10136), .B1(n15955), .B2(n11251), .ZN(
        n15918) );
  AOI21_X1 U19275 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15918), .ZN(n15920) );
  NAND2_X1 U19276 ( .A1(n19750), .A2(n16688), .ZN(n15919) );
  OAI211_X1 U19277 ( .C1(n20502), .C2(n15954), .A(n15920), .B(n15919), .ZN(
        n15921) );
  AOI21_X1 U19278 ( .B1(n17345), .B2(n19761), .A(n15921), .ZN(n15922) );
  OAI211_X1 U19279 ( .C1(n20169), .C2(n15959), .A(n15923), .B(n15922), .ZN(
        P2_U2852) );
  INV_X1 U19280 ( .A(n15924), .ZN(n15925) );
  NAND2_X1 U19281 ( .A1(n19753), .A2(n15925), .ZN(n15935) );
  XNOR2_X1 U19282 ( .A(n15935), .B(n15926), .ZN(n15934) );
  INV_X1 U19283 ( .A(n15959), .ZN(n15948) );
  OAI22_X1 U19284 ( .A1(n15955), .A2(n11247), .B1(n20431), .B2(n19748), .ZN(
        n15927) );
  AOI21_X1 U19285 ( .B1(n15951), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15927), .ZN(n15928) );
  OAI21_X1 U19286 ( .B1(n15929), .B2(n15941), .A(n15928), .ZN(n15930) );
  AOI21_X1 U19287 ( .B1(n19760), .B2(n20510), .A(n15930), .ZN(n15931) );
  OAI21_X1 U19288 ( .B1(n13240), .B2(n15945), .A(n15931), .ZN(n15932) );
  AOI21_X1 U19289 ( .B1(n20508), .B2(n15948), .A(n15932), .ZN(n15933) );
  OAI21_X1 U19290 ( .B1(n15934), .B2(n19734), .A(n15933), .ZN(P2_U2853) );
  INV_X1 U19291 ( .A(n15935), .ZN(n15938) );
  NAND2_X1 U19292 ( .A1(n15936), .A2(n16990), .ZN(n15937) );
  NAND2_X1 U19293 ( .A1(n15938), .A2(n15937), .ZN(n16998) );
  MUX2_X1 U19294 ( .A(n10546), .B(n19767), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15950) );
  NOR2_X1 U19295 ( .A1(n19748), .A2(n20429), .ZN(n15943) );
  OAI22_X1 U19296 ( .A1(n15941), .A2(n15940), .B1(n15955), .B2(n15939), .ZN(
        n15942) );
  AOI211_X1 U19297 ( .C1(n19760), .C2(n20513), .A(n15943), .B(n15942), .ZN(
        n15944) );
  OAI21_X1 U19298 ( .B1(n15946), .B2(n15945), .A(n15944), .ZN(n15947) );
  AOI21_X1 U19299 ( .B1(n20494), .B2(n15948), .A(n15947), .ZN(n15949) );
  OAI211_X1 U19300 ( .C1(n16998), .C2(n19734), .A(n15950), .B(n15949), .ZN(
        P2_U2854) );
  INV_X1 U19301 ( .A(n16990), .ZN(n15966) );
  OAI21_X1 U19302 ( .B1(n15952), .B2(n15951), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15964) );
  OAI22_X1 U19303 ( .A1(n15955), .A2(n11249), .B1(n15954), .B2(n15953), .ZN(
        n15956) );
  AOI21_X1 U19304 ( .B1(n19750), .B2(n15957), .A(n15956), .ZN(n15958) );
  OAI21_X1 U19305 ( .B1(n19722), .B2(n19748), .A(n15958), .ZN(n15961) );
  NOR2_X1 U19306 ( .A1(n20526), .A2(n15959), .ZN(n15960) );
  AOI211_X1 U19307 ( .C1(n19761), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        n15963) );
  OAI211_X1 U19308 ( .C1(n15966), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        P2_U2855) );
  AOI22_X1 U19309 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15971) );
  AOI22_X1 U19310 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15970) );
  AOI22_X1 U19311 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19312 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15968) );
  NAND4_X1 U19313 ( .A1(n15971), .A2(n15970), .A3(n15969), .A4(n15968), .ZN(
        n15977) );
  AOI22_X1 U19314 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14409), .ZN(n15975) );
  AOI22_X1 U19315 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15974) );
  AOI22_X1 U19316 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9589), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15973) );
  AOI22_X1 U19317 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15972) );
  NAND4_X1 U19318 ( .A1(n15975), .A2(n15974), .A3(n15973), .A4(n15972), .ZN(
        n15976) );
  OR2_X1 U19319 ( .A1(n15977), .A2(n15976), .ZN(n16278) );
  NAND3_X1 U19320 ( .A1(n15979), .A2(n15978), .A3(n16278), .ZN(n15981) );
  AOI22_X1 U19321 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15986) );
  AOI22_X1 U19322 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15985) );
  AOI22_X1 U19323 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15984) );
  AOI22_X1 U19324 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15983) );
  NAND4_X1 U19325 ( .A1(n15986), .A2(n15985), .A3(n15984), .A4(n15983), .ZN(
        n15992) );
  AOI22_X1 U19326 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n14409), .ZN(n15990) );
  AOI22_X1 U19327 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15989) );
  AOI22_X1 U19328 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n16048), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15988) );
  AOI22_X1 U19329 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15987) );
  NAND4_X1 U19330 ( .A1(n15990), .A2(n15989), .A3(n15988), .A4(n15987), .ZN(
        n15991) );
  NOR2_X1 U19331 ( .A1(n15992), .A2(n15991), .ZN(n16275) );
  AOI22_X1 U19332 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U19333 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15996) );
  AOI22_X1 U19334 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15995) );
  AOI22_X1 U19335 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15994) );
  NAND4_X1 U19336 ( .A1(n15997), .A2(n15996), .A3(n15995), .A4(n15994), .ZN(
        n16003) );
  AOI22_X1 U19337 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14409), .ZN(n16001) );
  AOI22_X1 U19338 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16000) );
  AOI22_X1 U19339 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9589), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19340 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15998) );
  NAND4_X1 U19341 ( .A1(n16001), .A2(n16000), .A3(n15999), .A4(n15998), .ZN(
        n16002) );
  AOI22_X1 U19342 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16007) );
  AOI22_X1 U19343 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U19344 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19345 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16004) );
  NAND4_X1 U19346 ( .A1(n16007), .A2(n16006), .A3(n16005), .A4(n16004), .ZN(
        n16013) );
  AOI22_X1 U19347 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n14409), .ZN(n16011) );
  AOI22_X1 U19348 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16010) );
  AOI22_X1 U19349 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n9589), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16009) );
  AOI22_X1 U19350 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16008) );
  NAND4_X1 U19351 ( .A1(n16011), .A2(n16010), .A3(n16009), .A4(n16008), .ZN(
        n16012) );
  NOR2_X1 U19352 ( .A1(n16013), .A2(n16012), .ZN(n16267) );
  AOI22_X1 U19353 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n16042), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16018) );
  AOI22_X1 U19354 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n16041), .B1(
        n14107), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16017) );
  AOI22_X1 U19355 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16016) );
  AOI22_X1 U19356 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16015) );
  NAND4_X1 U19357 ( .A1(n16018), .A2(n16017), .A3(n16016), .A4(n16015), .ZN(
        n16024) );
  AOI22_X1 U19358 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14409), .ZN(n16022) );
  AOI22_X1 U19359 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U19360 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9589), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16020) );
  AOI22_X1 U19361 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16019) );
  NAND4_X1 U19362 ( .A1(n16022), .A2(n16021), .A3(n16020), .A4(n16019), .ZN(
        n16023) );
  NOR2_X1 U19363 ( .A1(n16024), .A2(n16023), .ZN(n16261) );
  INV_X1 U19364 ( .A(n16261), .ZN(n16025) );
  AOI22_X1 U19365 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16028) );
  AOI22_X1 U19366 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16027) );
  AND2_X1 U19367 ( .A1(n16028), .A2(n16027), .ZN(n16031) );
  XNOR2_X1 U19368 ( .A(n14334), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16198) );
  AOI22_X1 U19369 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16090), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U19370 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16201), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16029) );
  NAND4_X1 U19371 ( .A1(n16031), .A2(n16198), .A3(n16030), .A4(n16029), .ZN(
        n16040) );
  NAND2_X1 U19372 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n16035) );
  NAND2_X1 U19373 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n16034) );
  NAND2_X1 U19374 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n16033) );
  NAND2_X1 U19375 ( .A1(n16195), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n16032) );
  AND4_X1 U19376 ( .A1(n16035), .A2(n16034), .A3(n16033), .A4(n16032), .ZN(
        n16038) );
  AOI22_X1 U19377 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U19378 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16036) );
  INV_X1 U19379 ( .A(n16198), .ZN(n16192) );
  NAND4_X1 U19380 ( .A1(n16038), .A2(n16037), .A3(n16036), .A4(n16192), .ZN(
        n16039) );
  NAND2_X1 U19381 ( .A1(n20549), .A2(n16077), .ZN(n16055) );
  AOI22_X1 U19382 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n16042), .B1(
        n16041), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16047) );
  AOI22_X1 U19383 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n14107), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U19384 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10990), .B1(
        n16043), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16045) );
  AOI22_X1 U19385 ( .A1(n11039), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15993), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16044) );
  NAND4_X1 U19386 ( .A1(n16047), .A2(n16046), .A3(n16045), .A4(n16044), .ZN(
        n16054) );
  AOI22_X1 U19387 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14409), .ZN(n16052) );
  AOI22_X1 U19388 ( .A1(n10995), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11044), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16051) );
  AOI22_X1 U19389 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16048), .B1(
        n11091), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U19390 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11069), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16049) );
  NAND4_X1 U19391 ( .A1(n16052), .A2(n16051), .A3(n16050), .A4(n16049), .ZN(
        n16053) );
  OR2_X1 U19392 ( .A1(n16054), .A2(n16053), .ZN(n16059) );
  XNOR2_X1 U19393 ( .A(n16055), .B(n16059), .ZN(n16078) );
  INV_X1 U19394 ( .A(n16077), .ZN(n16056) );
  NOR2_X1 U19395 ( .A1(n20549), .A2(n16056), .ZN(n16255) );
  INV_X1 U19396 ( .A(n16078), .ZN(n16057) );
  NAND2_X1 U19397 ( .A1(n16059), .A2(n16077), .ZN(n16081) );
  NAND2_X1 U19398 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n16063) );
  NAND2_X1 U19399 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n16062) );
  NAND2_X1 U19400 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n16061) );
  INV_X1 U19401 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21658) );
  NAND2_X1 U19402 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n16060) );
  AND4_X1 U19403 ( .A1(n16063), .A2(n16062), .A3(n16061), .A4(n16060), .ZN(
        n16066) );
  AOI22_X1 U19404 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U19405 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16064) );
  NAND4_X1 U19406 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n16192), .ZN(
        n16075) );
  NAND2_X1 U19407 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n16070) );
  NAND2_X1 U19408 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n16069) );
  NAND2_X1 U19409 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n16068) );
  NAND2_X1 U19410 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n16067) );
  AND4_X1 U19411 ( .A1(n16070), .A2(n16069), .A3(n16068), .A4(n16067), .ZN(
        n16073) );
  AOI22_X1 U19412 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16072) );
  AOI22_X1 U19413 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16071) );
  NAND4_X1 U19414 ( .A1(n16073), .A2(n16072), .A3(n16071), .A4(n16198), .ZN(
        n16074) );
  NAND2_X1 U19415 ( .A1(n16075), .A2(n16074), .ZN(n16080) );
  XNOR2_X1 U19416 ( .A(n16081), .B(n16080), .ZN(n16076) );
  NOR2_X1 U19417 ( .A1(n16076), .A2(n9595), .ZN(n16249) );
  NAND2_X1 U19418 ( .A1(n16248), .A2(n16249), .ZN(n16247) );
  NOR2_X1 U19419 ( .A1(n20549), .A2(n16080), .ZN(n16251) );
  NAND3_X1 U19420 ( .A1(n16078), .A2(n16077), .A3(n16251), .ZN(n16079) );
  NOR2_X1 U19421 ( .A1(n16081), .A2(n16080), .ZN(n16100) );
  NAND2_X1 U19422 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n16085) );
  NAND2_X1 U19423 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n16084) );
  NAND2_X1 U19424 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n16083) );
  NAND2_X1 U19425 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n16082) );
  AND4_X1 U19426 ( .A1(n16085), .A2(n16084), .A3(n16083), .A4(n16082), .ZN(
        n16089) );
  AOI22_X1 U19427 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16088) );
  INV_X1 U19428 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n20060) );
  AOI22_X1 U19429 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16087) );
  NAND4_X1 U19430 ( .A1(n16089), .A2(n16088), .A3(n16087), .A4(n16192), .ZN(
        n16099) );
  NAND2_X1 U19431 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n16094) );
  NAND2_X1 U19432 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n16093) );
  NAND2_X1 U19433 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n16092) );
  NAND2_X1 U19434 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n16091) );
  AND4_X1 U19435 ( .A1(n16094), .A2(n16093), .A3(n16092), .A4(n16091), .ZN(
        n16097) );
  AOI22_X1 U19436 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16096) );
  AOI22_X1 U19437 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16095) );
  NAND4_X1 U19438 ( .A1(n16097), .A2(n16096), .A3(n16095), .A4(n16198), .ZN(
        n16098) );
  AND2_X1 U19439 ( .A1(n16099), .A2(n16098), .ZN(n16117) );
  NAND2_X1 U19440 ( .A1(n16100), .A2(n16117), .ZN(n16122) );
  OAI211_X1 U19441 ( .C1(n16100), .C2(n16117), .A(n16122), .B(n16120), .ZN(
        n16119) );
  NAND2_X1 U19442 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n16104) );
  NAND2_X1 U19443 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n16103) );
  NAND2_X1 U19444 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n16102) );
  NAND2_X1 U19445 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n16101) );
  AND4_X1 U19446 ( .A1(n16104), .A2(n16103), .A3(n16102), .A4(n16101), .ZN(
        n16107) );
  AOI22_X1 U19447 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U19448 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16105) );
  NAND4_X1 U19449 ( .A1(n16107), .A2(n16106), .A3(n16105), .A4(n16192), .ZN(
        n16116) );
  NAND2_X1 U19450 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n16111) );
  NAND2_X1 U19451 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n16110) );
  NAND2_X1 U19452 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n16109) );
  NAND2_X1 U19453 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n16108) );
  AND4_X1 U19454 ( .A1(n16111), .A2(n16110), .A3(n16109), .A4(n16108), .ZN(
        n16114) );
  AOI22_X1 U19455 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16113) );
  AOI22_X1 U19456 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16112) );
  NAND4_X1 U19457 ( .A1(n16114), .A2(n16113), .A3(n16112), .A4(n16198), .ZN(
        n16115) );
  INV_X1 U19458 ( .A(n16117), .ZN(n16118) );
  NOR2_X1 U19459 ( .A1(n20549), .A2(n16118), .ZN(n16243) );
  XNOR2_X1 U19460 ( .A(n16122), .B(n16234), .ZN(n16121) );
  NAND2_X1 U19461 ( .A1(n16121), .A2(n16120), .ZN(n16236) );
  INV_X1 U19462 ( .A(n16122), .ZN(n16123) );
  AND2_X1 U19463 ( .A1(n16123), .A2(n16234), .ZN(n16140) );
  NAND2_X1 U19464 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n16127) );
  NAND2_X1 U19465 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n16126) );
  NAND2_X1 U19466 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n16125) );
  NAND2_X1 U19467 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n16124) );
  AND4_X1 U19468 ( .A1(n16127), .A2(n16126), .A3(n16125), .A4(n16124), .ZN(
        n16130) );
  AOI22_X1 U19469 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U19470 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16128) );
  NAND4_X1 U19471 ( .A1(n16130), .A2(n16129), .A3(n16128), .A4(n16192), .ZN(
        n16139) );
  NAND2_X1 U19472 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n16134) );
  NAND2_X1 U19473 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n16133) );
  NAND2_X1 U19474 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n16132) );
  NAND2_X1 U19475 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n16131) );
  AND4_X1 U19476 ( .A1(n16134), .A2(n16133), .A3(n16132), .A4(n16131), .ZN(
        n16137) );
  AOI22_X1 U19477 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16136) );
  AOI22_X1 U19478 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16135) );
  NAND4_X1 U19479 ( .A1(n16137), .A2(n16136), .A3(n16135), .A4(n16198), .ZN(
        n16138) );
  AND2_X1 U19480 ( .A1(n16139), .A2(n16138), .ZN(n16148) );
  NAND2_X1 U19481 ( .A1(n16140), .A2(n16148), .ZN(n16220) );
  INV_X1 U19482 ( .A(n16140), .ZN(n16143) );
  INV_X1 U19483 ( .A(n16148), .ZN(n16142) );
  AOI21_X1 U19484 ( .B1(n16143), .B2(n16142), .A(n9595), .ZN(n16144) );
  AND2_X1 U19485 ( .A1(n16220), .A2(n16144), .ZN(n16145) );
  NAND2_X1 U19486 ( .A1(n16146), .A2(n16145), .ZN(n16221) );
  NAND2_X1 U19487 ( .A1(n16147), .A2(n16221), .ZN(n16227) );
  NAND2_X1 U19488 ( .A1(n16235), .A2(n16148), .ZN(n16226) );
  INV_X1 U19489 ( .A(n16221), .ZN(n16166) );
  NAND2_X1 U19490 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n16152) );
  NAND2_X1 U19491 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n16151) );
  NAND2_X1 U19492 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n16150) );
  NAND2_X1 U19493 ( .A1(n16196), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n16149) );
  AND4_X1 U19494 ( .A1(n16152), .A2(n16151), .A3(n16150), .A4(n16149), .ZN(
        n16155) );
  AOI22_X1 U19495 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16154) );
  AOI22_X1 U19496 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16153) );
  NAND4_X1 U19497 ( .A1(n16155), .A2(n16154), .A3(n16153), .A4(n16192), .ZN(
        n16165) );
  NAND2_X1 U19498 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n16159) );
  NAND2_X1 U19499 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n16158) );
  NAND2_X1 U19500 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n16157) );
  NAND2_X1 U19501 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n16156) );
  AND4_X1 U19502 ( .A1(n16159), .A2(n16158), .A3(n16157), .A4(n16156), .ZN(
        n16163) );
  AOI22_X1 U19503 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16162) );
  AOI22_X1 U19504 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16161) );
  NAND4_X1 U19505 ( .A1(n16163), .A2(n16162), .A3(n16161), .A4(n16198), .ZN(
        n16164) );
  AND2_X1 U19506 ( .A1(n16165), .A2(n16164), .ZN(n16222) );
  INV_X1 U19507 ( .A(n16220), .ZN(n16168) );
  AND2_X1 U19508 ( .A1(n20549), .A2(n16222), .ZN(n16167) );
  AND2_X1 U19509 ( .A1(n16168), .A2(n16167), .ZN(n16186) );
  NAND2_X1 U19510 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16172) );
  NAND2_X1 U19511 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n16171) );
  NAND2_X1 U19512 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n16170) );
  NAND2_X1 U19513 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n16169) );
  AND4_X1 U19514 ( .A1(n16172), .A2(n16171), .A3(n16170), .A4(n16169), .ZN(
        n16175) );
  AOI22_X1 U19515 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16174) );
  AOI22_X1 U19516 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16173) );
  NAND4_X1 U19517 ( .A1(n16175), .A2(n16174), .A3(n16173), .A4(n16192), .ZN(
        n16184) );
  NAND2_X1 U19518 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n16179) );
  NAND2_X1 U19519 ( .A1(n16201), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n16178) );
  NAND2_X1 U19520 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n16177) );
  NAND2_X1 U19521 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n16176) );
  AND4_X1 U19522 ( .A1(n16179), .A2(n16178), .A3(n16177), .A4(n16176), .ZN(
        n16182) );
  AOI22_X1 U19523 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U19524 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16180) );
  NAND4_X1 U19525 ( .A1(n16182), .A2(n16181), .A3(n16180), .A4(n16198), .ZN(
        n16183) );
  AND2_X1 U19526 ( .A1(n16184), .A2(n16183), .ZN(n16185) );
  NAND2_X1 U19527 ( .A1(n16186), .A2(n16185), .ZN(n16187) );
  OAI21_X1 U19528 ( .B1(n16186), .B2(n16185), .A(n16187), .ZN(n16215) );
  NOR2_X1 U19529 ( .A1(n16216), .A2(n16215), .ZN(n16214) );
  INV_X1 U19530 ( .A(n16187), .ZN(n16188) );
  NOR2_X1 U19531 ( .A1(n16214), .A2(n16188), .ZN(n16210) );
  AOI22_X1 U19532 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16201), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16191) );
  AOI22_X1 U19533 ( .A1(n16189), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16090), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16190) );
  NAND2_X1 U19534 ( .A1(n16191), .A2(n16190), .ZN(n16208) );
  AOI22_X1 U19535 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16194) );
  AOI22_X1 U19536 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16193) );
  NAND3_X1 U19537 ( .A1(n16194), .A2(n16193), .A3(n16192), .ZN(n16207) );
  AOI22_X1 U19538 ( .A1(n16160), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16195), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U19539 ( .A1(n16197), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16196), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16199) );
  NAND3_X1 U19540 ( .A1(n16200), .A2(n16199), .A3(n16198), .ZN(n16206) );
  AOI22_X1 U19541 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16201), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U19542 ( .A1(n16090), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16203) );
  NAND2_X1 U19543 ( .A1(n16204), .A2(n16203), .ZN(n16205) );
  OAI22_X1 U19544 ( .A1(n16208), .A2(n16207), .B1(n16206), .B2(n16205), .ZN(
        n16209) );
  XNOR2_X1 U19545 ( .A(n16210), .B(n16209), .ZN(n16323) );
  NOR2_X1 U19546 ( .A1(n16211), .A2(n16287), .ZN(n16212) );
  OAI21_X1 U19547 ( .B1(n16323), .B2(n16301), .A(n16213), .ZN(P2_U2857) );
  INV_X1 U19548 ( .A(n16214), .ZN(n16325) );
  NAND2_X1 U19549 ( .A1(n16216), .A2(n16215), .ZN(n16324) );
  NAND3_X1 U19550 ( .A1(n16325), .A2(n16311), .A3(n16324), .ZN(n16218) );
  NAND2_X1 U19551 ( .A1(n16287), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16217) );
  OAI211_X1 U19552 ( .C1(n16219), .C2(n16287), .A(n16218), .B(n16217), .ZN(
        P2_U2858) );
  NAND2_X1 U19553 ( .A1(n16221), .A2(n16220), .ZN(n16223) );
  XNOR2_X1 U19554 ( .A(n16223), .B(n16222), .ZN(n16338) );
  NOR2_X1 U19555 ( .A1(n16739), .A2(n16287), .ZN(n16224) );
  AOI21_X1 U19556 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16287), .A(n16224), .ZN(
        n16225) );
  OAI21_X1 U19557 ( .B1(n16338), .B2(n16301), .A(n16225), .ZN(P2_U2859) );
  AND2_X1 U19558 ( .A1(n16227), .A2(n16226), .ZN(n16228) );
  NOR2_X1 U19559 ( .A1(n16229), .A2(n16228), .ZN(n16339) );
  NAND2_X1 U19560 ( .A1(n16339), .A2(n16311), .ZN(n16231) );
  NAND2_X1 U19561 ( .A1(n16287), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16230) );
  OAI211_X1 U19562 ( .C1(n16748), .C2(n16287), .A(n16231), .B(n16230), .ZN(
        P2_U2860) );
  NAND2_X1 U19563 ( .A1(n16232), .A2(n16243), .ZN(n16242) );
  NAND2_X1 U19564 ( .A1(n16242), .A2(n16233), .ZN(n16239) );
  NAND2_X1 U19565 ( .A1(n16235), .A2(n16234), .ZN(n16237) );
  XOR2_X1 U19566 ( .A(n16237), .B(n16236), .Z(n16238) );
  XNOR2_X1 U19567 ( .A(n16239), .B(n16238), .ZN(n16354) );
  MUX2_X1 U19568 ( .A(n16752), .B(n16240), .S(n16287), .Z(n16241) );
  OAI21_X1 U19569 ( .B1(n16354), .B2(n16301), .A(n16241), .ZN(P2_U2861) );
  OAI21_X1 U19570 ( .B1(n16232), .B2(n16243), .A(n16242), .ZN(n16362) );
  NAND2_X1 U19571 ( .A1(n16244), .A2(n16308), .ZN(n16246) );
  NAND2_X1 U19572 ( .A1(n16287), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16245) );
  OAI211_X1 U19573 ( .C1(n16362), .C2(n16301), .A(n16246), .B(n16245), .ZN(
        P2_U2862) );
  OAI21_X1 U19574 ( .B1(n16249), .B2(n16248), .A(n16247), .ZN(n16250) );
  XOR2_X1 U19575 ( .A(n16251), .B(n16250), .Z(n16369) );
  NAND2_X1 U19576 ( .A1(n16777), .A2(n16308), .ZN(n16253) );
  NAND2_X1 U19577 ( .A1(n16287), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16252) );
  OAI211_X1 U19578 ( .C1(n16369), .C2(n16301), .A(n16253), .B(n16252), .ZN(
        P2_U2863) );
  OAI21_X1 U19579 ( .B1(n16256), .B2(n16255), .A(n16254), .ZN(n16376) );
  INV_X1 U19580 ( .A(n16376), .ZN(n16257) );
  AOI22_X1 U19581 ( .A1(n16257), .A2(n16311), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n16287), .ZN(n16258) );
  OAI21_X1 U19582 ( .B1(n16259), .B2(n16287), .A(n16258), .ZN(P2_U2864) );
  INV_X1 U19583 ( .A(n16805), .ZN(n16265) );
  NAND2_X1 U19584 ( .A1(n16260), .A2(n16261), .ZN(n16262) );
  AND2_X1 U19585 ( .A1(n16263), .A2(n16262), .ZN(n16382) );
  AOI22_X1 U19586 ( .A1(n16382), .A2(n16311), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16287), .ZN(n16264) );
  OAI21_X1 U19587 ( .B1(n16265), .B2(n16287), .A(n16264), .ZN(P2_U2865) );
  INV_X1 U19588 ( .A(n16260), .ZN(n16266) );
  AOI21_X1 U19589 ( .B1(n16267), .B2(n16270), .A(n16266), .ZN(n16388) );
  AOI22_X1 U19590 ( .A1(n16388), .A2(n16311), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16287), .ZN(n16268) );
  OAI21_X1 U19591 ( .B1(n16269), .B2(n16287), .A(n16268), .ZN(P2_U2866) );
  OAI21_X1 U19592 ( .B1(n16274), .B2(n16271), .A(n16270), .ZN(n16399) );
  INV_X1 U19593 ( .A(n16399), .ZN(n16272) );
  AOI22_X1 U19594 ( .A1(n16272), .A2(n16311), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16287), .ZN(n16273) );
  OAI21_X1 U19595 ( .B1(n19730), .B2(n16287), .A(n16273), .ZN(P2_U2867) );
  INV_X1 U19596 ( .A(n16829), .ZN(n16277) );
  AOI21_X1 U19597 ( .B1(n16275), .B2(n16279), .A(n16274), .ZN(n16405) );
  AOI22_X1 U19598 ( .A1(n16405), .A2(n16311), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16287), .ZN(n16276) );
  OAI21_X1 U19599 ( .B1(n16277), .B2(n16287), .A(n16276), .ZN(P2_U2868) );
  INV_X1 U19600 ( .A(n16278), .ZN(n16281) );
  INV_X1 U19601 ( .A(n16279), .ZN(n16280) );
  AOI21_X1 U19602 ( .B1(n16282), .B2(n16281), .A(n16280), .ZN(n16415) );
  AOI22_X1 U19603 ( .A1(n16415), .A2(n16311), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16287), .ZN(n16283) );
  OAI21_X1 U19604 ( .B1(n16839), .B2(n16287), .A(n16283), .ZN(P2_U2869) );
  INV_X1 U19605 ( .A(n16284), .ZN(n16285) );
  AOI22_X1 U19606 ( .A1(n16285), .A2(n16311), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16287), .ZN(n16286) );
  OAI21_X1 U19607 ( .B1(n16855), .B2(n16287), .A(n16286), .ZN(P2_U2870) );
  MUX2_X1 U19608 ( .A(n16288), .B(n16866), .S(n16308), .Z(n16289) );
  OAI21_X1 U19609 ( .B1(n16301), .B2(n16290), .A(n16289), .ZN(P2_U2871) );
  NAND2_X1 U19610 ( .A1(n16291), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n16309) );
  NOR2_X1 U19611 ( .A1(n16309), .A2(n16292), .ZN(n16310) );
  NAND2_X1 U19612 ( .A1(n16310), .A2(n16304), .ZN(n16303) );
  NOR2_X1 U19613 ( .A1(n16303), .A2(n16298), .ZN(n16295) );
  INV_X1 U19614 ( .A(n14095), .ZN(n16293) );
  OAI211_X1 U19615 ( .C1(n16295), .C2(n16294), .A(n16293), .B(n16311), .ZN(
        n16297) );
  INV_X1 U19616 ( .A(n16603), .ZN(n16908) );
  NAND2_X1 U19617 ( .A1(n16908), .A2(n16308), .ZN(n16296) );
  OAI211_X1 U19618 ( .C1(n16308), .C2(n13273), .A(n16297), .B(n16296), .ZN(
        P2_U2876) );
  XNOR2_X1 U19619 ( .A(n16303), .B(n16298), .ZN(n16302) );
  MUX2_X1 U19620 ( .A(n16623), .B(n16299), .S(n16287), .Z(n16300) );
  OAI21_X1 U19621 ( .B1(n16302), .B2(n16301), .A(n16300), .ZN(P2_U2877) );
  OAI211_X1 U19622 ( .C1(n16310), .C2(n16304), .A(n16303), .B(n16311), .ZN(
        n16307) );
  INV_X1 U19623 ( .A(n16935), .ZN(n16305) );
  NAND2_X1 U19624 ( .A1(n16305), .A2(n16308), .ZN(n16306) );
  OAI211_X1 U19625 ( .C1(n16308), .C2(n10497), .A(n16307), .B(n16306), .ZN(
        P2_U2878) );
  INV_X1 U19626 ( .A(n16309), .ZN(n16314) );
  INV_X1 U19627 ( .A(n16310), .ZN(n16312) );
  OAI211_X1 U19628 ( .C1(n16314), .C2(n16313), .A(n16312), .B(n16311), .ZN(
        n16316) );
  NAND2_X1 U19629 ( .A1(n16287), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n16315) );
  OAI211_X1 U19630 ( .C1(n16949), .C2(n16287), .A(n16316), .B(n16315), .ZN(
        P2_U2879) );
  INV_X1 U19631 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16319) );
  AOI22_X1 U19632 ( .A1(n16408), .A2(n19829), .B1(n19785), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n16318) );
  NAND2_X1 U19633 ( .A1(n16395), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16317) );
  OAI211_X1 U19634 ( .C1(n16392), .C2(n16319), .A(n16318), .B(n16317), .ZN(
        n16320) );
  AOI21_X1 U19635 ( .B1(n16321), .B2(n19786), .A(n16320), .ZN(n16322) );
  OAI21_X1 U19636 ( .B1(n16323), .B2(n16398), .A(n16322), .ZN(P2_U2889) );
  NAND3_X1 U19637 ( .A1(n16325), .A2(n19790), .A3(n16324), .ZN(n16330) );
  AOI22_X1 U19638 ( .A1(n16408), .A2(n16326), .B1(n19785), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16327) );
  OAI21_X1 U19639 ( .B1(n16392), .B2(n19123), .A(n16327), .ZN(n16328) );
  AOI21_X1 U19640 ( .B1(n16395), .B2(BUF1_REG_29__SCAN_IN), .A(n16328), .ZN(
        n16329) );
  OAI211_X1 U19641 ( .C1(n16731), .C2(n19770), .A(n16330), .B(n16329), .ZN(
        P2_U2890) );
  INV_X1 U19642 ( .A(n16395), .ZN(n16413) );
  AOI22_X1 U19643 ( .A1(n16408), .A2(n16331), .B1(n19785), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16333) );
  NAND2_X1 U19644 ( .A1(n16409), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16332) );
  OAI211_X1 U19645 ( .C1(n16413), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16335) );
  AOI21_X1 U19646 ( .B1(n16336), .B2(n19786), .A(n16335), .ZN(n16337) );
  OAI21_X1 U19647 ( .B1(n16338), .B2(n16398), .A(n16337), .ZN(P2_U2891) );
  INV_X1 U19648 ( .A(n16339), .ZN(n16346) );
  NAND2_X1 U19649 ( .A1(n16395), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16343) );
  NAND2_X1 U19650 ( .A1(n16409), .A2(BUF2_REG_27__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U19651 ( .A1(n16408), .A2(n16340), .B1(n19785), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16341) );
  NAND3_X1 U19652 ( .A1(n16343), .A2(n16342), .A3(n16341), .ZN(n16344) );
  AOI21_X1 U19653 ( .B1(n16747), .B2(n19786), .A(n16344), .ZN(n16345) );
  OAI21_X1 U19654 ( .B1(n16398), .B2(n16346), .A(n16345), .ZN(P2_U2892) );
  AOI22_X1 U19655 ( .A1(n16408), .A2(n16347), .B1(n19785), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16349) );
  NAND2_X1 U19656 ( .A1(n16409), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16348) );
  OAI211_X1 U19657 ( .C1(n16413), .C2(n16350), .A(n16349), .B(n16348), .ZN(
        n16351) );
  AOI21_X1 U19658 ( .B1(n16352), .B2(n19786), .A(n16351), .ZN(n16353) );
  OAI21_X1 U19659 ( .B1(n16354), .B2(n16398), .A(n16353), .ZN(P2_U2893) );
  INV_X1 U19660 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16357) );
  AOI22_X1 U19661 ( .A1(n16408), .A2(n16355), .B1(n19785), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16356) );
  OAI21_X1 U19662 ( .B1(n16392), .B2(n16357), .A(n16356), .ZN(n16360) );
  NOR2_X1 U19663 ( .A1(n16358), .A2(n19770), .ZN(n16359) );
  AOI211_X1 U19664 ( .C1(n16395), .C2(BUF1_REG_25__SCAN_IN), .A(n16360), .B(
        n16359), .ZN(n16361) );
  OAI21_X1 U19665 ( .B1(n16398), .B2(n16362), .A(n16361), .ZN(P2_U2894) );
  NAND2_X1 U19666 ( .A1(n16395), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U19667 ( .A1(n16408), .A2(n16363), .B1(n19785), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16364) );
  NAND2_X1 U19668 ( .A1(n16365), .A2(n16364), .ZN(n16367) );
  NOR2_X1 U19669 ( .A1(n16775), .A2(n19770), .ZN(n16366) );
  AOI211_X1 U19670 ( .C1(n16409), .C2(BUF2_REG_24__SCAN_IN), .A(n16367), .B(
        n16366), .ZN(n16368) );
  OAI21_X1 U19671 ( .B1(n16398), .B2(n16369), .A(n16368), .ZN(P2_U2895) );
  AOI22_X1 U19672 ( .A1(n16408), .A2(n16370), .B1(n19785), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16371) );
  OAI21_X1 U19673 ( .B1(n16413), .B2(n16372), .A(n16371), .ZN(n16374) );
  NOR2_X1 U19674 ( .A1(n16787), .A2(n19770), .ZN(n16373) );
  AOI211_X1 U19675 ( .C1(n16409), .C2(BUF2_REG_23__SCAN_IN), .A(n16374), .B(
        n16373), .ZN(n16375) );
  OAI21_X1 U19676 ( .B1(n16398), .B2(n16376), .A(n16375), .ZN(P2_U2896) );
  NAND2_X1 U19677 ( .A1(n16409), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U19678 ( .A1(n16395), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16379) );
  AOI22_X1 U19679 ( .A1(n16408), .A2(n16377), .B1(n19785), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16378) );
  NAND3_X1 U19680 ( .A1(n16380), .A2(n16379), .A3(n16378), .ZN(n16381) );
  AOI21_X1 U19681 ( .B1(n16382), .B2(n19790), .A(n16381), .ZN(n16383) );
  OAI21_X1 U19682 ( .B1(n16803), .B2(n19770), .A(n16383), .ZN(P2_U2897) );
  INV_X1 U19683 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U19684 ( .A1(n16408), .A2(n19866), .B1(n19785), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16385) );
  NAND2_X1 U19685 ( .A1(n16395), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16384) );
  OAI211_X1 U19686 ( .C1(n16392), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        n16387) );
  AOI21_X1 U19687 ( .B1(n16388), .B2(n19790), .A(n16387), .ZN(n16389) );
  OAI21_X1 U19688 ( .B1(n16815), .B2(n19770), .A(n16389), .ZN(P2_U2898) );
  NAND2_X1 U19689 ( .A1(n19731), .A2(n19786), .ZN(n16397) );
  OAI22_X1 U19690 ( .A1(n16390), .A2(n19863), .B1(n13513), .B2(n19768), .ZN(
        n16394) );
  INV_X1 U19691 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16391) );
  NOR2_X1 U19692 ( .A1(n16392), .A2(n16391), .ZN(n16393) );
  AOI211_X1 U19693 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n16395), .A(n16394), .B(
        n16393), .ZN(n16396) );
  OAI211_X1 U19694 ( .C1(n16399), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        P2_U2899) );
  AOI22_X1 U19695 ( .A1(n16408), .A2(n16400), .B1(n19785), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16402) );
  NAND2_X1 U19696 ( .A1(n16409), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16401) );
  OAI211_X1 U19697 ( .C1(n16413), .C2(n16403), .A(n16402), .B(n16401), .ZN(
        n16404) );
  AOI21_X1 U19698 ( .B1(n16405), .B2(n19790), .A(n16404), .ZN(n16406) );
  OAI21_X1 U19699 ( .B1(n16823), .B2(n19770), .A(n16406), .ZN(P2_U2900) );
  INV_X1 U19700 ( .A(n16836), .ZN(n16417) );
  AOI22_X1 U19701 ( .A1(n16408), .A2(n16407), .B1(n19785), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16411) );
  NAND2_X1 U19702 ( .A1(n16409), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16410) );
  OAI211_X1 U19703 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        n16414) );
  AOI21_X1 U19704 ( .B1(n16415), .B2(n19790), .A(n16414), .ZN(n16416) );
  OAI21_X1 U19705 ( .B1(n16417), .B2(n19770), .A(n16416), .ZN(P2_U2901) );
  INV_X1 U19706 ( .A(n17328), .ZN(n16425) );
  INV_X1 U19707 ( .A(n20502), .ZN(n19778) );
  XOR2_X1 U19708 ( .A(n20502), .B(n20169), .Z(n19781) );
  OAI21_X1 U19709 ( .B1(n20508), .B2(n20510), .A(n16418), .ZN(n19780) );
  NAND2_X1 U19710 ( .A1(n19781), .A2(n19780), .ZN(n19779) );
  OAI21_X1 U19711 ( .B1(n20498), .B2(n19778), .A(n19779), .ZN(n16419) );
  NAND2_X1 U19712 ( .A1(n16419), .A2(n19771), .ZN(n19774) );
  INV_X1 U19713 ( .A(n19773), .ZN(n16420) );
  NAND3_X1 U19714 ( .A1(n19774), .A2(n16420), .A3(n19790), .ZN(n16423) );
  AOI22_X1 U19715 ( .A1(n16421), .A2(n19866), .B1(n19785), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n16422) );
  OAI211_X1 U19716 ( .C1(n16425), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        P2_U2914) );
  OAI21_X1 U19717 ( .B1(n16427), .B2(n16728), .A(n16727), .ZN(n16428) );
  NAND2_X1 U19718 ( .A1(n9902), .A2(n16428), .ZN(n16733) );
  NAND2_X1 U19719 ( .A1(n16431), .A2(n16430), .ZN(n16432) );
  XNOR2_X1 U19720 ( .A(n16429), .B(n16432), .ZN(n16732) );
  NAND2_X1 U19721 ( .A1(n16723), .A2(n16719), .ZN(n16434) );
  NOR2_X1 U19722 ( .A1(n17339), .A2(n20479), .ZN(n16730) );
  AOI21_X1 U19723 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16730), .ZN(n16433) );
  OAI211_X1 U19724 ( .C1(n16717), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        n16436) );
  OAI21_X1 U19725 ( .B1(n16722), .B2(n16733), .A(n16437), .ZN(P2_U2985) );
  XNOR2_X1 U19726 ( .A(n16442), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16443) );
  NOR2_X1 U19727 ( .A1(n17339), .A2(n16444), .ZN(n16736) );
  NOR2_X1 U19728 ( .A1(n16445), .A2(n16717), .ZN(n16446) );
  AOI211_X1 U19729 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n16714), .A(
        n16736), .B(n16446), .ZN(n16447) );
  OAI21_X1 U19730 ( .B1(n16739), .B2(n16682), .A(n16447), .ZN(n16448) );
  AOI21_X1 U19731 ( .B1(n16704), .B2(n16740), .A(n16448), .ZN(n16449) );
  INV_X1 U19732 ( .A(n16427), .ZN(n16452) );
  NOR2_X1 U19733 ( .A1(n17339), .A2(n20476), .ZN(n16743) );
  AOI21_X1 U19734 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16743), .ZN(n16453) );
  OAI21_X1 U19735 ( .B1(n16454), .B2(n16717), .A(n16453), .ZN(n16456) );
  NOR2_X1 U19736 ( .A1(n16748), .A2(n16682), .ZN(n16455) );
  INV_X1 U19737 ( .A(n16462), .ZN(n16463) );
  XNOR2_X1 U19738 ( .A(n16464), .B(n16463), .ZN(n16765) );
  NOR2_X1 U19739 ( .A1(n17339), .A2(n20473), .ZN(n16755) );
  NOR2_X1 U19740 ( .A1(n16465), .A2(n16717), .ZN(n16466) );
  AOI211_X1 U19741 ( .C1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n16714), .A(
        n16755), .B(n16466), .ZN(n16467) );
  OAI21_X1 U19742 ( .B1(n16752), .B2(n16682), .A(n16467), .ZN(n16468) );
  AOI21_X1 U19743 ( .B1(n16713), .B2(n16765), .A(n16468), .ZN(n16469) );
  OAI21_X1 U19744 ( .B1(n16768), .B2(n16722), .A(n16469), .ZN(P2_U2988) );
  OAI21_X1 U19745 ( .B1(n16483), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16470), .ZN(n16780) );
  NAND2_X1 U19746 ( .A1(n13136), .A2(n16493), .ZN(n16489) );
  XNOR2_X1 U19747 ( .A(n16471), .B(n21670), .ZN(n16488) );
  NAND2_X1 U19748 ( .A1(n16489), .A2(n16488), .ZN(n16790) );
  OAI21_X1 U19749 ( .B1(n16472), .B2(n21670), .A(n16790), .ZN(n16476) );
  NAND2_X1 U19750 ( .A1(n16474), .A2(n16473), .ZN(n16475) );
  NAND2_X1 U19751 ( .A1(n16777), .A2(n16719), .ZN(n16479) );
  INV_X1 U19752 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16477) );
  NOR2_X1 U19753 ( .A1(n17339), .A2(n16477), .ZN(n16770) );
  AOI21_X1 U19754 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16770), .ZN(n16478) );
  OAI211_X1 U19755 ( .C1(n16717), .C2(n16480), .A(n16479), .B(n16478), .ZN(
        n16481) );
  AOI21_X1 U19756 ( .B1(n16713), .B2(n16778), .A(n16481), .ZN(n16482) );
  OAI21_X1 U19757 ( .B1(n16722), .B2(n16780), .A(n16482), .ZN(P2_U2990) );
  NOR2_X1 U19758 ( .A1(n16511), .A2(n16798), .ZN(n16496) );
  INV_X1 U19759 ( .A(n16483), .ZN(n16484) );
  OAI21_X1 U19760 ( .B1(n16496), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16484), .ZN(n16794) );
  INV_X1 U19761 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20468) );
  NOR2_X1 U19762 ( .A1(n17339), .A2(n20468), .ZN(n16783) );
  AOI21_X1 U19763 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16783), .ZN(n16485) );
  OAI21_X1 U19764 ( .B1(n16486), .B2(n16717), .A(n16485), .ZN(n16487) );
  AOI21_X1 U19765 ( .B1(n16789), .B2(n16719), .A(n16487), .ZN(n16491) );
  OR2_X1 U19766 ( .A1(n16489), .A2(n16488), .ZN(n16791) );
  NAND3_X1 U19767 ( .A1(n16791), .A2(n16790), .A3(n16713), .ZN(n16490) );
  OAI211_X1 U19768 ( .C1(n16794), .C2(n16722), .A(n16491), .B(n16490), .ZN(
        P2_U2991) );
  NAND2_X1 U19769 ( .A1(n16493), .A2(n16492), .ZN(n16495) );
  XOR2_X1 U19770 ( .A(n16495), .B(n16494), .Z(n16808) );
  INV_X1 U19771 ( .A(n16496), .ZN(n16796) );
  NAND2_X1 U19772 ( .A1(n16511), .A2(n16798), .ZN(n16795) );
  NAND3_X1 U19773 ( .A1(n16796), .A2(n16704), .A3(n16795), .ZN(n16501) );
  NOR2_X1 U19774 ( .A1(n17339), .A2(n20466), .ZN(n16797) );
  AOI21_X1 U19775 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16797), .ZN(n16497) );
  OAI21_X1 U19776 ( .B1(n16498), .B2(n16717), .A(n16497), .ZN(n16499) );
  AOI21_X1 U19777 ( .B1(n16805), .B2(n16719), .A(n16499), .ZN(n16500) );
  OAI211_X1 U19778 ( .C1(n16808), .C2(n16707), .A(n16501), .B(n16500), .ZN(
        P2_U2992) );
  INV_X1 U19779 ( .A(n16502), .ZN(n16503) );
  NAND2_X1 U19780 ( .A1(n16507), .A2(n16506), .ZN(n16508) );
  NAND2_X1 U19781 ( .A1(n19745), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U19782 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16509) );
  OAI211_X1 U19783 ( .C1(n16510), .C2(n16717), .A(n16813), .B(n16509), .ZN(
        n16512) );
  INV_X1 U19784 ( .A(n16529), .ZN(n16514) );
  NAND2_X1 U19785 ( .A1(n16516), .A2(n16515), .ZN(n16517) );
  XNOR2_X1 U19786 ( .A(n16518), .B(n16517), .ZN(n16833) );
  INV_X1 U19787 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21594) );
  NOR2_X1 U19788 ( .A1(n17339), .A2(n21594), .ZN(n16821) );
  AOI21_X1 U19789 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16821), .ZN(n16519) );
  OAI21_X1 U19790 ( .B1(n16717), .B2(n16520), .A(n16519), .ZN(n16521) );
  AOI21_X1 U19791 ( .B1(n16829), .B2(n16719), .A(n16521), .ZN(n16523) );
  OAI211_X1 U19792 ( .C1(n16833), .C2(n16707), .A(n16523), .B(n16522), .ZN(
        P2_U2995) );
  INV_X1 U19793 ( .A(n16524), .ZN(n16525) );
  NAND2_X1 U19794 ( .A1(n16530), .A2(n16529), .ZN(n16531) );
  NAND2_X1 U19795 ( .A1(n19745), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16838) );
  OAI21_X1 U19796 ( .B1(n16700), .B2(n16532), .A(n16838), .ZN(n16533) );
  AOI21_X1 U19797 ( .B1(n16697), .B2(n16534), .A(n16533), .ZN(n16535) );
  OAI21_X1 U19798 ( .B1(n16839), .B2(n16682), .A(n16535), .ZN(n16536) );
  AOI21_X1 U19799 ( .B1(n16842), .B2(n16713), .A(n16536), .ZN(n16537) );
  XNOR2_X1 U19800 ( .A(n16846), .B(n16861), .ZN(n16546) );
  XOR2_X1 U19801 ( .A(n16539), .B(n16538), .Z(n16857) );
  NAND2_X1 U19802 ( .A1(n16540), .A2(n16719), .ZN(n16542) );
  NOR2_X1 U19803 ( .A1(n17339), .A2(n20459), .ZN(n16852) );
  AOI21_X1 U19804 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16852), .ZN(n16541) );
  OAI211_X1 U19805 ( .C1(n16717), .C2(n16543), .A(n16542), .B(n16541), .ZN(
        n16544) );
  AOI21_X1 U19806 ( .B1(n16857), .B2(n16713), .A(n16544), .ZN(n16545) );
  OAI21_X1 U19807 ( .B1(n16722), .B2(n16546), .A(n16545), .ZN(P2_U2997) );
  XNOR2_X1 U19808 ( .A(n16556), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16555) );
  XOR2_X1 U19809 ( .A(n16548), .B(n16547), .Z(n16862) );
  NAND2_X1 U19810 ( .A1(n16549), .A2(n16719), .ZN(n16551) );
  NOR2_X1 U19811 ( .A1(n17339), .A2(n20457), .ZN(n16863) );
  AOI21_X1 U19812 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16863), .ZN(n16550) );
  OAI211_X1 U19813 ( .C1(n16717), .C2(n16552), .A(n16551), .B(n16550), .ZN(
        n16553) );
  AOI21_X1 U19814 ( .B1(n16862), .B2(n16713), .A(n16553), .ZN(n16554) );
  OAI21_X1 U19815 ( .B1(n16555), .B2(n16722), .A(n16554), .ZN(P2_U2998) );
  OAI21_X1 U19816 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16557), .A(
        n16859), .ZN(n16880) );
  NAND2_X1 U19817 ( .A1(n16559), .A2(n16558), .ZN(n16561) );
  XOR2_X1 U19818 ( .A(n16561), .B(n16560), .Z(n16878) );
  NAND2_X1 U19819 ( .A1(n19745), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16869) );
  OAI21_X1 U19820 ( .B1(n16700), .B2(n16562), .A(n16869), .ZN(n16563) );
  AOI21_X1 U19821 ( .B1(n16697), .B2(n10543), .A(n16563), .ZN(n16564) );
  OAI21_X1 U19822 ( .B1(n16868), .B2(n16682), .A(n16564), .ZN(n16565) );
  AOI21_X1 U19823 ( .B1(n16878), .B2(n16713), .A(n16565), .ZN(n16566) );
  OAI21_X1 U19824 ( .B1(n16880), .B2(n16722), .A(n16566), .ZN(P2_U2999) );
  OAI21_X1 U19825 ( .B1(n16568), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16567), .ZN(n16893) );
  NAND2_X1 U19826 ( .A1(n16570), .A2(n16569), .ZN(n16571) );
  XNOR2_X1 U19827 ( .A(n16572), .B(n16571), .ZN(n16890) );
  NAND2_X1 U19828 ( .A1(n19745), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16883) );
  OAI21_X1 U19829 ( .B1(n16700), .B2(n16573), .A(n16883), .ZN(n16574) );
  AOI21_X1 U19830 ( .B1(n16697), .B2(n16575), .A(n16574), .ZN(n16576) );
  OAI21_X1 U19831 ( .B1(n16884), .B2(n16682), .A(n16576), .ZN(n16577) );
  AOI21_X1 U19832 ( .B1(n16890), .B2(n16713), .A(n16577), .ZN(n16578) );
  OAI21_X1 U19833 ( .B1(n16893), .B2(n16722), .A(n16578), .ZN(P2_U3000) );
  NAND2_X1 U19834 ( .A1(n16579), .A2(n16704), .ZN(n16586) );
  NAND2_X1 U19835 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16580) );
  OAI211_X1 U19836 ( .C1(n16717), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        n16583) );
  AOI21_X1 U19837 ( .B1(n16584), .B2(n16719), .A(n16583), .ZN(n16585) );
  OAI211_X1 U19838 ( .C1(n16707), .C2(n16587), .A(n16586), .B(n16585), .ZN(
        P2_U3001) );
  OAI21_X1 U19839 ( .B1(n16601), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16588), .ZN(n16906) );
  OAI21_X1 U19840 ( .B1(n16591), .B2(n16590), .A(n16589), .ZN(n16904) );
  NOR2_X1 U19841 ( .A1(n17339), .A2(n20449), .ZN(n16894) );
  NOR2_X1 U19842 ( .A1(n16717), .A2(n16592), .ZN(n16593) );
  AOI211_X1 U19843 ( .C1(n16714), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16894), .B(n16593), .ZN(n16594) );
  OAI21_X1 U19844 ( .B1(n16897), .B2(n16682), .A(n16594), .ZN(n16595) );
  AOI21_X1 U19845 ( .B1(n16904), .B2(n16713), .A(n16595), .ZN(n16596) );
  OAI21_X1 U19846 ( .B1(n16906), .B2(n16722), .A(n16596), .ZN(P2_U3002) );
  NAND2_X1 U19847 ( .A1(n16598), .A2(n16597), .ZN(n16599) );
  XNOR2_X1 U19848 ( .A(n16600), .B(n16599), .ZN(n16918) );
  NAND2_X1 U19849 ( .A1(n16907), .A2(n16704), .ZN(n16608) );
  OR2_X1 U19850 ( .A1(n17339), .A2(n20447), .ZN(n16909) );
  OAI21_X1 U19851 ( .B1(n16700), .B2(n16602), .A(n16909), .ZN(n16605) );
  NOR2_X1 U19852 ( .A1(n16603), .A2(n16682), .ZN(n16604) );
  AOI211_X1 U19853 ( .C1(n16697), .C2(n16606), .A(n16605), .B(n16604), .ZN(
        n16607) );
  INV_X1 U19854 ( .A(n16610), .ZN(n16613) );
  OAI21_X1 U19855 ( .B1(n16613), .B2(n16611), .A(n16612), .ZN(n16614) );
  NAND2_X1 U19856 ( .A1(n16614), .A2(n16627), .ZN(n16618) );
  NAND2_X1 U19857 ( .A1(n16616), .A2(n16615), .ZN(n16617) );
  XNOR2_X1 U19858 ( .A(n16618), .B(n16617), .ZN(n16927) );
  NOR2_X1 U19859 ( .A1(n17339), .A2(n20446), .ZN(n16920) );
  NOR2_X1 U19860 ( .A1(n16700), .A2(n16619), .ZN(n16620) );
  AOI211_X1 U19861 ( .C1(n16621), .C2(n16697), .A(n16920), .B(n16620), .ZN(
        n16622) );
  OAI21_X1 U19862 ( .B1(n16623), .B2(n16682), .A(n16622), .ZN(n16624) );
  AOI21_X1 U19863 ( .B1(n16927), .B2(n16713), .A(n16624), .ZN(n16625) );
  OAI21_X1 U19864 ( .B1(n16929), .B2(n16722), .A(n16625), .ZN(P2_U3004) );
  NAND2_X1 U19865 ( .A1(n16628), .A2(n16627), .ZN(n16633) );
  NAND2_X1 U19866 ( .A1(n16610), .A2(n16629), .ZN(n16659) );
  OAI21_X1 U19867 ( .B1(n16659), .B2(n10266), .A(n16631), .ZN(n16632) );
  XOR2_X1 U19868 ( .A(n16633), .B(n16632), .Z(n16938) );
  NOR2_X1 U19869 ( .A1(n17339), .A2(n20444), .ZN(n16931) );
  NOR2_X1 U19870 ( .A1(n16717), .A2(n16634), .ZN(n16635) );
  AOI211_X1 U19871 ( .C1(n16714), .C2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16931), .B(n16635), .ZN(n16636) );
  OAI21_X1 U19872 ( .B1(n16935), .B2(n16682), .A(n16636), .ZN(n16637) );
  AOI21_X1 U19873 ( .B1(n16938), .B2(n16713), .A(n16637), .ZN(n16638) );
  OAI21_X1 U19874 ( .B1(n16941), .B2(n16722), .A(n16638), .ZN(P2_U3005) );
  INV_X1 U19875 ( .A(n16656), .ZN(n16639) );
  AOI21_X1 U19876 ( .B1(n16659), .B2(n16657), .A(n16639), .ZN(n16643) );
  NAND2_X1 U19877 ( .A1(n16641), .A2(n16640), .ZN(n16642) );
  XNOR2_X1 U19878 ( .A(n16643), .B(n16642), .ZN(n16953) );
  OR2_X1 U19879 ( .A1(n16645), .A2(n16644), .ZN(n16942) );
  NAND3_X1 U19880 ( .A1(n16942), .A2(n16704), .A3(n16646), .ZN(n16652) );
  INV_X1 U19881 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20442) );
  NOR2_X1 U19882 ( .A1(n17339), .A2(n20442), .ZN(n16945) );
  AOI21_X1 U19883 ( .B1(n16714), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16945), .ZN(n16647) );
  OAI21_X1 U19884 ( .B1(n16717), .B2(n16648), .A(n16647), .ZN(n16649) );
  AOI21_X1 U19885 ( .B1(n16650), .B2(n16719), .A(n16649), .ZN(n16651) );
  OAI211_X1 U19886 ( .C1(n16953), .C2(n16707), .A(n16652), .B(n16651), .ZN(
        P2_U3006) );
  XNOR2_X1 U19887 ( .A(n16654), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16655) );
  XNOR2_X1 U19888 ( .A(n16653), .B(n16655), .ZN(n16966) );
  NAND2_X1 U19889 ( .A1(n16657), .A2(n16656), .ZN(n16658) );
  XNOR2_X1 U19890 ( .A(n16659), .B(n16658), .ZN(n16964) );
  NAND2_X1 U19891 ( .A1(n19745), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16956) );
  OAI21_X1 U19892 ( .B1(n16700), .B2(n16660), .A(n16956), .ZN(n16661) );
  AOI21_X1 U19893 ( .B1(n16697), .B2(n16662), .A(n16661), .ZN(n16663) );
  OAI21_X1 U19894 ( .B1(n16955), .B2(n16682), .A(n16663), .ZN(n16664) );
  AOI21_X1 U19895 ( .B1(n16964), .B2(n16713), .A(n16664), .ZN(n16665) );
  OAI21_X1 U19896 ( .B1(n16966), .B2(n16722), .A(n16665), .ZN(P2_U3007) );
  OAI21_X1 U19897 ( .B1(n16666), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16667), .ZN(n16976) );
  NAND2_X1 U19898 ( .A1(n16697), .A2(n19755), .ZN(n16668) );
  NAND2_X1 U19899 ( .A1(n19745), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16968) );
  OAI211_X1 U19900 ( .C1(n16700), .C2(n16669), .A(n16668), .B(n16968), .ZN(
        n16673) );
  XNOR2_X1 U19901 ( .A(n16671), .B(n16670), .ZN(n16970) );
  NOR2_X1 U19902 ( .A1(n16970), .A2(n16707), .ZN(n16672) );
  AOI211_X1 U19903 ( .C1(n16719), .C2(n19762), .A(n16673), .B(n16672), .ZN(
        n16674) );
  OAI21_X1 U19904 ( .B1(n16722), .B2(n16976), .A(n16674), .ZN(P2_U3008) );
  OAI21_X1 U19905 ( .B1(n16678), .B2(n16676), .A(n16675), .ZN(n16677) );
  INV_X1 U19906 ( .A(n16679), .ZN(n16681) );
  XNOR2_X1 U19907 ( .A(n16681), .B(n16680), .ZN(n17335) );
  NOR2_X1 U19908 ( .A1(n17331), .A2(n16682), .ZN(n16686) );
  AOI22_X1 U19909 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19745), .ZN(n16683) );
  OAI21_X1 U19910 ( .B1(n16717), .B2(n16684), .A(n16683), .ZN(n16685) );
  AOI211_X1 U19911 ( .C1(n17335), .C2(n16713), .A(n16686), .B(n16685), .ZN(
        n16687) );
  OAI21_X1 U19912 ( .B1(n17332), .B2(n16722), .A(n16687), .ZN(P2_U3009) );
  INV_X1 U19913 ( .A(n16688), .ZN(n16689) );
  OAI21_X1 U19914 ( .B1(n10329), .B2(n16690), .A(n16689), .ZN(n16712) );
  INV_X1 U19915 ( .A(n16712), .ZN(n16691) );
  NAND2_X1 U19916 ( .A1(n16691), .A2(n17354), .ZN(n16692) );
  AOI22_X1 U19917 ( .A1(n16712), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16692), .B2(n16710), .ZN(n16695) );
  XNOR2_X1 U19918 ( .A(n16693), .B(n16703), .ZN(n16694) );
  XNOR2_X1 U19919 ( .A(n16695), .B(n16694), .ZN(n16989) );
  NAND2_X1 U19920 ( .A1(n16697), .A2(n16696), .ZN(n16698) );
  INV_X1 U19921 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20434) );
  NAND2_X1 U19922 ( .A1(n19745), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n16977) );
  OAI211_X1 U19923 ( .C1(n16700), .C2(n16699), .A(n16698), .B(n16977), .ZN(
        n16701) );
  AOI21_X1 U19924 ( .B1(n16983), .B2(n16719), .A(n16701), .ZN(n16706) );
  NAND2_X1 U19925 ( .A1(n16985), .A2(n16704), .ZN(n16705) );
  OAI211_X1 U19926 ( .C1(n16989), .C2(n16707), .A(n16706), .B(n16705), .ZN(
        P2_U3010) );
  XNOR2_X1 U19927 ( .A(n16709), .B(n16708), .ZN(n17349) );
  XNOR2_X1 U19928 ( .A(n16710), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16711) );
  XNOR2_X1 U19929 ( .A(n16712), .B(n16711), .ZN(n17352) );
  NAND2_X1 U19930 ( .A1(n17352), .A2(n16713), .ZN(n16721) );
  AOI22_X1 U19931 ( .A1(n16714), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19745), .ZN(n16715) );
  OAI21_X1 U19932 ( .B1(n16717), .B2(n16716), .A(n16715), .ZN(n16718) );
  AOI21_X1 U19933 ( .B1(n17345), .B2(n16719), .A(n16718), .ZN(n16720) );
  OAI211_X1 U19934 ( .C1(n17349), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        P2_U3011) );
  NAND2_X1 U19935 ( .A1(n16724), .A2(n16745), .ZN(n16744) );
  AOI21_X1 U19936 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16727), .A(
        n16728), .ZN(n16726) );
  INV_X1 U19937 ( .A(n16724), .ZN(n16725) );
  NOR2_X1 U19938 ( .A1(n16734), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16735) );
  OAI21_X1 U19939 ( .B1(n16742), .B2(n16988), .A(n16741), .ZN(P2_U3018) );
  OAI21_X1 U19940 ( .B1(n16751), .B2(n16988), .A(n16750), .ZN(P2_U3019) );
  INV_X1 U19941 ( .A(n16752), .ZN(n16764) );
  OAI21_X1 U19942 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16753), .ZN(n16754) );
  INV_X1 U19943 ( .A(n16754), .ZN(n16756) );
  AOI21_X1 U19944 ( .B1(n16757), .B2(n16756), .A(n16755), .ZN(n16761) );
  OR2_X1 U19945 ( .A1(n16759), .A2(n16758), .ZN(n16760) );
  OAI211_X1 U19946 ( .C1(n16762), .C2(n17340), .A(n16761), .B(n16760), .ZN(
        n16763) );
  AOI21_X1 U19947 ( .B1(n16764), .B2(n17346), .A(n16763), .ZN(n16767) );
  NAND2_X1 U19948 ( .A1(n16765), .A2(n17351), .ZN(n16766) );
  OAI211_X1 U19949 ( .C1(n16768), .C2(n17348), .A(n16767), .B(n16766), .ZN(
        P2_U3020) );
  INV_X1 U19950 ( .A(n16781), .ZN(n16799) );
  NOR2_X1 U19951 ( .A1(n16769), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16771) );
  AOI21_X1 U19952 ( .B1(n16799), .B2(n16771), .A(n16770), .ZN(n16774) );
  NAND3_X1 U19953 ( .A1(n16772), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16800), .ZN(n16773) );
  OAI211_X1 U19954 ( .C1(n16775), .C2(n17340), .A(n16774), .B(n16773), .ZN(
        n16776) );
  AOI21_X1 U19955 ( .B1(n16777), .B2(n17346), .A(n16776), .ZN(n16779) );
  AOI211_X1 U19956 ( .C1(n21670), .C2(n16798), .A(n16782), .B(n16781), .ZN(
        n16784) );
  NOR2_X1 U19957 ( .A1(n16784), .A2(n16783), .ZN(n16786) );
  NAND3_X1 U19958 ( .A1(n16812), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16800), .ZN(n16785) );
  OAI211_X1 U19959 ( .C1(n16787), .C2(n17340), .A(n16786), .B(n16785), .ZN(
        n16788) );
  AOI21_X1 U19960 ( .B1(n17346), .B2(n16789), .A(n16788), .ZN(n16793) );
  NAND3_X1 U19961 ( .A1(n16791), .A2(n16790), .A3(n17351), .ZN(n16792) );
  OAI211_X1 U19962 ( .C1(n16794), .C2(n17348), .A(n16793), .B(n16792), .ZN(
        P2_U3023) );
  NAND3_X1 U19963 ( .A1(n16796), .A2(n16984), .A3(n16795), .ZN(n16807) );
  AOI21_X1 U19964 ( .B1(n16799), .B2(n16798), .A(n16797), .ZN(n16802) );
  NAND3_X1 U19965 ( .A1(n16812), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n16800), .ZN(n16801) );
  OAI211_X1 U19966 ( .C1(n16803), .C2(n17340), .A(n16802), .B(n16801), .ZN(
        n16804) );
  AOI21_X1 U19967 ( .B1(n16805), .B2(n17346), .A(n16804), .ZN(n16806) );
  OAI211_X1 U19968 ( .C1(n16808), .C2(n16988), .A(n16807), .B(n16806), .ZN(
        P2_U3024) );
  OAI21_X1 U19969 ( .B1(n16824), .B2(n16810), .A(n16809), .ZN(n16811) );
  NAND2_X1 U19970 ( .A1(n16812), .A2(n16811), .ZN(n16814) );
  OAI211_X1 U19971 ( .C1(n17340), .C2(n16815), .A(n16814), .B(n16813), .ZN(
        n16817) );
  INV_X1 U19972 ( .A(n16821), .ZN(n16822) );
  OAI21_X1 U19973 ( .B1(n16823), .B2(n17340), .A(n16822), .ZN(n16828) );
  INV_X1 U19974 ( .A(n16824), .ZN(n16826) );
  MUX2_X1 U19975 ( .A(n16834), .B(n16826), .S(n16825), .Z(n16827) );
  AOI211_X1 U19976 ( .C1(n16829), .C2(n17346), .A(n16828), .B(n16827), .ZN(
        n16832) );
  NAND2_X1 U19977 ( .A1(n16873), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16858) );
  INV_X1 U19978 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16851) );
  NOR3_X1 U19979 ( .A1(n16858), .A2(n16861), .A3(n16851), .ZN(n16835) );
  MUX2_X1 U19980 ( .A(n16835), .B(n16834), .S(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Z(n16841) );
  NAND2_X1 U19981 ( .A1(n16836), .A2(n17327), .ZN(n16837) );
  OAI211_X1 U19982 ( .C1(n16839), .C2(n17330), .A(n16838), .B(n16837), .ZN(
        n16840) );
  OR2_X1 U19983 ( .A1(n16984), .A2(n16844), .ZN(n16845) );
  INV_X1 U19984 ( .A(n16847), .ZN(n16876) );
  AOI21_X1 U19985 ( .B1(n16853), .B2(n17327), .A(n16852), .ZN(n16854) );
  OAI21_X1 U19986 ( .B1(n16855), .B2(n17330), .A(n16854), .ZN(n16856) );
  AOI21_X1 U19987 ( .B1(n16857), .B2(n17351), .A(n16856), .ZN(n16860) );
  AOI21_X1 U19988 ( .B1(n16864), .B2(n17327), .A(n16863), .ZN(n16865) );
  NOR2_X1 U19989 ( .A1(n16868), .A2(n17330), .ZN(n16872) );
  OAI21_X1 U19990 ( .B1(n16870), .B2(n17340), .A(n16869), .ZN(n16871) );
  AOI211_X1 U19991 ( .C1(n16873), .C2(n16875), .A(n16872), .B(n16871), .ZN(
        n16874) );
  OAI21_X1 U19992 ( .B1(n16876), .B2(n16875), .A(n16874), .ZN(n16877) );
  AOI21_X1 U19993 ( .B1(n16878), .B2(n17351), .A(n16877), .ZN(n16879) );
  OAI21_X1 U19994 ( .B1(n16880), .B2(n17348), .A(n16879), .ZN(P2_U3031) );
  NAND2_X1 U19995 ( .A1(n16881), .A2(n17327), .ZN(n16882) );
  OAI211_X1 U19996 ( .C1(n16884), .C2(n17330), .A(n16883), .B(n16882), .ZN(
        n16888) );
  NOR3_X1 U19997 ( .A1(n16886), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16885), .ZN(n16887) );
  AOI211_X1 U19998 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16889), .A(
        n16888), .B(n16887), .ZN(n16892) );
  NAND2_X1 U19999 ( .A1(n16890), .A2(n17351), .ZN(n16891) );
  OAI211_X1 U20000 ( .C1(n16893), .C2(n17348), .A(n16892), .B(n16891), .ZN(
        P2_U3032) );
  AOI21_X1 U20001 ( .B1(n16895), .B2(n17327), .A(n16894), .ZN(n16896) );
  OAI21_X1 U20002 ( .B1(n16897), .B2(n17330), .A(n16896), .ZN(n16898) );
  AOI21_X1 U20003 ( .B1(n16899), .B2(n16901), .A(n16898), .ZN(n16900) );
  OAI21_X1 U20004 ( .B1(n16902), .B2(n16901), .A(n16900), .ZN(n16903) );
  AOI21_X1 U20005 ( .B1(n16904), .B2(n17351), .A(n16903), .ZN(n16905) );
  OAI21_X1 U20006 ( .B1(n16906), .B2(n17348), .A(n16905), .ZN(P2_U3034) );
  NAND2_X1 U20007 ( .A1(n16908), .A2(n17346), .ZN(n16910) );
  OAI211_X1 U20008 ( .C1(n17340), .C2(n16911), .A(n16910), .B(n16909), .ZN(
        n16913) );
  NAND3_X1 U20009 ( .A1(n9727), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16919), .ZN(n16923) );
  AOI21_X1 U20010 ( .B1(n9662), .B2(n16923), .A(n16914), .ZN(n16912) );
  AOI211_X1 U20011 ( .C1(n16915), .C2(n16914), .A(n16913), .B(n16912), .ZN(
        n16916) );
  OAI211_X1 U20012 ( .C1(n16918), .C2(n16988), .A(n16917), .B(n16916), .ZN(
        P2_U3035) );
  NOR2_X1 U20013 ( .A1(n9662), .A2(n16919), .ZN(n16926) );
  AOI21_X1 U20014 ( .B1(n16921), .B2(n17346), .A(n16920), .ZN(n16922) );
  OAI211_X1 U20015 ( .C1(n16924), .C2(n17340), .A(n16923), .B(n16922), .ZN(
        n16925) );
  AOI211_X1 U20016 ( .C1(n16927), .C2(n17351), .A(n16926), .B(n16925), .ZN(
        n16928) );
  OAI21_X1 U20017 ( .B1(n16929), .B2(n17348), .A(n16928), .ZN(P2_U3036) );
  NAND2_X1 U20018 ( .A1(n9727), .A2(n16930), .ZN(n16934) );
  AOI21_X1 U20019 ( .B1(n16932), .B2(n17327), .A(n16931), .ZN(n16933) );
  OAI211_X1 U20020 ( .C1(n16935), .C2(n17330), .A(n16934), .B(n16933), .ZN(
        n16936) );
  AOI21_X1 U20021 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16937), .A(
        n16936), .ZN(n16940) );
  NAND2_X1 U20022 ( .A1(n16938), .A2(n17351), .ZN(n16939) );
  OAI211_X1 U20023 ( .C1(n16941), .C2(n17348), .A(n16940), .B(n16939), .ZN(
        P2_U3037) );
  NAND3_X1 U20024 ( .A1(n16942), .A2(n16984), .A3(n16646), .ZN(n16952) );
  INV_X1 U20025 ( .A(n16962), .ZN(n16944) );
  OAI211_X1 U20026 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16944), .B(n16943), .ZN(n16948) );
  AOI21_X1 U20027 ( .B1(n16946), .B2(n17327), .A(n16945), .ZN(n16947) );
  OAI211_X1 U20028 ( .C1(n16949), .C2(n17330), .A(n16948), .B(n16947), .ZN(
        n16950) );
  AOI21_X1 U20029 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16954), .A(
        n16950), .ZN(n16951) );
  OAI211_X1 U20030 ( .C1(n16953), .C2(n16988), .A(n16952), .B(n16951), .ZN(
        P2_U3038) );
  NAND2_X1 U20031 ( .A1(n16954), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16961) );
  INV_X1 U20032 ( .A(n16955), .ZN(n16959) );
  OAI21_X1 U20033 ( .B1(n16957), .B2(n17340), .A(n16956), .ZN(n16958) );
  AOI21_X1 U20034 ( .B1(n16959), .B2(n17346), .A(n16958), .ZN(n16960) );
  OAI211_X1 U20035 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16962), .A(
        n16961), .B(n16960), .ZN(n16963) );
  AOI21_X1 U20036 ( .B1(n16964), .B2(n17351), .A(n16963), .ZN(n16965) );
  OAI21_X1 U20037 ( .B1(n16966), .B2(n17348), .A(n16965), .ZN(P2_U3039) );
  AOI22_X1 U20038 ( .A1(n19762), .A2(n17346), .B1(n17327), .B2(n19759), .ZN(
        n16969) );
  OAI211_X1 U20039 ( .C1(n16967), .C2(n16973), .A(n16969), .B(n16968), .ZN(
        n16972) );
  NOR2_X1 U20040 ( .A1(n16970), .A2(n16988), .ZN(n16971) );
  AOI211_X1 U20041 ( .C1(n16974), .C2(n16973), .A(n16972), .B(n16971), .ZN(
        n16975) );
  OAI21_X1 U20042 ( .B1(n17348), .B2(n16976), .A(n16975), .ZN(P2_U3040) );
  OAI21_X1 U20043 ( .B1(n19771), .B2(n17340), .A(n16977), .ZN(n16982) );
  INV_X1 U20044 ( .A(n16978), .ZN(n16979) );
  MUX2_X1 U20045 ( .A(n16980), .B(n16979), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n16981) );
  AOI211_X1 U20046 ( .C1(n16983), .C2(n17346), .A(n16982), .B(n16981), .ZN(
        n16987) );
  NAND2_X1 U20047 ( .A1(n16985), .A2(n16984), .ZN(n16986) );
  OAI211_X1 U20048 ( .C1(n16989), .C2(n16988), .A(n16987), .B(n16986), .ZN(
        P2_U3042) );
  INV_X1 U20049 ( .A(n17016), .ZN(n16994) );
  MUX2_X1 U20050 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16990), .S(
        n19753), .Z(n16999) );
  OAI222_X1 U20051 ( .A1(n16994), .A2(n16993), .B1(n16992), .B2(n16999), .C1(
        n20493), .C2(n16991), .ZN(n16995) );
  MUX2_X1 U20052 ( .A(n16995), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n17010), .Z(P2_U3601) );
  NAND2_X1 U20053 ( .A1(n16996), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16997) );
  NAND2_X1 U20054 ( .A1(n16998), .A2(n16997), .ZN(n17007) );
  NAND2_X1 U20055 ( .A1(n16999), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20056 ( .A1(n20494), .A2(n17016), .B1(n17050), .B2(n17000), .ZN(
        n17001) );
  OAI21_X1 U20057 ( .B1(n17007), .B2(n17005), .A(n17001), .ZN(n17003) );
  MUX2_X1 U20058 ( .A(n17004), .B(n17003), .S(n17002), .Z(P2_U3600) );
  INV_X1 U20059 ( .A(n17005), .ZN(n17006) );
  AOI222_X1 U20060 ( .A1(n17008), .A2(n17050), .B1(n20508), .B2(n17016), .C1(
        n17007), .C2(n17006), .ZN(n17011) );
  NAND2_X1 U20061 ( .A1(n17010), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17009) );
  OAI21_X1 U20062 ( .B1(n17011), .B2(n17010), .A(n17009), .ZN(P2_U3599) );
  OAI21_X1 U20063 ( .B1(n20018), .B2(n20008), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17012) );
  NAND2_X1 U20064 ( .A1(n17012), .A2(n19948), .ZN(n17021) );
  INV_X1 U20065 ( .A(n17013), .ZN(n20302) );
  NOR2_X1 U20066 ( .A1(n17014), .A2(n20302), .ZN(n20231) );
  NAND2_X1 U20067 ( .A1(n20231), .A2(n20505), .ZN(n17026) );
  NAND2_X1 U20068 ( .A1(n20505), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20079) );
  INV_X1 U20069 ( .A(n20079), .ZN(n20076) );
  NAND2_X1 U20070 ( .A1(n20076), .A2(n20521), .ZN(n17043) );
  NOR2_X1 U20071 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17043), .ZN(
        n20002) );
  OAI21_X1 U20072 ( .B1(n17022), .B2(n20002), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17015) );
  INV_X1 U20073 ( .A(n20009), .ZN(n17036) );
  OR2_X1 U20074 ( .A1(n20522), .A2(n20551), .ZN(n17017) );
  INV_X1 U20075 ( .A(n17019), .ZN(n17020) );
  NOR2_X2 U20076 ( .A1(n20265), .A2(n17020), .ZN(n20353) );
  INV_X1 U20077 ( .A(n20353), .ZN(n17035) );
  INV_X1 U20078 ( .A(n17021), .ZN(n17027) );
  INV_X1 U20079 ( .A(n17022), .ZN(n17023) );
  AOI21_X1 U20080 ( .B1(n17023), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n17024) );
  OAI21_X1 U20081 ( .B1(n17024), .B2(n20002), .A(n20361), .ZN(n17025) );
  AOI21_X2 U20082 ( .B1(n17027), .B2(n17026), .A(n17025), .ZN(n20013) );
  INV_X1 U20083 ( .A(n20013), .ZN(n17033) );
  AOI22_X1 U20084 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19883), .ZN(n20366) );
  NOR2_X1 U20085 ( .A1(n19978), .A2(n20366), .ZN(n17032) );
  AOI22_X1 U20086 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19883), .ZN(n20297) );
  NAND2_X1 U20087 ( .A1(n19880), .A2(n17030), .ZN(n20296) );
  INV_X1 U20088 ( .A(n20002), .ZN(n20006) );
  OAI22_X1 U20089 ( .A1(n20040), .A2(n20297), .B1(n20296), .B2(n20006), .ZN(
        n17031) );
  AOI211_X1 U20090 ( .C1(n17033), .C2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17032), .B(n17031), .ZN(n17034) );
  OAI21_X1 U20091 ( .B1(n17036), .B2(n17035), .A(n17034), .ZN(P2_U3080) );
  AOI21_X1 U20092 ( .B1(n17045), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20543), 
        .ZN(n17041) );
  NAND2_X1 U20093 ( .A1(n17041), .A2(n17043), .ZN(n17040) );
  NAND2_X1 U20094 ( .A1(n11082), .A2(n20501), .ZN(n17038) );
  NOR2_X1 U20095 ( .A1(n20260), .A2(n20079), .ZN(n20032) );
  INV_X1 U20096 ( .A(n20032), .ZN(n20043) );
  AND2_X1 U20097 ( .A1(n20543), .A2(n20043), .ZN(n17037) );
  AOI21_X1 U20098 ( .B1(n17038), .B2(n17037), .A(n20265), .ZN(n17039) );
  INV_X1 U20099 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17049) );
  INV_X1 U20100 ( .A(n17041), .ZN(n17044) );
  OAI21_X1 U20101 ( .B1(n11082), .B2(n20032), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17042) );
  INV_X1 U20102 ( .A(n20366), .ZN(n20241) );
  AOI22_X1 U20103 ( .A1(n20018), .A2(n20241), .B1(n20352), .B2(n20032), .ZN(
        n17046) );
  OAI21_X1 U20104 ( .B1(n20297), .B2(n20041), .A(n17046), .ZN(n17047) );
  AOI21_X1 U20105 ( .B1(n20036), .B2(n20353), .A(n17047), .ZN(n17048) );
  OAI21_X1 U20106 ( .B1(n20022), .B2(n17049), .A(n17048), .ZN(P2_U3088) );
  NAND2_X1 U20107 ( .A1(n17054), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17357) );
  NAND2_X1 U20108 ( .A1(n20547), .A2(n17050), .ZN(n17057) );
  NAND2_X1 U20109 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20553), .ZN(n17051) );
  AOI21_X1 U20110 ( .B1(n17054), .B2(n17052), .A(n17051), .ZN(n17053) );
  AOI211_X1 U20111 ( .C1(n17055), .C2(n17054), .A(n19757), .B(n17053), .ZN(
        n17056) );
  OAI21_X1 U20112 ( .B1(n17357), .B2(n17057), .A(n17056), .ZN(P2_U3177) );
  INV_X1 U20113 ( .A(n17182), .ZN(n17059) );
  INV_X1 U20114 ( .A(n17180), .ZN(n17058) );
  NOR2_X1 U20115 ( .A1(n18696), .A2(n17058), .ZN(n17086) );
  AOI21_X1 U20116 ( .B1(n17059), .B2(n18812), .A(n17086), .ZN(n17077) );
  AOI21_X1 U20117 ( .B1(n17061), .B2(n18663), .A(n17060), .ZN(n17062) );
  XNOR2_X1 U20118 ( .A(n17062), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17179) );
  NAND2_X1 U20119 ( .A1(n17179), .A2(n18714), .ZN(n17073) );
  NOR2_X1 U20120 ( .A1(n17063), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17070) );
  OR2_X1 U20121 ( .A1(n18745), .A2(n18985), .ZN(n17064) );
  OAI21_X2 U20122 ( .B1(n18696), .B2(n18664), .A(n17064), .ZN(n18724) );
  NAND2_X1 U20123 ( .A1(n13950), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17191) );
  OAI211_X1 U20124 ( .C1(n17068), .C2(n10310), .A(n17067), .B(n17191), .ZN(
        n17069) );
  AOI211_X1 U20125 ( .C1(n18730), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        n17072) );
  OAI211_X1 U20126 ( .C1(n17077), .C2(n17188), .A(n17073), .B(n17072), .ZN(
        P3_U2800) );
  XNOR2_X1 U20127 ( .A(n18663), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17224) );
  INV_X1 U20128 ( .A(n17114), .ZN(n17074) );
  NAND2_X1 U20129 ( .A1(n17074), .A2(n18644), .ZN(n17112) );
  INV_X1 U20130 ( .A(n17112), .ZN(n17075) );
  AOI211_X1 U20131 ( .C1(n18663), .C2(n17225), .A(n17224), .B(n17075), .ZN(
        n17076) );
  XNOR2_X1 U20132 ( .A(n17076), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17203) );
  INV_X1 U20133 ( .A(n17077), .ZN(n17092) );
  NAND2_X1 U20134 ( .A1(n17104), .A2(n17185), .ZN(n17213) );
  NOR3_X1 U20135 ( .A1(n17182), .A2(n17213), .A3(n18745), .ZN(n17091) );
  INV_X1 U20136 ( .A(n17472), .ZN(n17089) );
  OAI21_X1 U20137 ( .B1(n17079), .B2(n19136), .A(n17478), .ZN(n17084) );
  NOR2_X1 U20138 ( .A1(n19075), .A2(n19644), .ZN(n17194) );
  INV_X1 U20139 ( .A(n17080), .ZN(n17082) );
  NOR2_X1 U20140 ( .A1(n17082), .A2(n17081), .ZN(n17083) );
  AOI211_X1 U20141 ( .C1(n17085), .C2(n17084), .A(n17194), .B(n17083), .ZN(
        n17088) );
  NAND3_X1 U20142 ( .A1(n17086), .A2(n17185), .A3(n17237), .ZN(n17087) );
  OAI211_X1 U20143 ( .C1(n17089), .C2(n18706), .A(n17088), .B(n17087), .ZN(
        n17090) );
  AOI211_X1 U20144 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17092), .A(
        n17091), .B(n17090), .ZN(n17093) );
  OAI21_X1 U20145 ( .B1(n17203), .B2(n18732), .A(n17093), .ZN(P3_U2801) );
  NAND2_X1 U20146 ( .A1(n17112), .A2(n17225), .ZN(n17115) );
  NAND2_X1 U20147 ( .A1(n17115), .A2(n17224), .ZN(n17217) );
  OAI211_X1 U20148 ( .C1(n17115), .C2(n17224), .A(n17217), .B(n18714), .ZN(
        n17110) );
  INV_X1 U20149 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17094) );
  NAND3_X1 U20150 ( .A1(n17233), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17094), .ZN(n17102) );
  OAI21_X1 U20151 ( .B1(n14477), .B2(n9899), .A(n18807), .ZN(n17098) );
  INV_X1 U20152 ( .A(n17095), .ZN(n17096) );
  NOR2_X1 U20153 ( .A1(n17096), .A2(n19570), .ZN(n17097) );
  NOR2_X1 U20154 ( .A1(n17098), .A2(n17097), .ZN(n18532) );
  NAND2_X1 U20155 ( .A1(n18573), .A2(n10578), .ZN(n17099) );
  NAND2_X1 U20156 ( .A1(n18532), .A2(n17099), .ZN(n17116) );
  AND2_X1 U20157 ( .A1(n19022), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17226) );
  AOI21_X1 U20158 ( .B1(n17116), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17226), .ZN(n17101) );
  NAND2_X1 U20159 ( .A1(n18730), .A2(n17483), .ZN(n17100) );
  OAI211_X1 U20160 ( .C1(n18555), .C2(n17102), .A(n17101), .B(n17100), .ZN(
        n17103) );
  INV_X1 U20161 ( .A(n17103), .ZN(n17109) );
  OAI22_X1 U20162 ( .A1(n17104), .A2(n18745), .B1(n17237), .B2(n18696), .ZN(
        n18527) );
  OR2_X1 U20163 ( .A1(n18527), .A2(n17240), .ZN(n17120) );
  NAND2_X1 U20164 ( .A1(n18696), .A2(n18745), .ZN(n18594) );
  NAND3_X1 U20165 ( .A1(n17120), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18594), .ZN(n17108) );
  INV_X1 U20166 ( .A(n14477), .ZN(n17105) );
  NOR2_X1 U20167 ( .A1(n18649), .A2(n17105), .ZN(n17121) );
  OAI211_X1 U20168 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17121), .B(n17106), .ZN(n17107) );
  NAND4_X1 U20169 ( .A1(n17110), .A2(n17109), .A3(n17108), .A4(n17107), .ZN(
        P3_U2802) );
  INV_X1 U20170 ( .A(n17225), .ZN(n17111) );
  OAI21_X1 U20171 ( .B1(n17112), .B2(n17111), .A(n18644), .ZN(n17113) );
  OAI21_X1 U20172 ( .B1(n17115), .B2(n17114), .A(n17113), .ZN(n17246) );
  OR2_X1 U20173 ( .A1(n17246), .A2(n18732), .ZN(n17125) );
  INV_X1 U20174 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19640) );
  OAI22_X1 U20175 ( .A1(n19075), .A2(n19640), .B1(n18706), .B2(n10302), .ZN(
        n17118) );
  AND2_X1 U20176 ( .A1(n17116), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17117) );
  NOR2_X1 U20177 ( .A1(n17118), .A2(n17117), .ZN(n17124) );
  OAI21_X1 U20178 ( .B1(n18555), .B2(n17241), .A(n17240), .ZN(n17119) );
  NAND2_X1 U20179 ( .A1(n17120), .A2(n17119), .ZN(n17123) );
  NAND2_X1 U20180 ( .A1(n17121), .A2(n21668), .ZN(n17122) );
  NAND4_X1 U20181 ( .A1(n17125), .A2(n17124), .A3(n17123), .A4(n17122), .ZN(
        P3_U2803) );
  AOI22_X1 U20182 ( .A1(n18698), .A2(n18664), .B1(n18985), .B2(n18812), .ZN(
        n17161) );
  INV_X1 U20183 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17135) );
  INV_X1 U20184 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U20185 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17150), .ZN(
        n17662) );
  AOI21_X1 U20186 ( .B1(n17673), .B2(n17662), .A(n17623), .ZN(n17664) );
  NOR2_X1 U20187 ( .A1(n19136), .A2(n17126), .ZN(n18752) );
  AND2_X1 U20188 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18752), .ZN(
        n18738) );
  AND2_X1 U20189 ( .A1(n17626), .A2(n18738), .ZN(n17152) );
  NAND2_X1 U20190 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17152), .ZN(
        n17136) );
  NOR2_X1 U20191 ( .A1(n17673), .A2(n17136), .ZN(n18683) );
  AOI211_X1 U20192 ( .C1(n17136), .C2(n17673), .A(n18817), .B(n18683), .ZN(
        n17128) );
  INV_X1 U20193 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19606) );
  NOR2_X1 U20194 ( .A1(n19075), .A2(n19606), .ZN(n17127) );
  AOI211_X1 U20195 ( .C1(n17664), .C2(n18813), .A(n17128), .B(n17127), .ZN(
        n17134) );
  INV_X1 U20196 ( .A(n17129), .ZN(n18990) );
  OR2_X1 U20197 ( .A1(n18990), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18998) );
  OAI21_X1 U20198 ( .B1(n17135), .B2(n17129), .A(n18998), .ZN(n17132) );
  OR2_X1 U20199 ( .A1(n17130), .A2(n18644), .ZN(n18667) );
  INV_X1 U20200 ( .A(n18667), .ZN(n17154) );
  NAND2_X1 U20201 ( .A1(n17154), .A2(n19010), .ZN(n17139) );
  NAND2_X1 U20202 ( .A1(n18988), .A2(n18644), .ZN(n18687) );
  OAI22_X1 U20203 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17139), .B1(
        n18990), .B2(n18687), .ZN(n17131) );
  XOR2_X1 U20204 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17131), .Z(
        n18980) );
  AOI22_X1 U20205 ( .A1(n18724), .A2(n17132), .B1(n18714), .B2(n18980), .ZN(
        n17133) );
  OAI211_X1 U20206 ( .C1(n17161), .C2(n17135), .A(n17134), .B(n17133), .ZN(
        P3_U2819) );
  INV_X1 U20207 ( .A(n17136), .ZN(n17138) );
  INV_X1 U20208 ( .A(n18817), .ZN(n17147) );
  AOI21_X1 U20209 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17147), .A(
        n17152), .ZN(n17137) );
  OAI21_X1 U20210 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17150), .A(
        n17662), .ZN(n17674) );
  OAI22_X1 U20211 ( .A1(n17138), .A2(n17137), .B1(n18803), .B2(n17674), .ZN(
        n17146) );
  OAI21_X1 U20212 ( .B1(n19010), .B2(n18687), .A(n17139), .ZN(n17140) );
  XNOR2_X1 U20213 ( .A(n17144), .B(n17140), .ZN(n19002) );
  INV_X1 U20214 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19604) );
  NOR2_X1 U20215 ( .A1(n19075), .A2(n19604), .ZN(n17141) );
  AOI21_X1 U20216 ( .B1(n18714), .B2(n19002), .A(n17141), .ZN(n17143) );
  OAI211_X1 U20217 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n18724), .B(n18990), .ZN(
        n17142) );
  OAI211_X1 U20218 ( .C1(n17161), .C2(n17144), .A(n17143), .B(n17142), .ZN(
        n17145) );
  OR2_X1 U20219 ( .A1(n17146), .A2(n17145), .ZN(P3_U2820) );
  INV_X1 U20220 ( .A(n17163), .ZN(n17148) );
  AOI22_X1 U20221 ( .A1(n17148), .A2(n18738), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17147), .ZN(n17151) );
  NAND2_X1 U20222 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17149), .ZN(
        n17725) );
  OR2_X1 U20223 ( .A1(n17163), .A2(n17725), .ZN(n17162) );
  AOI21_X1 U20224 ( .B1(n17687), .B2(n17162), .A(n17150), .ZN(n17689) );
  INV_X1 U20225 ( .A(n17689), .ZN(n17686) );
  OAI22_X1 U20226 ( .A1(n17152), .A2(n17151), .B1(n18803), .B2(n17686), .ZN(
        n17153) );
  INV_X1 U20227 ( .A(n17153), .ZN(n17160) );
  INV_X1 U20228 ( .A(n18687), .ZN(n18719) );
  NOR2_X1 U20229 ( .A1(n17154), .A2(n18719), .ZN(n17155) );
  XOR2_X1 U20230 ( .A(n17155), .B(n19010), .Z(n19006) );
  INV_X1 U20231 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19602) );
  NOR2_X1 U20232 ( .A1(n19075), .A2(n19602), .ZN(n17158) );
  INV_X1 U20233 ( .A(n18724), .ZN(n17156) );
  NOR2_X1 U20234 ( .A1(n17156), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17157) );
  AOI211_X1 U20235 ( .C1(n18714), .C2(n19006), .A(n17158), .B(n17157), .ZN(
        n17159) );
  OAI211_X1 U20236 ( .C1(n17161), .C2(n19010), .A(n17160), .B(n17159), .ZN(
        P3_U2821) );
  OAI21_X1 U20237 ( .B1(n17149), .B2(n9899), .A(n18807), .ZN(n18736) );
  NOR2_X1 U20238 ( .A1(n19075), .A2(n19601), .ZN(n17166) );
  INV_X1 U20239 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18737) );
  NOR2_X1 U20240 ( .A1(n18737), .A2(n17725), .ZN(n17710) );
  OAI21_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17710), .A(
        n17162), .ZN(n17701) );
  OAI211_X1 U20242 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17149), .B(n17163), .ZN(n17164)
         );
  OAI22_X1 U20243 ( .A1(n18803), .A2(n17701), .B1(n19136), .B2(n17164), .ZN(
        n17165) );
  AOI211_X1 U20244 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18736), .A(
        n17166), .B(n17165), .ZN(n17171) );
  INV_X1 U20245 ( .A(n17167), .ZN(n17169) );
  AOI22_X1 U20246 ( .A1(n18698), .A2(n17169), .B1(n18812), .B2(n17168), .ZN(
        n17170) );
  OAI211_X1 U20247 ( .C1(n17172), .C2(n18732), .A(n17171), .B(n17170), .ZN(
        P3_U2822) );
  INV_X1 U20248 ( .A(n17173), .ZN(n17175) );
  NAND2_X1 U20249 ( .A1(n17175), .A2(n17174), .ZN(n19078) );
  NAND2_X1 U20250 ( .A1(n18812), .A2(n19078), .ZN(n17178) );
  NAND3_X1 U20251 ( .A1(n19559), .A2(n19570), .A3(n18807), .ZN(n17176) );
  AOI22_X1 U20252 ( .A1(n13950), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17176), .ZN(n17177) );
  OAI211_X1 U20253 ( .C1(n19078), .C2(n18801), .A(n17178), .B(n17177), .ZN(
        P3_U2830) );
  NAND2_X1 U20254 ( .A1(n17179), .A2(n19007), .ZN(n17193) );
  NAND3_X1 U20255 ( .A1(n17180), .A2(n19074), .A3(n18394), .ZN(n17181) );
  OAI21_X1 U20256 ( .B1(n17182), .B2(n19021), .A(n17181), .ZN(n17200) );
  OAI21_X1 U20257 ( .B1(n17200), .B2(n17183), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17192) );
  AOI21_X1 U20258 ( .B1(n17237), .B2(n18961), .A(n17184), .ZN(n17187) );
  NAND2_X1 U20259 ( .A1(n19070), .A2(n17185), .ZN(n17186) );
  OAI22_X1 U20260 ( .A1(n17213), .A2(n19021), .B1(n17187), .B2(n17186), .ZN(
        n17196) );
  NAND3_X1 U20261 ( .A1(n17196), .A2(n17189), .A3(n17188), .ZN(n17190) );
  NAND4_X1 U20262 ( .A1(n17193), .A2(n17192), .A3(n17191), .A4(n17190), .ZN(
        P3_U2832) );
  INV_X1 U20263 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17195) );
  AOI21_X1 U20264 ( .B1(n17196), .B2(n17195), .A(n17194), .ZN(n17202) );
  NAND2_X1 U20265 ( .A1(n18943), .A2(n19061), .ZN(n18999) );
  INV_X1 U20266 ( .A(n18999), .ZN(n18992) );
  OAI21_X1 U20267 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18992), .A(
        n17197), .ZN(n17219) );
  AOI21_X1 U20268 ( .B1(n17219), .B2(n19070), .A(n19042), .ZN(n17198) );
  OAI21_X1 U20269 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n19035), .A(
        n17198), .ZN(n17199) );
  OAI21_X1 U20270 ( .B1(n17200), .B2(n17199), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17201) );
  OAI211_X1 U20271 ( .C1(n17203), .C2(n18956), .A(n17202), .B(n17201), .ZN(
        P3_U2833) );
  INV_X1 U20272 ( .A(n17214), .ZN(n17212) );
  OR2_X1 U20273 ( .A1(n18985), .A2(n10205), .ZN(n17205) );
  NAND2_X1 U20274 ( .A1(n18988), .A2(n18961), .ZN(n17204) );
  NAND2_X1 U20275 ( .A1(n17205), .A2(n17204), .ZN(n17250) );
  INV_X1 U20276 ( .A(n17206), .ZN(n17207) );
  OAI21_X1 U20277 ( .B1(n17208), .B2(n19052), .A(n17207), .ZN(n18826) );
  AOI21_X1 U20278 ( .B1(n17250), .B2(n17209), .A(n18826), .ZN(n18870) );
  NOR2_X1 U20279 ( .A1(n18870), .A2(n19080), .ZN(n18879) );
  NAND2_X1 U20280 ( .A1(n18879), .A2(n18828), .ZN(n18850) );
  INV_X1 U20281 ( .A(n18850), .ZN(n17210) );
  AOI22_X1 U20282 ( .A1(n17212), .A2(n19074), .B1(n17211), .B2(n17210), .ZN(
        n17230) );
  INV_X1 U20283 ( .A(n17213), .ZN(n17222) );
  NAND4_X1 U20284 ( .A1(n17217), .A2(n17216), .A3(n17215), .A4(n17214), .ZN(
        n17221) );
  AOI21_X1 U20285 ( .B1(n17237), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18987), .ZN(n17218) );
  NOR3_X1 U20286 ( .A1(n17219), .A2(n19042), .A3(n17218), .ZN(n17220) );
  OAI211_X1 U20287 ( .C1(n17222), .C2(n10205), .A(n17221), .B(n17220), .ZN(
        n17223) );
  NAND3_X1 U20288 ( .A1(n17223), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n19075), .ZN(n17229) );
  NOR3_X1 U20289 ( .A1(n17225), .A2(n17224), .A3(n18956), .ZN(n17227) );
  NOR2_X1 U20290 ( .A1(n17227), .A2(n17226), .ZN(n17228) );
  OAI211_X1 U20291 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n17230), .A(
        n17229), .B(n17228), .ZN(P3_U2834) );
  AOI21_X1 U20292 ( .B1(n18971), .B2(n18857), .A(n18872), .ZN(n17231) );
  AOI21_X1 U20293 ( .B1(n17232), .B2(n17231), .A(n19062), .ZN(n18840) );
  OAI22_X1 U20294 ( .A1(n18943), .A2(n18827), .B1(n18994), .B2(n17233), .ZN(
        n17234) );
  AOI211_X1 U20295 ( .C1(n19081), .C2(n14436), .A(n17235), .B(n17234), .ZN(
        n17236) );
  OAI211_X1 U20296 ( .C1(n17237), .C2(n18987), .A(n19070), .B(n17236), .ZN(
        n17238) );
  AOI211_X1 U20297 ( .C1(n19519), .C2(n17239), .A(n18840), .B(n17238), .ZN(
        n18819) );
  AOI221_X1 U20298 ( .B1(n18943), .B2(n18819), .C1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n18819), .A(n17240), .ZN(
        n17243) );
  NOR3_X1 U20299 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17241), .A3(
        n18850), .ZN(n17242) );
  AOI21_X1 U20300 ( .B1(n19075), .B2(n17243), .A(n17242), .ZN(n17245) );
  NAND2_X1 U20301 ( .A1(n13950), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17244) );
  OAI211_X1 U20302 ( .C1(n17246), .C2(n18956), .A(n17245), .B(n17244), .ZN(
        P3_U2835) );
  XNOR2_X1 U20303 ( .A(n17247), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18633) );
  NOR3_X1 U20304 ( .A1(n19064), .A2(n18883), .A3(n14427), .ZN(n17248) );
  NOR2_X1 U20305 ( .A1(n19519), .A2(n18961), .ZN(n18896) );
  INV_X1 U20306 ( .A(n18896), .ZN(n18989) );
  AOI22_X1 U20307 ( .A1(n19519), .A2(n18927), .B1(n18961), .B2(n18645), .ZN(
        n18873) );
  NAND3_X1 U20308 ( .A1(n18910), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n19075), .ZN(n17253) );
  NAND2_X1 U20309 ( .A1(n19070), .A2(n18973), .ZN(n19011) );
  NOR2_X1 U20310 ( .A1(n17251), .A2(n19011), .ZN(n18922) );
  NOR2_X1 U20311 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n14427), .ZN(
        n18636) );
  AOI22_X1 U20312 ( .A1(n18922), .A2(n18636), .B1(n13950), .B2(
        P3_REIP_REG_17__SCAN_IN), .ZN(n17252) );
  OAI211_X1 U20313 ( .C1(n18633), .C2(n18956), .A(n17253), .B(n17252), .ZN(
        P3_U2845) );
  MUX2_X1 U20314 ( .A(n17254), .B(n18943), .S(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n19530) );
  AOI22_X1 U20315 ( .A1(n19553), .A2(n9882), .B1(n18884), .B2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20316 ( .B1(n19530), .B2(n17256), .A(n17255), .ZN(n17257) );
  MUX2_X1 U20317 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17257), .S(
        n17280), .Z(P3_U3290) );
  INV_X1 U20318 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17525) );
  NAND2_X1 U20319 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n17258) );
  NAND2_X1 U20320 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17937) );
  NOR4_X1 U20321 ( .A1(n17525), .A2(n17936), .A3(n17258), .A4(n17937), .ZN(
        n17941) );
  INV_X1 U20322 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17610) );
  INV_X1 U20323 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18135) );
  INV_X1 U20324 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n18112) );
  INV_X1 U20325 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18200) );
  NAND2_X1 U20326 ( .A1(n19102), .A2(n19675), .ZN(n17261) );
  INV_X1 U20327 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18253) );
  NAND3_X1 U20328 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18252) );
  NOR4_X1 U20329 ( .A1(n17744), .A2(n18253), .A3(n18257), .A4(n18252), .ZN(
        n18244) );
  NAND2_X1 U20330 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n9686), .ZN(n18110) );
  AND3_X1 U20331 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n18073), .ZN(n18037) );
  NAND3_X1 U20332 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n18037), .ZN(n17987) );
  NOR2_X1 U20333 ( .A1(n17943), .A2(n17987), .ZN(n17262) );
  NAND4_X1 U20334 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17941), .A4(n17262), .ZN(n17813) );
  NOR2_X1 U20335 ( .A1(n17814), .A2(n17813), .ZN(n17934) );
  NAND2_X1 U20336 ( .A1(n18266), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17264) );
  NAND2_X1 U20337 ( .A1(n17934), .A2(n17935), .ZN(n17263) );
  OAI22_X1 U20338 ( .A1(n17934), .A2(n17264), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17263), .ZN(P3_U2672) );
  NAND2_X1 U20339 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19528), .ZN(n19270) );
  NOR2_X1 U20340 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17265), .ZN(
        n17277) );
  NAND2_X1 U20341 ( .A1(n17277), .A2(n17266), .ZN(n19085) );
  INV_X1 U20342 ( .A(n19659), .ZN(n17269) );
  INV_X1 U20343 ( .A(n17267), .ZN(n17268) );
  AOI21_X1 U20344 ( .B1(n19085), .B2(n17269), .A(n17268), .ZN(n17270) );
  AND2_X1 U20345 ( .A1(n19184), .A2(n17270), .ZN(n19092) );
  INV_X1 U20346 ( .A(n19092), .ZN(n17275) );
  NAND2_X1 U20347 ( .A1(n19270), .A2(n17275), .ZN(n17273) );
  INV_X1 U20348 ( .A(n17273), .ZN(n17272) );
  INV_X1 U20349 ( .A(n19087), .ZN(n19674) );
  OAI22_X1 U20350 ( .A1(n19674), .A2(n18790), .B1(n19528), .B2(n19660), .ZN(
        n17276) );
  NAND3_X1 U20351 ( .A1(n10732), .A2(n17275), .A3(n17276), .ZN(n17271) );
  OAI221_X1 U20352 ( .B1(n10732), .B2(n17272), .C1(n10732), .C2(n19205), .A(
        n17271), .ZN(P3_U2864) );
  NAND2_X1 U20353 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19273) );
  NOR2_X1 U20354 ( .A1(n19674), .A2(n18790), .ZN(n17274) );
  AOI221_X1 U20355 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19273), .C1(n17274), 
        .C2(n19273), .A(n17273), .ZN(n19091) );
  INV_X1 U20356 ( .A(n19205), .ZN(n19435) );
  OAI221_X1 U20357 ( .B1(n19435), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19435), .C2(n17276), .A(n17275), .ZN(n19089) );
  AOI22_X1 U20358 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19091), .B1(
        n19089), .B2(n19095), .ZN(P3_U2865) );
  NOR2_X1 U20359 ( .A1(n17278), .A2(n17277), .ZN(n19521) );
  NAND3_X1 U20360 ( .A1(n17280), .A2(n19693), .A3(n19521), .ZN(n17279) );
  OAI21_X1 U20361 ( .B1(n17280), .B2(n17752), .A(n17279), .ZN(P3_U3284) );
  NOR3_X1 U20362 ( .A1(n17282), .A2(n17281), .A3(n21327), .ZN(n17287) );
  AOI211_X1 U20363 ( .C1(n17287), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17284), .B(n17283), .ZN(n17285) );
  INV_X1 U20364 ( .A(n17285), .ZN(n17286) );
  OAI21_X1 U20365 ( .B1(n17287), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17286), .ZN(n17288) );
  AOI222_X1 U20366 ( .A1(n17289), .A2(n21276), .B1(n17289), .B2(n17288), .C1(
        n21276), .C2(n17288), .ZN(n17290) );
  AOI222_X1 U20367 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17291), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17290), .C1(n17291), 
        .C2(n17290), .ZN(n17299) );
  OAI21_X1 U20368 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17292), .ZN(n17293) );
  NAND4_X1 U20369 ( .A1(n17296), .A2(n17295), .A3(n17294), .A4(n17293), .ZN(
        n17297) );
  AOI211_X1 U20370 ( .C1(n17299), .C2(n21623), .A(n17298), .B(n17297), .ZN(
        n17314) );
  NAND3_X1 U20371 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n17309), .A3(n21501), 
        .ZN(n17300) );
  AOI22_X1 U20372 ( .A1(n17303), .A2(n17302), .B1(n17301), .B2(n17300), .ZN(
        n17320) );
  OAI221_X1 U20373 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n17314), 
        .A(n17320), .ZN(n17326) );
  NOR2_X1 U20374 ( .A1(n17305), .A2(n17304), .ZN(n17306) );
  NOR2_X1 U20375 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17306), .ZN(n17312) );
  AOI211_X1 U20376 ( .C1(n17309), .C2(n21503), .A(n17308), .B(n17307), .ZN(
        n17310) );
  NAND2_X1 U20377 ( .A1(n17326), .A2(n17310), .ZN(n17311) );
  AOI22_X1 U20378 ( .A1(n17326), .A2(n17312), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n17311), .ZN(n17313) );
  OAI21_X1 U20379 ( .B1(n17314), .B2(n20568), .A(n17313), .ZN(P1_U3161) );
  INV_X1 U20380 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17438) );
  NOR2_X1 U20381 ( .A1(n20667), .A2(n17438), .ZN(P1_U2905) );
  INV_X1 U20382 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19709) );
  INV_X1 U20383 ( .A(n20538), .ZN(n17315) );
  OAI221_X1 U20384 ( .B1(n19709), .B2(n17316), .C1(n17315), .C2(n17316), .A(
        n20265), .ZN(n20530) );
  NOR2_X1 U20385 ( .A1(n17317), .A2(n20530), .ZN(P2_U3047) );
  NAND2_X1 U20386 ( .A1(n21282), .A2(n21590), .ZN(n17324) );
  AOI21_X1 U20387 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n17326), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17323) );
  NAND4_X1 U20388 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21503), .A4(n21590), .ZN(n17318) );
  AND2_X1 U20389 ( .A1(n17319), .A2(n17318), .ZN(n21502) );
  AOI21_X1 U20390 ( .B1(n21502), .B2(n17321), .A(n17320), .ZN(n17322) );
  AOI211_X1 U20391 ( .C1(n21587), .C2(n17324), .A(n17323), .B(n17322), .ZN(
        P1_U3162) );
  OAI221_X1 U20392 ( .B1(n21282), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n21282), 
        .C2(n17326), .A(n17325), .ZN(P1_U3466) );
  AOI22_X1 U20393 ( .A1(n17328), .A2(n17327), .B1(n19745), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n17329) );
  OAI21_X1 U20394 ( .B1(n17331), .B2(n17330), .A(n17329), .ZN(n17334) );
  NOR2_X1 U20395 ( .A1(n17332), .A2(n17348), .ZN(n17333) );
  AOI211_X1 U20396 ( .C1(n17351), .C2(n17335), .A(n17334), .B(n17333), .ZN(
        n17336) );
  OAI221_X1 U20397 ( .B1(n16967), .B2(n17338), .C1(n16967), .C2(n17337), .A(
        n17336), .ZN(P2_U3041) );
  OAI22_X1 U20398 ( .A1(n17340), .A2(n20502), .B1(n10136), .B2(n17339), .ZN(
        n17344) );
  NOR2_X1 U20399 ( .A1(n17342), .A2(n17341), .ZN(n17343) );
  AOI211_X1 U20400 ( .C1(n17346), .C2(n17345), .A(n17344), .B(n17343), .ZN(
        n17347) );
  OAI21_X1 U20401 ( .B1(n17349), .B2(n17348), .A(n17347), .ZN(n17350) );
  AOI21_X1 U20402 ( .B1(n17352), .B2(n17351), .A(n17350), .ZN(n17353) );
  OAI21_X1 U20403 ( .B1(n17355), .B2(n17354), .A(n17353), .ZN(P2_U3043) );
  AOI21_X1 U20404 ( .B1(n17357), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17356), 
        .ZN(n17358) );
  INV_X1 U20405 ( .A(n17358), .ZN(P2_U3593) );
  NOR3_X1 U20406 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n17360) );
  NOR4_X1 U20407 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17359) );
  INV_X2 U20408 ( .A(n17425), .ZN(U215) );
  NAND4_X1 U20409 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17360), .A3(n17359), .A4(
        U215), .ZN(U213) );
  INV_X1 U20410 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17362) );
  INV_X1 U20411 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21684) );
  OAI222_X1 U20412 ( .A1(U214), .A2(n17438), .B1(n17406), .B2(n17362), .C1(
        U212), .C2(n21684), .ZN(U216) );
  AOI222_X1 U20413 ( .A1(n17403), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17401), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17404), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17363) );
  INV_X1 U20414 ( .A(n17363), .ZN(U217) );
  AOI22_X1 U20415 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17403), .ZN(n17364) );
  OAI21_X1 U20416 ( .B1(n14942), .B2(n17406), .A(n17364), .ZN(U218) );
  AOI22_X1 U20417 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17403), .ZN(n17365) );
  OAI21_X1 U20418 ( .B1(n16334), .B2(n17406), .A(n17365), .ZN(U219) );
  AOI22_X1 U20419 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17403), .ZN(n17366) );
  OAI21_X1 U20420 ( .B1(n14955), .B2(n17406), .A(n17366), .ZN(U220) );
  AOI22_X1 U20421 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17403), .ZN(n17367) );
  OAI21_X1 U20422 ( .B1(n16350), .B2(n17406), .A(n17367), .ZN(U221) );
  AOI222_X1 U20423 ( .A1(n17403), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n17401), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n17404), .C2(P1_DATAO_REG_25__SCAN_IN), 
        .ZN(n17368) );
  INV_X1 U20424 ( .A(n17368), .ZN(U222) );
  AOI222_X1 U20425 ( .A1(n17403), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n17401), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n17404), .C2(P1_DATAO_REG_24__SCAN_IN), 
        .ZN(n17369) );
  INV_X1 U20426 ( .A(n17369), .ZN(U223) );
  AOI22_X1 U20427 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17403), .ZN(n17370) );
  OAI21_X1 U20428 ( .B1(n16372), .B2(n17406), .A(n17370), .ZN(U224) );
  AOI22_X1 U20429 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17403), .ZN(n17371) );
  OAI21_X1 U20430 ( .B1(n14983), .B2(n17406), .A(n17371), .ZN(U225) );
  INV_X1 U20431 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U20432 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17403), .ZN(n17372) );
  OAI21_X1 U20433 ( .B1(n17373), .B2(n17406), .A(n17372), .ZN(U226) );
  INV_X1 U20434 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21665) );
  AOI22_X1 U20435 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17403), .ZN(n17374) );
  OAI21_X1 U20436 ( .B1(n21665), .B2(n17406), .A(n17374), .ZN(U227) );
  AOI22_X1 U20437 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n17404), .ZN(n17375) );
  OAI21_X1 U20438 ( .B1(n21728), .B2(U212), .A(n17375), .ZN(U228) );
  AOI22_X1 U20439 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17403), .ZN(n17376) );
  OAI21_X1 U20440 ( .B1(n16412), .B2(n17406), .A(n17376), .ZN(U229) );
  INV_X1 U20441 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U20442 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17403), .ZN(n17377) );
  OAI21_X1 U20443 ( .B1(n19851), .B2(n17406), .A(n17377), .ZN(U230) );
  INV_X1 U20444 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20445 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17403), .ZN(n17378) );
  OAI21_X1 U20446 ( .B1(n17379), .B2(n17406), .A(n17378), .ZN(U231) );
  INV_X1 U20447 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20448 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17404), .ZN(n17380) );
  OAI21_X1 U20449 ( .B1(n17381), .B2(U212), .A(n17380), .ZN(U232) );
  INV_X1 U20450 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20451 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17404), .ZN(n17382) );
  OAI21_X1 U20452 ( .B1(n17383), .B2(U212), .A(n17382), .ZN(U233) );
  INV_X1 U20453 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20454 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17404), .ZN(n17384) );
  OAI21_X1 U20455 ( .B1(n17420), .B2(U212), .A(n17384), .ZN(U234) );
  AOI22_X1 U20456 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17403), .ZN(n17385) );
  OAI21_X1 U20457 ( .B1(n21639), .B2(n17406), .A(n17385), .ZN(U235) );
  INV_X1 U20458 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20459 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17404), .ZN(n17386) );
  OAI21_X1 U20460 ( .B1(n17387), .B2(U212), .A(n17386), .ZN(U236) );
  AOI22_X1 U20461 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17403), .ZN(n17388) );
  OAI21_X1 U20462 ( .B1(n17389), .B2(n17406), .A(n17388), .ZN(U237) );
  AOI22_X1 U20463 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17403), .ZN(n17390) );
  OAI21_X1 U20464 ( .B1(n17391), .B2(n17406), .A(n17390), .ZN(U238) );
  AOI22_X1 U20465 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17403), .ZN(n17392) );
  OAI21_X1 U20466 ( .B1(n17393), .B2(n17406), .A(n17392), .ZN(U239) );
  INV_X1 U20467 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20468 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17404), .ZN(n17394) );
  OAI21_X1 U20469 ( .B1(n17414), .B2(U212), .A(n17394), .ZN(U240) );
  INV_X1 U20470 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20471 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17404), .ZN(n17395) );
  OAI21_X1 U20472 ( .B1(n17413), .B2(U212), .A(n17395), .ZN(U241) );
  INV_X1 U20473 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20474 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17404), .ZN(n17396) );
  OAI21_X1 U20475 ( .B1(n17412), .B2(U212), .A(n17396), .ZN(U242) );
  AOI22_X1 U20476 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17403), .ZN(n17397) );
  OAI21_X1 U20477 ( .B1(n13774), .B2(n17406), .A(n17397), .ZN(U243) );
  AOI22_X1 U20478 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17403), .ZN(n17398) );
  OAI21_X1 U20479 ( .B1(n17399), .B2(n17406), .A(n17398), .ZN(U244) );
  AOI22_X1 U20480 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17403), .ZN(n17400) );
  OAI21_X1 U20481 ( .B1(n13779), .B2(n17406), .A(n17400), .ZN(U245) );
  INV_X1 U20482 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20483 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17401), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17404), .ZN(n17402) );
  OAI21_X1 U20484 ( .B1(n17408), .B2(U212), .A(n17402), .ZN(U246) );
  AOI22_X1 U20485 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17404), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17403), .ZN(n17405) );
  OAI21_X1 U20486 ( .B1(n13706), .B2(n17406), .A(n17405), .ZN(U247) );
  OAI22_X1 U20487 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17425), .ZN(n17407) );
  INV_X1 U20488 ( .A(n17407), .ZN(U251) );
  INV_X1 U20489 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19103) );
  AOI22_X1 U20490 ( .A1(n17425), .A2(n17408), .B1(n19103), .B2(U215), .ZN(U252) );
  OAI22_X1 U20491 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17425), .ZN(n17409) );
  INV_X1 U20492 ( .A(n17409), .ZN(U253) );
  OAI22_X1 U20493 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17425), .ZN(n17410) );
  INV_X1 U20494 ( .A(n17410), .ZN(U254) );
  OAI22_X1 U20495 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17425), .ZN(n17411) );
  INV_X1 U20496 ( .A(n17411), .ZN(U255) );
  AOI22_X1 U20497 ( .A1(n17425), .A2(n17412), .B1(n19124), .B2(U215), .ZN(U256) );
  INV_X1 U20498 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19128) );
  AOI22_X1 U20499 ( .A1(n17425), .A2(n17413), .B1(n19128), .B2(U215), .ZN(U257) );
  AOI22_X1 U20500 ( .A1(n17425), .A2(n17414), .B1(n19133), .B2(U215), .ZN(U258) );
  OAI22_X1 U20501 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17425), .ZN(n17415) );
  INV_X1 U20502 ( .A(n17415), .ZN(U259) );
  OAI22_X1 U20503 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17425), .ZN(n17416) );
  INV_X1 U20504 ( .A(n17416), .ZN(U260) );
  OAI22_X1 U20505 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17425), .ZN(n17417) );
  INV_X1 U20506 ( .A(n17417), .ZN(U261) );
  OAI22_X1 U20507 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17425), .ZN(n17418) );
  INV_X1 U20508 ( .A(n17418), .ZN(U262) );
  OAI22_X1 U20509 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17425), .ZN(n17419) );
  INV_X1 U20510 ( .A(n17419), .ZN(U263) );
  INV_X1 U20511 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18516) );
  AOI22_X1 U20512 ( .A1(n17425), .A2(n17420), .B1(n18516), .B2(U215), .ZN(U264) );
  OAI22_X1 U20513 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17425), .ZN(n17421) );
  INV_X1 U20514 ( .A(n17421), .ZN(U265) );
  OAI22_X1 U20515 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17425), .ZN(n17422) );
  INV_X1 U20516 ( .A(n17422), .ZN(U266) );
  OAI22_X1 U20517 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17425), .ZN(n17423) );
  INV_X1 U20518 ( .A(n17423), .ZN(U267) );
  OAI22_X1 U20519 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17425), .ZN(n17424) );
  INV_X1 U20520 ( .A(n17424), .ZN(U268) );
  OAI22_X1 U20521 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17425), .ZN(n17426) );
  INV_X1 U20522 ( .A(n17426), .ZN(U269) );
  INV_X1 U20523 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19114) );
  AOI22_X1 U20524 ( .A1(n17425), .A2(n21728), .B1(n19114), .B2(U215), .ZN(U270) );
  OAI22_X1 U20525 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17425), .ZN(n17428) );
  INV_X1 U20526 ( .A(n17428), .ZN(U271) );
  OAI22_X1 U20527 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17425), .ZN(n17429) );
  INV_X1 U20528 ( .A(n17429), .ZN(U272) );
  OAI22_X1 U20529 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17425), .ZN(n17430) );
  INV_X1 U20530 ( .A(n17430), .ZN(U273) );
  OAI22_X1 U20531 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17425), .ZN(n17431) );
  INV_X1 U20532 ( .A(n17431), .ZN(U274) );
  OAI22_X1 U20533 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17425), .ZN(n17432) );
  INV_X1 U20534 ( .A(n17432), .ZN(U275) );
  OAI22_X1 U20535 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17425), .ZN(n17433) );
  INV_X1 U20536 ( .A(n17433), .ZN(U276) );
  OAI22_X1 U20537 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17425), .ZN(n17434) );
  INV_X1 U20538 ( .A(n17434), .ZN(U277) );
  OAI22_X1 U20539 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17425), .ZN(n17435) );
  INV_X1 U20540 ( .A(n17435), .ZN(U278) );
  OAI22_X1 U20541 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17425), .ZN(n17436) );
  INV_X1 U20542 ( .A(n17436), .ZN(U279) );
  OAI22_X1 U20543 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17425), .ZN(n17437) );
  INV_X1 U20544 ( .A(n17437), .ZN(U280) );
  INV_X1 U20545 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19797) );
  AOI22_X1 U20546 ( .A1(n17425), .A2(n19797), .B1(n16319), .B2(U215), .ZN(U281) );
  INV_X1 U20547 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19135) );
  AOI22_X1 U20548 ( .A1(n17425), .A2(n21684), .B1(n19135), .B2(U215), .ZN(U282) );
  INV_X1 U20549 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17439) );
  AOI222_X1 U20550 ( .A1(n17439), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n17438), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n21684), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n17440) );
  INV_X2 U20551 ( .A(n17442), .ZN(n17441) );
  INV_X1 U20552 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19605) );
  AOI22_X1 U20553 ( .A1(n17441), .A2(n19605), .B1(n21626), .B2(n17442), .ZN(
        U347) );
  INV_X1 U20554 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19603) );
  INV_X1 U20555 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20445) );
  AOI22_X1 U20556 ( .A1(n17441), .A2(n19603), .B1(n20445), .B2(n17442), .ZN(
        U348) );
  INV_X1 U20557 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19600) );
  INV_X1 U20558 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20443) );
  AOI22_X1 U20559 ( .A1(n17441), .A2(n19600), .B1(n20443), .B2(n17442), .ZN(
        U349) );
  INV_X1 U20560 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19599) );
  INV_X1 U20561 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20441) );
  AOI22_X1 U20562 ( .A1(n17441), .A2(n19599), .B1(n20441), .B2(n17442), .ZN(
        U350) );
  INV_X1 U20563 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19598) );
  INV_X1 U20564 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U20565 ( .A1(n17441), .A2(n19598), .B1(n20439), .B2(n17442), .ZN(
        U351) );
  INV_X1 U20566 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19596) );
  INV_X1 U20567 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20437) );
  AOI22_X1 U20568 ( .A1(n17441), .A2(n19596), .B1(n20437), .B2(n17442), .ZN(
        U352) );
  INV_X1 U20569 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19595) );
  INV_X1 U20570 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20435) );
  AOI22_X1 U20571 ( .A1(n17441), .A2(n19595), .B1(n20435), .B2(n17442), .ZN(
        U353) );
  INV_X1 U20572 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19592) );
  INV_X1 U20573 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20433) );
  AOI22_X1 U20574 ( .A1(n17441), .A2(n19592), .B1(n20433), .B2(n17442), .ZN(
        U354) );
  INV_X1 U20575 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19648) );
  INV_X1 U20576 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20482) );
  AOI22_X1 U20577 ( .A1(n17441), .A2(n19648), .B1(n20482), .B2(n17442), .ZN(
        U355) );
  INV_X1 U20578 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19645) );
  INV_X1 U20579 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20480) );
  AOI22_X1 U20580 ( .A1(n17441), .A2(n19645), .B1(n20480), .B2(n17442), .ZN(
        U356) );
  INV_X1 U20581 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19642) );
  INV_X1 U20582 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20478) );
  AOI22_X1 U20583 ( .A1(n17441), .A2(n19642), .B1(n20478), .B2(n17442), .ZN(
        U357) );
  INV_X1 U20584 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19641) );
  INV_X1 U20585 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20475) );
  AOI22_X1 U20586 ( .A1(n17441), .A2(n19641), .B1(n20475), .B2(n17442), .ZN(
        U358) );
  INV_X1 U20587 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19639) );
  INV_X1 U20588 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20474) );
  AOI22_X1 U20589 ( .A1(n17441), .A2(n19639), .B1(n20474), .B2(n17442), .ZN(
        U359) );
  INV_X1 U20590 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19636) );
  INV_X1 U20591 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20472) );
  AOI22_X1 U20592 ( .A1(n17441), .A2(n19636), .B1(n20472), .B2(n17442), .ZN(
        U360) );
  INV_X1 U20593 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19634) );
  INV_X1 U20594 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20470) );
  AOI22_X1 U20595 ( .A1(n17441), .A2(n19634), .B1(n20470), .B2(n17442), .ZN(
        U361) );
  INV_X1 U20596 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19630) );
  INV_X1 U20597 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20469) );
  AOI22_X1 U20598 ( .A1(n17441), .A2(n19630), .B1(n20469), .B2(n17442), .ZN(
        U362) );
  INV_X1 U20599 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19629) );
  INV_X1 U20600 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U20601 ( .A1(n17441), .A2(n19629), .B1(n20467), .B2(n17442), .ZN(
        U363) );
  INV_X1 U20602 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19627) );
  INV_X1 U20603 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20465) );
  AOI22_X1 U20604 ( .A1(n17441), .A2(n19627), .B1(n20465), .B2(n17442), .ZN(
        U364) );
  INV_X1 U20605 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19591) );
  INV_X1 U20606 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U20607 ( .A1(n17441), .A2(n19591), .B1(n20432), .B2(n17442), .ZN(
        U365) );
  INV_X1 U20608 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19624) );
  INV_X1 U20609 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20463) );
  AOI22_X1 U20610 ( .A1(n17441), .A2(n19624), .B1(n20463), .B2(n17442), .ZN(
        U366) );
  INV_X1 U20611 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19623) );
  INV_X1 U20612 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20462) );
  AOI22_X1 U20613 ( .A1(n17441), .A2(n19623), .B1(n20462), .B2(n17442), .ZN(
        U367) );
  INV_X1 U20614 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19621) );
  INV_X1 U20615 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20461) );
  AOI22_X1 U20616 ( .A1(n17441), .A2(n19621), .B1(n20461), .B2(n17442), .ZN(
        U368) );
  INV_X1 U20617 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19618) );
  INV_X1 U20618 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20460) );
  AOI22_X1 U20619 ( .A1(n17441), .A2(n19618), .B1(n20460), .B2(n17442), .ZN(
        U369) );
  INV_X1 U20620 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19617) );
  INV_X1 U20621 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20458) );
  AOI22_X1 U20622 ( .A1(n17441), .A2(n19617), .B1(n20458), .B2(n17442), .ZN(
        U370) );
  INV_X1 U20623 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19615) );
  INV_X1 U20624 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20456) );
  AOI22_X1 U20625 ( .A1(n17440), .A2(n19615), .B1(n20456), .B2(n17442), .ZN(
        U371) );
  INV_X1 U20626 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19612) );
  INV_X1 U20627 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20454) );
  AOI22_X1 U20628 ( .A1(n17441), .A2(n19612), .B1(n20454), .B2(n17442), .ZN(
        U372) );
  INV_X1 U20629 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19611) );
  INV_X1 U20630 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20452) );
  AOI22_X1 U20631 ( .A1(n17440), .A2(n19611), .B1(n20452), .B2(n17442), .ZN(
        U373) );
  INV_X1 U20632 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19609) );
  INV_X1 U20633 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20450) );
  AOI22_X1 U20634 ( .A1(n17440), .A2(n19609), .B1(n20450), .B2(n17442), .ZN(
        U374) );
  INV_X1 U20635 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19607) );
  INV_X1 U20636 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20448) );
  AOI22_X1 U20637 ( .A1(n17440), .A2(n19607), .B1(n20448), .B2(n17442), .ZN(
        U375) );
  INV_X1 U20638 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19588) );
  INV_X1 U20639 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U20640 ( .A1(n17441), .A2(n19588), .B1(n20430), .B2(n17442), .ZN(
        U376) );
  INV_X1 U20641 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19587) );
  NAND2_X1 U20642 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19587), .ZN(n19575) );
  INV_X1 U20643 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19585) );
  AOI22_X1 U20644 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19575), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19585), .ZN(n19656) );
  AOI21_X1 U20645 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19656), .ZN(n17443) );
  INV_X1 U20646 ( .A(n17443), .ZN(P3_U2633) );
  OAI21_X1 U20647 ( .B1(n17450), .B2(n18473), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17444) );
  OAI21_X1 U20648 ( .B1(n17446), .B2(n17445), .A(n17444), .ZN(P3_U2634) );
  AOI21_X1 U20649 ( .B1(n19585), .B2(n19587), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17447) );
  AOI22_X1 U20650 ( .A1(n19647), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17447), 
        .B2(n19690), .ZN(P3_U2635) );
  OAI21_X1 U20651 ( .B1(n19572), .B2(BS16), .A(n19656), .ZN(n19654) );
  OAI21_X1 U20652 ( .B1(n19656), .B2(n19680), .A(n19654), .ZN(P3_U2636) );
  INV_X1 U20653 ( .A(n19516), .ZN(n17449) );
  NOR3_X1 U20654 ( .A1(n17450), .A2(n17449), .A3(n17448), .ZN(n19545) );
  INV_X1 U20655 ( .A(n19675), .ZN(n19549) );
  NOR2_X1 U20656 ( .A1(n19545), .A2(n19549), .ZN(n19670) );
  OAI21_X1 U20657 ( .B1(n19670), .B2(n17452), .A(n17451), .ZN(P3_U2637) );
  NOR4_X1 U20658 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n17456) );
  NOR4_X1 U20659 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n17455) );
  NOR4_X1 U20660 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17454) );
  NOR4_X1 U20661 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17453) );
  NAND4_X1 U20662 ( .A1(n17456), .A2(n17455), .A3(n17454), .A4(n17453), .ZN(
        n17462) );
  NOR4_X1 U20663 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n17460) );
  AOI211_X1 U20664 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_25__SCAN_IN), .B(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17459) );
  NOR4_X1 U20665 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17458) );
  NOR4_X1 U20666 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17457) );
  NAND4_X1 U20667 ( .A1(n17460), .A2(n17459), .A3(n17458), .A4(n17457), .ZN(
        n17461) );
  NOR2_X1 U20668 ( .A1(n17462), .A2(n17461), .ZN(n17466) );
  INV_X1 U20669 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21651) );
  INV_X1 U20670 ( .A(n17466), .ZN(n19667) );
  NOR2_X1 U20671 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(n19667), .ZN(n17464)
         );
  INV_X1 U20672 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19666) );
  INV_X1 U20673 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17463) );
  NAND3_X1 U20674 ( .A1(n17464), .A2(n19666), .A3(n17463), .ZN(n17465) );
  OAI221_X1 U20675 ( .B1(n17466), .B2(n21651), .C1(n19667), .C2(n13988), .A(
        n17465), .ZN(P3_U2638) );
  INV_X1 U20676 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19650) );
  NAND2_X1 U20677 ( .A1(n17464), .A2(n13988), .ZN(n19664) );
  OAI211_X1 U20678 ( .C1(n17466), .C2(n19650), .A(n19664), .B(n17465), .ZN(
        P3_U2639) );
  AOI22_X1 U20679 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17467), .B1(n17800), 
        .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n17477) );
  NOR2_X1 U20680 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17487), .ZN(n17475) );
  INV_X1 U20681 ( .A(n17484), .ZN(n17469) );
  AOI21_X1 U20682 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17469), .A(n17468), .ZN(
        n17474) );
  AOI211_X1 U20683 ( .C1(n17472), .C2(n17471), .A(n17470), .B(n19566), .ZN(
        n17473) );
  AOI211_X1 U20684 ( .C1(n17480), .C2(n17475), .A(n17474), .B(n17473), .ZN(
        n17476) );
  INV_X1 U20685 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17491) );
  NOR2_X1 U20686 ( .A1(n17592), .A2(n17479), .ZN(n17502) );
  AOI22_X1 U20687 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17502), .B1(n17800), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17490) );
  INV_X1 U20688 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19643) );
  INV_X1 U20689 ( .A(n17480), .ZN(n17500) );
  AOI21_X1 U20690 ( .B1(n19643), .B2(n19640), .A(n17500), .ZN(n17488) );
  AOI211_X1 U20691 ( .C1(n17483), .C2(n17481), .A(n17482), .B(n19566), .ZN(
        n17486) );
  AOI211_X1 U20692 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17496), .A(n17484), .B(
        n17805), .ZN(n17485) );
  AOI211_X1 U20693 ( .C1(n17488), .C2(n17487), .A(n17486), .B(n17485), .ZN(
        n17489) );
  OAI211_X1 U20694 ( .C1(n17491), .C2(n17801), .A(n17490), .B(n17489), .ZN(
        P3_U2643) );
  AOI211_X1 U20695 ( .C1(n17493), .C2(n17492), .A(n9644), .B(n19566), .ZN(
        n17495) );
  OAI22_X1 U20696 ( .A1(n21668), .A2(n17801), .B1(n17768), .B2(n17497), .ZN(
        n17494) );
  AOI211_X1 U20697 ( .C1(n17502), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17495), 
        .B(n17494), .ZN(n17499) );
  OAI211_X1 U20698 ( .C1(n17503), .C2(n17497), .A(n17774), .B(n17496), .ZN(
        n17498) );
  OAI211_X1 U20699 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17500), .A(n17499), 
        .B(n17498), .ZN(P3_U2644) );
  INV_X1 U20700 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19633) );
  NOR2_X1 U20701 ( .A1(n19633), .A2(n17501), .ZN(n17516) );
  AOI21_X1 U20702 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n17516), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17511) );
  INV_X1 U20703 ( .A(n17502), .ZN(n17510) );
  AOI22_X1 U20704 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17716), .B1(
        n17800), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17509) );
  AOI211_X1 U20705 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17517), .A(n17503), .B(
        n17805), .ZN(n17507) );
  AOI211_X1 U20706 ( .C1(n18524), .C2(n17504), .A(n17505), .B(n19566), .ZN(
        n17506) );
  NOR2_X1 U20707 ( .A1(n17507), .A2(n17506), .ZN(n17508) );
  OAI211_X1 U20708 ( .C1(n17511), .C2(n17510), .A(n17509), .B(n17508), .ZN(
        P3_U2645) );
  AOI22_X1 U20709 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17716), .B1(
        n17800), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n17523) );
  INV_X1 U20710 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19635) );
  AOI211_X1 U20711 ( .C1(n17514), .C2(n17513), .A(n17512), .B(n19566), .ZN(
        n17515) );
  AOI21_X1 U20712 ( .B1(n17516), .B2(n19635), .A(n17515), .ZN(n17522) );
  OAI211_X1 U20713 ( .C1(n17524), .C2(n17518), .A(n17774), .B(n17517), .ZN(
        n17521) );
  AND2_X1 U20714 ( .A1(n17594), .A2(n17519), .ZN(n17538) );
  NOR2_X1 U20715 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17806), .ZN(n17532) );
  OAI21_X1 U20716 ( .B1(n17538), .B2(n17532), .A(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n17520) );
  NAND4_X1 U20717 ( .A1(n17523), .A2(n17522), .A3(n17521), .A4(n17520), .ZN(
        P3_U2646) );
  AOI211_X1 U20718 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17539), .A(n17524), .B(
        n17805), .ZN(n17527) );
  OAI22_X1 U20719 ( .A1(n18550), .A2(n17801), .B1(n17768), .B2(n17525), .ZN(
        n17526) );
  AOI211_X1 U20720 ( .C1(n17538), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17527), 
        .B(n17526), .ZN(n17534) );
  AOI211_X1 U20721 ( .C1(n18546), .C2(n17529), .A(n17528), .B(n19566), .ZN(
        n17530) );
  AOI21_X1 U20722 ( .B1(n17532), .B2(n17531), .A(n17530), .ZN(n17533) );
  NAND2_X1 U20723 ( .A1(n17534), .A2(n17533), .ZN(P3_U2647) );
  AOI22_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17716), .B1(
        n17800), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n17543) );
  AOI211_X1 U20725 ( .C1(n18560), .C2(n17536), .A(n17535), .B(n19566), .ZN(
        n17537) );
  AOI21_X1 U20726 ( .B1(n17538), .B2(P3_REIP_REG_23__SCAN_IN), .A(n17537), 
        .ZN(n17542) );
  NAND4_X1 U20727 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n17551), .A4(n19631), .ZN(n17541) );
  OAI211_X1 U20728 ( .C1(n17545), .C2(n17936), .A(n17774), .B(n17539), .ZN(
        n17540) );
  NAND4_X1 U20729 ( .A1(n17543), .A2(n17542), .A3(n17541), .A4(n17540), .ZN(
        P3_U2648) );
  AOI211_X1 U20730 ( .C1(n18580), .C2(n9758), .A(n17544), .B(n19566), .ZN(
        n17549) );
  AOI211_X1 U20731 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17556), .A(n17545), .B(
        n17805), .ZN(n17548) );
  AOI22_X1 U20732 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17716), .B1(
        n17800), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n17546) );
  INV_X1 U20733 ( .A(n17546), .ZN(n17547) );
  NOR3_X1 U20734 ( .A1(n17549), .A2(n17548), .A3(n17547), .ZN(n17553) );
  NAND2_X1 U20735 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17550) );
  OAI211_X1 U20736 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17551), .B(n17550), .ZN(n17552) );
  OAI211_X1 U20737 ( .C1(n19628), .C2(n17562), .A(n17553), .B(n17552), .ZN(
        P3_U2649) );
  AOI211_X1 U20738 ( .C1(n18590), .C2(n17555), .A(n17554), .B(n19566), .ZN(
        n17560) );
  OAI211_X1 U20739 ( .C1(n17557), .C2(n18005), .A(n17774), .B(n17556), .ZN(
        n17558) );
  OAI21_X1 U20740 ( .B1(n18005), .B2(n17768), .A(n17558), .ZN(n17559) );
  AOI211_X1 U20741 ( .C1(n17716), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17560), .B(n17559), .ZN(n17561) );
  OAI221_X1 U20742 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17563), .C1(n19626), 
        .C2(n17562), .A(n17561), .ZN(P3_U2650) );
  INV_X1 U20743 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19622) );
  NAND2_X1 U20744 ( .A1(n17594), .A2(n17564), .ZN(n17584) );
  NOR2_X1 U20745 ( .A1(n18816), .A2(n18609), .ZN(n18608) );
  NAND2_X1 U20746 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18608), .ZN(
        n17576) );
  INV_X1 U20747 ( .A(n17576), .ZN(n17565) );
  OAI21_X1 U20748 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17565), .A(
        n18571), .ZN(n18613) );
  OAI21_X1 U20749 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17576), .A(
        n17748), .ZN(n17567) );
  OAI21_X1 U20750 ( .B1(n18613), .B2(n17567), .A(n17781), .ZN(n17566) );
  AOI21_X1 U20751 ( .B1(n18613), .B2(n17567), .A(n17566), .ZN(n17571) );
  OAI211_X1 U20752 ( .C1(n17579), .C2(n18038), .A(n17774), .B(n17568), .ZN(
        n17569) );
  OAI211_X1 U20753 ( .C1(n17768), .C2(n18038), .A(n19075), .B(n17569), .ZN(
        n17570) );
  AOI211_X1 U20754 ( .C1(n17716), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17571), .B(n17570), .ZN(n17575) );
  OAI211_X1 U20755 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17573), .B(n17572), .ZN(n17574) );
  OAI211_X1 U20756 ( .C1(n19622), .C2(n17584), .A(n17575), .B(n17574), .ZN(
        P3_U2652) );
  INV_X1 U20757 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19620) );
  OAI21_X1 U20758 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18608), .A(
        n17576), .ZN(n18619) );
  INV_X1 U20759 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17587) );
  NAND2_X1 U20760 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17603), .ZN(
        n17602) );
  OR2_X1 U20761 ( .A1(n17602), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17586) );
  OAI21_X1 U20762 ( .B1(n17587), .B2(n17586), .A(n17748), .ZN(n17578) );
  OAI21_X1 U20763 ( .B1(n18619), .B2(n17578), .A(n17781), .ZN(n17577) );
  AOI21_X1 U20764 ( .B1(n18619), .B2(n17578), .A(n17577), .ZN(n17582) );
  AOI211_X1 U20765 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17589), .A(n17579), .B(
        n17805), .ZN(n17581) );
  INV_X1 U20766 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18622) );
  OAI22_X1 U20767 ( .A1(n18622), .A2(n17801), .B1(n17768), .B2(n18054), .ZN(
        n17580) );
  NOR4_X1 U20768 ( .A1(n19022), .A2(n17582), .A3(n17581), .A4(n17580), .ZN(
        n17583) );
  OAI221_X1 U20769 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17585), .C1(n19620), 
        .C2(n17584), .A(n17583), .ZN(P3_U2653) );
  NAND2_X1 U20770 ( .A1(n17748), .A2(n17586), .ZN(n17588) );
  AOI21_X1 U20771 ( .B1(n17587), .B2(n17602), .A(n18608), .ZN(n18632) );
  XOR2_X1 U20772 ( .A(n17588), .B(n18632), .Z(n17600) );
  OAI211_X1 U20773 ( .C1(n17601), .C2(n18075), .A(n17774), .B(n17589), .ZN(
        n17590) );
  OAI211_X1 U20774 ( .C1(n17768), .C2(n18075), .A(n19075), .B(n17590), .ZN(
        n17598) );
  NAND2_X1 U20775 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17593) );
  NOR2_X1 U20776 ( .A1(n17593), .A2(n17591), .ZN(n17596) );
  NOR2_X1 U20777 ( .A1(n17592), .A2(n17635), .ZN(n17631) );
  AOI21_X1 U20778 ( .B1(n17594), .B2(n17593), .A(n17631), .ZN(n17606) );
  INV_X1 U20779 ( .A(n17606), .ZN(n17595) );
  MUX2_X1 U20780 ( .A(n17596), .B(n17595), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n17597) );
  AOI211_X1 U20781 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n17716), .A(
        n17598), .B(n17597), .ZN(n17599) );
  OAI21_X1 U20782 ( .B1(n17600), .B2(n19566), .A(n17599), .ZN(P3_U2654) );
  AOI211_X1 U20783 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17617), .A(n17601), .B(
        n17805), .ZN(n17608) );
  AOI21_X1 U20784 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17616), .A(
        P3_REIP_REG_16__SCAN_IN), .ZN(n17605) );
  OAI21_X1 U20785 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17603), .A(
        n17602), .ZN(n18653) );
  XOR2_X1 U20786 ( .A(n17613), .B(n18653), .Z(n17604) );
  OAI22_X1 U20787 ( .A1(n17606), .A2(n17605), .B1(n19566), .B2(n17604), .ZN(
        n17607) );
  AOI211_X1 U20788 ( .C1(n17716), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17608), .B(n17607), .ZN(n17609) );
  OAI211_X1 U20789 ( .C1(n17768), .C2(n17610), .A(n17609), .B(n19075), .ZN(
        P3_U2655) );
  OAI21_X1 U20790 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18647), .A(
        n17611), .ZN(n18658) );
  AOI21_X1 U20791 ( .B1(n17748), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19566), .ZN(n17809) );
  INV_X1 U20792 ( .A(n17809), .ZN(n17639) );
  AOI211_X1 U20793 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17748), .A(
        n18658), .B(n17639), .ZN(n17612) );
  AOI21_X1 U20794 ( .B1(n17716), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17612), .ZN(n17620) );
  NAND3_X1 U20795 ( .A1(n17613), .A2(n17781), .A3(n18658), .ZN(n17614) );
  OAI211_X1 U20796 ( .C1(n17768), .C2(n21713), .A(n19075), .B(n17614), .ZN(
        n17615) );
  AOI221_X1 U20797 ( .B1(n17631), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n17616), 
        .C2(n19614), .A(n17615), .ZN(n17619) );
  OAI211_X1 U20798 ( .C1(n17621), .C2(n21713), .A(n17774), .B(n17617), .ZN(
        n17618) );
  NAND3_X1 U20799 ( .A1(n17620), .A2(n17619), .A3(n17618), .ZN(P3_U2656) );
  AOI211_X1 U20800 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17644), .A(n17621), .B(
        n17805), .ZN(n17622) );
  NOR2_X1 U20801 ( .A1(n19022), .A2(n17622), .ZN(n17633) );
  INV_X1 U20802 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17625) );
  OAI22_X1 U20803 ( .A1(n17625), .A2(n17801), .B1(n17768), .B2(n18135), .ZN(
        n17630) );
  NAND2_X1 U20804 ( .A1(n18700), .A2(n17623), .ZN(n17624) );
  AOI21_X1 U20805 ( .B1(n17625), .B2(n17624), .A(n18647), .ZN(n18694) );
  NOR2_X1 U20806 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18816), .ZN(
        n17789) );
  NAND2_X1 U20807 ( .A1(n17149), .A2(n17789), .ZN(n17711) );
  INV_X1 U20808 ( .A(n17711), .ZN(n17717) );
  AOI21_X1 U20809 ( .B1(n17626), .B2(n17717), .A(n10301), .ZN(n17688) );
  AOI21_X1 U20810 ( .B1(n17748), .B2(n17627), .A(n17688), .ZN(n17655) );
  OAI21_X1 U20811 ( .B1(n18700), .B2(n10301), .A(n17655), .ZN(n17643) );
  OAI21_X1 U20812 ( .B1(n18694), .B2(n17643), .A(n17781), .ZN(n17628) );
  AOI21_X1 U20813 ( .B1(n18694), .B2(n17643), .A(n17628), .ZN(n17629) );
  AOI211_X1 U20814 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17631), .A(n17630), 
        .B(n17629), .ZN(n17632) );
  OAI211_X1 U20815 ( .C1(n17635), .C2(n17634), .A(n17633), .B(n17632), .ZN(
        P3_U2657) );
  NOR2_X1 U20816 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17806), .ZN(n17636) );
  AOI21_X1 U20817 ( .B1(n17637), .B2(n17636), .A(n19022), .ZN(n17648) );
  AOI21_X1 U20818 ( .B1(n17796), .B2(n17650), .A(n17785), .ZN(n17666) );
  OAI21_X1 U20819 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17806), .A(n17666), 
        .ZN(n17642) );
  INV_X1 U20820 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18722) );
  NOR2_X1 U20821 ( .A1(n18722), .A2(n18703), .ZN(n17654) );
  OAI22_X1 U20822 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17654), .B1(
        n18703), .B2(n17638), .ZN(n18705) );
  AOI211_X1 U20823 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17748), .A(
        n18705), .B(n17639), .ZN(n17641) );
  INV_X1 U20824 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18707) );
  OAI22_X1 U20825 ( .A1(n18707), .A2(n17801), .B1(n17768), .B2(n18113), .ZN(
        n17640) );
  AOI211_X1 U20826 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17642), .A(n17641), 
        .B(n17640), .ZN(n17647) );
  NAND3_X1 U20827 ( .A1(n17781), .A2(n18705), .A3(n17643), .ZN(n17646) );
  OAI211_X1 U20828 ( .C1(n17649), .C2(n18113), .A(n17774), .B(n17644), .ZN(
        n17645) );
  NAND4_X1 U20829 ( .A1(n17648), .A2(n17647), .A3(n17646), .A4(n17645), .ZN(
        P3_U2658) );
  AOI211_X1 U20830 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17669), .A(n17649), .B(
        n17805), .ZN(n17653) );
  NOR3_X1 U20831 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17806), .A3(n17650), 
        .ZN(n17652) );
  OAI22_X1 U20832 ( .A1(n18722), .A2(n17801), .B1(n17768), .B2(n18112), .ZN(
        n17651) );
  NOR4_X1 U20833 ( .A1(n19022), .A2(n17653), .A3(n17652), .A4(n17651), .ZN(
        n17659) );
  AOI21_X1 U20834 ( .B1(n18722), .B2(n18703), .A(n17654), .ZN(n18729) );
  INV_X1 U20835 ( .A(n17655), .ZN(n17657) );
  INV_X1 U20836 ( .A(n18729), .ZN(n17656) );
  OAI221_X1 U20837 ( .B1(n18729), .B2(n17657), .C1(n17656), .C2(n17655), .A(
        n17781), .ZN(n17658) );
  OAI211_X1 U20838 ( .C1(n17666), .C2(n19608), .A(n17659), .B(n17658), .ZN(
        P3_U2659) );
  NOR2_X1 U20839 ( .A1(n19604), .A2(n19602), .ZN(n17661) );
  NAND2_X1 U20840 ( .A1(n17796), .A2(n17678), .ZN(n17675) );
  INV_X1 U20841 ( .A(n17675), .ZN(n17660) );
  AOI21_X1 U20842 ( .B1(n17661), .B2(n17660), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17667) );
  OAI21_X1 U20843 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17662), .A(
        n17748), .ZN(n17663) );
  XOR2_X1 U20844 ( .A(n17664), .B(n17663), .Z(n17665) );
  OAI22_X1 U20845 ( .A1(n17667), .A2(n17666), .B1(n19566), .B2(n17665), .ZN(
        n17668) );
  AOI211_X1 U20846 ( .C1(n17800), .C2(P3_EBX_REG_11__SCAN_IN), .A(n13950), .B(
        n17668), .ZN(n17672) );
  OAI211_X1 U20847 ( .C1(n17679), .C2(n17670), .A(n17774), .B(n17669), .ZN(
        n17671) );
  OAI211_X1 U20848 ( .C1(n17801), .C2(n17673), .A(n17672), .B(n17671), .ZN(
        P3_U2660) );
  XOR2_X1 U20849 ( .A(n17688), .B(n17674), .Z(n17685) );
  NOR3_X1 U20850 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n19602), .A3(n17675), 
        .ZN(n17676) );
  AOI211_X1 U20851 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n17716), .A(
        n13950), .B(n17676), .ZN(n17684) );
  NOR2_X1 U20852 ( .A1(n17678), .A2(n17806), .ZN(n17677) );
  NOR2_X1 U20853 ( .A1(n17785), .A2(n17677), .ZN(n17702) );
  NAND3_X1 U20854 ( .A1(n17678), .A2(n17796), .A3(n19602), .ZN(n17693) );
  AOI21_X1 U20855 ( .B1(n17702), .B2(n17693), .A(n19604), .ZN(n17682) );
  AOI211_X1 U20856 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17680), .A(n17679), .B(
        n17805), .ZN(n17681) );
  AOI211_X1 U20857 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17800), .A(n17682), .B(
        n17681), .ZN(n17683) );
  OAI211_X1 U20858 ( .C1(n19566), .C2(n17685), .A(n17684), .B(n17683), .ZN(
        P3_U2661) );
  AOI21_X1 U20859 ( .B1(n17687), .B2(n17803), .A(n17686), .ZN(n17691) );
  NOR2_X1 U20860 ( .A1(n17689), .A2(n17688), .ZN(n17690) );
  AOI211_X1 U20861 ( .C1(n17748), .C2(n17691), .A(n17690), .B(n19566), .ZN(
        n17692) );
  AOI211_X1 U20862 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17716), .A(
        n13950), .B(n17692), .ZN(n17699) );
  AOI21_X1 U20863 ( .B1(n17774), .B2(n17704), .A(n17800), .ZN(n17696) );
  OR2_X1 U20864 ( .A1(n17704), .A2(n17805), .ZN(n17694) );
  OAI221_X1 U20865 ( .B1(n17696), .B2(n17695), .C1(n17694), .C2(
        P3_EBX_REG_9__SCAN_IN), .A(n17693), .ZN(n17697) );
  INV_X1 U20866 ( .A(n17697), .ZN(n17698) );
  OAI211_X1 U20867 ( .C1(n17702), .C2(n19602), .A(n17699), .B(n17698), .ZN(
        P3_U2662) );
  OAI21_X1 U20868 ( .B1(n18737), .B2(n17711), .A(n17748), .ZN(n17700) );
  XNOR2_X1 U20869 ( .A(n17701), .B(n17700), .ZN(n17709) );
  AOI21_X1 U20870 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17716), .A(
        n19022), .ZN(n17708) );
  AOI221_X1 U20871 ( .B1(n17806), .B2(n19601), .C1(n17703), .C2(n19601), .A(
        n17702), .ZN(n17706) );
  AOI211_X1 U20872 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17718), .A(n17704), .B(
        n17805), .ZN(n17705) );
  AOI211_X1 U20873 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17800), .A(n17706), .B(
        n17705), .ZN(n17707) );
  OAI211_X1 U20874 ( .C1(n19566), .C2(n17709), .A(n17708), .B(n17707), .ZN(
        P3_U2663) );
  AOI21_X1 U20875 ( .B1(n18737), .B2(n17725), .A(n17710), .ZN(n18742) );
  NAND2_X1 U20876 ( .A1(n17788), .A2(n17711), .ZN(n17726) );
  OAI22_X1 U20877 ( .A1(n18742), .A2(n17726), .B1(n17768), .B2(n17719), .ZN(
        n17715) );
  NAND4_X1 U20878 ( .A1(n17796), .A2(n17755), .A3(P3_REIP_REG_5__SCAN_IN), 
        .A4(P3_REIP_REG_4__SCAN_IN), .ZN(n17733) );
  INV_X1 U20879 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19597) );
  XOR2_X1 U20880 ( .A(P3_REIP_REG_7__SCAN_IN), .B(n19597), .Z(n17713) );
  INV_X1 U20881 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21686) );
  OAI21_X1 U20882 ( .B1(n17755), .B2(n17806), .A(n17812), .ZN(n17772) );
  AOI21_X1 U20883 ( .B1(n17796), .B2(n17712), .A(n17772), .ZN(n17735) );
  OAI22_X1 U20884 ( .A1(n17733), .A2(n17713), .B1(n21686), .B2(n17735), .ZN(
        n17714) );
  AOI211_X1 U20885 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17716), .A(
        n17715), .B(n17714), .ZN(n17722) );
  OAI211_X1 U20886 ( .C1(n17717), .C2(n10301), .A(n17781), .B(n18742), .ZN(
        n17721) );
  OAI211_X1 U20887 ( .C1(n17723), .C2(n17719), .A(n17774), .B(n17718), .ZN(
        n17720) );
  NAND4_X1 U20888 ( .A1(n17722), .A2(n19075), .A3(n17721), .A4(n17720), .ZN(
        P3_U2664) );
  AOI211_X1 U20889 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17737), .A(n17723), .B(
        n17805), .ZN(n17731) );
  INV_X1 U20890 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17739) );
  NAND2_X1 U20891 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17724), .ZN(
        n17746) );
  NOR2_X1 U20892 ( .A1(n17739), .A2(n17746), .ZN(n17734) );
  OAI21_X1 U20893 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17734), .A(
        n17725), .ZN(n18754) );
  INV_X1 U20894 ( .A(n18754), .ZN(n17728) );
  OAI21_X1 U20895 ( .B1(n17734), .B2(n10301), .A(n17809), .ZN(n17727) );
  AOI22_X1 U20896 ( .A1(n17728), .A2(n17727), .B1(n17726), .B2(n18754), .ZN(
        n17730) );
  INV_X1 U20897 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18245) );
  OAI22_X1 U20898 ( .A1(n18753), .A2(n17801), .B1(n17768), .B2(n18245), .ZN(
        n17729) );
  NOR4_X1 U20899 ( .A1(n19022), .A2(n17731), .A3(n17730), .A4(n17729), .ZN(
        n17732) );
  OAI221_X1 U20900 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17733), .C1(n19597), 
        .C2(n17735), .A(n17732), .ZN(P3_U2665) );
  AOI21_X1 U20901 ( .B1(n17739), .B2(n17746), .A(n17734), .ZN(n18760) );
  OAI21_X1 U20902 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17746), .A(
        n17748), .ZN(n17747) );
  XNOR2_X1 U20903 ( .A(n18760), .B(n17747), .ZN(n17742) );
  NAND3_X1 U20904 ( .A1(n17796), .A2(n17755), .A3(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n17736) );
  AOI21_X1 U20905 ( .B1(n13980), .B2(n17736), .A(n17735), .ZN(n17741) );
  OAI211_X1 U20906 ( .C1(n17754), .C2(n17744), .A(n17774), .B(n17737), .ZN(
        n17738) );
  OAI21_X1 U20907 ( .B1(n17801), .B2(n17739), .A(n17738), .ZN(n17740) );
  AOI211_X1 U20908 ( .C1(n17742), .C2(n17781), .A(n17741), .B(n17740), .ZN(
        n17743) );
  OAI211_X1 U20909 ( .C1(n17768), .C2(n17744), .A(n17743), .B(n19075), .ZN(
        P3_U2666) );
  NOR2_X1 U20910 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17745), .ZN(
        n18770) );
  NOR2_X1 U20911 ( .A1(n18816), .A2(n17745), .ZN(n17763) );
  OAI21_X1 U20912 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17763), .A(
        n17746), .ZN(n18777) );
  INV_X1 U20913 ( .A(n18777), .ZN(n17749) );
  AOI22_X1 U20914 ( .A1(n17749), .A2(n17748), .B1(n17747), .B2(n18777), .ZN(
        n17750) );
  AOI21_X1 U20915 ( .B1(n18770), .B2(n17789), .A(n17750), .ZN(n17762) );
  AOI21_X1 U20916 ( .B1(n17752), .B2(n17878), .A(n17783), .ZN(n17753) );
  AOI211_X1 U20917 ( .C1(n17800), .C2(P3_EBX_REG_4__SCAN_IN), .A(n13950), .B(
        n17753), .ZN(n17761) );
  AOI211_X1 U20918 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17773), .A(n17754), .B(
        n17805), .ZN(n17759) );
  NAND2_X1 U20919 ( .A1(n17796), .A2(n17755), .ZN(n17757) );
  OAI22_X1 U20920 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17757), .B1(n17756), 
        .B2(n17801), .ZN(n17758) );
  AOI211_X1 U20921 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n17772), .A(n17759), .B(
        n17758), .ZN(n17760) );
  OAI211_X1 U20922 ( .C1(n17762), .C2(n19566), .A(n17761), .B(n17760), .ZN(
        P3_U2667) );
  INV_X1 U20923 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17777) );
  OAI21_X1 U20924 ( .B1(n17806), .B2(n17795), .A(n19593), .ZN(n17771) );
  NAND2_X1 U20925 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17782) );
  AOI21_X1 U20926 ( .B1(n17777), .B2(n17782), .A(n17763), .ZN(n18788) );
  NOR2_X1 U20927 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17782), .ZN(
        n17786) );
  NOR2_X1 U20928 ( .A1(n17786), .A2(n10301), .ZN(n17765) );
  OAI21_X1 U20929 ( .B1(n18788), .B2(n17765), .A(n17781), .ZN(n17764) );
  AOI21_X1 U20930 ( .B1(n18788), .B2(n17765), .A(n17764), .ZN(n17770) );
  AOI21_X1 U20931 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17766), .A(
        n9601), .ZN(n17767) );
  OAI22_X1 U20932 ( .A1(n17768), .A2(n18257), .B1(n17783), .B2(n17767), .ZN(
        n17769) );
  AOI211_X1 U20933 ( .C1(n17772), .C2(n17771), .A(n17770), .B(n17769), .ZN(
        n17776) );
  OAI211_X1 U20934 ( .C1(n17778), .C2(n18257), .A(n17774), .B(n17773), .ZN(
        n17775) );
  OAI211_X1 U20935 ( .C1(n17801), .C2(n17777), .A(n17776), .B(n17775), .ZN(
        P3_U2668) );
  INV_X1 U20936 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18808) );
  NAND2_X1 U20937 ( .A1(n9868), .A2(n9870), .ZN(n17779) );
  AOI211_X1 U20938 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17779), .A(n17778), .B(
        n17805), .ZN(n17794) );
  NAND2_X1 U20939 ( .A1(n17781), .A2(n10301), .ZN(n17792) );
  OAI21_X1 U20940 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17782), .ZN(n18802) );
  INV_X1 U20941 ( .A(n17783), .ZN(n19697) );
  AOI22_X1 U20942 ( .A1(n17785), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19697), 
        .B2(n17784), .ZN(n17791) );
  INV_X1 U20943 ( .A(n17786), .ZN(n17787) );
  OAI211_X1 U20944 ( .C1(n17789), .C2(n18802), .A(n17788), .B(n17787), .ZN(
        n17790) );
  OAI211_X1 U20945 ( .C1(n17792), .C2(n18802), .A(n17791), .B(n17790), .ZN(
        n17793) );
  AOI211_X1 U20946 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17800), .A(n17794), .B(
        n17793), .ZN(n17798) );
  OAI211_X1 U20947 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17796), .B(n17795), .ZN(n17797) );
  OAI211_X1 U20948 ( .C1(n17801), .C2(n18808), .A(n17798), .B(n17797), .ZN(
        P3_U2669) );
  AOI22_X1 U20949 ( .A1(n17800), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17799), .B2(
        n19697), .ZN(n17811) );
  OAI21_X1 U20950 ( .B1(n17803), .B2(n17802), .A(n17801), .ZN(n17808) );
  NOR2_X1 U20951 ( .A1(n9868), .A2(n9870), .ZN(n18262) );
  INV_X1 U20952 ( .A(n18262), .ZN(n17804) );
  OAI21_X1 U20953 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17804), .ZN(n18268) );
  OAI22_X1 U20954 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17806), .B1(n17805), 
        .B2(n18268), .ZN(n17807) );
  AOI221_X1 U20955 ( .B1(n17809), .B2(n18816), .C1(n17808), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17807), .ZN(n17810) );
  OAI211_X1 U20956 ( .C1(n17812), .C2(n13988), .A(n17811), .B(n17810), .ZN(
        P3_U2670) );
  NAND2_X1 U20957 ( .A1(n17814), .A2(n17813), .ZN(n17815) );
  NAND2_X1 U20958 ( .A1(n17815), .A2(n18266), .ZN(n17933) );
  INV_X1 U20959 ( .A(n18227), .ZN(n18122) );
  INV_X1 U20960 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17817) );
  AOI22_X1 U20961 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17816) );
  OAI21_X1 U20962 ( .B1(n9588), .B2(n17817), .A(n17816), .ZN(n17818) );
  AOI21_X1 U20963 ( .B1(n18122), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17818), .ZN(n17821) );
  AOI22_X1 U20964 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U20965 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17819) );
  NAND3_X1 U20966 ( .A1(n17821), .A2(n17820), .A3(n17819), .ZN(n17827) );
  AOI22_X1 U20967 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U20968 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17824) );
  AOI22_X1 U20969 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17823) );
  AOI22_X1 U20970 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17822) );
  NAND4_X1 U20971 ( .A1(n17825), .A2(n17824), .A3(n17823), .A4(n17822), .ZN(
        n17826) );
  NOR2_X1 U20972 ( .A1(n17827), .A2(n17826), .ZN(n17939) );
  INV_X1 U20973 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18007) );
  INV_X1 U20974 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17828) );
  OAI22_X1 U20975 ( .A1(n17919), .A2(n18014), .B1(n18060), .B2(n17828), .ZN(
        n17832) );
  INV_X1 U20976 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17830) );
  INV_X1 U20977 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17829) );
  OAI22_X1 U20978 ( .A1(n9588), .A2(n17830), .B1(n10620), .B2(n17829), .ZN(
        n17831) );
  AOI211_X1 U20979 ( .C1(n18043), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17832), .B(n17831), .ZN(n17834) );
  AOI22_X1 U20980 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17833) );
  OAI211_X1 U20981 ( .C1(n18227), .C2(n18007), .A(n17834), .B(n17833), .ZN(
        n17840) );
  AOI22_X1 U20982 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U20983 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U20984 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U20985 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17835) );
  NAND4_X1 U20986 ( .A1(n17838), .A2(n17837), .A3(n17836), .A4(n17835), .ZN(
        n17839) );
  NOR2_X1 U20987 ( .A1(n17840), .A2(n17839), .ZN(n17948) );
  INV_X1 U20988 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17847) );
  AOI22_X1 U20989 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U20990 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17841) );
  OAI211_X1 U20991 ( .C1(n9603), .C2(n17843), .A(n17842), .B(n17841), .ZN(
        n17844) );
  INV_X1 U20992 ( .A(n17844), .ZN(n17846) );
  AOI22_X1 U20993 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17845) );
  OAI211_X1 U20994 ( .C1(n18227), .C2(n17847), .A(n17846), .B(n17845), .ZN(
        n17853) );
  AOI22_X1 U20995 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U20996 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U20997 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17849) );
  AOI22_X1 U20998 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17848) );
  NAND4_X1 U20999 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n17848), .ZN(
        n17852) );
  NOR2_X1 U21000 ( .A1(n17853), .A2(n17852), .ZN(n17959) );
  INV_X1 U21001 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U21002 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17854) );
  OAI21_X1 U21003 ( .B1(n9588), .B2(n17855), .A(n17854), .ZN(n17856) );
  AOI21_X1 U21004 ( .B1(n18122), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17856), .ZN(n17859) );
  AOI22_X1 U21005 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17858) );
  AOI22_X1 U21006 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17857) );
  NAND3_X1 U21007 ( .A1(n17859), .A2(n17858), .A3(n17857), .ZN(n17865) );
  AOI22_X1 U21008 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17863) );
  AOI22_X1 U21009 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U21010 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17861) );
  AOI22_X1 U21011 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9610), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17860) );
  NAND4_X1 U21012 ( .A1(n17863), .A2(n17862), .A3(n17861), .A4(n17860), .ZN(
        n17864) );
  NOR2_X1 U21013 ( .A1(n17865), .A2(n17864), .ZN(n17969) );
  INV_X1 U21014 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18097) );
  INV_X1 U21015 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17916) );
  AOI22_X1 U21016 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9591), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17867) );
  AOI22_X1 U21017 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17866) );
  OAI211_X1 U21018 ( .C1(n9603), .C2(n17916), .A(n17867), .B(n17866), .ZN(
        n17868) );
  INV_X1 U21019 ( .A(n17868), .ZN(n17870) );
  AOI22_X1 U21020 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17869) );
  OAI211_X1 U21021 ( .C1(n18097), .C2(n18227), .A(n17870), .B(n17869), .ZN(
        n17876) );
  AOI22_X1 U21022 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n18235), .ZN(n17874) );
  AOI22_X1 U21023 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17873) );
  AOI22_X1 U21024 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17872) );
  AOI22_X1 U21025 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17871) );
  NAND4_X1 U21026 ( .A1(n17874), .A2(n17873), .A3(n17872), .A4(n17871), .ZN(
        n17875) );
  NOR2_X1 U21027 ( .A1(n17876), .A2(n17875), .ZN(n17968) );
  NOR2_X1 U21028 ( .A1(n17969), .A2(n17968), .ZN(n17964) );
  INV_X1 U21029 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17879) );
  INV_X1 U21030 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17877) );
  OAI22_X1 U21031 ( .A1(n9588), .A2(n17879), .B1(n17878), .B2(n17877), .ZN(
        n17884) );
  AOI22_X1 U21032 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U21033 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17880) );
  OAI211_X1 U21034 ( .C1(n9602), .C2(n17882), .A(n17881), .B(n17880), .ZN(
        n17883) );
  AOI211_X1 U21035 ( .C1(n18122), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n17884), .B(n17883), .ZN(n17892) );
  INV_X1 U21036 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18203) );
  NOR2_X1 U21037 ( .A1(n18125), .A2(n18203), .ZN(n17888) );
  OAI22_X1 U21038 ( .A1(n17919), .A2(n17886), .B1(n18123), .B2(n17885), .ZN(
        n17887) );
  AOI211_X1 U21039 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n18233), .A(
        n17888), .B(n17887), .ZN(n17891) );
  AOI22_X1 U21040 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17890) );
  AOI22_X1 U21041 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17889) );
  NAND4_X1 U21042 ( .A1(n17892), .A2(n17891), .A3(n17890), .A4(n17889), .ZN(
        n17963) );
  NAND2_X1 U21043 ( .A1(n17964), .A2(n17963), .ZN(n17962) );
  NOR2_X1 U21044 ( .A1(n17959), .A2(n17962), .ZN(n17954) );
  INV_X1 U21045 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17893) );
  INV_X1 U21046 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n21657) );
  OAI22_X1 U21047 ( .A1(n9588), .A2(n17893), .B1(n21657), .B2(n17878), .ZN(
        n17898) );
  AOI22_X1 U21048 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17895) );
  AOI22_X1 U21049 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U21050 ( .C1(n9602), .C2(n17896), .A(n17895), .B(n17894), .ZN(
        n17897) );
  AOI211_X1 U21051 ( .C1(n18122), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n17898), .B(n17897), .ZN(n17905) );
  NOR2_X1 U21052 ( .A1(n18123), .A2(n17899), .ZN(n17901) );
  INV_X1 U21053 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18170) );
  INV_X1 U21054 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18172) );
  OAI22_X1 U21055 ( .A1(n9761), .A2(n18170), .B1(n18125), .B2(n18172), .ZN(
        n17900) );
  AOI211_X1 U21056 ( .C1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .C2(n9597), .A(
        n17901), .B(n17900), .ZN(n17904) );
  AOI22_X1 U21057 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U21058 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17902) );
  NAND4_X1 U21059 ( .A1(n17905), .A2(n17904), .A3(n17903), .A4(n17902), .ZN(
        n17953) );
  NAND2_X1 U21060 ( .A1(n17954), .A2(n17953), .ZN(n17952) );
  NOR2_X1 U21061 ( .A1(n17948), .A2(n17952), .ZN(n18289) );
  AOI22_X1 U21062 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U21063 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17908) );
  AOI22_X1 U21064 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U21065 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17906) );
  NAND4_X1 U21066 ( .A1(n17909), .A2(n17908), .A3(n17907), .A4(n17906), .ZN(
        n17915) );
  AOI22_X1 U21067 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U21068 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17910) );
  OAI211_X1 U21069 ( .C1(n21633), .C2(n9603), .A(n17911), .B(n17910), .ZN(
        n17914) );
  INV_X1 U21070 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17988) );
  AOI22_X1 U21071 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17912) );
  OAI21_X1 U21072 ( .B1(n18227), .B2(n17988), .A(n17912), .ZN(n17913) );
  OR3_X1 U21073 ( .A1(n17915), .A2(n17914), .A3(n17913), .ZN(n18288) );
  NAND2_X1 U21074 ( .A1(n18289), .A2(n18288), .ZN(n18287) );
  NOR2_X1 U21075 ( .A1(n17939), .A2(n18287), .ZN(n17938) );
  INV_X1 U21076 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17925) );
  INV_X1 U21077 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17917) );
  OAI22_X1 U21078 ( .A1(n17917), .A2(n13880), .B1(n18095), .B2(n17916), .ZN(
        n17922) );
  INV_X1 U21079 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17920) );
  OAI22_X1 U21080 ( .A1(n9588), .A2(n17920), .B1(n17919), .B2(n17918), .ZN(
        n17921) );
  AOI211_X1 U21081 ( .C1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n9590), .A(
        n17922), .B(n17921), .ZN(n17924) );
  AOI22_X1 U21082 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18234), .B1(
        n9612), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17923) );
  OAI211_X1 U21083 ( .C1(n18227), .C2(n17925), .A(n17924), .B(n17923), .ZN(
        n17931) );
  AOI22_X1 U21084 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U21085 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U21086 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17927) );
  AOI22_X1 U21087 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17926) );
  NAND4_X1 U21088 ( .A1(n17929), .A2(n17928), .A3(n17927), .A4(n17926), .ZN(
        n17930) );
  NOR2_X1 U21089 ( .A1(n17931), .A2(n17930), .ZN(n17932) );
  XOR2_X1 U21090 ( .A(n17938), .B(n17932), .Z(n18282) );
  OAI22_X1 U21091 ( .A1(n17934), .A2(n17933), .B1(n18282), .B2(n18266), .ZN(
        P3_U2673) );
  NAND2_X1 U21092 ( .A1(n17935), .A2(n18272), .ZN(n18267) );
  INV_X1 U21093 ( .A(n18267), .ZN(n18269) );
  NAND2_X1 U21094 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17971), .ZN(n17961) );
  AOI21_X1 U21095 ( .B1(n17939), .B2(n18287), .A(n17938), .ZN(n18283) );
  NOR2_X1 U21096 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17967), .ZN(n17940) );
  AOI22_X1 U21097 ( .A1(n18270), .A2(n18283), .B1(n17941), .B2(n17940), .ZN(
        n17942) );
  OAI21_X1 U21098 ( .B1(n17945), .B2(n17943), .A(n17942), .ZN(P3_U2674) );
  INV_X1 U21099 ( .A(n17951), .ZN(n17957) );
  NAND2_X1 U21100 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17957), .ZN(n17947) );
  INV_X1 U21101 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17946) );
  OAI211_X1 U21102 ( .C1(n18289), .C2(n18288), .A(n18270), .B(n18287), .ZN(
        n17944) );
  OAI221_X1 U21103 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17947), .C1(n17946), 
        .C2(n17945), .A(n17944), .ZN(P3_U2675) );
  AOI21_X1 U21104 ( .B1(n17948), .B2(n17952), .A(n18289), .ZN(n18295) );
  AOI22_X1 U21105 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17949), .B1(n18270), 
        .B2(n18295), .ZN(n17950) );
  OAI21_X1 U21106 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17951), .A(n17950), .ZN(
        P3_U2676) );
  OAI21_X1 U21107 ( .B1(n17954), .B2(n17953), .A(n17952), .ZN(n18302) );
  NAND2_X1 U21108 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17966), .ZN(n17958) );
  INV_X1 U21109 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17956) );
  OAI222_X1 U21110 ( .A1(n18302), .A2(n18184), .B1(n17958), .B2(n17957), .C1(
        n17956), .C2(n17955), .ZN(P3_U2677) );
  XNOR2_X1 U21111 ( .A(n17959), .B(n17962), .ZN(n18307) );
  NAND3_X1 U21112 ( .A1(n17961), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n18266), 
        .ZN(n17960) );
  OAI221_X1 U21113 ( .B1(n17961), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n18184), 
        .C2(n18307), .A(n17960), .ZN(P3_U2678) );
  AOI21_X1 U21114 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18266), .A(n17971), .ZN(
        n17965) );
  OAI21_X1 U21115 ( .B1(n17964), .B2(n17963), .A(n17962), .ZN(n18312) );
  OAI22_X1 U21116 ( .A1(n17966), .A2(n17965), .B1(n18184), .B2(n18312), .ZN(
        P3_U2679) );
  INV_X1 U21117 ( .A(n17967), .ZN(n17986) );
  AOI21_X1 U21118 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18266), .A(n17986), .ZN(
        n17970) );
  XNOR2_X1 U21119 ( .A(n17969), .B(n17968), .ZN(n18317) );
  OAI22_X1 U21120 ( .A1(n17971), .A2(n17970), .B1(n18266), .B2(n18317), .ZN(
        P3_U2680) );
  AOI21_X1 U21121 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18266), .A(n17972), .ZN(
        n17985) );
  INV_X1 U21122 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U21123 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17973) );
  OAI21_X1 U21124 ( .B1(n9588), .B2(n17974), .A(n17973), .ZN(n17975) );
  AOI21_X1 U21125 ( .B1(n18122), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17975), .ZN(n17978) );
  AOI22_X1 U21126 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21127 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17976) );
  NAND3_X1 U21128 ( .A1(n17978), .A2(n17977), .A3(n17976), .ZN(n17984) );
  AOI22_X1 U21129 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U21130 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U21131 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17980) );
  AOI22_X1 U21132 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17979) );
  NAND4_X1 U21133 ( .A1(n17982), .A2(n17981), .A3(n17980), .A4(n17979), .ZN(
        n17983) );
  NOR2_X1 U21134 ( .A1(n17984), .A2(n17983), .ZN(n18321) );
  OAI22_X1 U21135 ( .A1(n17986), .A2(n17985), .B1(n18321), .B2(n18266), .ZN(
        P3_U2681) );
  NAND2_X1 U21136 ( .A1(n18266), .A2(n17987), .ZN(n18024) );
  INV_X1 U21137 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17989) );
  OAI22_X1 U21138 ( .A1(n9588), .A2(n17989), .B1(n17878), .B2(n17988), .ZN(
        n17994) );
  INV_X1 U21139 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U21140 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21141 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17990) );
  OAI211_X1 U21142 ( .C1(n9602), .C2(n17992), .A(n17991), .B(n17990), .ZN(
        n17993) );
  AOI211_X1 U21143 ( .C1(n18122), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17994), .B(n17993), .ZN(n18003) );
  NOR2_X1 U21144 ( .A1(n18123), .A2(n17995), .ZN(n17999) );
  OAI22_X1 U21145 ( .A1(n9761), .A2(n17997), .B1(n18125), .B2(n17996), .ZN(
        n17998) );
  AOI211_X1 U21146 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n17999), .B(n17998), .ZN(n18002) );
  AOI22_X1 U21147 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U21148 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18000) );
  NAND4_X1 U21149 ( .A1(n18003), .A2(n18002), .A3(n18001), .A4(n18000), .ZN(
        n18326) );
  NAND2_X1 U21150 ( .A1(n18270), .A2(n18326), .ZN(n18004) );
  OAI221_X1 U21151 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18006), .C1(n18005), 
        .C2(n18024), .A(n18004), .ZN(P3_U2682) );
  INV_X1 U21152 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18008) );
  OAI22_X1 U21153 ( .A1(n9588), .A2(n18008), .B1(n17878), .B2(n18007), .ZN(
        n18012) );
  AOI22_X1 U21154 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U21155 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18009) );
  OAI211_X1 U21156 ( .C1(n21664), .C2(n9603), .A(n18010), .B(n18009), .ZN(
        n18011) );
  AOI211_X1 U21157 ( .C1(n18122), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n18012), .B(n18011), .ZN(n18021) );
  NOR2_X1 U21158 ( .A1(n18123), .A2(n18013), .ZN(n18017) );
  OAI22_X1 U21159 ( .A1(n9761), .A2(n18015), .B1(n18125), .B2(n18014), .ZN(
        n18016) );
  AOI211_X1 U21160 ( .C1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .C2(n14134), .A(
        n18017), .B(n18016), .ZN(n18020) );
  AOI22_X1 U21161 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U21162 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18018) );
  NAND4_X1 U21163 ( .A1(n18021), .A2(n18020), .A3(n18019), .A4(n18018), .ZN(
        n18330) );
  NOR2_X1 U21164 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18038), .ZN(n18022) );
  AOI22_X1 U21165 ( .A1(n18270), .A2(n18330), .B1(n9647), .B2(n18022), .ZN(
        n18023) );
  OAI21_X1 U21166 ( .B1(n10320), .B2(n18024), .A(n18023), .ZN(P3_U2683) );
  INV_X1 U21167 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U21168 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18025) );
  OAI21_X1 U21169 ( .B1(n9588), .B2(n18026), .A(n18025), .ZN(n18027) );
  AOI21_X1 U21170 ( .B1(n18122), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18027), .ZN(n18030) );
  AOI22_X1 U21171 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U21172 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18028) );
  NAND3_X1 U21173 ( .A1(n18030), .A2(n18029), .A3(n18028), .ZN(n18036) );
  AOI22_X1 U21174 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U21175 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U21176 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18032) );
  AOI22_X1 U21177 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9612), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18031) );
  NAND4_X1 U21178 ( .A1(n18034), .A2(n18033), .A3(n18032), .A4(n18031), .ZN(
        n18035) );
  NOR2_X1 U21179 ( .A1(n18036), .A2(n18035), .ZN(n18339) );
  NOR2_X1 U21180 ( .A1(n18270), .A2(n18037), .ZN(n18055) );
  AOI22_X1 U21181 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18055), .B1(n9647), .B2(
        n18038), .ZN(n18039) );
  OAI21_X1 U21182 ( .B1(n18339), .B2(n18184), .A(n18039), .ZN(P3_U2684) );
  INV_X1 U21183 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18040) );
  OAI22_X1 U21184 ( .A1(n18123), .A2(n18041), .B1(n13880), .B2(n18040), .ZN(
        n18042) );
  AOI21_X1 U21185 ( .B1(n18043), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n18042), .ZN(n18047) );
  AOI22_X1 U21186 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18046) );
  AOI22_X1 U21187 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18045) );
  NAND2_X1 U21188 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n18044) );
  NAND4_X1 U21189 ( .A1(n18047), .A2(n18046), .A3(n18045), .A4(n18044), .ZN(
        n18053) );
  AOI22_X1 U21190 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U21191 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U21192 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U21193 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18048) );
  NAND4_X1 U21194 ( .A1(n18051), .A2(n18050), .A3(n18049), .A4(n18048), .ZN(
        n18052) );
  NOR2_X1 U21195 ( .A1(n18053), .A2(n18052), .ZN(n18344) );
  OAI21_X1 U21196 ( .B1(n18075), .B2(n18074), .A(n18054), .ZN(n18056) );
  NAND2_X1 U21197 ( .A1(n18056), .A2(n18055), .ZN(n18057) );
  OAI21_X1 U21198 ( .B1(n18344), .B2(n18184), .A(n18057), .ZN(P3_U2685) );
  INV_X1 U21199 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18066) );
  INV_X1 U21200 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n21655) );
  INV_X1 U21201 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18058) );
  OAI22_X1 U21202 ( .A1(n18123), .A2(n21655), .B1(n18095), .B2(n18058), .ZN(
        n18063) );
  INV_X1 U21203 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18061) );
  INV_X1 U21204 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18059) );
  OAI22_X1 U21205 ( .A1(n9588), .A2(n18061), .B1(n18060), .B2(n18059), .ZN(
        n18062) );
  AOI211_X1 U21206 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n18063), .B(n18062), .ZN(n18065) );
  AOI22_X1 U21207 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18064) );
  OAI211_X1 U21208 ( .C1(n18227), .C2(n18066), .A(n18065), .B(n18064), .ZN(
        n18072) );
  AOI22_X1 U21209 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U21210 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18069) );
  AOI22_X1 U21211 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U21212 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18067) );
  NAND4_X1 U21213 ( .A1(n18070), .A2(n18069), .A3(n18068), .A4(n18067), .ZN(
        n18071) );
  NOR2_X1 U21214 ( .A1(n18072), .A2(n18071), .ZN(n18349) );
  NOR2_X1 U21215 ( .A1(n18270), .A2(n18073), .ZN(n18091) );
  INV_X1 U21216 ( .A(n18074), .ZN(n18076) );
  AOI22_X1 U21217 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18091), .B1(n18076), 
        .B2(n18075), .ZN(n18077) );
  OAI21_X1 U21218 ( .B1(n18349), .B2(n18184), .A(n18077), .ZN(P3_U2686) );
  INV_X1 U21219 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U21220 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U21221 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18078) );
  OAI211_X1 U21222 ( .C1(n9602), .C2(n18080), .A(n18079), .B(n18078), .ZN(
        n18081) );
  INV_X1 U21223 ( .A(n18081), .ZN(n18083) );
  AOI22_X1 U21224 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18082) );
  OAI211_X1 U21225 ( .C1(n18227), .C2(n18084), .A(n18083), .B(n18082), .ZN(
        n18090) );
  AOI22_X1 U21226 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18088) );
  AOI22_X1 U21227 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18087) );
  AOI22_X1 U21228 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18086) );
  AOI22_X1 U21229 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18085) );
  NAND4_X1 U21230 ( .A1(n18088), .A2(n18087), .A3(n18086), .A4(n18085), .ZN(
        n18089) );
  NOR2_X1 U21231 ( .A1(n18090), .A2(n18089), .ZN(n18355) );
  INV_X1 U21232 ( .A(n18110), .ZN(n18092) );
  OAI21_X1 U21233 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18092), .A(n18091), .ZN(
        n18093) );
  OAI21_X1 U21234 ( .B1(n18355), .B2(n18184), .A(n18093), .ZN(P3_U2687) );
  INV_X1 U21235 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18103) );
  INV_X1 U21236 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18096) );
  OAI22_X1 U21237 ( .A1(n18096), .A2(n13880), .B1(n18095), .B2(n18094), .ZN(
        n18100) );
  INV_X1 U21238 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18098) );
  OAI22_X1 U21239 ( .A1(n9588), .A2(n18098), .B1(n18097), .B2(n17878), .ZN(
        n18099) );
  AOI211_X1 U21240 ( .C1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .C2(n18043), .A(
        n18100), .B(n18099), .ZN(n18102) );
  AOI22_X1 U21241 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18101) );
  OAI211_X1 U21242 ( .C1(n18227), .C2(n18103), .A(n18102), .B(n18101), .ZN(
        n18109) );
  AOI22_X1 U21243 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U21244 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18106) );
  AOI22_X1 U21245 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U21246 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18104) );
  NAND4_X1 U21247 ( .A1(n18107), .A2(n18106), .A3(n18105), .A4(n18104), .ZN(
        n18108) );
  NOR2_X1 U21248 ( .A1(n18109), .A2(n18108), .ZN(n18360) );
  OAI21_X1 U21249 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n9686), .A(n18110), .ZN(
        n18111) );
  AOI22_X1 U21250 ( .A1(n18270), .A2(n18360), .B1(n18111), .B2(n18184), .ZN(
        P3_U2688) );
  NOR3_X1 U21251 ( .A1(n19131), .A2(n18112), .A3(n18183), .ZN(n18150) );
  NAND2_X1 U21252 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18150), .ZN(n18149) );
  NOR2_X1 U21253 ( .A1(n18270), .A2(n18150), .ZN(n18165) );
  AOI21_X1 U21254 ( .B1(n18269), .B2(n18113), .A(n18165), .ZN(n18134) );
  INV_X1 U21255 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18115) );
  INV_X1 U21256 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18114) );
  OAI22_X1 U21257 ( .A1(n9588), .A2(n18115), .B1(n17878), .B2(n18114), .ZN(
        n18121) );
  INV_X1 U21258 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U21259 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U21260 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18117) );
  OAI211_X1 U21261 ( .C1(n9602), .C2(n18119), .A(n18118), .B(n18117), .ZN(
        n18120) );
  AOI211_X1 U21262 ( .C1(n18122), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18121), .B(n18120), .ZN(n18132) );
  INV_X1 U21263 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21667) );
  NOR2_X1 U21264 ( .A1(n18123), .A2(n21667), .ZN(n18128) );
  OAI22_X1 U21265 ( .A1(n9761), .A2(n18126), .B1(n18125), .B2(n18124), .ZN(
        n18127) );
  AOI211_X1 U21266 ( .C1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .C2(n9597), .A(
        n18128), .B(n18127), .ZN(n18131) );
  AOI22_X1 U21267 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U21268 ( .A1(n9612), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18129) );
  NAND4_X1 U21269 ( .A1(n18132), .A2(n18131), .A3(n18130), .A4(n18129), .ZN(
        n18362) );
  NAND2_X1 U21270 ( .A1(n18270), .A2(n18362), .ZN(n18133) );
  OAI221_X1 U21271 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18149), .C1(n18135), 
        .C2(n18134), .A(n18133), .ZN(P3_U2689) );
  INV_X1 U21272 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18142) );
  INV_X1 U21273 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U21274 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U21275 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18136) );
  OAI211_X1 U21276 ( .C1(n9602), .C2(n18138), .A(n18137), .B(n18136), .ZN(
        n18139) );
  INV_X1 U21277 ( .A(n18139), .ZN(n18141) );
  AOI22_X1 U21278 ( .A1(n13898), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18140) );
  OAI211_X1 U21279 ( .C1(n18227), .C2(n18142), .A(n18141), .B(n18140), .ZN(
        n18148) );
  AOI22_X1 U21280 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18146) );
  AOI22_X1 U21281 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18145) );
  AOI22_X1 U21282 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U21283 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18143) );
  NAND4_X1 U21284 ( .A1(n18146), .A2(n18145), .A3(n18144), .A4(n18143), .ZN(
        n18147) );
  NOR2_X1 U21285 ( .A1(n18148), .A2(n18147), .ZN(n18366) );
  OAI211_X1 U21286 ( .C1(n18150), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18266), .B(
        n18149), .ZN(n18151) );
  OAI21_X1 U21287 ( .B1(n18366), .B2(n18184), .A(n18151), .ZN(P3_U2690) );
  INV_X1 U21288 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18158) );
  INV_X1 U21289 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18154) );
  AOI22_X1 U21290 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U21291 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18210), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18152) );
  OAI211_X1 U21292 ( .C1(n9603), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        n18155) );
  INV_X1 U21293 ( .A(n18155), .ZN(n18157) );
  AOI22_X1 U21294 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18156) );
  OAI211_X1 U21295 ( .C1(n18227), .C2(n18158), .A(n18157), .B(n18156), .ZN(
        n18164) );
  AOI22_X1 U21296 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U21297 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21298 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U21299 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18159) );
  NAND4_X1 U21300 ( .A1(n18162), .A2(n18161), .A3(n18160), .A4(n18159), .ZN(
        n18163) );
  NOR2_X1 U21301 ( .A1(n18164), .A2(n18163), .ZN(n18370) );
  INV_X1 U21302 ( .A(n18183), .ZN(n18166) );
  OAI21_X1 U21303 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18166), .A(n18165), .ZN(
        n18167) );
  OAI21_X1 U21304 ( .B1(n18370), .B2(n18184), .A(n18167), .ZN(P3_U2691) );
  AOI22_X1 U21305 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U21306 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18175) );
  NAND2_X1 U21307 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n18169) );
  NAND2_X1 U21308 ( .A1(n10621), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n18168) );
  OAI211_X1 U21309 ( .C1(n9603), .C2(n18170), .A(n18169), .B(n18168), .ZN(
        n18171) );
  INV_X1 U21310 ( .A(n18171), .ZN(n18174) );
  OR2_X1 U21311 ( .A1(n18227), .A2(n18172), .ZN(n18173) );
  NAND4_X1 U21312 ( .A1(n18176), .A2(n18175), .A3(n18174), .A4(n18173), .ZN(
        n18182) );
  AOI22_X1 U21313 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U21314 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U21315 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18178) );
  AOI22_X1 U21316 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18177) );
  NAND4_X1 U21317 ( .A1(n18180), .A2(n18179), .A3(n18178), .A4(n18177), .ZN(
        n18181) );
  NOR2_X1 U21318 ( .A1(n18182), .A2(n18181), .ZN(n18373) );
  OAI21_X1 U21319 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n9754), .A(n18183), .ZN(
        n18185) );
  AOI22_X1 U21320 ( .A1(n18270), .A2(n18373), .B1(n18185), .B2(n18184), .ZN(
        P3_U2692) );
  NAND2_X1 U21321 ( .A1(n18266), .A2(n18197), .ZN(n18217) );
  AOI22_X1 U21322 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18189) );
  AOI22_X1 U21323 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U21324 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U21325 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18186) );
  NAND4_X1 U21326 ( .A1(n18189), .A2(n18188), .A3(n18187), .A4(n18186), .ZN(
        n18196) );
  INV_X1 U21327 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U21328 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U21329 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18190) );
  OAI211_X1 U21330 ( .C1(n9602), .C2(n18192), .A(n18191), .B(n18190), .ZN(
        n18195) );
  AOI22_X1 U21331 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18193) );
  OAI21_X1 U21332 ( .B1(n18265), .B2(n18227), .A(n18193), .ZN(n18194) );
  OR3_X1 U21333 ( .A1(n18196), .A2(n18195), .A3(n18194), .ZN(n18377) );
  NOR3_X1 U21334 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n19131), .A3(n18197), .ZN(
        n18198) );
  AOI21_X1 U21335 ( .B1(n18270), .B2(n18377), .A(n18198), .ZN(n18199) );
  OAI21_X1 U21336 ( .B1(n18200), .B2(n18217), .A(n18199), .ZN(P3_U2693) );
  AOI22_X1 U21337 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18202) );
  NAND2_X1 U21338 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n18201) );
  OAI211_X1 U21339 ( .C1(n18203), .C2(n18227), .A(n18202), .B(n18201), .ZN(
        n18204) );
  INV_X1 U21340 ( .A(n18204), .ZN(n18208) );
  AOI22_X1 U21341 ( .A1(n14134), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U21342 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18205), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18206) );
  NAND3_X1 U21343 ( .A1(n18208), .A2(n18207), .A3(n18206), .ZN(n18216) );
  AOI22_X1 U21344 ( .A1(n18209), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U21345 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10621), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U21346 ( .A1(n18232), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U21347 ( .A1(n9604), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9611), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18211) );
  NAND4_X1 U21348 ( .A1(n18214), .A2(n18213), .A3(n18212), .A4(n18211), .ZN(
        n18215) );
  NOR2_X1 U21349 ( .A1(n18216), .A2(n18215), .ZN(n18384) );
  NOR2_X1 U21350 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n18243), .ZN(n18218) );
  OAI22_X1 U21351 ( .A1(n18384), .A2(n18184), .B1(n18218), .B2(n18217), .ZN(
        P3_U2694) );
  OAI21_X1 U21352 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18247), .A(n18266), .ZN(
        n18242) );
  AOI22_X1 U21353 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U21354 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17751), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18230) );
  INV_X1 U21355 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18223) );
  NAND2_X1 U21356 ( .A1(n18210), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n18222) );
  NAND2_X1 U21357 ( .A1(n10621), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n18221) );
  OAI211_X1 U21358 ( .C1(n9603), .C2(n18223), .A(n18222), .B(n18221), .ZN(
        n18225) );
  INV_X1 U21359 ( .A(n18225), .ZN(n18229) );
  INV_X1 U21360 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18226) );
  OR2_X1 U21361 ( .A1(n18227), .A2(n18226), .ZN(n18228) );
  NAND4_X1 U21362 ( .A1(n18231), .A2(n18230), .A3(n18229), .A4(n18228), .ZN(
        n18241) );
  AOI22_X1 U21363 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U21364 ( .A1(n18233), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18232), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18238) );
  AOI22_X1 U21365 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13898), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U21366 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18236) );
  NAND4_X1 U21367 ( .A1(n18239), .A2(n18238), .A3(n18237), .A4(n18236), .ZN(
        n18240) );
  NOR2_X1 U21368 ( .A1(n18241), .A2(n18240), .ZN(n18387) );
  OAI22_X1 U21369 ( .A1(n18243), .A2(n18242), .B1(n18387), .B2(n18266), .ZN(
        P3_U2695) );
  NAND2_X1 U21370 ( .A1(n18244), .A2(n18269), .ZN(n18248) );
  NOR2_X1 U21371 ( .A1(n18245), .A2(n18248), .ZN(n18251) );
  AOI21_X1 U21372 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18266), .A(n18251), .ZN(
        n18246) );
  OAI22_X1 U21373 ( .A1(n18247), .A2(n18246), .B1(n18103), .B2(n18184), .ZN(
        P3_U2696) );
  INV_X1 U21374 ( .A(n18248), .ZN(n18255) );
  AOI21_X1 U21375 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18266), .A(n18255), .ZN(
        n18250) );
  INV_X1 U21376 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18249) );
  OAI22_X1 U21377 ( .A1(n18251), .A2(n18250), .B1(n18249), .B2(n18184), .ZN(
        P3_U2697) );
  NOR2_X1 U21378 ( .A1(n18252), .A2(n18267), .ZN(n18263) );
  INV_X1 U21379 ( .A(n18263), .ZN(n18256) );
  NOR3_X1 U21380 ( .A1(n18253), .A2(n18257), .A3(n18256), .ZN(n18259) );
  AOI21_X1 U21381 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18266), .A(n18259), .ZN(
        n18254) );
  OAI22_X1 U21382 ( .A1(n18255), .A2(n18254), .B1(n18142), .B2(n18184), .ZN(
        P3_U2698) );
  NOR2_X1 U21383 ( .A1(n18257), .A2(n18256), .ZN(n18261) );
  AOI21_X1 U21384 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18266), .A(n18261), .ZN(
        n18258) );
  OAI22_X1 U21385 ( .A1(n18259), .A2(n18258), .B1(n18158), .B2(n18184), .ZN(
        P3_U2699) );
  AOI21_X1 U21386 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18266), .A(n18263), .ZN(
        n18260) );
  OAI22_X1 U21387 ( .A1(n18261), .A2(n18260), .B1(n18172), .B2(n18184), .ZN(
        P3_U2700) );
  AOI221_X1 U21388 ( .B1(n18262), .B2(n18272), .C1(n19131), .C2(n18272), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18264) );
  AOI211_X1 U21389 ( .C1(n18270), .C2(n18265), .A(n18264), .B(n18263), .ZN(
        P3_U2701) );
  OAI222_X1 U21390 ( .A1(n18268), .A2(n18267), .B1(n9870), .B2(n18272), .C1(
        n18203), .C2(n18266), .ZN(P3_U2702) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18270), .B1(
        n18269), .B2(n9868), .ZN(n18271) );
  OAI21_X1 U21392 ( .B1(n18272), .B2(n9868), .A(n18271), .ZN(P3_U2703) );
  INV_X1 U21393 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18419) );
  INV_X1 U21394 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18422) );
  INV_X1 U21395 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18456) );
  INV_X1 U21396 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18459) );
  NAND3_X1 U21397 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .ZN(n18393) );
  NOR4_X1 U21398 ( .A1(n18456), .A2(n18459), .A3(n18273), .A4(n18393), .ZN(
        n18383) );
  NAND4_X1 U21399 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n18274)
         );
  NAND4_X1 U21400 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n18275), .ZN(n18361) );
  NAND4_X1 U21401 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n18318)
         );
  NAND2_X1 U21402 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18290), .ZN(n18284) );
  NAND2_X1 U21403 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18279), .ZN(n18278) );
  NAND2_X1 U21404 ( .A1(n18278), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n18277) );
  NAND2_X1 U21405 ( .A1(n19127), .A2(n18357), .ZN(n18320) );
  NAND2_X1 U21406 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18350), .ZN(n18276) );
  OAI221_X1 U21407 ( .B1(n18278), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n18277), 
        .C2(n18357), .A(n18276), .ZN(P3_U2704) );
  NOR2_X2 U21408 ( .A1(n19122), .A2(n18408), .ZN(n18351) );
  AOI22_X1 U21409 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18350), .ZN(n18281) );
  OAI211_X1 U21410 ( .C1(n18279), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18408), .B(
        n18278), .ZN(n18280) );
  OAI211_X1 U21411 ( .C1(n18282), .C2(n18410), .A(n18281), .B(n18280), .ZN(
        P3_U2705) );
  INV_X1 U21412 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19123) );
  AOI22_X1 U21413 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18351), .B1(n18389), .B2(
        n18283), .ZN(n18286) );
  OAI211_X1 U21414 ( .C1(n18290), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18408), .B(
        n18284), .ZN(n18285) );
  OAI211_X1 U21415 ( .C1(n18320), .C2(n19123), .A(n18286), .B(n18285), .ZN(
        P3_U2706) );
  OAI21_X1 U21416 ( .B1(n18289), .B2(n18288), .A(n18287), .ZN(n18294) );
  AOI22_X1 U21417 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18350), .ZN(n18293) );
  AOI211_X1 U21418 ( .C1(n18419), .C2(n18296), .A(n18290), .B(n18357), .ZN(
        n18291) );
  INV_X1 U21419 ( .A(n18291), .ZN(n18292) );
  OAI211_X1 U21420 ( .C1(n18294), .C2(n18410), .A(n18293), .B(n18292), .ZN(
        P3_U2707) );
  INV_X1 U21421 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19112) );
  AOI22_X1 U21422 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18351), .B1(n18389), .B2(
        n18295), .ZN(n18298) );
  OAI211_X1 U21423 ( .C1(n9664), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18408), .B(
        n18296), .ZN(n18297) );
  OAI211_X1 U21424 ( .C1(n18320), .C2(n19112), .A(n18298), .B(n18297), .ZN(
        P3_U2708) );
  AOI22_X1 U21425 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18350), .ZN(n18301) );
  AOI211_X1 U21426 ( .C1(n18422), .C2(n18303), .A(n9664), .B(n18357), .ZN(
        n18299) );
  INV_X1 U21427 ( .A(n18299), .ZN(n18300) );
  OAI211_X1 U21428 ( .C1(n18302), .C2(n18410), .A(n18301), .B(n18300), .ZN(
        P3_U2709) );
  AOI22_X1 U21429 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18350), .ZN(n18306) );
  OAI211_X1 U21430 ( .C1(n18304), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18408), .B(
        n18303), .ZN(n18305) );
  OAI211_X1 U21431 ( .C1(n18307), .C2(n18410), .A(n18306), .B(n18305), .ZN(
        P3_U2710) );
  AOI22_X1 U21432 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18350), .ZN(n18311) );
  OAI211_X1 U21433 ( .C1(n18309), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18408), .B(
        n18308), .ZN(n18310) );
  OAI211_X1 U21434 ( .C1(n18312), .C2(n18410), .A(n18311), .B(n18310), .ZN(
        P3_U2711) );
  AOI22_X1 U21435 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18350), .ZN(n18316) );
  OAI211_X1 U21436 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18314), .A(n18408), .B(
        n18313), .ZN(n18315) );
  OAI211_X1 U21437 ( .C1(n18317), .C2(n18410), .A(n18316), .B(n18315), .ZN(
        P3_U2712) );
  NOR3_X1 U21438 ( .A1(n19131), .A2(n18352), .A3(n18318), .ZN(n18334) );
  NAND2_X1 U21439 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18334), .ZN(n18325) );
  NOR2_X1 U21440 ( .A1(n18357), .A2(n18334), .ZN(n18331) );
  AOI21_X1 U21441 ( .B1(n18382), .B2(n18431), .A(n18331), .ZN(n18324) );
  OAI22_X1 U21442 ( .A1(n18321), .A2(n18410), .B1(n19872), .B2(n18320), .ZN(
        n18322) );
  AOI21_X1 U21443 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n18351), .A(n18322), .ZN(
        n18323) );
  OAI221_X1 U21444 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n18325), .C1(n18429), 
        .C2(n18324), .A(n18323), .ZN(P3_U2713) );
  INV_X1 U21445 ( .A(n18351), .ZN(n18329) );
  AOI22_X1 U21446 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18350), .B1(n18389), .B2(
        n18326), .ZN(n18328) );
  AOI22_X1 U21447 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18331), .B1(n18334), 
        .B2(n18431), .ZN(n18327) );
  OAI211_X1 U21448 ( .C1(n19124), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2714) );
  INV_X1 U21449 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18477) );
  NOR3_X1 U21450 ( .A1(n19131), .A2(n18352), .A3(n18477), .ZN(n18335) );
  NAND3_X1 U21451 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(n18335), .ZN(n18336) );
  AOI22_X1 U21452 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18350), .B1(n18389), .B2(
        n18330), .ZN(n18333) );
  AOI22_X1 U21453 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18351), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n18331), .ZN(n18332) );
  OAI211_X1 U21454 ( .C1(n18334), .C2(n18336), .A(n18333), .B(n18332), .ZN(
        P3_U2715) );
  AOI22_X1 U21455 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18350), .ZN(n18338) );
  INV_X1 U21456 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18437) );
  INV_X1 U21457 ( .A(n18335), .ZN(n18345) );
  NOR2_X1 U21458 ( .A1(n18437), .A2(n18345), .ZN(n18340) );
  OAI211_X1 U21459 ( .C1(n18340), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18408), .B(
        n18336), .ZN(n18337) );
  OAI211_X1 U21460 ( .C1(n18339), .C2(n18410), .A(n18338), .B(n18337), .ZN(
        P3_U2716) );
  AOI22_X1 U21461 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18350), .ZN(n18343) );
  AOI211_X1 U21462 ( .C1(n18437), .C2(n18345), .A(n18340), .B(n18357), .ZN(
        n18341) );
  INV_X1 U21463 ( .A(n18341), .ZN(n18342) );
  OAI211_X1 U21464 ( .C1(n18344), .C2(n18410), .A(n18343), .B(n18342), .ZN(
        P3_U2717) );
  AOI22_X1 U21465 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18350), .ZN(n18348) );
  INV_X1 U21466 ( .A(n18352), .ZN(n18346) );
  OAI211_X1 U21467 ( .C1(n18346), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18408), .B(
        n18345), .ZN(n18347) );
  OAI211_X1 U21468 ( .C1(n18349), .C2(n18410), .A(n18348), .B(n18347), .ZN(
        P3_U2718) );
  AOI22_X1 U21469 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18351), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18350), .ZN(n18354) );
  OAI211_X1 U21470 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18356), .A(n18408), .B(
        n18352), .ZN(n18353) );
  OAI211_X1 U21471 ( .C1(n18355), .C2(n18410), .A(n18354), .B(n18353), .ZN(
        P3_U2719) );
  AOI211_X1 U21472 ( .C1(n18522), .C2(n18361), .A(n18357), .B(n18356), .ZN(
        n18358) );
  AOI21_X1 U21473 ( .B1(n18378), .B2(BUF2_REG_15__SCAN_IN), .A(n18358), .ZN(
        n18359) );
  OAI21_X1 U21474 ( .B1(n18360), .B2(n18410), .A(n18359), .ZN(P3_U2720) );
  INV_X1 U21475 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18509) );
  NAND4_X1 U21476 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18383), .A3(
        P3_EAX_REG_8__SCAN_IN), .A4(n18382), .ZN(n18380) );
  INV_X1 U21477 ( .A(n18380), .ZN(n18386) );
  NAND2_X1 U21478 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18386), .ZN(n18376) );
  NOR2_X1 U21479 ( .A1(n18509), .A2(n18376), .ZN(n18369) );
  NAND2_X1 U21480 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18372), .ZN(n18365) );
  INV_X1 U21481 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21692) );
  NAND2_X1 U21482 ( .A1(n18408), .A2(n18361), .ZN(n18364) );
  AOI22_X1 U21483 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18378), .B1(n18389), .B2(
        n18362), .ZN(n18363) );
  OAI221_X1 U21484 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18365), .C1(n21692), 
        .C2(n18364), .A(n18363), .ZN(P3_U2721) );
  INV_X1 U21485 ( .A(n18365), .ZN(n18368) );
  AOI21_X1 U21486 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18408), .A(n18372), .ZN(
        n18367) );
  OAI222_X1 U21487 ( .A1(n18413), .A2(n18516), .B1(n18368), .B2(n18367), .C1(
        n18410), .C2(n18366), .ZN(P3_U2722) );
  INV_X1 U21488 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18511) );
  AOI21_X1 U21489 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18408), .A(n18369), .ZN(
        n18371) );
  OAI222_X1 U21490 ( .A1(n18413), .A2(n18511), .B1(n18372), .B2(n18371), .C1(
        n18410), .C2(n18370), .ZN(P3_U2723) );
  NAND2_X1 U21491 ( .A1(n18408), .A2(n18376), .ZN(n18381) );
  INV_X1 U21492 ( .A(n18373), .ZN(n18374) );
  AOI22_X1 U21493 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18378), .B1(n18389), .B2(
        n18374), .ZN(n18375) );
  OAI221_X1 U21494 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18376), .C1(n18509), 
        .C2(n18381), .A(n18375), .ZN(P3_U2724) );
  INV_X1 U21495 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18451) );
  AOI22_X1 U21496 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18378), .B1(n18389), .B2(
        n18377), .ZN(n18379) );
  OAI221_X1 U21497 ( .B1(n18381), .B2(n18451), .C1(n18381), .C2(n18380), .A(
        n18379), .ZN(P3_U2725) );
  INV_X1 U21498 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18505) );
  AND2_X1 U21499 ( .A1(n18383), .A2(n18382), .ZN(n18396) );
  AOI22_X1 U21500 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18408), .B1(
        P3_EAX_REG_8__SCAN_IN), .B2(n18396), .ZN(n18385) );
  OAI222_X1 U21501 ( .A1(n18413), .A2(n18505), .B1(n18386), .B2(n18385), .C1(
        n18410), .C2(n18384), .ZN(P3_U2726) );
  INV_X1 U21502 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18503) );
  INV_X1 U21503 ( .A(n18387), .ZN(n18388) );
  INV_X1 U21504 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U21505 ( .A1(n18389), .A2(n18388), .B1(n18396), .B2(n18454), .ZN(
        n18392) );
  NAND3_X1 U21506 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18408), .A3(n18390), .ZN(
        n18391) );
  OAI211_X1 U21507 ( .C1(n18413), .C2(n18503), .A(n18392), .B(n18391), .ZN(
        P3_U2727) );
  INV_X1 U21508 ( .A(n18407), .ZN(n18400) );
  NOR2_X1 U21509 ( .A1(n18393), .A2(n18400), .ZN(n18403) );
  AND2_X1 U21510 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18403), .ZN(n18399) );
  AOI21_X1 U21511 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18408), .A(n18399), .ZN(
        n18395) );
  OAI222_X1 U21512 ( .A1(n19133), .A2(n18413), .B1(n18396), .B2(n18395), .C1(
        n18410), .C2(n18394), .ZN(P3_U2728) );
  AOI21_X1 U21513 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18408), .A(n18403), .ZN(
        n18398) );
  OAI222_X1 U21514 ( .A1(n19128), .A2(n18413), .B1(n18399), .B2(n18398), .C1(
        n18410), .C2(n18397), .ZN(P3_U2729) );
  INV_X1 U21515 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18465) );
  NOR2_X1 U21516 ( .A1(n18465), .A2(n18400), .ZN(n18412) );
  AND2_X1 U21517 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18412), .ZN(n18406) );
  AOI21_X1 U21518 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18408), .A(n18406), .ZN(
        n18402) );
  OAI222_X1 U21519 ( .A1(n19124), .A2(n18413), .B1(n18403), .B2(n18402), .C1(
        n18410), .C2(n18401), .ZN(P3_U2730) );
  INV_X1 U21520 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19118) );
  AOI21_X1 U21521 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18408), .A(n18412), .ZN(
        n18405) );
  OAI222_X1 U21522 ( .A1(n19118), .A2(n18413), .B1(n18406), .B2(n18405), .C1(
        n18410), .C2(n18404), .ZN(P3_U2731) );
  INV_X1 U21523 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19113) );
  AOI21_X1 U21524 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18408), .A(n18407), .ZN(
        n18411) );
  OAI222_X1 U21525 ( .A1(n19113), .A2(n18413), .B1(n18412), .B2(n18411), .C1(
        n18410), .C2(n18409), .ZN(P3_U2732) );
  NOR2_X4 U21526 ( .A1(n18469), .A2(n18442), .ZN(n18457) );
  AND2_X1 U21527 ( .A1(n18457), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21528 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18492) );
  AOI22_X1 U21529 ( .A1(n18469), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18415) );
  OAI21_X1 U21530 ( .B1(n18492), .B2(n18440), .A(n18415), .ZN(P3_U2737) );
  INV_X1 U21531 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18417) );
  AOI22_X1 U21532 ( .A1(n18469), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18416) );
  OAI21_X1 U21533 ( .B1(n18417), .B2(n18440), .A(n18416), .ZN(P3_U2738) );
  AOI22_X1 U21534 ( .A1(n18469), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18418) );
  OAI21_X1 U21535 ( .B1(n18419), .B2(n18440), .A(n18418), .ZN(P3_U2739) );
  INV_X1 U21536 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U21537 ( .A1(n18469), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18420) );
  OAI21_X1 U21538 ( .B1(n18488), .B2(n18440), .A(n18420), .ZN(P3_U2740) );
  AOI22_X1 U21539 ( .A1(n18469), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18421) );
  OAI21_X1 U21540 ( .B1(n18422), .B2(n18440), .A(n18421), .ZN(P3_U2741) );
  AOI22_X1 U21541 ( .A1(n18469), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18423) );
  OAI21_X1 U21542 ( .B1(n10358), .B2(n18440), .A(n18423), .ZN(P3_U2742) );
  INV_X1 U21543 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U21544 ( .A1(n18469), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18424) );
  OAI21_X1 U21545 ( .B1(n18425), .B2(n18440), .A(n18424), .ZN(P3_U2743) );
  INV_X1 U21546 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18427) );
  INV_X2 U21547 ( .A(n19676), .ZN(n18469) );
  AOI22_X1 U21548 ( .A1(n18469), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18426) );
  OAI21_X1 U21549 ( .B1(n18427), .B2(n18440), .A(n18426), .ZN(P3_U2744) );
  AOI22_X1 U21550 ( .A1(n18469), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18428) );
  OAI21_X1 U21551 ( .B1(n18429), .B2(n18440), .A(n18428), .ZN(P3_U2745) );
  AOI22_X1 U21552 ( .A1(n18469), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18430) );
  OAI21_X1 U21553 ( .B1(n18431), .B2(n18440), .A(n18430), .ZN(P3_U2746) );
  INV_X1 U21554 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18433) );
  AOI22_X1 U21555 ( .A1(n18469), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18432) );
  OAI21_X1 U21556 ( .B1(n18433), .B2(n18440), .A(n18432), .ZN(P3_U2747) );
  INV_X1 U21557 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18435) );
  AOI22_X1 U21558 ( .A1(n18469), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18434) );
  OAI21_X1 U21559 ( .B1(n18435), .B2(n18440), .A(n18434), .ZN(P3_U2748) );
  AOI22_X1 U21560 ( .A1(n18469), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18436) );
  OAI21_X1 U21561 ( .B1(n18437), .B2(n18440), .A(n18436), .ZN(P3_U2749) );
  AOI22_X1 U21562 ( .A1(n18469), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18438) );
  OAI21_X1 U21563 ( .B1(n18477), .B2(n18440), .A(n18438), .ZN(P3_U2750) );
  INV_X1 U21564 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18441) );
  AOI22_X1 U21565 ( .A1(n18469), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18439) );
  OAI21_X1 U21566 ( .B1(n18441), .B2(n18440), .A(n18439), .ZN(P3_U2751) );
  AOI22_X1 U21567 ( .A1(n18469), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18443) );
  OAI21_X1 U21568 ( .B1(n18522), .B2(n18471), .A(n18443), .ZN(P3_U2752) );
  AOI22_X1 U21569 ( .A1(n18469), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18444) );
  OAI21_X1 U21570 ( .B1(n21692), .B2(n18471), .A(n18444), .ZN(P3_U2753) );
  INV_X1 U21571 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18446) );
  AOI22_X1 U21572 ( .A1(n18469), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18445) );
  OAI21_X1 U21573 ( .B1(n18446), .B2(n18471), .A(n18445), .ZN(P3_U2754) );
  INV_X1 U21574 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18448) );
  AOI22_X1 U21575 ( .A1(n18469), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18447) );
  OAI21_X1 U21576 ( .B1(n18448), .B2(n18471), .A(n18447), .ZN(P3_U2755) );
  AOI22_X1 U21577 ( .A1(n18469), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18449) );
  OAI21_X1 U21578 ( .B1(n18509), .B2(n18471), .A(n18449), .ZN(P3_U2756) );
  AOI22_X1 U21579 ( .A1(n18469), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18450) );
  OAI21_X1 U21580 ( .B1(n18451), .B2(n18471), .A(n18450), .ZN(P3_U2757) );
  INV_X1 U21581 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21619) );
  AOI22_X1 U21582 ( .A1(n18469), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18452) );
  OAI21_X1 U21583 ( .B1(n21619), .B2(n18471), .A(n18452), .ZN(P3_U2758) );
  AOI22_X1 U21584 ( .A1(n18469), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18453) );
  OAI21_X1 U21585 ( .B1(n18454), .B2(n18471), .A(n18453), .ZN(P3_U2759) );
  AOI22_X1 U21586 ( .A1(n18469), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18455) );
  OAI21_X1 U21587 ( .B1(n18456), .B2(n18471), .A(n18455), .ZN(P3_U2760) );
  AOI22_X1 U21588 ( .A1(n18469), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18458) );
  OAI21_X1 U21589 ( .B1(n18459), .B2(n18471), .A(n18458), .ZN(P3_U2761) );
  INV_X1 U21590 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18461) );
  AOI22_X1 U21591 ( .A1(n18469), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18460) );
  OAI21_X1 U21592 ( .B1(n18461), .B2(n18471), .A(n18460), .ZN(P3_U2762) );
  INV_X1 U21593 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18463) );
  AOI22_X1 U21594 ( .A1(n18469), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18462) );
  OAI21_X1 U21595 ( .B1(n18463), .B2(n18471), .A(n18462), .ZN(P3_U2763) );
  AOI22_X1 U21596 ( .A1(n18469), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18464) );
  OAI21_X1 U21597 ( .B1(n18465), .B2(n18471), .A(n18464), .ZN(P3_U2764) );
  INV_X1 U21598 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18467) );
  AOI22_X1 U21599 ( .A1(n18469), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18466) );
  OAI21_X1 U21600 ( .B1(n18467), .B2(n18471), .A(n18466), .ZN(P3_U2765) );
  AOI22_X1 U21601 ( .A1(n18469), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18468) );
  OAI21_X1 U21602 ( .B1(n18495), .B2(n18471), .A(n18468), .ZN(P3_U2766) );
  AOI22_X1 U21603 ( .A1(n18469), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18457), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18470) );
  OAI21_X1 U21604 ( .B1(n18472), .B2(n18471), .A(n18470), .ZN(P3_U2767) );
  AOI22_X1 U21605 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18518), .ZN(n18475) );
  OAI21_X1 U21606 ( .B1(n19096), .B2(n18515), .A(n18475), .ZN(P3_U2768) );
  AOI22_X1 U21607 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18519), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18518), .ZN(n18476) );
  OAI21_X1 U21608 ( .B1(n18477), .B2(n18521), .A(n18476), .ZN(P3_U2769) );
  AOI22_X1 U21609 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18518), .ZN(n18478) );
  OAI21_X1 U21610 ( .B1(n19107), .B2(n18515), .A(n18478), .ZN(P3_U2770) );
  AOI22_X1 U21611 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18518), .ZN(n18479) );
  OAI21_X1 U21612 ( .B1(n19113), .B2(n18515), .A(n18479), .ZN(P3_U2771) );
  AOI22_X1 U21613 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18518), .ZN(n18480) );
  OAI21_X1 U21614 ( .B1(n19118), .B2(n18515), .A(n18480), .ZN(P3_U2772) );
  AOI22_X1 U21615 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18518), .ZN(n18481) );
  OAI21_X1 U21616 ( .B1(n19124), .B2(n18515), .A(n18481), .ZN(P3_U2773) );
  AOI22_X1 U21617 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18518), .ZN(n18482) );
  OAI21_X1 U21618 ( .B1(n19128), .B2(n18515), .A(n18482), .ZN(P3_U2774) );
  AOI22_X1 U21619 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18518), .ZN(n18483) );
  OAI21_X1 U21620 ( .B1(n19133), .B2(n18515), .A(n18483), .ZN(P3_U2775) );
  AOI22_X1 U21621 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18518), .ZN(n18484) );
  OAI21_X1 U21622 ( .B1(n18503), .B2(n18515), .A(n18484), .ZN(P3_U2776) );
  AOI22_X1 U21623 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18518), .ZN(n18485) );
  OAI21_X1 U21624 ( .B1(n18505), .B2(n18515), .A(n18485), .ZN(P3_U2777) );
  INV_X1 U21625 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18507) );
  AOI22_X1 U21626 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18518), .ZN(n18486) );
  OAI21_X1 U21627 ( .B1(n18507), .B2(n18515), .A(n18486), .ZN(P3_U2778) );
  AOI22_X1 U21628 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18519), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18518), .ZN(n18487) );
  OAI21_X1 U21629 ( .B1(n18488), .B2(n18521), .A(n18487), .ZN(P3_U2779) );
  AOI22_X1 U21630 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18518), .ZN(n18489) );
  OAI21_X1 U21631 ( .B1(n18511), .B2(n18515), .A(n18489), .ZN(P3_U2780) );
  AOI22_X1 U21632 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18513), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18518), .ZN(n18490) );
  OAI21_X1 U21633 ( .B1(n18516), .B2(n18515), .A(n18490), .ZN(P3_U2781) );
  AOI22_X1 U21634 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18519), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18518), .ZN(n18491) );
  OAI21_X1 U21635 ( .B1(n18492), .B2(n18521), .A(n18491), .ZN(P3_U2782) );
  AOI22_X1 U21636 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18518), .ZN(n18493) );
  OAI21_X1 U21637 ( .B1(n19096), .B2(n18515), .A(n18493), .ZN(P3_U2783) );
  AOI22_X1 U21638 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18519), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18518), .ZN(n18494) );
  OAI21_X1 U21639 ( .B1(n18495), .B2(n18521), .A(n18494), .ZN(P3_U2784) );
  AOI22_X1 U21640 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18518), .ZN(n18496) );
  OAI21_X1 U21641 ( .B1(n19107), .B2(n18515), .A(n18496), .ZN(P3_U2785) );
  AOI22_X1 U21642 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18512), .ZN(n18497) );
  OAI21_X1 U21643 ( .B1(n19113), .B2(n18515), .A(n18497), .ZN(P3_U2786) );
  AOI22_X1 U21644 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18512), .ZN(n18498) );
  OAI21_X1 U21645 ( .B1(n19118), .B2(n18515), .A(n18498), .ZN(P3_U2787) );
  AOI22_X1 U21646 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18512), .ZN(n18499) );
  OAI21_X1 U21647 ( .B1(n19124), .B2(n18515), .A(n18499), .ZN(P3_U2788) );
  AOI22_X1 U21648 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18512), .ZN(n18500) );
  OAI21_X1 U21649 ( .B1(n19128), .B2(n18515), .A(n18500), .ZN(P3_U2789) );
  AOI22_X1 U21650 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18512), .ZN(n18501) );
  OAI21_X1 U21651 ( .B1(n19133), .B2(n18515), .A(n18501), .ZN(P3_U2790) );
  AOI22_X1 U21652 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18512), .ZN(n18502) );
  OAI21_X1 U21653 ( .B1(n18503), .B2(n18515), .A(n18502), .ZN(P3_U2791) );
  AOI22_X1 U21654 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18512), .ZN(n18504) );
  OAI21_X1 U21655 ( .B1(n18505), .B2(n18515), .A(n18504), .ZN(P3_U2792) );
  AOI22_X1 U21656 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18512), .ZN(n18506) );
  OAI21_X1 U21657 ( .B1(n18507), .B2(n18515), .A(n18506), .ZN(P3_U2793) );
  AOI22_X1 U21658 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18519), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18518), .ZN(n18508) );
  OAI21_X1 U21659 ( .B1(n18509), .B2(n18521), .A(n18508), .ZN(P3_U2794) );
  AOI22_X1 U21660 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18512), .ZN(n18510) );
  OAI21_X1 U21661 ( .B1(n18511), .B2(n18515), .A(n18510), .ZN(P3_U2795) );
  AOI22_X1 U21662 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18513), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18512), .ZN(n18514) );
  OAI21_X1 U21663 ( .B1(n18516), .B2(n18515), .A(n18514), .ZN(P3_U2796) );
  AOI22_X1 U21664 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18519), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18518), .ZN(n18517) );
  OAI21_X1 U21665 ( .B1(n21692), .B2(n18521), .A(n18517), .ZN(P3_U2797) );
  AOI22_X1 U21666 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18519), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18518), .ZN(n18520) );
  OAI21_X1 U21667 ( .B1(n18522), .B2(n18521), .A(n18520), .ZN(P3_U2798) );
  AOI21_X1 U21668 ( .B1(n18523), .B2(n17078), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18531) );
  AOI22_X1 U21669 ( .A1(n13950), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18524), 
        .B2(n18813), .ZN(n18530) );
  OAI21_X1 U21670 ( .B1(n18526), .B2(n18818), .A(n18525), .ZN(n18821) );
  NAND3_X1 U21671 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18827), .A3(
        n18818), .ZN(n18824) );
  INV_X1 U21672 ( .A(n18824), .ZN(n18528) );
  AOI222_X1 U21673 ( .A1(n18821), .A2(n18714), .B1(n18528), .B2(n18566), .C1(
        n18527), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18529) );
  OAI211_X1 U21674 ( .C1(n18532), .C2(n18531), .A(n18530), .B(n18529), .ZN(
        P3_U2804) );
  NOR2_X1 U21675 ( .A1(n18927), .A2(n18539), .ZN(n18839) );
  NAND2_X1 U21676 ( .A1(n18839), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18533) );
  XOR2_X1 U21677 ( .A(n18533), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18831) );
  AND2_X1 U21678 ( .A1(n10577), .A2(n17078), .ZN(n18561) );
  AOI211_X1 U21679 ( .C1(n18704), .C2(n18534), .A(n18776), .B(n18561), .ZN(
        n18563) );
  OAI21_X1 U21680 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18598), .A(
        n18563), .ZN(n18549) );
  NOR2_X1 U21681 ( .A1(n18649), .A2(n10577), .ZN(n18551) );
  OAI211_X1 U21682 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18551), .B(n18535), .ZN(n18536) );
  NAND2_X1 U21683 ( .A1(n19022), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18835) );
  OAI211_X1 U21684 ( .C1(n18706), .C2(n18537), .A(n18536), .B(n18835), .ZN(
        n18538) );
  AOI21_X1 U21685 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18549), .A(
        n18538), .ZN(n18545) );
  NOR2_X1 U21686 ( .A1(n18645), .A2(n18539), .ZN(n18843) );
  NAND2_X1 U21687 ( .A1(n18843), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18540) );
  XOR2_X1 U21688 ( .A(n18540), .B(n14436), .Z(n18833) );
  OAI21_X1 U21689 ( .B1(n18542), .B2(n18663), .A(n18541), .ZN(n18543) );
  XNOR2_X1 U21690 ( .A(n18543), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18834) );
  AOI22_X1 U21691 ( .A1(n18698), .A2(n18833), .B1(n18714), .B2(n18834), .ZN(
        n18544) );
  OAI211_X1 U21692 ( .C1(n18745), .C2(n18831), .A(n18545), .B(n18544), .ZN(
        P3_U2805) );
  NAND2_X1 U21693 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14434), .ZN(
        n18851) );
  AOI22_X1 U21694 ( .A1(n13950), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18730), 
        .B2(n18546), .ZN(n18547) );
  INV_X1 U21695 ( .A(n18547), .ZN(n18548) );
  AOI221_X1 U21696 ( .B1(n18551), .B2(n18550), .C1(n18549), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18548), .ZN(n18554) );
  OAI22_X1 U21697 ( .A1(n18839), .A2(n18745), .B1(n18843), .B2(n18696), .ZN(
        n18565) );
  XNOR2_X1 U21698 ( .A(n18552), .B(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18838) );
  AOI22_X1 U21699 ( .A1(n18565), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n18714), .B2(n18838), .ZN(n18553) );
  OAI211_X1 U21700 ( .C1(n18555), .C2(n18851), .A(n18554), .B(n18553), .ZN(
        P3_U2806) );
  NAND2_X1 U21701 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18557) );
  OAI211_X1 U21702 ( .C1(n18558), .C2(n18569), .A(n18556), .B(n18557), .ZN(
        n18559) );
  XNOR2_X1 U21703 ( .A(n18559), .B(n18844), .ZN(n18856) );
  AOI22_X1 U21704 ( .A1(n9725), .A2(n18561), .B1(n18560), .B2(n18813), .ZN(
        n18562) );
  NAND2_X1 U21705 ( .A1(n19022), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18855) );
  OAI211_X1 U21706 ( .C1(n18563), .C2(n10299), .A(n18562), .B(n18855), .ZN(
        n18564) );
  AOI221_X1 U21707 ( .B1(n18566), .B2(n18844), .C1(n18565), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18564), .ZN(n18567) );
  OAI21_X1 U21708 ( .B1(n18732), .B2(n18856), .A(n18567), .ZN(P3_U2807) );
  NOR2_X1 U21709 ( .A1(n9659), .A2(n18869), .ZN(n18568) );
  OAI21_X1 U21710 ( .B1(n18569), .B2(n18568), .A(n18556), .ZN(n18570) );
  XNOR2_X1 U21711 ( .A(n18570), .B(n18872), .ZN(n18878) );
  AOI22_X1 U21712 ( .A1(n18704), .A2(n18571), .B1(n18790), .B2(n18574), .ZN(
        n18572) );
  NAND2_X1 U21713 ( .A1(n18572), .A2(n18807), .ZN(n18596) );
  AOI21_X1 U21714 ( .B1(n18573), .B2(n10298), .A(n18596), .ZN(n18582) );
  NAND2_X1 U21715 ( .A1(n19022), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18876) );
  NOR2_X1 U21716 ( .A1(n18574), .A2(n18649), .ZN(n18581) );
  OAI211_X1 U21717 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18581), .B(n18575), .ZN(n18576) );
  OAI211_X1 U21718 ( .C1(n18582), .C2(n18577), .A(n18876), .B(n18576), .ZN(
        n18579) );
  INV_X1 U21719 ( .A(n18637), .ZN(n18657) );
  NOR2_X1 U21720 ( .A1(n18628), .A2(n18862), .ZN(n18885) );
  NAND3_X1 U21721 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18866), .A3(
        n18885), .ZN(n18863) );
  NOR2_X1 U21722 ( .A1(n18657), .A2(n18863), .ZN(n18578) );
  INV_X1 U21723 ( .A(n18656), .ZN(n18618) );
  AOI21_X1 U21724 ( .B1(n18594), .B2(n18863), .A(n18618), .ZN(n18587) );
  INV_X1 U21725 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18887) );
  NAND2_X1 U21726 ( .A1(n18866), .A2(n18887), .ZN(n18893) );
  NAND2_X1 U21727 ( .A1(n18637), .A2(n18885), .ZN(n18617) );
  INV_X1 U21728 ( .A(n18581), .ZN(n18584) );
  INV_X1 U21729 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18583) );
  NAND2_X1 U21730 ( .A1(n19022), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18891) );
  OAI221_X1 U21731 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18584), .C1(
        n18583), .C2(n18582), .A(n18891), .ZN(n18589) );
  OR2_X1 U21732 ( .A1(n18663), .A2(n18862), .ZN(n18624) );
  OAI22_X1 U21733 ( .A1(n18626), .A2(n18585), .B1(n18882), .B2(n18603), .ZN(
        n18586) );
  XNOR2_X1 U21734 ( .A(n18586), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18880) );
  OAI22_X1 U21735 ( .A1(n18587), .A2(n18887), .B1(n18880), .B2(n18732), .ZN(
        n18588) );
  AOI211_X1 U21736 ( .C1(n18730), .C2(n18590), .A(n18589), .B(n18588), .ZN(
        n18591) );
  OAI21_X1 U21737 ( .B1(n18893), .B2(n18617), .A(n18591), .ZN(P3_U2809) );
  INV_X1 U21738 ( .A(n18625), .ZN(n18592) );
  NAND2_X1 U21739 ( .A1(n18603), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18605) );
  OAI211_X1 U21740 ( .C1(n18592), .C2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n18556), .B(n18605), .ZN(n18593) );
  XNOR2_X1 U21741 ( .A(n18593), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18900) );
  NAND2_X1 U21742 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18885), .ZN(
        n18858) );
  AOI21_X1 U21743 ( .B1(n18594), .B2(n18858), .A(n18618), .ZN(n18616) );
  NAND2_X1 U21744 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18864), .ZN(
        n18904) );
  OAI22_X1 U21745 ( .A1(n18616), .A2(n18864), .B1(n18617), .B2(n18904), .ZN(
        n18595) );
  AOI21_X1 U21746 ( .B1(n18714), .B2(n18900), .A(n18595), .ZN(n18602) );
  NAND2_X1 U21747 ( .A1(n19022), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18902) );
  OAI221_X1 U21748 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18597), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n17078), .A(n18596), .ZN(
        n18601) );
  OAI21_X1 U21749 ( .B1(n18730), .B2(n18573), .A(n18599), .ZN(n18600) );
  NAND4_X1 U21750 ( .A1(n18602), .A2(n18902), .A3(n18601), .A4(n18600), .ZN(
        P3_U2810) );
  INV_X1 U21751 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18908) );
  NOR2_X1 U21752 ( .A1(n18626), .A2(n18625), .ZN(n18606) );
  INV_X1 U21753 ( .A(n18603), .ZN(n18604) );
  NOR2_X1 U21754 ( .A1(n18606), .A2(n18604), .ZN(n18607) );
  OAI22_X1 U21755 ( .A1(n18607), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n18606), .B2(n18605), .ZN(n18905) );
  AOI21_X1 U21756 ( .B1(n18790), .B2(n18609), .A(n18776), .ZN(n18640) );
  OAI21_X1 U21757 ( .B1(n18608), .B2(n19570), .A(n18640), .ZN(n18621) );
  AOI22_X1 U21758 ( .A1(n13950), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18621), .ZN(n18612) );
  NOR2_X1 U21759 ( .A1(n18649), .A2(n18609), .ZN(n18623) );
  OAI211_X1 U21760 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18623), .B(n18610), .ZN(n18611) );
  OAI211_X1 U21761 ( .C1(n18706), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        n18614) );
  AOI21_X1 U21762 ( .B1(n18714), .B2(n18905), .A(n18614), .ZN(n18615) );
  OAI221_X1 U21763 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18617), 
        .C1(n18908), .C2(n18616), .A(n18615), .ZN(P3_U2811) );
  AOI21_X1 U21764 ( .B1(n18637), .B2(n18628), .A(n18618), .ZN(n18634) );
  OAI22_X1 U21765 ( .A1(n19075), .A2(n19620), .B1(n18706), .B2(n18619), .ZN(
        n18620) );
  AOI221_X1 U21766 ( .B1(n18623), .B2(n18622), .C1(n18621), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18620), .ZN(n18630) );
  NAND2_X1 U21767 ( .A1(n18625), .A2(n18624), .ZN(n18627) );
  XOR2_X1 U21768 ( .A(n18627), .B(n18626), .Z(n18912) );
  NOR2_X1 U21769 ( .A1(n18628), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18911) );
  AOI22_X1 U21770 ( .A1(n18912), .A2(n18714), .B1(n18637), .B2(n18911), .ZN(
        n18629) );
  OAI211_X1 U21771 ( .C1(n18634), .C2(n18862), .A(n18630), .B(n18629), .ZN(
        P3_U2812) );
  AOI21_X1 U21772 ( .B1(n17078), .B2(n18631), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18641) );
  AOI22_X1 U21773 ( .A1(n13950), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18632), 
        .B2(n18813), .ZN(n18639) );
  OAI22_X1 U21774 ( .A1(n18634), .A2(n14430), .B1(n18732), .B2(n18633), .ZN(
        n18635) );
  AOI21_X1 U21775 ( .B1(n18637), .B2(n18636), .A(n18635), .ZN(n18638) );
  OAI211_X1 U21776 ( .C1(n18641), .C2(n18640), .A(n18639), .B(n18638), .ZN(
        P3_U2813) );
  INV_X1 U21777 ( .A(n18642), .ZN(n18643) );
  AOI21_X1 U21778 ( .B1(n18645), .B2(n18644), .A(n18643), .ZN(n18646) );
  XOR2_X1 U21779 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18646), .Z(
        n18923) );
  AOI21_X1 U21780 ( .B1(n18790), .B2(n18648), .A(n18776), .ZN(n18685) );
  OAI21_X1 U21781 ( .B1(n18647), .B2(n19570), .A(n18685), .ZN(n18660) );
  AOI22_X1 U21782 ( .A1(n19022), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18660), .ZN(n18652) );
  NOR2_X1 U21783 ( .A1(n18649), .A2(n18648), .ZN(n18662) );
  OAI211_X1 U21784 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18662), .B(n18650), .ZN(n18651) );
  OAI211_X1 U21785 ( .C1(n18706), .C2(n18653), .A(n18652), .B(n18651), .ZN(
        n18654) );
  AOI21_X1 U21786 ( .B1(n18714), .B2(n18923), .A(n18654), .ZN(n18655) );
  OAI221_X1 U21787 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18657), 
        .C1(n14427), .C2(n18656), .A(n18655), .ZN(P3_U2814) );
  INV_X1 U21788 ( .A(n18944), .ZN(n18710) );
  OR3_X1 U21789 ( .A1(n18985), .A2(n18710), .A3(n18668), .ZN(n18691) );
  NAND2_X1 U21790 ( .A1(n18675), .A2(n18691), .ZN(n18933) );
  INV_X1 U21791 ( .A(n18933), .ZN(n18680) );
  NAND2_X1 U21792 ( .A1(n18812), .A2(n18927), .ZN(n18679) );
  INV_X1 U21793 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18661) );
  OAI22_X1 U21794 ( .A1(n19075), .A2(n19614), .B1(n18706), .B2(n18658), .ZN(
        n18659) );
  AOI221_X1 U21795 ( .B1(n18662), .B2(n18661), .C1(n18660), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18659), .ZN(n18678) );
  NOR2_X1 U21796 ( .A1(n18663), .A2(n18969), .ZN(n18711) );
  NOR2_X1 U21797 ( .A1(n18664), .A2(n18717), .ZN(n18712) );
  INV_X1 U21798 ( .A(n18712), .ZN(n18669) );
  INV_X1 U21799 ( .A(n18665), .ZN(n18666) );
  NOR2_X1 U21800 ( .A1(n18667), .A2(n18666), .ZN(n18718) );
  INV_X1 U21801 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18948) );
  NAND2_X1 U21802 ( .A1(n18718), .A2(n18948), .ZN(n18688) );
  OAI21_X1 U21803 ( .B1(n18669), .B2(n18668), .A(n18688), .ZN(n18670) );
  OAI21_X1 U21804 ( .B1(n18671), .B2(n18711), .A(n18670), .ZN(n18672) );
  XOR2_X1 U21805 ( .A(n18675), .B(n18672), .Z(n18936) );
  NOR2_X1 U21806 ( .A1(n18929), .A2(n18696), .ZN(n18676) );
  NAND2_X1 U21807 ( .A1(n18988), .A2(n18944), .ZN(n18960) );
  INV_X1 U21808 ( .A(n18960), .ZN(n18674) );
  NAND2_X1 U21809 ( .A1(n18674), .A2(n18673), .ZN(n18681) );
  NAND2_X1 U21810 ( .A1(n18681), .A2(n18675), .ZN(n18931) );
  AOI22_X1 U21811 ( .A1(n18714), .A2(n18936), .B1(n18676), .B2(n18931), .ZN(
        n18677) );
  OAI211_X1 U21812 ( .C1(n18680), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        P3_U2815) );
  NOR2_X1 U21813 ( .A1(n18960), .A2(n18948), .ZN(n18682) );
  OAI21_X1 U21814 ( .B1(n18682), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18681), .ZN(n18952) );
  AOI21_X1 U21815 ( .B1(n18700), .B2(n18683), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18684) );
  NAND2_X1 U21816 ( .A1(n19022), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U21817 ( .B1(n18685), .B2(n18684), .A(n18954), .ZN(n18693) );
  NOR2_X1 U21818 ( .A1(n18710), .A2(n18948), .ZN(n18940) );
  INV_X1 U21819 ( .A(n18940), .ZN(n18686) );
  OAI22_X1 U21820 ( .A1(n18688), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18687), .B2(n18686), .ZN(n18689) );
  INV_X1 U21821 ( .A(n18689), .ZN(n18690) );
  XOR2_X1 U21822 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18690), .Z(
        n18957) );
  OAI221_X1 U21823 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18940), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18697), .A(n18691), .ZN(
        n18949) );
  OAI22_X1 U21824 ( .A1(n18957), .A2(n18732), .B1(n18745), .B2(n18949), .ZN(
        n18692) );
  AOI211_X1 U21825 ( .C1(n18694), .C2(n18813), .A(n18693), .B(n18692), .ZN(
        n18695) );
  OAI21_X1 U21826 ( .B1(n18696), .B2(n18952), .A(n18695), .ZN(P3_U2816) );
  NAND2_X1 U21827 ( .A1(n18944), .A2(n18697), .ZN(n18962) );
  AOI22_X1 U21828 ( .A1(n18698), .A2(n18960), .B1(n18812), .B2(n18962), .ZN(
        n18726) );
  NAND2_X1 U21829 ( .A1(n18701), .A2(n18699), .ZN(n18723) );
  AOI211_X1 U21830 ( .C1(n18722), .C2(n18707), .A(n18700), .B(n18723), .ZN(
        n18709) );
  OAI21_X1 U21831 ( .B1(n18701), .B2(n9899), .A(n18807), .ZN(n18702) );
  AOI21_X1 U21832 ( .B1(n18704), .B2(n18703), .A(n18702), .ZN(n18721) );
  OAI22_X1 U21833 ( .A1(n18721), .A2(n18707), .B1(n18706), .B2(n18705), .ZN(
        n18708) );
  AOI211_X1 U21834 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n19022), .A(n18709), 
        .B(n18708), .ZN(n18716) );
  NOR2_X1 U21835 ( .A1(n18710), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18958) );
  OAI22_X1 U21836 ( .A1(n18712), .A2(n18969), .B1(n18711), .B2(n18718), .ZN(
        n18713) );
  XNOR2_X1 U21837 ( .A(n18713), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18959) );
  AOI22_X1 U21838 ( .A1(n18724), .A2(n18958), .B1(n18714), .B2(n18959), .ZN(
        n18715) );
  OAI211_X1 U21839 ( .C1(n18726), .C2(n18948), .A(n18716), .B(n18715), .ZN(
        P3_U2817) );
  INV_X1 U21840 ( .A(n18717), .ZN(n18993) );
  AOI21_X1 U21841 ( .B1(n18719), .B2(n18993), .A(n18718), .ZN(n18720) );
  XNOR2_X1 U21842 ( .A(n18969), .B(n18720), .ZN(n18974) );
  NAND2_X1 U21843 ( .A1(n19022), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18976) );
  OAI221_X1 U21844 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18723), .C1(
        n18722), .C2(n18721), .A(n18976), .ZN(n18728) );
  NAND3_X1 U21845 ( .A1(n18724), .A2(n18993), .A3(n18969), .ZN(n18725) );
  OAI21_X1 U21846 ( .B1(n18726), .B2(n18969), .A(n18725), .ZN(n18727) );
  AOI211_X1 U21847 ( .C1(n18730), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        n18731) );
  OAI21_X1 U21848 ( .B1(n18974), .B2(n18732), .A(n18731), .ZN(P3_U2818) );
  NAND2_X1 U21849 ( .A1(n18734), .A2(n18733), .ZN(n18735) );
  XOR2_X1 U21850 ( .A(n18735), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19020) );
  NOR2_X1 U21851 ( .A1(n19075), .A2(n21686), .ZN(n19012) );
  AOI221_X1 U21852 ( .B1(n18738), .B2(n18737), .C1(n18736), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n19012), .ZN(n18744) );
  OAI21_X1 U21853 ( .B1(n18740), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18739), .ZN(n18741) );
  INV_X1 U21854 ( .A(n18741), .ZN(n19016) );
  AOI22_X1 U21855 ( .A1(n18813), .A2(n18742), .B1(n10202), .B2(n19016), .ZN(
        n18743) );
  OAI211_X1 U21856 ( .C1(n18745), .C2(n19020), .A(n18744), .B(n18743), .ZN(
        P3_U2823) );
  OAI21_X1 U21857 ( .B1(n18748), .B2(n18747), .A(n18746), .ZN(n18749) );
  INV_X1 U21858 ( .A(n18749), .ZN(n19024) );
  AOI22_X1 U21859 ( .A1(n10202), .A2(n19024), .B1(n18753), .B2(n18752), .ZN(
        n18757) );
  AOI21_X1 U21860 ( .B1(n18751), .B2(n19026), .A(n18750), .ZN(n19025) );
  OR2_X1 U21861 ( .A1(n18817), .A2(n18752), .ZN(n18764) );
  OAI22_X1 U21862 ( .A1(n18803), .A2(n18754), .B1(n18753), .B2(n18764), .ZN(
        n18755) );
  AOI21_X1 U21863 ( .B1(n18812), .B2(n19025), .A(n18755), .ZN(n18756) );
  OAI211_X1 U21864 ( .C1(n19075), .C2(n19597), .A(n18757), .B(n18756), .ZN(
        P3_U2824) );
  AOI21_X1 U21865 ( .B1(n17724), .B2(n18807), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18765) );
  AOI21_X1 U21866 ( .B1(n10202), .B2(n18759), .A(n18758), .ZN(n18763) );
  AOI22_X1 U21867 ( .A1(n18812), .A2(n18761), .B1(n18760), .B2(n18813), .ZN(
        n18762) );
  OAI211_X1 U21868 ( .C1(n18765), .C2(n18764), .A(n18763), .B(n18762), .ZN(
        P3_U2825) );
  INV_X1 U21869 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19594) );
  OAI21_X1 U21870 ( .B1(n18768), .B2(n18767), .A(n18766), .ZN(n18769) );
  INV_X1 U21871 ( .A(n18769), .ZN(n19031) );
  AOI22_X1 U21872 ( .A1(n10202), .A2(n19031), .B1(n17078), .B2(n18770), .ZN(
        n18780) );
  OAI21_X1 U21873 ( .B1(n18773), .B2(n18772), .A(n18771), .ZN(n18775) );
  XOR2_X1 U21874 ( .A(n18775), .B(n18774), .Z(n19036) );
  AOI21_X1 U21875 ( .B1(n18790), .B2(n17745), .A(n18776), .ZN(n18787) );
  OAI22_X1 U21876 ( .A1(n18803), .A2(n18777), .B1(n18787), .B2(n17756), .ZN(
        n18778) );
  AOI21_X1 U21877 ( .B1(n18812), .B2(n19036), .A(n18778), .ZN(n18779) );
  OAI211_X1 U21878 ( .C1(n19075), .C2(n19594), .A(n18780), .B(n18779), .ZN(
        P3_U2826) );
  AOI21_X1 U21879 ( .B1(n18783), .B2(n18782), .A(n18781), .ZN(n19041) );
  OR2_X1 U21880 ( .A1(n18784), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18785) );
  AND2_X1 U21881 ( .A1(n18786), .A2(n18785), .ZN(n19046) );
  AOI22_X1 U21882 ( .A1(n18812), .A2(n19041), .B1(n10202), .B2(n19046), .ZN(
        n18793) );
  INV_X1 U21883 ( .A(n18787), .ZN(n18789) );
  AOI22_X1 U21884 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n18789), .B1(
        n18788), .B2(n18813), .ZN(n18792) );
  NAND4_X1 U21885 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18790), .A3(
        n18807), .A4(n17745), .ZN(n18791) );
  NAND2_X1 U21886 ( .A1(n19022), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19049) );
  NAND4_X1 U21887 ( .A1(n18793), .A2(n18792), .A3(n18791), .A4(n19049), .ZN(
        P3_U2827) );
  AOI21_X1 U21888 ( .B1(n18796), .B2(n18795), .A(n18794), .ZN(n19051) );
  OAI21_X1 U21889 ( .B1(n18799), .B2(n18798), .A(n18797), .ZN(n19055) );
  AND2_X1 U21890 ( .A1(n19022), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19068) );
  INV_X1 U21891 ( .A(n19068), .ZN(n18800) );
  OAI21_X1 U21892 ( .B1(n18801), .B2(n19055), .A(n18800), .ZN(n18805) );
  NOR2_X1 U21893 ( .A1(n18803), .A2(n18802), .ZN(n18804) );
  AOI211_X1 U21894 ( .C1(n18812), .C2(n19051), .A(n18805), .B(n18804), .ZN(
        n18806) );
  OAI221_X1 U21895 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19136), .C1(
        n18808), .C2(n18807), .A(n18806), .ZN(P3_U2828) );
  AOI21_X1 U21896 ( .B1(n10202), .B2(n18810), .A(n18809), .ZN(n18815) );
  AOI22_X1 U21897 ( .A1(n18813), .A2(n18816), .B1(n18812), .B2(n18811), .ZN(
        n18814) );
  OAI211_X1 U21898 ( .C1(n18817), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        P3_U2829) );
  NOR3_X1 U21899 ( .A1(n18819), .A2(n13950), .A3(n18818), .ZN(n18820) );
  AOI21_X1 U21900 ( .B1(n19007), .B2(n18821), .A(n18820), .ZN(n18823) );
  NAND2_X1 U21901 ( .A1(n19022), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18822) );
  OAI211_X1 U21902 ( .C1(n18824), .C2(n18850), .A(n18823), .B(n18822), .ZN(
        P3_U2836) );
  NAND2_X1 U21903 ( .A1(n18827), .A2(n18846), .ZN(n18825) );
  OAI211_X1 U21904 ( .C1(n18840), .C2(n18825), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18920), .ZN(n18830) );
  NAND4_X1 U21905 ( .A1(n18828), .A2(n18827), .A3(n14436), .A4(n18826), .ZN(
        n18829) );
  OAI211_X1 U21906 ( .C1(n18831), .C2(n10205), .A(n18830), .B(n18829), .ZN(
        n18832) );
  AOI21_X1 U21907 ( .B1(n18961), .B2(n18833), .A(n18832), .ZN(n18837) );
  AOI22_X1 U21908 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19042), .B1(
        n19007), .B2(n18834), .ZN(n18836) );
  OAI211_X1 U21909 ( .C1(n18837), .C2(n19080), .A(n18836), .B(n18835), .ZN(
        P3_U2837) );
  AOI22_X1 U21910 ( .A1(n18838), .A2(n19007), .B1(n13950), .B2(
        P3_REIP_REG_24__SCAN_IN), .ZN(n18849) );
  INV_X1 U21911 ( .A(n18839), .ZN(n18841) );
  AOI211_X1 U21912 ( .C1(n19519), .C2(n18841), .A(n18840), .B(n19042), .ZN(
        n18842) );
  OAI21_X1 U21913 ( .B1(n18843), .B2(n18987), .A(n18842), .ZN(n18847) );
  NOR2_X1 U21914 ( .A1(n18844), .A2(n18847), .ZN(n18845) );
  AOI21_X1 U21915 ( .B1(n18846), .B2(n18845), .A(n19022), .ZN(n18852) );
  OAI211_X1 U21916 ( .C1(n18920), .C2(n18847), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18852), .ZN(n18848) );
  OAI211_X1 U21917 ( .C1(n18851), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        P3_U2838) );
  NOR4_X1 U21918 ( .A1(n19042), .A2(n18870), .A3(n18869), .A4(n18872), .ZN(
        n18853) );
  OAI21_X1 U21919 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18853), .A(
        n18852), .ZN(n18854) );
  OAI211_X1 U21920 ( .C1(n18856), .C2(n18956), .A(n18855), .B(n18854), .ZN(
        P3_U2839) );
  AND2_X1 U21921 ( .A1(n18971), .A2(n18857), .ZN(n18868) );
  INV_X1 U21922 ( .A(n18883), .ZN(n18859) );
  INV_X1 U21923 ( .A(n18858), .ZN(n18897) );
  AOI21_X1 U21924 ( .B1(n18859), .B2(n18897), .A(n18943), .ZN(n18860) );
  AOI211_X1 U21925 ( .C1(n9887), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        n18895) );
  AOI22_X1 U21926 ( .A1(n19081), .A2(n18864), .B1(n18863), .B2(n18989), .ZN(
        n18865) );
  NAND2_X1 U21927 ( .A1(n18895), .A2(n18865), .ZN(n18881) );
  OAI22_X1 U21928 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18992), .B1(
        n18866), .B2(n19061), .ZN(n18867) );
  NOR4_X1 U21929 ( .A1(n18868), .A2(n18872), .A3(n18881), .A4(n18867), .ZN(
        n18874) );
  OR2_X1 U21930 ( .A1(n18870), .A2(n18869), .ZN(n18871) );
  AOI22_X1 U21931 ( .A1(n18874), .A2(n18873), .B1(n18872), .B2(n18871), .ZN(
        n18875) );
  AOI22_X1 U21932 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19042), .B1(
        n19070), .B2(n18875), .ZN(n18877) );
  OAI211_X1 U21933 ( .C1(n18878), .C2(n18956), .A(n18877), .B(n18876), .ZN(
        P3_U2840) );
  NAND2_X1 U21934 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18879), .ZN(
        n18909) );
  INV_X1 U21935 ( .A(n18880), .ZN(n18890) );
  AOI21_X1 U21936 ( .B1(n18882), .B2(n18947), .A(n18881), .ZN(n18888) );
  NOR2_X1 U21937 ( .A1(n18884), .A2(n18883), .ZN(n18917) );
  AOI21_X1 U21938 ( .B1(n18885), .B2(n18917), .A(n18994), .ZN(n18886) );
  NOR2_X1 U21939 ( .A1(n18886), .A2(n18921), .ZN(n18894) );
  AOI211_X1 U21940 ( .C1(n18888), .C2(n18894), .A(n13950), .B(n18887), .ZN(
        n18889) );
  AOI21_X1 U21941 ( .B1(n19007), .B2(n18890), .A(n18889), .ZN(n18892) );
  OAI211_X1 U21942 ( .C1(n18893), .C2(n18909), .A(n18892), .B(n18891), .ZN(
        P3_U2841) );
  NAND3_X1 U21943 ( .A1(n18908), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18947), 
        .ZN(n18899) );
  OAI211_X1 U21944 ( .C1(n18897), .C2(n18896), .A(n18895), .B(n18894), .ZN(
        n18898) );
  NAND2_X1 U21945 ( .A1(n19075), .A2(n18898), .ZN(n18907) );
  NAND2_X1 U21946 ( .A1(n18899), .A2(n18907), .ZN(n18901) );
  AOI22_X1 U21947 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18901), .B1(
        n19007), .B2(n18900), .ZN(n18903) );
  OAI211_X1 U21948 ( .C1(n18904), .C2(n18909), .A(n18903), .B(n18902), .ZN(
        P3_U2842) );
  AOI22_X1 U21949 ( .A1(n13950), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n19007), 
        .B2(n18905), .ZN(n18906) );
  OAI221_X1 U21950 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18909), 
        .C1(n18908), .C2(n18907), .A(n18906), .ZN(P3_U2843) );
  AOI22_X1 U21951 ( .A1(n18912), .A2(n19007), .B1(n18911), .B2(n18922), .ZN(
        n18913) );
  OAI221_X1 U21952 ( .B1(n19022), .B2(n18914), .C1(n19075), .C2(n19620), .A(
        n18913), .ZN(P3_U2844) );
  OAI22_X1 U21953 ( .A1(n19061), .A2(n18915), .B1(n18943), .B2(n18981), .ZN(
        n18916) );
  INV_X1 U21954 ( .A(n18916), .ZN(n18982) );
  AOI21_X1 U21955 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18994), .A(
        n18917), .ZN(n18918) );
  INV_X1 U21956 ( .A(n18918), .ZN(n18919) );
  OAI211_X1 U21957 ( .C1(n18942), .C2(n18992), .A(n18982), .B(n18919), .ZN(
        n18934) );
  OAI221_X1 U21958 ( .B1(n18921), .B2(n18920), .C1(n18921), .C2(n18934), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18925) );
  AOI22_X1 U21959 ( .A1(n18923), .A2(n19007), .B1(n18922), .B2(n14427), .ZN(
        n18924) );
  OAI221_X1 U21960 ( .B1(n19022), .B2(n18925), .C1(n19075), .C2(n19616), .A(
        n18924), .ZN(P3_U2846) );
  AOI21_X1 U21961 ( .B1(n18942), .B2(n18941), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18926) );
  INV_X1 U21962 ( .A(n18926), .ZN(n18935) );
  INV_X1 U21963 ( .A(n18927), .ZN(n18928) );
  NOR2_X1 U21964 ( .A1(n18928), .A2(n10205), .ZN(n18932) );
  NOR2_X1 U21965 ( .A1(n18929), .A2(n18987), .ZN(n18930) );
  AOI222_X1 U21966 ( .A1(n18935), .A2(n18934), .B1(n18933), .B2(n18932), .C1(
        n18931), .C2(n18930), .ZN(n18939) );
  AOI22_X1 U21967 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19042), .B1(
        n19007), .B2(n18936), .ZN(n18938) );
  NAND2_X1 U21968 ( .A1(n19022), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18937) );
  OAI211_X1 U21969 ( .C1(n18939), .C2(n19080), .A(n18938), .B(n18937), .ZN(
        P3_U2847) );
  AOI21_X1 U21970 ( .B1(n18941), .B2(n18940), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18951) );
  AOI21_X1 U21971 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18943), .A(
        n18942), .ZN(n18946) );
  NAND3_X1 U21972 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18944), .A3(
        n18981), .ZN(n18972) );
  NAND2_X1 U21973 ( .A1(n18971), .A2(n18972), .ZN(n18964) );
  OAI211_X1 U21974 ( .C1(n18944), .C2(n19061), .A(n18982), .B(n18964), .ZN(
        n18945) );
  AOI211_X1 U21975 ( .C1(n18948), .C2(n18947), .A(n18946), .B(n18945), .ZN(
        n18950) );
  OAI222_X1 U21976 ( .A1(n18952), .A2(n18987), .B1(n18951), .B2(n18950), .C1(
        n10205), .C2(n18949), .ZN(n18953) );
  AOI22_X1 U21977 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19042), .B1(
        n19070), .B2(n18953), .ZN(n18955) );
  OAI211_X1 U21978 ( .C1(n18957), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        P3_U2848) );
  INV_X1 U21979 ( .A(n18958), .ZN(n18968) );
  AOI22_X1 U21980 ( .A1(n13950), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19007), 
        .B2(n18959), .ZN(n18967) );
  AOI22_X1 U21981 ( .A1(n19519), .A2(n18962), .B1(n18961), .B2(n18960), .ZN(
        n18963) );
  OAI211_X1 U21982 ( .C1(n18993), .C2(n18992), .A(n18982), .B(n18963), .ZN(
        n18970) );
  OAI211_X1 U21983 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18992), .A(
        n19070), .B(n18964), .ZN(n18965) );
  OAI211_X1 U21984 ( .C1(n18970), .C2(n18965), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19075), .ZN(n18966) );
  OAI211_X1 U21985 ( .C1(n18968), .C2(n19011), .A(n18967), .B(n18966), .ZN(
        P3_U2849) );
  AOI211_X1 U21986 ( .C1(n18972), .C2(n18971), .A(n18970), .B(n18969), .ZN(
        n18979) );
  OAI221_X1 U21987 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18993), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18973), .A(n19070), .ZN(
        n18978) );
  INV_X1 U21988 ( .A(n18974), .ZN(n18975) );
  AOI22_X1 U21989 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19042), .B1(
        n19007), .B2(n18975), .ZN(n18977) );
  OAI211_X1 U21990 ( .C1(n18979), .C2(n18978), .A(n18977), .B(n18976), .ZN(
        P3_U2850) );
  AOI22_X1 U21991 ( .A1(n13950), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19007), 
        .B2(n18980), .ZN(n18997) );
  AOI21_X1 U21992 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18981), .A(
        n18994), .ZN(n18984) );
  NAND2_X1 U21993 ( .A1(n18982), .A2(n19070), .ZN(n18983) );
  AOI211_X1 U21994 ( .C1(n19519), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        n18986) );
  OAI21_X1 U21995 ( .B1(n18988), .B2(n18987), .A(n18986), .ZN(n19005) );
  AOI21_X1 U21996 ( .B1(n18990), .B2(n18989), .A(n19005), .ZN(n18991) );
  OAI21_X1 U21997 ( .B1(n18994), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18991), .ZN(n19000) );
  OAI22_X1 U21998 ( .A1(n18994), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18993), .B2(n18992), .ZN(n18995) );
  OAI211_X1 U21999 ( .C1(n19000), .C2(n18995), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19075), .ZN(n18996) );
  OAI211_X1 U22000 ( .C1(n18998), .C2(n19011), .A(n18997), .B(n18996), .ZN(
        P3_U2851) );
  OAI221_X1 U22001 ( .B1(n19000), .B2(n19010), .C1(n19000), .C2(n18999), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19004) );
  NOR3_X1 U22002 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n19010), .A3(
        n19011), .ZN(n19001) );
  AOI21_X1 U22003 ( .B1(n19007), .B2(n19002), .A(n19001), .ZN(n19003) );
  OAI221_X1 U22004 ( .B1(n19022), .B2(n19004), .C1(n19075), .C2(n19604), .A(
        n19003), .ZN(P3_U2852) );
  NAND2_X1 U22005 ( .A1(n19075), .A2(n19005), .ZN(n19009) );
  AOI22_X1 U22006 ( .A1(n13950), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19007), 
        .B2(n19006), .ZN(n19008) );
  OAI221_X1 U22007 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19011), .C1(
        n19010), .C2(n19009), .A(n19008), .ZN(P3_U2853) );
  AOI21_X1 U22008 ( .B1(n19042), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19012), .ZN(n19019) );
  AOI221_X1 U22009 ( .B1(n19026), .B2(n19015), .C1(n19014), .C2(n19015), .A(
        n19013), .ZN(n19017) );
  AOI22_X1 U22010 ( .A1(n19017), .A2(n19070), .B1(n19074), .B2(n19016), .ZN(
        n19018) );
  OAI211_X1 U22011 ( .C1(n19021), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        P3_U2855) );
  AOI22_X1 U22012 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n19030) );
  AOI22_X1 U22013 ( .A1(n19079), .A2(n19025), .B1(n19074), .B2(n19024), .ZN(
        n19029) );
  NAND3_X1 U22014 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19027), .A3(
        n19026), .ZN(n19028) );
  NAND3_X1 U22015 ( .A1(n19030), .A2(n19029), .A3(n19028), .ZN(P3_U2856) );
  AOI22_X1 U22016 ( .A1(n19074), .A2(n19031), .B1(n13950), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n19039) );
  OAI21_X1 U22017 ( .B1(n19061), .B2(n19054), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19032) );
  AOI211_X1 U22018 ( .C1(n19034), .C2(n19033), .A(n19064), .B(n19032), .ZN(
        n19043) );
  OAI21_X1 U22019 ( .B1(n19043), .B2(n19035), .A(n19072), .ZN(n19037) );
  AOI22_X1 U22020 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19037), .B1(
        n19079), .B2(n19036), .ZN(n19038) );
  OAI211_X1 U22021 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n19040), .A(
        n19039), .B(n19038), .ZN(P3_U2858) );
  AOI22_X1 U22022 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19042), .B1(
        n19079), .B2(n19041), .ZN(n19050) );
  INV_X1 U22023 ( .A(n19043), .ZN(n19044) );
  OAI211_X1 U22024 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19045), .A(
        n19070), .B(n19044), .ZN(n19048) );
  NAND2_X1 U22025 ( .A1(n19074), .A2(n19046), .ZN(n19047) );
  NAND4_X1 U22026 ( .A1(n19050), .A2(n19049), .A3(n19048), .A4(n19047), .ZN(
        P3_U2859) );
  INV_X1 U22027 ( .A(n19051), .ZN(n19067) );
  NOR3_X1 U22028 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19053), .A3(
        n19052), .ZN(n19059) );
  NOR2_X1 U22029 ( .A1(n19061), .A2(n19054), .ZN(n19057) );
  NOR2_X1 U22030 ( .A1(n19514), .A2(n19055), .ZN(n19056) );
  OR2_X1 U22031 ( .A1(n19057), .A2(n19056), .ZN(n19058) );
  NOR2_X1 U22032 ( .A1(n19059), .A2(n19058), .ZN(n19066) );
  NAND2_X1 U22033 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19060) );
  OAI22_X1 U22034 ( .A1(n19062), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19061), .B2(n19060), .ZN(n19063) );
  OAI21_X1 U22035 ( .B1(n19064), .B2(n19063), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19065) );
  OAI211_X1 U22036 ( .C1(n19067), .C2(n10205), .A(n19066), .B(n19065), .ZN(
        n19069) );
  AOI21_X1 U22037 ( .B1(n19070), .B2(n19069), .A(n19068), .ZN(n19071) );
  OAI21_X1 U22038 ( .B1(n19073), .B2(n19072), .A(n19071), .ZN(P3_U2860) );
  INV_X1 U22039 ( .A(n19074), .ZN(n19076) );
  OAI22_X1 U22040 ( .A1(n19076), .A2(n19078), .B1(n19666), .B2(n19075), .ZN(
        n19077) );
  AOI21_X1 U22041 ( .B1(n19079), .B2(n19078), .A(n19077), .ZN(n19084) );
  OAI211_X1 U22042 ( .C1(n19081), .C2(n19080), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n19075), .ZN(n19082) );
  NAND3_X1 U22043 ( .A1(n19084), .A2(n19083), .A3(n19082), .ZN(P3_U2862) );
  INV_X1 U22044 ( .A(n19085), .ZN(n19086) );
  OAI211_X1 U22045 ( .C1(n19086), .C2(P3_FLUSH_REG_SCAN_IN), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n19558)
         );
  OAI21_X1 U22046 ( .B1(n19092), .B2(n19087), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19088) );
  OAI221_X1 U22047 ( .B1(n19092), .B2(n19558), .C1(n19092), .C2(n19270), .A(
        n19088), .ZN(P3_U2863) );
  NAND2_X1 U22048 ( .A1(n19541), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19227) );
  NAND2_X1 U22049 ( .A1(n19095), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19362) );
  NAND2_X1 U22050 ( .A1(n19435), .A2(n19364), .ZN(n19385) );
  AND2_X1 U22051 ( .A1(n19227), .A2(n19385), .ZN(n19090) );
  OAI22_X1 U22052 ( .A1(n19091), .A2(n19541), .B1(n19090), .B2(n19089), .ZN(
        P3_U2866) );
  AND2_X1 U22053 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19092), .ZN(
        P3_U2867) );
  NAND2_X1 U22054 ( .A1(n19095), .A2(n19541), .ZN(n19183) );
  INV_X1 U22055 ( .A(n19183), .ZN(n19185) );
  NAND2_X1 U22056 ( .A1(n19533), .A2(n19185), .ZN(n19162) );
  NOR2_X1 U22057 ( .A1(n19094), .A2(n19093), .ZN(n19132) );
  AND2_X1 U22058 ( .A1(n17078), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19462) );
  NOR2_X1 U22059 ( .A1(n19095), .A2(n19541), .ZN(n19097) );
  NAND2_X1 U22060 ( .A1(n19097), .A2(n19339), .ZN(n19456) );
  NOR2_X2 U22061 ( .A1(n19184), .A2(n19096), .ZN(n19457) );
  NOR2_X1 U22062 ( .A1(n19541), .A2(n19273), .ZN(n19460) );
  NAND2_X1 U22063 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19460), .ZN(
        n19512) );
  NAND2_X1 U22064 ( .A1(n19512), .A2(n19162), .ZN(n19098) );
  INV_X1 U22065 ( .A(n19098), .ZN(n19160) );
  NOR2_X1 U22066 ( .A1(n19409), .A2(n19160), .ZN(n19134) );
  AOI22_X1 U22067 ( .A1(n19462), .A2(n19155), .B1(n19457), .B2(n19134), .ZN(
        n19101) );
  NOR2_X1 U22068 ( .A1(n19339), .A2(n19316), .ZN(n19386) );
  INV_X1 U22069 ( .A(n19097), .ZN(n19099) );
  NOR2_X1 U22070 ( .A1(n19386), .A2(n19099), .ZN(n19436) );
  AOI21_X1 U22071 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19184), .ZN(n19433) );
  AOI22_X1 U22072 ( .A1(n17078), .A2(n19436), .B1(n19433), .B2(n19098), .ZN(
        n19137) );
  NAND2_X1 U22073 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19461), .ZN(
        n19430) );
  INV_X1 U22074 ( .A(n19430), .ZN(n19507) );
  AND2_X1 U22075 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17078), .ZN(n19458) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19137), .B1(
        n19507), .B2(n19458), .ZN(n19100) );
  OAI211_X1 U22077 ( .C1(n19162), .C2(n19465), .A(n19101), .B(n19100), .ZN(
        P3_U2868) );
  NAND2_X1 U22078 ( .A1(n19132), .A2(n19102), .ZN(n19471) );
  AND2_X1 U22079 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17078), .ZN(n19467) );
  NOR2_X2 U22080 ( .A1(n19184), .A2(n19103), .ZN(n19466) );
  AOI22_X1 U22081 ( .A1(n19507), .A2(n19467), .B1(n19134), .B2(n19466), .ZN(
        n19105) );
  NOR2_X2 U22082 ( .A1(n19136), .A2(n21618), .ZN(n19468) );
  AOI22_X1 U22083 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19137), .B1(
        n19155), .B2(n19468), .ZN(n19104) );
  OAI211_X1 U22084 ( .C1(n19162), .C2(n19471), .A(n19105), .B(n19104), .ZN(
        P3_U2869) );
  AND2_X1 U22085 ( .A1(n17078), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19474) );
  NOR2_X2 U22086 ( .A1(n19184), .A2(n19107), .ZN(n19472) );
  AOI22_X1 U22087 ( .A1(n19155), .A2(n19474), .B1(n19134), .B2(n19472), .ZN(
        n19110) );
  INV_X1 U22088 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19108) );
  NOR2_X2 U22089 ( .A1(n19108), .A2(n19136), .ZN(n19473) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19137), .B1(
        n19507), .B2(n19473), .ZN(n19109) );
  OAI211_X1 U22091 ( .C1(n19162), .C2(n19477), .A(n19110), .B(n19109), .ZN(
        P3_U2870) );
  NOR2_X2 U22092 ( .A1(n19112), .A2(n19136), .ZN(n19478) );
  NOR2_X2 U22093 ( .A1(n19184), .A2(n19113), .ZN(n19479) );
  AOI22_X1 U22094 ( .A1(n19507), .A2(n19478), .B1(n19134), .B2(n19479), .ZN(
        n19116) );
  NOR2_X2 U22095 ( .A1(n19136), .A2(n19114), .ZN(n19480) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19137), .B1(
        n19155), .B2(n19480), .ZN(n19115) );
  OAI211_X1 U22097 ( .C1(n19162), .C2(n19483), .A(n19116), .B(n19115), .ZN(
        P3_U2871) );
  AND2_X1 U22098 ( .A1(n17078), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19486) );
  NOR2_X2 U22099 ( .A1(n19184), .A2(n19118), .ZN(n19484) );
  AOI22_X1 U22100 ( .A1(n19155), .A2(n19486), .B1(n19134), .B2(n19484), .ZN(
        n19121) );
  INV_X1 U22101 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19119) );
  NOR2_X2 U22102 ( .A1(n19119), .A2(n19136), .ZN(n19485) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19137), .B1(
        n19507), .B2(n19485), .ZN(n19120) );
  OAI211_X1 U22104 ( .C1(n19162), .C2(n19489), .A(n19121), .B(n19120), .ZN(
        P3_U2872) );
  NOR2_X2 U22105 ( .A1(n19123), .A2(n19136), .ZN(n19492) );
  NOR2_X2 U22106 ( .A1(n19184), .A2(n19124), .ZN(n19490) );
  AOI22_X1 U22107 ( .A1(n19507), .A2(n19492), .B1(n19134), .B2(n19490), .ZN(
        n19126) );
  AND2_X1 U22108 ( .A1(n17078), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19491) );
  AOI22_X1 U22109 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19137), .B1(
        n19155), .B2(n19491), .ZN(n19125) );
  OAI211_X1 U22110 ( .C1(n19162), .C2(n19495), .A(n19126), .B(n19125), .ZN(
        P3_U2873) );
  NOR2_X2 U22111 ( .A1(n19136), .A2(n19872), .ZN(n19498) );
  NOR2_X2 U22112 ( .A1(n19184), .A2(n19128), .ZN(n19496) );
  AOI22_X1 U22113 ( .A1(n19155), .A2(n19498), .B1(n19134), .B2(n19496), .ZN(
        n19130) );
  NOR2_X2 U22114 ( .A1(n16319), .A2(n19136), .ZN(n19497) );
  AOI22_X1 U22115 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19137), .B1(
        n19507), .B2(n19497), .ZN(n19129) );
  OAI211_X1 U22116 ( .C1(n19162), .C2(n19501), .A(n19130), .B(n19129), .ZN(
        P3_U2874) );
  AND2_X1 U22117 ( .A1(n17078), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19506) );
  NOR2_X2 U22118 ( .A1(n19184), .A2(n19133), .ZN(n19503) );
  AOI22_X1 U22119 ( .A1(n19155), .A2(n19506), .B1(n19134), .B2(n19503), .ZN(
        n19139) );
  NOR2_X2 U22120 ( .A1(n19136), .A2(n19135), .ZN(n19505) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19137), .B1(
        n19507), .B2(n19505), .ZN(n19138) );
  OAI211_X1 U22122 ( .C1(n19162), .C2(n19511), .A(n19139), .B(n19138), .ZN(
        P3_U2875) );
  NAND2_X1 U22123 ( .A1(n19185), .A2(n19316), .ZN(n19159) );
  NAND2_X1 U22124 ( .A1(n10732), .A2(n19560), .ZN(n19317) );
  NOR2_X1 U22125 ( .A1(n19183), .A2(n19317), .ZN(n19154) );
  AOI22_X1 U22126 ( .A1(n19178), .A2(n19462), .B1(n19457), .B2(n19154), .ZN(
        n19141) );
  AND2_X1 U22127 ( .A1(n19387), .A2(n19270), .ZN(n19459) );
  AND2_X1 U22128 ( .A1(n10732), .A2(n19459), .ZN(n19318) );
  AOI22_X1 U22129 ( .A1(n17078), .A2(n19460), .B1(n19185), .B2(n19318), .ZN(
        n19156) );
  AOI22_X1 U22130 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19156), .B1(
        n19458), .B2(n19155), .ZN(n19140) );
  OAI211_X1 U22131 ( .C1(n19465), .C2(n19159), .A(n19141), .B(n19140), .ZN(
        P3_U2876) );
  AOI22_X1 U22132 ( .A1(n19178), .A2(n19468), .B1(n19466), .B2(n19154), .ZN(
        n19143) );
  AOI22_X1 U22133 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19467), .ZN(n19142) );
  OAI211_X1 U22134 ( .C1(n19471), .C2(n19159), .A(n19143), .B(n19142), .ZN(
        P3_U2877) );
  AOI22_X1 U22135 ( .A1(n19178), .A2(n19474), .B1(n19472), .B2(n19154), .ZN(
        n19145) );
  AOI22_X1 U22136 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19473), .ZN(n19144) );
  OAI211_X1 U22137 ( .C1(n19477), .C2(n19159), .A(n19145), .B(n19144), .ZN(
        P3_U2878) );
  AOI22_X1 U22138 ( .A1(n19155), .A2(n19478), .B1(n19479), .B2(n19154), .ZN(
        n19147) );
  AOI22_X1 U22139 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19156), .B1(
        n19178), .B2(n19480), .ZN(n19146) );
  OAI211_X1 U22140 ( .C1(n19483), .C2(n19159), .A(n19147), .B(n19146), .ZN(
        P3_U2879) );
  AOI22_X1 U22141 ( .A1(n19155), .A2(n19485), .B1(n19484), .B2(n19154), .ZN(
        n19149) );
  AOI22_X1 U22142 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19156), .B1(
        n19178), .B2(n19486), .ZN(n19148) );
  OAI211_X1 U22143 ( .C1(n19489), .C2(n19159), .A(n19149), .B(n19148), .ZN(
        P3_U2880) );
  AOI22_X1 U22144 ( .A1(n19178), .A2(n19491), .B1(n19490), .B2(n19154), .ZN(
        n19151) );
  AOI22_X1 U22145 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19492), .ZN(n19150) );
  OAI211_X1 U22146 ( .C1(n19495), .C2(n19159), .A(n19151), .B(n19150), .ZN(
        P3_U2881) );
  AOI22_X1 U22147 ( .A1(n19178), .A2(n19498), .B1(n19496), .B2(n19154), .ZN(
        n19153) );
  AOI22_X1 U22148 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19497), .ZN(n19152) );
  OAI211_X1 U22149 ( .C1(n19501), .C2(n19159), .A(n19153), .B(n19152), .ZN(
        P3_U2882) );
  AOI22_X1 U22150 ( .A1(n19178), .A2(n19506), .B1(n19503), .B2(n19154), .ZN(
        n19158) );
  AOI22_X1 U22151 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19156), .B1(
        n19155), .B2(n19505), .ZN(n19157) );
  OAI211_X1 U22152 ( .C1(n19511), .C2(n19159), .A(n19158), .B(n19157), .ZN(
        P3_U2883) );
  NAND2_X1 U22153 ( .A1(n19185), .A2(n19339), .ZN(n19182) );
  INV_X1 U22154 ( .A(n19182), .ZN(n19244) );
  NOR2_X1 U22155 ( .A1(n19223), .A2(n19244), .ZN(n19206) );
  NOR2_X1 U22156 ( .A1(n19409), .A2(n19206), .ZN(n19177) );
  AOI22_X1 U22157 ( .A1(n19178), .A2(n19458), .B1(n19457), .B2(n19177), .ZN(
        n19164) );
  OAI21_X1 U22158 ( .B1(n19160), .B2(n19205), .A(n19206), .ZN(n19161) );
  OAI211_X1 U22159 ( .C1(n19244), .C2(n19660), .A(n19387), .B(n19161), .ZN(
        n19179) );
  AOI22_X1 U22160 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19462), .ZN(n19163) );
  OAI211_X1 U22161 ( .C1(n19465), .C2(n19182), .A(n19164), .B(n19163), .ZN(
        P3_U2884) );
  AOI22_X1 U22162 ( .A1(n19178), .A2(n19467), .B1(n19466), .B2(n19177), .ZN(
        n19166) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19468), .ZN(n19165) );
  OAI211_X1 U22164 ( .C1(n19471), .C2(n19182), .A(n19166), .B(n19165), .ZN(
        P3_U2885) );
  AOI22_X1 U22165 ( .A1(n19201), .A2(n19474), .B1(n19472), .B2(n19177), .ZN(
        n19168) );
  AOI22_X1 U22166 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n19473), .ZN(n19167) );
  OAI211_X1 U22167 ( .C1(n19477), .C2(n19182), .A(n19168), .B(n19167), .ZN(
        P3_U2886) );
  AOI22_X1 U22168 ( .A1(n19201), .A2(n19480), .B1(n19479), .B2(n19177), .ZN(
        n19170) );
  AOI22_X1 U22169 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n19478), .ZN(n19169) );
  OAI211_X1 U22170 ( .C1(n19483), .C2(n19182), .A(n19170), .B(n19169), .ZN(
        P3_U2887) );
  AOI22_X1 U22171 ( .A1(n19178), .A2(n19485), .B1(n19484), .B2(n19177), .ZN(
        n19172) );
  AOI22_X1 U22172 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19486), .ZN(n19171) );
  OAI211_X1 U22173 ( .C1(n19489), .C2(n19182), .A(n19172), .B(n19171), .ZN(
        P3_U2888) );
  AOI22_X1 U22174 ( .A1(n19178), .A2(n19492), .B1(n19490), .B2(n19177), .ZN(
        n19174) );
  AOI22_X1 U22175 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19491), .ZN(n19173) );
  OAI211_X1 U22176 ( .C1(n19495), .C2(n19182), .A(n19174), .B(n19173), .ZN(
        P3_U2889) );
  AOI22_X1 U22177 ( .A1(n19178), .A2(n19497), .B1(n19496), .B2(n19177), .ZN(
        n19176) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19498), .ZN(n19175) );
  OAI211_X1 U22179 ( .C1(n19501), .C2(n19182), .A(n19176), .B(n19175), .ZN(
        P3_U2890) );
  AOI22_X1 U22180 ( .A1(n19178), .A2(n19505), .B1(n19503), .B2(n19177), .ZN(
        n19181) );
  AOI22_X1 U22181 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19179), .B1(
        n19201), .B2(n19506), .ZN(n19180) );
  OAI211_X1 U22182 ( .C1(n19511), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        P3_U2891) );
  NOR2_X1 U22183 ( .A1(n10732), .A2(n19183), .ZN(n19228) );
  AND2_X1 U22184 ( .A1(n19560), .A2(n19228), .ZN(n19200) );
  AOI22_X1 U22185 ( .A1(n19201), .A2(n19458), .B1(n19457), .B2(n19200), .ZN(
        n19187) );
  AOI21_X1 U22186 ( .B1(n10732), .B2(n19205), .A(n19184), .ZN(n19272) );
  OAI211_X1 U22187 ( .C1(n19266), .C2(n19660), .A(n19185), .B(n19272), .ZN(
        n19202) );
  AOI22_X1 U22188 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19202), .B1(
        n19462), .B2(n19223), .ZN(n19186) );
  OAI211_X1 U22189 ( .C1(n19465), .C2(n19249), .A(n19187), .B(n19186), .ZN(
        P3_U2892) );
  AOI22_X1 U22190 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19202), .B1(
        n19466), .B2(n19200), .ZN(n19189) );
  AOI22_X1 U22191 ( .A1(n19201), .A2(n19467), .B1(n19468), .B2(n19223), .ZN(
        n19188) );
  OAI211_X1 U22192 ( .C1(n19471), .C2(n19249), .A(n19189), .B(n19188), .ZN(
        P3_U2893) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19202), .B1(
        n19472), .B2(n19200), .ZN(n19191) );
  AOI22_X1 U22194 ( .A1(n19201), .A2(n19473), .B1(n19474), .B2(n19223), .ZN(
        n19190) );
  OAI211_X1 U22195 ( .C1(n19477), .C2(n19249), .A(n19191), .B(n19190), .ZN(
        P3_U2894) );
  AOI22_X1 U22196 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19202), .B1(
        n19479), .B2(n19200), .ZN(n19193) );
  AOI22_X1 U22197 ( .A1(n19201), .A2(n19478), .B1(n19480), .B2(n19223), .ZN(
        n19192) );
  OAI211_X1 U22198 ( .C1(n19483), .C2(n19249), .A(n19193), .B(n19192), .ZN(
        P3_U2895) );
  AOI22_X1 U22199 ( .A1(n19486), .A2(n19223), .B1(n19484), .B2(n19200), .ZN(
        n19195) );
  AOI22_X1 U22200 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19202), .B1(
        n19201), .B2(n19485), .ZN(n19194) );
  OAI211_X1 U22201 ( .C1(n19489), .C2(n19249), .A(n19195), .B(n19194), .ZN(
        P3_U2896) );
  AOI22_X1 U22202 ( .A1(n19201), .A2(n19492), .B1(n19490), .B2(n19200), .ZN(
        n19197) );
  AOI22_X1 U22203 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19202), .B1(
        n19491), .B2(n19223), .ZN(n19196) );
  OAI211_X1 U22204 ( .C1(n19495), .C2(n19249), .A(n19197), .B(n19196), .ZN(
        P3_U2897) );
  AOI22_X1 U22205 ( .A1(n19201), .A2(n19497), .B1(n19496), .B2(n19200), .ZN(
        n19199) );
  AOI22_X1 U22206 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19202), .B1(
        n19498), .B2(n19223), .ZN(n19198) );
  OAI211_X1 U22207 ( .C1(n19501), .C2(n19249), .A(n19199), .B(n19198), .ZN(
        P3_U2898) );
  AOI22_X1 U22208 ( .A1(n19201), .A2(n19505), .B1(n19503), .B2(n19200), .ZN(
        n19204) );
  AOI22_X1 U22209 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19202), .B1(
        n19506), .B2(n19223), .ZN(n19203) );
  OAI211_X1 U22210 ( .C1(n19511), .C2(n19249), .A(n19204), .B(n19203), .ZN(
        P3_U2899) );
  INV_X1 U22211 ( .A(n19227), .ZN(n19271) );
  NAND2_X1 U22212 ( .A1(n19533), .A2(n19271), .ZN(n19248) );
  AOI21_X1 U22213 ( .B1(n19249), .B2(n19248), .A(n19409), .ZN(n19222) );
  AOI22_X1 U22214 ( .A1(n19462), .A2(n19244), .B1(n19457), .B2(n19222), .ZN(
        n19209) );
  INV_X1 U22215 ( .A(n19248), .ZN(n19290) );
  AOI221_X1 U22216 ( .B1(n19206), .B2(n19249), .C1(n19205), .C2(n19249), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22217 ( .B1(n19290), .B2(n19207), .A(n19387), .ZN(n19224) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19224), .B1(
        n19458), .B2(n19223), .ZN(n19208) );
  OAI211_X1 U22219 ( .C1(n19465), .C2(n19248), .A(n19209), .B(n19208), .ZN(
        P3_U2900) );
  AOI22_X1 U22220 ( .A1(n19468), .A2(n19244), .B1(n19466), .B2(n19222), .ZN(
        n19211) );
  AOI22_X1 U22221 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19224), .B1(
        n19467), .B2(n19223), .ZN(n19210) );
  OAI211_X1 U22222 ( .C1(n19471), .C2(n19248), .A(n19211), .B(n19210), .ZN(
        P3_U2901) );
  AOI22_X1 U22223 ( .A1(n19473), .A2(n19223), .B1(n19472), .B2(n19222), .ZN(
        n19213) );
  AOI22_X1 U22224 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19224), .B1(
        n19474), .B2(n19244), .ZN(n19212) );
  OAI211_X1 U22225 ( .C1(n19477), .C2(n19248), .A(n19213), .B(n19212), .ZN(
        P3_U2902) );
  AOI22_X1 U22226 ( .A1(n19480), .A2(n19244), .B1(n19479), .B2(n19222), .ZN(
        n19215) );
  AOI22_X1 U22227 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19224), .B1(
        n19478), .B2(n19223), .ZN(n19214) );
  OAI211_X1 U22228 ( .C1(n19483), .C2(n19248), .A(n19215), .B(n19214), .ZN(
        P3_U2903) );
  AOI22_X1 U22229 ( .A1(n19485), .A2(n19223), .B1(n19484), .B2(n19222), .ZN(
        n19217) );
  AOI22_X1 U22230 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19224), .B1(
        n19486), .B2(n19244), .ZN(n19216) );
  OAI211_X1 U22231 ( .C1(n19489), .C2(n19248), .A(n19217), .B(n19216), .ZN(
        P3_U2904) );
  AOI22_X1 U22232 ( .A1(n19492), .A2(n19223), .B1(n19490), .B2(n19222), .ZN(
        n19219) );
  AOI22_X1 U22233 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19224), .B1(
        n19491), .B2(n19244), .ZN(n19218) );
  OAI211_X1 U22234 ( .C1(n19495), .C2(n19248), .A(n19219), .B(n19218), .ZN(
        P3_U2905) );
  AOI22_X1 U22235 ( .A1(n19498), .A2(n19244), .B1(n19496), .B2(n19222), .ZN(
        n19221) );
  AOI22_X1 U22236 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19224), .B1(
        n19497), .B2(n19223), .ZN(n19220) );
  OAI211_X1 U22237 ( .C1(n19501), .C2(n19248), .A(n19221), .B(n19220), .ZN(
        P3_U2906) );
  AOI22_X1 U22238 ( .A1(n19505), .A2(n19223), .B1(n19503), .B2(n19222), .ZN(
        n19226) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19224), .B1(
        n19506), .B2(n19244), .ZN(n19225) );
  OAI211_X1 U22240 ( .C1(n19511), .C2(n19248), .A(n19226), .B(n19225), .ZN(
        P3_U2907) );
  NAND2_X1 U22241 ( .A1(n19316), .A2(n19271), .ZN(n19274) );
  NOR2_X1 U22242 ( .A1(n19317), .A2(n19227), .ZN(n19243) );
  AOI22_X1 U22243 ( .A1(n19458), .A2(n19244), .B1(n19457), .B2(n19243), .ZN(
        n19230) );
  AOI22_X1 U22244 ( .A1(n17078), .A2(n19228), .B1(n19318), .B2(n19271), .ZN(
        n19245) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19245), .B1(
        n19462), .B2(n19266), .ZN(n19229) );
  OAI211_X1 U22246 ( .C1(n19465), .C2(n19274), .A(n19230), .B(n19229), .ZN(
        P3_U2908) );
  AOI22_X1 U22247 ( .A1(n19467), .A2(n19244), .B1(n19466), .B2(n19243), .ZN(
        n19232) );
  AOI22_X1 U22248 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19245), .B1(
        n19468), .B2(n19266), .ZN(n19231) );
  OAI211_X1 U22249 ( .C1(n19471), .C2(n19274), .A(n19232), .B(n19231), .ZN(
        P3_U2909) );
  AOI22_X1 U22250 ( .A1(n19474), .A2(n19266), .B1(n19472), .B2(n19243), .ZN(
        n19234) );
  AOI22_X1 U22251 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19245), .B1(
        n19473), .B2(n19244), .ZN(n19233) );
  OAI211_X1 U22252 ( .C1(n19477), .C2(n19274), .A(n19234), .B(n19233), .ZN(
        P3_U2910) );
  AOI22_X1 U22253 ( .A1(n19480), .A2(n19266), .B1(n19479), .B2(n19243), .ZN(
        n19236) );
  AOI22_X1 U22254 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19245), .B1(
        n19478), .B2(n19244), .ZN(n19235) );
  OAI211_X1 U22255 ( .C1(n19483), .C2(n19274), .A(n19236), .B(n19235), .ZN(
        P3_U2911) );
  AOI22_X1 U22256 ( .A1(n19485), .A2(n19244), .B1(n19484), .B2(n19243), .ZN(
        n19238) );
  AOI22_X1 U22257 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19245), .B1(
        n19486), .B2(n19266), .ZN(n19237) );
  OAI211_X1 U22258 ( .C1(n19489), .C2(n19274), .A(n19238), .B(n19237), .ZN(
        P3_U2912) );
  AOI22_X1 U22259 ( .A1(n19492), .A2(n19244), .B1(n19490), .B2(n19243), .ZN(
        n19240) );
  AOI22_X1 U22260 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19245), .B1(
        n19491), .B2(n19266), .ZN(n19239) );
  OAI211_X1 U22261 ( .C1(n19495), .C2(n19274), .A(n19240), .B(n19239), .ZN(
        P3_U2913) );
  AOI22_X1 U22262 ( .A1(n19498), .A2(n19266), .B1(n19496), .B2(n19243), .ZN(
        n19242) );
  AOI22_X1 U22263 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19245), .B1(
        n19497), .B2(n19244), .ZN(n19241) );
  OAI211_X1 U22264 ( .C1(n19501), .C2(n19274), .A(n19242), .B(n19241), .ZN(
        P3_U2914) );
  AOI22_X1 U22265 ( .A1(n19506), .A2(n19266), .B1(n19503), .B2(n19243), .ZN(
        n19247) );
  AOI22_X1 U22266 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19245), .B1(
        n19505), .B2(n19244), .ZN(n19246) );
  OAI211_X1 U22267 ( .C1(n19511), .C2(n19274), .A(n19247), .B(n19246), .ZN(
        P3_U2915) );
  NAND2_X1 U22268 ( .A1(n19339), .A2(n19271), .ZN(n19296) );
  NAND2_X1 U22269 ( .A1(n19274), .A2(n19296), .ZN(n19295) );
  AND2_X1 U22270 ( .A1(n19560), .A2(n19295), .ZN(n19265) );
  AOI22_X1 U22271 ( .A1(n19458), .A2(n19266), .B1(n19457), .B2(n19265), .ZN(
        n19252) );
  NAND2_X1 U22272 ( .A1(n19249), .A2(n19248), .ZN(n19250) );
  OAI221_X1 U22273 ( .B1(n19295), .B2(n19435), .C1(n19295), .C2(n19250), .A(
        n19433), .ZN(n19267) );
  AOI22_X1 U22274 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19267), .B1(
        n19462), .B2(n19290), .ZN(n19251) );
  OAI211_X1 U22275 ( .C1(n19465), .C2(n19296), .A(n19252), .B(n19251), .ZN(
        P3_U2916) );
  AOI22_X1 U22276 ( .A1(n19467), .A2(n19266), .B1(n19466), .B2(n19265), .ZN(
        n19254) );
  AOI22_X1 U22277 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19267), .B1(
        n19468), .B2(n19290), .ZN(n19253) );
  OAI211_X1 U22278 ( .C1(n19471), .C2(n19296), .A(n19254), .B(n19253), .ZN(
        P3_U2917) );
  AOI22_X1 U22279 ( .A1(n19474), .A2(n19290), .B1(n19472), .B2(n19265), .ZN(
        n19256) );
  AOI22_X1 U22280 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19267), .B1(
        n19473), .B2(n19266), .ZN(n19255) );
  OAI211_X1 U22281 ( .C1(n19477), .C2(n19296), .A(n19256), .B(n19255), .ZN(
        P3_U2918) );
  AOI22_X1 U22282 ( .A1(n19479), .A2(n19265), .B1(n19478), .B2(n19266), .ZN(
        n19258) );
  AOI22_X1 U22283 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19267), .B1(
        n19480), .B2(n19290), .ZN(n19257) );
  OAI211_X1 U22284 ( .C1(n19483), .C2(n19296), .A(n19258), .B(n19257), .ZN(
        P3_U2919) );
  AOI22_X1 U22285 ( .A1(n19486), .A2(n19290), .B1(n19484), .B2(n19265), .ZN(
        n19260) );
  AOI22_X1 U22286 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19267), .B1(
        n19485), .B2(n19266), .ZN(n19259) );
  OAI211_X1 U22287 ( .C1(n19489), .C2(n19296), .A(n19260), .B(n19259), .ZN(
        P3_U2920) );
  AOI22_X1 U22288 ( .A1(n19492), .A2(n19266), .B1(n19490), .B2(n19265), .ZN(
        n19262) );
  AOI22_X1 U22289 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19267), .B1(
        n19491), .B2(n19290), .ZN(n19261) );
  OAI211_X1 U22290 ( .C1(n19495), .C2(n19296), .A(n19262), .B(n19261), .ZN(
        P3_U2921) );
  AOI22_X1 U22291 ( .A1(n19497), .A2(n19266), .B1(n19496), .B2(n19265), .ZN(
        n19264) );
  AOI22_X1 U22292 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19267), .B1(
        n19498), .B2(n19290), .ZN(n19263) );
  OAI211_X1 U22293 ( .C1(n19501), .C2(n19296), .A(n19264), .B(n19263), .ZN(
        P3_U2922) );
  AOI22_X1 U22294 ( .A1(n19506), .A2(n19290), .B1(n19503), .B2(n19265), .ZN(
        n19269) );
  AOI22_X1 U22295 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19267), .B1(
        n19505), .B2(n19266), .ZN(n19268) );
  OAI211_X1 U22296 ( .C1(n19511), .C2(n19296), .A(n19269), .B(n19268), .ZN(
        P3_U2923) );
  NOR3_X4 U22297 ( .A1(n19528), .A2(n19273), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19358) );
  NAND3_X1 U22298 ( .A1(n19272), .A2(n19271), .A3(n19270), .ZN(n19291) );
  NOR2_X1 U22299 ( .A1(n19273), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19319) );
  AOI22_X1 U22300 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19291), .B1(
        n19457), .B2(n19289), .ZN(n19276) );
  AOI22_X1 U22301 ( .A1(n19458), .A2(n19290), .B1(n19462), .B2(n19313), .ZN(
        n19275) );
  OAI211_X1 U22302 ( .C1(n19465), .C2(n19294), .A(n19276), .B(n19275), .ZN(
        P3_U2924) );
  AOI22_X1 U22303 ( .A1(n19468), .A2(n19313), .B1(n19466), .B2(n19289), .ZN(
        n19278) );
  AOI22_X1 U22304 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19291), .B1(
        n19467), .B2(n19290), .ZN(n19277) );
  OAI211_X1 U22305 ( .C1(n19471), .C2(n19294), .A(n19278), .B(n19277), .ZN(
        P3_U2925) );
  AOI22_X1 U22306 ( .A1(n19474), .A2(n19313), .B1(n19472), .B2(n19289), .ZN(
        n19280) );
  AOI22_X1 U22307 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19291), .B1(
        n19473), .B2(n19290), .ZN(n19279) );
  OAI211_X1 U22308 ( .C1(n19477), .C2(n19294), .A(n19280), .B(n19279), .ZN(
        P3_U2926) );
  AOI22_X1 U22309 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19291), .B1(
        n19479), .B2(n19289), .ZN(n19282) );
  AOI22_X1 U22310 ( .A1(n19480), .A2(n19313), .B1(n19478), .B2(n19290), .ZN(
        n19281) );
  OAI211_X1 U22311 ( .C1(n19483), .C2(n19294), .A(n19282), .B(n19281), .ZN(
        P3_U2927) );
  AOI22_X1 U22312 ( .A1(n19486), .A2(n19313), .B1(n19484), .B2(n19289), .ZN(
        n19284) );
  AOI22_X1 U22313 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19291), .B1(
        n19485), .B2(n19290), .ZN(n19283) );
  OAI211_X1 U22314 ( .C1(n19489), .C2(n19294), .A(n19284), .B(n19283), .ZN(
        P3_U2928) );
  AOI22_X1 U22315 ( .A1(n19492), .A2(n19290), .B1(n19490), .B2(n19289), .ZN(
        n19286) );
  AOI22_X1 U22316 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19291), .B1(
        n19491), .B2(n19313), .ZN(n19285) );
  OAI211_X1 U22317 ( .C1(n19495), .C2(n19294), .A(n19286), .B(n19285), .ZN(
        P3_U2929) );
  AOI22_X1 U22318 ( .A1(n19498), .A2(n19313), .B1(n19496), .B2(n19289), .ZN(
        n19288) );
  AOI22_X1 U22319 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19291), .B1(
        n19497), .B2(n19290), .ZN(n19287) );
  OAI211_X1 U22320 ( .C1(n19501), .C2(n19294), .A(n19288), .B(n19287), .ZN(
        P3_U2930) );
  AOI22_X1 U22321 ( .A1(n19505), .A2(n19290), .B1(n19503), .B2(n19289), .ZN(
        n19293) );
  AOI22_X1 U22322 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19291), .B1(
        n19506), .B2(n19313), .ZN(n19292) );
  OAI211_X1 U22323 ( .C1(n19511), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        P3_U2931) );
  NAND2_X1 U22324 ( .A1(n19533), .A2(n19364), .ZN(n19342) );
  NAND2_X1 U22325 ( .A1(n19294), .A2(n19342), .ZN(n19340) );
  OAI221_X1 U22326 ( .B1(n19340), .B2(n19435), .C1(n19340), .C2(n19295), .A(
        n19433), .ZN(n19312) );
  AND2_X1 U22327 ( .A1(n19560), .A2(n19340), .ZN(n19311) );
  AOI22_X1 U22328 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19312), .B1(
        n19457), .B2(n19311), .ZN(n19298) );
  INV_X1 U22329 ( .A(n19296), .ZN(n19335) );
  AOI22_X1 U22330 ( .A1(n19458), .A2(n19313), .B1(n19462), .B2(n19335), .ZN(
        n19297) );
  OAI211_X1 U22331 ( .C1(n19465), .C2(n19342), .A(n19298), .B(n19297), .ZN(
        P3_U2932) );
  AOI22_X1 U22332 ( .A1(n19467), .A2(n19313), .B1(n19466), .B2(n19311), .ZN(
        n19300) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19312), .B1(
        n19468), .B2(n19335), .ZN(n19299) );
  OAI211_X1 U22334 ( .C1(n19471), .C2(n19342), .A(n19300), .B(n19299), .ZN(
        P3_U2933) );
  AOI22_X1 U22335 ( .A1(n19474), .A2(n19335), .B1(n19472), .B2(n19311), .ZN(
        n19302) );
  AOI22_X1 U22336 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19312), .B1(
        n19473), .B2(n19313), .ZN(n19301) );
  OAI211_X1 U22337 ( .C1(n19477), .C2(n19342), .A(n19302), .B(n19301), .ZN(
        P3_U2934) );
  AOI22_X1 U22338 ( .A1(n19479), .A2(n19311), .B1(n19478), .B2(n19313), .ZN(
        n19304) );
  AOI22_X1 U22339 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19312), .B1(
        n19480), .B2(n19335), .ZN(n19303) );
  OAI211_X1 U22340 ( .C1(n19483), .C2(n19342), .A(n19304), .B(n19303), .ZN(
        P3_U2935) );
  AOI22_X1 U22341 ( .A1(n19486), .A2(n19335), .B1(n19484), .B2(n19311), .ZN(
        n19306) );
  AOI22_X1 U22342 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19312), .B1(
        n19485), .B2(n19313), .ZN(n19305) );
  OAI211_X1 U22343 ( .C1(n19489), .C2(n19342), .A(n19306), .B(n19305), .ZN(
        P3_U2936) );
  AOI22_X1 U22344 ( .A1(n19491), .A2(n19335), .B1(n19490), .B2(n19311), .ZN(
        n19308) );
  AOI22_X1 U22345 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19312), .B1(
        n19492), .B2(n19313), .ZN(n19307) );
  OAI211_X1 U22346 ( .C1(n19495), .C2(n19342), .A(n19308), .B(n19307), .ZN(
        P3_U2937) );
  AOI22_X1 U22347 ( .A1(n19498), .A2(n19335), .B1(n19496), .B2(n19311), .ZN(
        n19310) );
  AOI22_X1 U22348 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19312), .B1(
        n19497), .B2(n19313), .ZN(n19309) );
  OAI211_X1 U22349 ( .C1(n19501), .C2(n19342), .A(n19310), .B(n19309), .ZN(
        P3_U2938) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19312), .B1(
        n19503), .B2(n19311), .ZN(n19315) );
  AOI22_X1 U22351 ( .A1(n19505), .A2(n19313), .B1(n19506), .B2(n19335), .ZN(
        n19314) );
  OAI211_X1 U22352 ( .C1(n19511), .C2(n19342), .A(n19315), .B(n19314), .ZN(
        P3_U2939) );
  NAND2_X1 U22353 ( .A1(n19316), .A2(n19364), .ZN(n19363) );
  NOR2_X1 U22354 ( .A1(n19317), .A2(n19362), .ZN(n19334) );
  AOI22_X1 U22355 ( .A1(n19462), .A2(n19358), .B1(n19457), .B2(n19334), .ZN(
        n19321) );
  AOI22_X1 U22356 ( .A1(n17078), .A2(n19319), .B1(n19318), .B2(n19364), .ZN(
        n19336) );
  AOI22_X1 U22357 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19336), .B1(
        n19458), .B2(n19335), .ZN(n19320) );
  OAI211_X1 U22358 ( .C1(n19465), .C2(n19363), .A(n19321), .B(n19320), .ZN(
        P3_U2940) );
  AOI22_X1 U22359 ( .A1(n19468), .A2(n19358), .B1(n19466), .B2(n19334), .ZN(
        n19323) );
  AOI22_X1 U22360 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19336), .B1(
        n19467), .B2(n19335), .ZN(n19322) );
  OAI211_X1 U22361 ( .C1(n19471), .C2(n19363), .A(n19323), .B(n19322), .ZN(
        P3_U2941) );
  AOI22_X1 U22362 ( .A1(n19474), .A2(n19358), .B1(n19472), .B2(n19334), .ZN(
        n19325) );
  AOI22_X1 U22363 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19336), .B1(
        n19473), .B2(n19335), .ZN(n19324) );
  OAI211_X1 U22364 ( .C1(n19477), .C2(n19363), .A(n19325), .B(n19324), .ZN(
        P3_U2942) );
  AOI22_X1 U22365 ( .A1(n19480), .A2(n19358), .B1(n19479), .B2(n19334), .ZN(
        n19327) );
  AOI22_X1 U22366 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19336), .B1(
        n19478), .B2(n19335), .ZN(n19326) );
  OAI211_X1 U22367 ( .C1(n19483), .C2(n19363), .A(n19327), .B(n19326), .ZN(
        P3_U2943) );
  AOI22_X1 U22368 ( .A1(n19486), .A2(n19358), .B1(n19484), .B2(n19334), .ZN(
        n19329) );
  AOI22_X1 U22369 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19336), .B1(
        n19485), .B2(n19335), .ZN(n19328) );
  OAI211_X1 U22370 ( .C1(n19489), .C2(n19363), .A(n19329), .B(n19328), .ZN(
        P3_U2944) );
  AOI22_X1 U22371 ( .A1(n19491), .A2(n19358), .B1(n19490), .B2(n19334), .ZN(
        n19331) );
  AOI22_X1 U22372 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19336), .B1(
        n19492), .B2(n19335), .ZN(n19330) );
  OAI211_X1 U22373 ( .C1(n19495), .C2(n19363), .A(n19331), .B(n19330), .ZN(
        P3_U2945) );
  AOI22_X1 U22374 ( .A1(n19497), .A2(n19335), .B1(n19496), .B2(n19334), .ZN(
        n19333) );
  AOI22_X1 U22375 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19336), .B1(
        n19498), .B2(n19358), .ZN(n19332) );
  OAI211_X1 U22376 ( .C1(n19501), .C2(n19363), .A(n19333), .B(n19332), .ZN(
        P3_U2946) );
  AOI22_X1 U22377 ( .A1(n19506), .A2(n19358), .B1(n19503), .B2(n19334), .ZN(
        n19338) );
  AOI22_X1 U22378 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19336), .B1(
        n19505), .B2(n19335), .ZN(n19337) );
  OAI211_X1 U22379 ( .C1(n19511), .C2(n19363), .A(n19338), .B(n19337), .ZN(
        P3_U2947) );
  NAND2_X1 U22380 ( .A1(n19339), .A2(n19364), .ZN(n19384) );
  AOI21_X1 U22381 ( .B1(n19363), .B2(n19384), .A(n19409), .ZN(n19357) );
  AOI22_X1 U22382 ( .A1(n19458), .A2(n19358), .B1(n19457), .B2(n19357), .ZN(
        n19344) );
  NAND2_X1 U22383 ( .A1(n19363), .A2(n19384), .ZN(n19341) );
  OAI221_X1 U22384 ( .B1(n19341), .B2(n19435), .C1(n19341), .C2(n19340), .A(
        n19433), .ZN(n19359) );
  INV_X1 U22385 ( .A(n19342), .ZN(n19380) );
  AOI22_X1 U22386 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19359), .B1(
        n19462), .B2(n19380), .ZN(n19343) );
  OAI211_X1 U22387 ( .C1(n19465), .C2(n19384), .A(n19344), .B(n19343), .ZN(
        P3_U2948) );
  AOI22_X1 U22388 ( .A1(n19468), .A2(n19380), .B1(n19466), .B2(n19357), .ZN(
        n19346) );
  AOI22_X1 U22389 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19359), .B1(
        n19467), .B2(n19358), .ZN(n19345) );
  OAI211_X1 U22390 ( .C1(n19471), .C2(n19384), .A(n19346), .B(n19345), .ZN(
        P3_U2949) );
  AOI22_X1 U22391 ( .A1(n19473), .A2(n19358), .B1(n19472), .B2(n19357), .ZN(
        n19348) );
  AOI22_X1 U22392 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19359), .B1(
        n19474), .B2(n19380), .ZN(n19347) );
  OAI211_X1 U22393 ( .C1(n19477), .C2(n19384), .A(n19348), .B(n19347), .ZN(
        P3_U2950) );
  AOI22_X1 U22394 ( .A1(n19479), .A2(n19357), .B1(n19478), .B2(n19358), .ZN(
        n19350) );
  AOI22_X1 U22395 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19359), .B1(
        n19480), .B2(n19380), .ZN(n19349) );
  OAI211_X1 U22396 ( .C1(n19483), .C2(n19384), .A(n19350), .B(n19349), .ZN(
        P3_U2951) );
  AOI22_X1 U22397 ( .A1(n19486), .A2(n19380), .B1(n19484), .B2(n19357), .ZN(
        n19352) );
  AOI22_X1 U22398 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19359), .B1(
        n19485), .B2(n19358), .ZN(n19351) );
  OAI211_X1 U22399 ( .C1(n19489), .C2(n19384), .A(n19352), .B(n19351), .ZN(
        P3_U2952) );
  AOI22_X1 U22400 ( .A1(n19491), .A2(n19380), .B1(n19490), .B2(n19357), .ZN(
        n19354) );
  AOI22_X1 U22401 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19359), .B1(
        n19492), .B2(n19358), .ZN(n19353) );
  OAI211_X1 U22402 ( .C1(n19495), .C2(n19384), .A(n19354), .B(n19353), .ZN(
        P3_U2953) );
  AOI22_X1 U22403 ( .A1(n19497), .A2(n19358), .B1(n19496), .B2(n19357), .ZN(
        n19356) );
  AOI22_X1 U22404 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19359), .B1(
        n19498), .B2(n19380), .ZN(n19355) );
  OAI211_X1 U22405 ( .C1(n19501), .C2(n19384), .A(n19356), .B(n19355), .ZN(
        P3_U2954) );
  AOI22_X1 U22406 ( .A1(n19505), .A2(n19358), .B1(n19503), .B2(n19357), .ZN(
        n19361) );
  AOI22_X1 U22407 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19359), .B1(
        n19506), .B2(n19380), .ZN(n19360) );
  OAI211_X1 U22408 ( .C1(n19511), .C2(n19384), .A(n19361), .B(n19360), .ZN(
        P3_U2955) );
  NOR2_X1 U22409 ( .A1(n10732), .A2(n19362), .ZN(n19410) );
  AND2_X1 U22410 ( .A1(n19560), .A2(n19410), .ZN(n19379) );
  AOI22_X1 U22411 ( .A1(n19462), .A2(n19404), .B1(n19457), .B2(n19379), .ZN(
        n19366) );
  AOI22_X1 U22412 ( .A1(n17078), .A2(n19364), .B1(n19459), .B2(n19410), .ZN(
        n19381) );
  AOI22_X1 U22413 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19381), .B1(
        n19458), .B2(n19380), .ZN(n19365) );
  OAI211_X1 U22414 ( .C1(n19465), .C2(n19432), .A(n19366), .B(n19365), .ZN(
        P3_U2956) );
  AOI22_X1 U22415 ( .A1(n19468), .A2(n19404), .B1(n19466), .B2(n19379), .ZN(
        n19368) );
  AOI22_X1 U22416 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19381), .B1(
        n19467), .B2(n19380), .ZN(n19367) );
  OAI211_X1 U22417 ( .C1(n19471), .C2(n19432), .A(n19368), .B(n19367), .ZN(
        P3_U2957) );
  AOI22_X1 U22418 ( .A1(n19474), .A2(n19404), .B1(n19472), .B2(n19379), .ZN(
        n19370) );
  AOI22_X1 U22419 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19381), .B1(
        n19473), .B2(n19380), .ZN(n19369) );
  OAI211_X1 U22420 ( .C1(n19477), .C2(n19432), .A(n19370), .B(n19369), .ZN(
        P3_U2958) );
  AOI22_X1 U22421 ( .A1(n19480), .A2(n19404), .B1(n19479), .B2(n19379), .ZN(
        n19372) );
  AOI22_X1 U22422 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19381), .B1(
        n19478), .B2(n19380), .ZN(n19371) );
  OAI211_X1 U22423 ( .C1(n19483), .C2(n19432), .A(n19372), .B(n19371), .ZN(
        P3_U2959) );
  AOI22_X1 U22424 ( .A1(n19485), .A2(n19380), .B1(n19484), .B2(n19379), .ZN(
        n19374) );
  AOI22_X1 U22425 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19381), .B1(
        n19486), .B2(n19404), .ZN(n19373) );
  OAI211_X1 U22426 ( .C1(n19489), .C2(n19432), .A(n19374), .B(n19373), .ZN(
        P3_U2960) );
  AOI22_X1 U22427 ( .A1(n19491), .A2(n19404), .B1(n19490), .B2(n19379), .ZN(
        n19376) );
  AOI22_X1 U22428 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19381), .B1(
        n19492), .B2(n19380), .ZN(n19375) );
  OAI211_X1 U22429 ( .C1(n19495), .C2(n19432), .A(n19376), .B(n19375), .ZN(
        P3_U2961) );
  AOI22_X1 U22430 ( .A1(n19497), .A2(n19380), .B1(n19496), .B2(n19379), .ZN(
        n19378) );
  AOI22_X1 U22431 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19381), .B1(
        n19498), .B2(n19404), .ZN(n19377) );
  OAI211_X1 U22432 ( .C1(n19501), .C2(n19432), .A(n19378), .B(n19377), .ZN(
        P3_U2962) );
  AOI22_X1 U22433 ( .A1(n19505), .A2(n19380), .B1(n19503), .B2(n19379), .ZN(
        n19383) );
  AOI22_X1 U22434 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19381), .B1(
        n19506), .B2(n19404), .ZN(n19382) );
  OAI211_X1 U22435 ( .C1(n19511), .C2(n19432), .A(n19383), .B(n19382), .ZN(
        P3_U2963) );
  INV_X1 U22436 ( .A(n19461), .ZN(n19408) );
  NOR2_X2 U22437 ( .A1(n19408), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19504) );
  AOI21_X1 U22438 ( .B1(n19432), .B2(n19431), .A(n19409), .ZN(n19403) );
  AOI22_X1 U22439 ( .A1(n19462), .A2(n19426), .B1(n19457), .B2(n19403), .ZN(
        n19390) );
  AOI221_X1 U22440 ( .B1(n19386), .B2(n19432), .C1(n19385), .C2(n19432), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19388) );
  OAI21_X1 U22441 ( .B1(n19504), .B2(n19388), .A(n19387), .ZN(n19405) );
  AOI22_X1 U22442 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19405), .B1(
        n19458), .B2(n19404), .ZN(n19389) );
  OAI211_X1 U22443 ( .C1(n19465), .C2(n19431), .A(n19390), .B(n19389), .ZN(
        P3_U2964) );
  AOI22_X1 U22444 ( .A1(n19468), .A2(n19426), .B1(n19466), .B2(n19403), .ZN(
        n19392) );
  AOI22_X1 U22445 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19405), .B1(
        n19467), .B2(n19404), .ZN(n19391) );
  OAI211_X1 U22446 ( .C1(n19471), .C2(n19431), .A(n19392), .B(n19391), .ZN(
        P3_U2965) );
  AOI22_X1 U22447 ( .A1(n19474), .A2(n19426), .B1(n19472), .B2(n19403), .ZN(
        n19394) );
  AOI22_X1 U22448 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19405), .B1(
        n19473), .B2(n19404), .ZN(n19393) );
  OAI211_X1 U22449 ( .C1(n19477), .C2(n19431), .A(n19394), .B(n19393), .ZN(
        P3_U2966) );
  AOI22_X1 U22450 ( .A1(n19479), .A2(n19403), .B1(n19478), .B2(n19404), .ZN(
        n19396) );
  AOI22_X1 U22451 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19405), .B1(
        n19480), .B2(n19426), .ZN(n19395) );
  OAI211_X1 U22452 ( .C1(n19483), .C2(n19431), .A(n19396), .B(n19395), .ZN(
        P3_U2967) );
  AOI22_X1 U22453 ( .A1(n19485), .A2(n19404), .B1(n19484), .B2(n19403), .ZN(
        n19398) );
  AOI22_X1 U22454 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19405), .B1(
        n19486), .B2(n19426), .ZN(n19397) );
  OAI211_X1 U22455 ( .C1(n19489), .C2(n19431), .A(n19398), .B(n19397), .ZN(
        P3_U2968) );
  AOI22_X1 U22456 ( .A1(n19491), .A2(n19426), .B1(n19490), .B2(n19403), .ZN(
        n19400) );
  AOI22_X1 U22457 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19405), .B1(
        n19492), .B2(n19404), .ZN(n19399) );
  OAI211_X1 U22458 ( .C1(n19495), .C2(n19431), .A(n19400), .B(n19399), .ZN(
        P3_U2969) );
  AOI22_X1 U22459 ( .A1(n19498), .A2(n19426), .B1(n19496), .B2(n19403), .ZN(
        n19402) );
  AOI22_X1 U22460 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19405), .B1(
        n19497), .B2(n19404), .ZN(n19401) );
  OAI211_X1 U22461 ( .C1(n19501), .C2(n19431), .A(n19402), .B(n19401), .ZN(
        P3_U2970) );
  AOI22_X1 U22462 ( .A1(n19505), .A2(n19404), .B1(n19503), .B2(n19403), .ZN(
        n19407) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19405), .B1(
        n19506), .B2(n19426), .ZN(n19406) );
  OAI211_X1 U22464 ( .C1(n19511), .C2(n19431), .A(n19407), .B(n19406), .ZN(
        P3_U2971) );
  INV_X1 U22465 ( .A(n19432), .ZN(n19452) );
  NOR2_X1 U22466 ( .A1(n19409), .A2(n19408), .ZN(n19425) );
  AOI22_X1 U22467 ( .A1(n19462), .A2(n19452), .B1(n19457), .B2(n19425), .ZN(
        n19412) );
  AOI22_X1 U22468 ( .A1(n17078), .A2(n19410), .B1(n19461), .B2(n19459), .ZN(
        n19427) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19427), .B1(
        n19458), .B2(n19426), .ZN(n19411) );
  OAI211_X1 U22470 ( .C1(n19430), .C2(n19465), .A(n19412), .B(n19411), .ZN(
        P3_U2972) );
  AOI22_X1 U22471 ( .A1(n19467), .A2(n19426), .B1(n19466), .B2(n19425), .ZN(
        n19414) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19427), .B1(
        n19468), .B2(n19452), .ZN(n19413) );
  OAI211_X1 U22473 ( .C1(n19430), .C2(n19471), .A(n19414), .B(n19413), .ZN(
        P3_U2973) );
  AOI22_X1 U22474 ( .A1(n19474), .A2(n19452), .B1(n19472), .B2(n19425), .ZN(
        n19416) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19427), .B1(
        n19473), .B2(n19426), .ZN(n19415) );
  OAI211_X1 U22476 ( .C1(n19430), .C2(n19477), .A(n19416), .B(n19415), .ZN(
        P3_U2974) );
  AOI22_X1 U22477 ( .A1(n19479), .A2(n19425), .B1(n19478), .B2(n19426), .ZN(
        n19418) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19427), .B1(
        n19480), .B2(n19452), .ZN(n19417) );
  OAI211_X1 U22479 ( .C1(n19430), .C2(n19483), .A(n19418), .B(n19417), .ZN(
        P3_U2975) );
  AOI22_X1 U22480 ( .A1(n19486), .A2(n19452), .B1(n19484), .B2(n19425), .ZN(
        n19420) );
  AOI22_X1 U22481 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19427), .B1(
        n19485), .B2(n19426), .ZN(n19419) );
  OAI211_X1 U22482 ( .C1(n19430), .C2(n19489), .A(n19420), .B(n19419), .ZN(
        P3_U2976) );
  AOI22_X1 U22483 ( .A1(n19491), .A2(n19452), .B1(n19490), .B2(n19425), .ZN(
        n19422) );
  AOI22_X1 U22484 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19427), .B1(
        n19492), .B2(n19426), .ZN(n19421) );
  OAI211_X1 U22485 ( .C1(n19430), .C2(n19495), .A(n19422), .B(n19421), .ZN(
        P3_U2977) );
  AOI22_X1 U22486 ( .A1(n19497), .A2(n19426), .B1(n19496), .B2(n19425), .ZN(
        n19424) );
  AOI22_X1 U22487 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19427), .B1(
        n19498), .B2(n19452), .ZN(n19423) );
  OAI211_X1 U22488 ( .C1(n19430), .C2(n19501), .A(n19424), .B(n19423), .ZN(
        P3_U2978) );
  AOI22_X1 U22489 ( .A1(n19505), .A2(n19426), .B1(n19503), .B2(n19425), .ZN(
        n19429) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19427), .B1(
        n19506), .B2(n19452), .ZN(n19428) );
  OAI211_X1 U22491 ( .C1(n19430), .C2(n19511), .A(n19429), .B(n19428), .ZN(
        P3_U2979) );
  AOI22_X1 U22492 ( .A1(n19458), .A2(n19452), .B1(n19457), .B2(n19451), .ZN(
        n19438) );
  NAND2_X1 U22493 ( .A1(n19432), .A2(n19431), .ZN(n19434) );
  OAI221_X1 U22494 ( .B1(n19436), .B2(n19435), .C1(n19436), .C2(n19434), .A(
        n19433), .ZN(n19453) );
  AOI22_X1 U22495 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19453), .B1(
        n19462), .B2(n19504), .ZN(n19437) );
  OAI211_X1 U22496 ( .C1(n19465), .C2(n19456), .A(n19438), .B(n19437), .ZN(
        P3_U2980) );
  AOI22_X1 U22497 ( .A1(n19467), .A2(n19452), .B1(n19466), .B2(n19451), .ZN(
        n19440) );
  AOI22_X1 U22498 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19453), .B1(
        n19468), .B2(n19504), .ZN(n19439) );
  OAI211_X1 U22499 ( .C1(n19456), .C2(n19471), .A(n19440), .B(n19439), .ZN(
        P3_U2981) );
  AOI22_X1 U22500 ( .A1(n19473), .A2(n19452), .B1(n19472), .B2(n19451), .ZN(
        n19442) );
  AOI22_X1 U22501 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19453), .B1(
        n19474), .B2(n19504), .ZN(n19441) );
  OAI211_X1 U22502 ( .C1(n19456), .C2(n19477), .A(n19442), .B(n19441), .ZN(
        P3_U2982) );
  AOI22_X1 U22503 ( .A1(n19479), .A2(n19451), .B1(n19478), .B2(n19452), .ZN(
        n19444) );
  AOI22_X1 U22504 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19453), .B1(
        n19480), .B2(n19504), .ZN(n19443) );
  OAI211_X1 U22505 ( .C1(n19456), .C2(n19483), .A(n19444), .B(n19443), .ZN(
        P3_U2983) );
  AOI22_X1 U22506 ( .A1(n19485), .A2(n19452), .B1(n19484), .B2(n19451), .ZN(
        n19446) );
  AOI22_X1 U22507 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19453), .B1(
        n19486), .B2(n19504), .ZN(n19445) );
  OAI211_X1 U22508 ( .C1(n19456), .C2(n19489), .A(n19446), .B(n19445), .ZN(
        P3_U2984) );
  AOI22_X1 U22509 ( .A1(n19492), .A2(n19452), .B1(n19490), .B2(n19451), .ZN(
        n19448) );
  AOI22_X1 U22510 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19453), .B1(
        n19491), .B2(n19504), .ZN(n19447) );
  OAI211_X1 U22511 ( .C1(n19456), .C2(n19495), .A(n19448), .B(n19447), .ZN(
        P3_U2985) );
  AOI22_X1 U22512 ( .A1(n19497), .A2(n19452), .B1(n19496), .B2(n19451), .ZN(
        n19450) );
  AOI22_X1 U22513 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19453), .B1(
        n19498), .B2(n19504), .ZN(n19449) );
  OAI211_X1 U22514 ( .C1(n19456), .C2(n19501), .A(n19450), .B(n19449), .ZN(
        P3_U2986) );
  AOI22_X1 U22515 ( .A1(n19505), .A2(n19452), .B1(n19503), .B2(n19451), .ZN(
        n19455) );
  AOI22_X1 U22516 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19453), .B1(
        n19506), .B2(n19504), .ZN(n19454) );
  OAI211_X1 U22517 ( .C1(n19456), .C2(n19511), .A(n19455), .B(n19454), .ZN(
        P3_U2987) );
  AND2_X1 U22518 ( .A1(n19560), .A2(n19460), .ZN(n19502) );
  AOI22_X1 U22519 ( .A1(n19458), .A2(n19504), .B1(n19457), .B2(n19502), .ZN(
        n19464) );
  AOI22_X1 U22520 ( .A1(n17078), .A2(n19461), .B1(n19460), .B2(n19459), .ZN(
        n19508) );
  AOI22_X1 U22521 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19462), .ZN(n19463) );
  OAI211_X1 U22522 ( .C1(n19512), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P3_U2988) );
  AOI22_X1 U22523 ( .A1(n19467), .A2(n19504), .B1(n19466), .B2(n19502), .ZN(
        n19470) );
  AOI22_X1 U22524 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19468), .ZN(n19469) );
  OAI211_X1 U22525 ( .C1(n19512), .C2(n19471), .A(n19470), .B(n19469), .ZN(
        P3_U2989) );
  AOI22_X1 U22526 ( .A1(n19473), .A2(n19504), .B1(n19472), .B2(n19502), .ZN(
        n19476) );
  AOI22_X1 U22527 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19474), .ZN(n19475) );
  OAI211_X1 U22528 ( .C1(n19512), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P3_U2990) );
  AOI22_X1 U22529 ( .A1(n19479), .A2(n19502), .B1(n19478), .B2(n19504), .ZN(
        n19482) );
  AOI22_X1 U22530 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19480), .ZN(n19481) );
  OAI211_X1 U22531 ( .C1(n19512), .C2(n19483), .A(n19482), .B(n19481), .ZN(
        P3_U2991) );
  AOI22_X1 U22532 ( .A1(n19485), .A2(n19504), .B1(n19484), .B2(n19502), .ZN(
        n19488) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19486), .ZN(n19487) );
  OAI211_X1 U22534 ( .C1(n19512), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        P3_U2992) );
  AOI22_X1 U22535 ( .A1(n19507), .A2(n19491), .B1(n19490), .B2(n19502), .ZN(
        n19494) );
  AOI22_X1 U22536 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19508), .B1(
        n19492), .B2(n19504), .ZN(n19493) );
  OAI211_X1 U22537 ( .C1(n19512), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P3_U2993) );
  AOI22_X1 U22538 ( .A1(n19497), .A2(n19504), .B1(n19496), .B2(n19502), .ZN(
        n19500) );
  AOI22_X1 U22539 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19498), .ZN(n19499) );
  OAI211_X1 U22540 ( .C1(n19512), .C2(n19501), .A(n19500), .B(n19499), .ZN(
        P3_U2994) );
  AOI22_X1 U22541 ( .A1(n19505), .A2(n19504), .B1(n19503), .B2(n19502), .ZN(
        n19510) );
  AOI22_X1 U22542 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19506), .ZN(n19509) );
  OAI211_X1 U22543 ( .C1(n19512), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P3_U2995) );
  OAI22_X1 U22544 ( .A1(n19517), .A2(n19516), .B1(n19515), .B2(n19514), .ZN(
        n19518) );
  AOI221_X1 U22545 ( .B1(n9887), .B2(n10204), .C1(n19519), .C2(n10204), .A(
        n19518), .ZN(n19672) );
  INV_X1 U22546 ( .A(n19535), .ZN(n19537) );
  AOI211_X1 U22547 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19537), .A(
        n19521), .B(n19520), .ZN(n19548) );
  NAND2_X1 U22548 ( .A1(n19535), .A2(n19522), .ZN(n19526) );
  NOR2_X1 U22549 ( .A1(n19537), .A2(n19523), .ZN(n19525) );
  MUX2_X1 U22550 ( .A(n19526), .B(n19525), .S(n19524), .Z(n19544) );
  INV_X1 U22551 ( .A(n19527), .ZN(n19532) );
  INV_X1 U22552 ( .A(n19530), .ZN(n19529) );
  NOR3_X1 U22553 ( .A1(n19529), .A2(n10732), .A3(n19528), .ZN(n19531) );
  OAI22_X1 U22554 ( .A1(n19532), .A2(n19531), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19530), .ZN(n19534) );
  AOI21_X1 U22555 ( .B1(n19534), .B2(n19535), .A(n19533), .ZN(n19539) );
  AOI22_X1 U22556 ( .A1(n19537), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19536), .B2(n19535), .ZN(n19540) );
  OR2_X1 U22557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19540), .ZN(
        n19538) );
  AOI221_X1 U22558 ( .B1(n19539), .B2(n19538), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n19540), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19543) );
  OAI21_X1 U22559 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n19540), .ZN(n19542) );
  AOI222_X1 U22560 ( .A1(n19544), .A2(n19543), .B1(n19544), .B2(n19542), .C1(
        n19543), .C2(n19541), .ZN(n19547) );
  OAI21_X1 U22561 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19545), .ZN(n19546) );
  NAND4_X1 U22562 ( .A1(n19672), .A2(n19548), .A3(n19547), .A4(n19546), .ZN(
        n19556) );
  AOI211_X1 U22563 ( .C1(n19551), .C2(n19550), .A(n19549), .B(n19556), .ZN(
        n19658) );
  AOI21_X1 U22564 ( .B1(n19677), .B2(n19692), .A(n19658), .ZN(n19561) );
  NAND2_X1 U22565 ( .A1(n19677), .A2(n18469), .ZN(n19565) );
  INV_X1 U22566 ( .A(n19565), .ZN(n19552) );
  AOI211_X1 U22567 ( .C1(n19553), .C2(n19685), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n19552), .ZN(n19554) );
  AOI211_X1 U22568 ( .C1(n19675), .C2(n19556), .A(n19555), .B(n19554), .ZN(
        n19557) );
  OAI221_X1 U22569 ( .B1(n19657), .B2(n19561), .C1(n19657), .C2(n19558), .A(
        n19557), .ZN(P3_U2996) );
  NOR4_X1 U22570 ( .A1(n19657), .A2(n19559), .A3(n19682), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19568) );
  INV_X1 U22571 ( .A(n19568), .ZN(n19564) );
  NAND3_X1 U22572 ( .A1(n19562), .A2(n19561), .A3(n19560), .ZN(n19563) );
  NAND4_X1 U22573 ( .A1(n19566), .A2(n19565), .A3(n19564), .A4(n19563), .ZN(
        P3_U2997) );
  OAI21_X1 U22574 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19567), .ZN(n19569) );
  AOI21_X1 U22575 ( .B1(n19570), .B2(n19569), .A(n19568), .ZN(P3_U2998) );
  AND2_X1 U22576 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19571), .ZN(
        P3_U2999) );
  AND2_X1 U22577 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19571), .ZN(
        P3_U3000) );
  AND2_X1 U22578 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19571), .ZN(
        P3_U3001) );
  AND2_X1 U22579 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19571), .ZN(
        P3_U3002) );
  AND2_X1 U22580 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19571), .ZN(
        P3_U3003) );
  AND2_X1 U22581 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19571), .ZN(
        P3_U3004) );
  INV_X1 U22582 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21705) );
  NOR2_X1 U22583 ( .A1(n21705), .A2(n19656), .ZN(P3_U3005) );
  AND2_X1 U22584 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19571), .ZN(
        P3_U3006) );
  AND2_X1 U22585 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19571), .ZN(
        P3_U3007) );
  INV_X1 U22586 ( .A(P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n21687) );
  NOR2_X1 U22587 ( .A1(n21687), .A2(n19656), .ZN(P3_U3008) );
  AND2_X1 U22588 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19571), .ZN(
        P3_U3009) );
  AND2_X1 U22589 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19571), .ZN(
        P3_U3010) );
  AND2_X1 U22590 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19571), .ZN(
        P3_U3011) );
  AND2_X1 U22591 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19571), .ZN(
        P3_U3012) );
  AND2_X1 U22592 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19571), .ZN(
        P3_U3013) );
  AND2_X1 U22593 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19571), .ZN(
        P3_U3014) );
  AND2_X1 U22594 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19571), .ZN(
        P3_U3015) );
  AND2_X1 U22595 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19571), .ZN(
        P3_U3016) );
  AND2_X1 U22596 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19571), .ZN(
        P3_U3017) );
  AND2_X1 U22597 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19571), .ZN(
        P3_U3018) );
  AND2_X1 U22598 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19571), .ZN(
        P3_U3019) );
  AND2_X1 U22599 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19571), .ZN(
        P3_U3020) );
  AND2_X1 U22600 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19571), .ZN(P3_U3021) );
  AND2_X1 U22601 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19571), .ZN(P3_U3022) );
  AND2_X1 U22602 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19571), .ZN(P3_U3023) );
  AND2_X1 U22603 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19571), .ZN(P3_U3024) );
  AND2_X1 U22604 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19571), .ZN(P3_U3025) );
  AND2_X1 U22605 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19571), .ZN(P3_U3026) );
  AND2_X1 U22606 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19571), .ZN(P3_U3027) );
  AND2_X1 U22607 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19571), .ZN(P3_U3028) );
  OAI21_X1 U22608 ( .B1(n19572), .B2(n21512), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19573) );
  AOI22_X1 U22609 ( .A1(n19585), .A2(n19587), .B1(n19690), .B2(n19573), .ZN(
        n19574) );
  NAND3_X1 U22610 ( .A1(NA), .A2(n19585), .A3(n21652), .ZN(n19580) );
  OAI211_X1 U22611 ( .C1(n19575), .C2(n19682), .A(n19574), .B(n19580), .ZN(
        P3_U3029) );
  AOI21_X1 U22612 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19576) );
  AOI21_X1 U22613 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n19576), .ZN(
        n19577) );
  AOI22_X1 U22614 ( .A1(n19677), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19577), .ZN(n19578) );
  NAND2_X1 U22615 ( .A1(n19578), .A2(n19679), .ZN(P3_U3030) );
  NAND2_X1 U22616 ( .A1(n19677), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19581) );
  INV_X1 U22617 ( .A(n19581), .ZN(n19579) );
  AOI21_X1 U22618 ( .B1(n19585), .B2(n19580), .A(n19579), .ZN(n19586) );
  NOR2_X1 U22619 ( .A1(n19587), .A2(n21512), .ZN(n19583) );
  OAI22_X1 U22620 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19581), .ZN(n19582) );
  OAI22_X1 U22621 ( .A1(n19583), .A2(n19582), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19584) );
  OAI22_X1 U22622 ( .A1(n19586), .A2(n19587), .B1(n19585), .B2(n19584), .ZN(
        P3_U3031) );
  INV_X1 U22623 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19590) );
  NAND2_X2 U22624 ( .A1(n19647), .A2(n19587), .ZN(n19637) );
  OAI222_X1 U22625 ( .A1(n13988), .A2(n19632), .B1(n19588), .B2(n19647), .C1(
        n19590), .C2(n19637), .ZN(P3_U3032) );
  INV_X2 U22626 ( .A(n19589), .ZN(n19632) );
  OAI222_X1 U22627 ( .A1(n19637), .A2(n19593), .B1(n19591), .B2(n19647), .C1(
        n19590), .C2(n19632), .ZN(P3_U3033) );
  OAI222_X1 U22628 ( .A1(n19593), .A2(n19632), .B1(n19592), .B2(n19647), .C1(
        n19594), .C2(n19637), .ZN(P3_U3034) );
  OAI222_X1 U22629 ( .A1(n19637), .A2(n13980), .B1(n19595), .B2(n19647), .C1(
        n19594), .C2(n19632), .ZN(P3_U3035) );
  OAI222_X1 U22630 ( .A1(n19637), .A2(n19597), .B1(n19596), .B2(n19647), .C1(
        n13980), .C2(n19632), .ZN(P3_U3036) );
  OAI222_X1 U22631 ( .A1(n19637), .A2(n21686), .B1(n19598), .B2(n19647), .C1(
        n19597), .C2(n19632), .ZN(P3_U3037) );
  OAI222_X1 U22632 ( .A1(n19637), .A2(n19601), .B1(n19599), .B2(n19647), .C1(
        n21686), .C2(n19632), .ZN(P3_U3038) );
  OAI222_X1 U22633 ( .A1(n19601), .A2(n19632), .B1(n19600), .B2(n19647), .C1(
        n19602), .C2(n19637), .ZN(P3_U3039) );
  OAI222_X1 U22634 ( .A1(n19637), .A2(n19604), .B1(n19603), .B2(n19647), .C1(
        n19602), .C2(n19632), .ZN(P3_U3040) );
  OAI222_X1 U22635 ( .A1(n19637), .A2(n19606), .B1(n19605), .B2(n19647), .C1(
        n19604), .C2(n19632), .ZN(P3_U3041) );
  OAI222_X1 U22636 ( .A1(n19637), .A2(n19608), .B1(n19607), .B2(n19647), .C1(
        n19606), .C2(n19632), .ZN(P3_U3042) );
  INV_X1 U22637 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19610) );
  OAI222_X1 U22638 ( .A1(n19637), .A2(n19610), .B1(n19609), .B2(n19647), .C1(
        n19608), .C2(n19632), .ZN(P3_U3043) );
  OAI222_X1 U22639 ( .A1(n19637), .A2(n19613), .B1(n19611), .B2(n19647), .C1(
        n19610), .C2(n19632), .ZN(P3_U3044) );
  OAI222_X1 U22640 ( .A1(n19613), .A2(n19632), .B1(n19612), .B2(n19647), .C1(
        n19614), .C2(n19637), .ZN(P3_U3045) );
  OAI222_X1 U22641 ( .A1(n19637), .A2(n19616), .B1(n19615), .B2(n19647), .C1(
        n19614), .C2(n19632), .ZN(P3_U3046) );
  OAI222_X1 U22642 ( .A1(n19637), .A2(n19619), .B1(n19617), .B2(n19647), .C1(
        n19616), .C2(n19632), .ZN(P3_U3047) );
  OAI222_X1 U22643 ( .A1(n19619), .A2(n19632), .B1(n19618), .B2(n19647), .C1(
        n19620), .C2(n19637), .ZN(P3_U3048) );
  OAI222_X1 U22644 ( .A1(n19637), .A2(n19622), .B1(n19621), .B2(n19647), .C1(
        n19620), .C2(n19632), .ZN(P3_U3049) );
  INV_X1 U22645 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19625) );
  OAI222_X1 U22646 ( .A1(n19637), .A2(n19625), .B1(n19623), .B2(n19647), .C1(
        n19622), .C2(n19632), .ZN(P3_U3050) );
  OAI222_X1 U22647 ( .A1(n19625), .A2(n19632), .B1(n19624), .B2(n19647), .C1(
        n19626), .C2(n19637), .ZN(P3_U3051) );
  OAI222_X1 U22648 ( .A1(n19637), .A2(n19628), .B1(n19627), .B2(n19647), .C1(
        n19626), .C2(n19632), .ZN(P3_U3052) );
  OAI222_X1 U22649 ( .A1(n19637), .A2(n19631), .B1(n19629), .B2(n19647), .C1(
        n19628), .C2(n19632), .ZN(P3_U3053) );
  OAI222_X1 U22650 ( .A1(n19631), .A2(n19632), .B1(n19630), .B2(n19647), .C1(
        n19633), .C2(n19637), .ZN(P3_U3054) );
  OAI222_X1 U22651 ( .A1(n19637), .A2(n19635), .B1(n19634), .B2(n19647), .C1(
        n19633), .C2(n19632), .ZN(P3_U3055) );
  INV_X1 U22652 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19638) );
  OAI222_X1 U22653 ( .A1(n19637), .A2(n19638), .B1(n19636), .B2(n19647), .C1(
        n19635), .C2(n19632), .ZN(P3_U3056) );
  OAI222_X1 U22654 ( .A1(n19637), .A2(n19640), .B1(n19639), .B2(n19647), .C1(
        n19638), .C2(n19632), .ZN(P3_U3057) );
  OAI222_X1 U22655 ( .A1(n19637), .A2(n19643), .B1(n19641), .B2(n19647), .C1(
        n19640), .C2(n19632), .ZN(P3_U3058) );
  OAI222_X1 U22656 ( .A1(n19643), .A2(n19632), .B1(n19642), .B2(n19647), .C1(
        n19644), .C2(n19637), .ZN(P3_U3059) );
  OAI222_X1 U22657 ( .A1(n19637), .A2(n19649), .B1(n19645), .B2(n19647), .C1(
        n19644), .C2(n19632), .ZN(P3_U3060) );
  OAI222_X1 U22658 ( .A1(n19632), .A2(n19649), .B1(n19648), .B2(n19647), .C1(
        n19646), .C2(n19637), .ZN(P3_U3061) );
  INV_X1 U22659 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n21718) );
  AOI22_X1 U22660 ( .A1(n19647), .A2(n19650), .B1(n21718), .B2(n19690), .ZN(
        P3_U3274) );
  MUX2_X1 U22661 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n19690), .Z(P3_U3275) );
  OAI22_X1 U22662 ( .A1(n19690), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19647), .ZN(n19651) );
  INV_X1 U22663 ( .A(n19651), .ZN(P3_U3276) );
  OAI22_X1 U22664 ( .A1(n19690), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19647), .ZN(n19652) );
  INV_X1 U22665 ( .A(n19652), .ZN(P3_U3277) );
  OAI21_X1 U22666 ( .B1(n19656), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19654), 
        .ZN(n19653) );
  INV_X1 U22667 ( .A(n19653), .ZN(P3_U3280) );
  INV_X1 U22668 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19655) );
  OAI21_X1 U22669 ( .B1(n19656), .B2(n19655), .A(n19654), .ZN(P3_U3281) );
  NOR2_X1 U22670 ( .A1(n19658), .A2(n19657), .ZN(n19661) );
  OAI21_X1 U22671 ( .B1(n19661), .B2(n19660), .A(n19659), .ZN(P3_U3282) );
  NOR2_X1 U22672 ( .A1(n13988), .A2(n19667), .ZN(n19662) );
  AOI22_X1 U22673 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n19662), .B1(
        P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n19667), .ZN(n19663) );
  OAI221_X1 U22674 ( .B1(n19664), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .C1(n19664), .C2(P3_REIP_REG_0__SCAN_IN), .A(n19663), .ZN(P3_U3292) );
  INV_X1 U22675 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19668) );
  NOR2_X1 U22676 ( .A1(n19667), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U22677 ( .A1(n19668), .A2(n19667), .B1(n19666), .B2(n19665), .ZN(
        P3_U3293) );
  INV_X1 U22678 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19696) );
  OAI22_X1 U22679 ( .A1(n19690), .A2(n19696), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19647), .ZN(n19669) );
  INV_X1 U22680 ( .A(n19669), .ZN(P3_U3294) );
  INV_X1 U22681 ( .A(n19670), .ZN(n19673) );
  NAND2_X1 U22682 ( .A1(n19673), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19671) );
  OAI21_X1 U22683 ( .B1(n19673), .B2(n19672), .A(n19671), .ZN(P3_U3295) );
  OAI22_X1 U22684 ( .A1(n19677), .A2(n19676), .B1(n19675), .B2(n19674), .ZN(
        n19678) );
  NOR2_X1 U22685 ( .A1(n19695), .A2(n19678), .ZN(n19689) );
  AOI21_X1 U22686 ( .B1(n19681), .B2(n19680), .A(n19679), .ZN(n19683) );
  OAI211_X1 U22687 ( .C1(n19684), .C2(n19683), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19682), .ZN(n19686) );
  AOI21_X1 U22688 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19686), .A(n19685), 
        .ZN(n19688) );
  NAND2_X1 U22689 ( .A1(n19689), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19687) );
  OAI21_X1 U22690 ( .B1(n19689), .B2(n19688), .A(n19687), .ZN(P3_U3296) );
  OAI22_X1 U22691 ( .A1(n19690), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19647), .ZN(n19691) );
  INV_X1 U22692 ( .A(n19691), .ZN(P3_U3297) );
  AOI21_X1 U22693 ( .B1(n19693), .B2(n19692), .A(n19695), .ZN(n19699) );
  AOI22_X1 U22694 ( .A1(n19699), .A2(n19696), .B1(n19695), .B2(n19694), .ZN(
        P3_U3298) );
  INV_X1 U22695 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19698) );
  AOI21_X1 U22696 ( .B1(n19699), .B2(n19698), .A(n19697), .ZN(P3_U3299) );
  NAND2_X1 U22697 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20428), .ZN(n20420) );
  NOR2_X1 U22698 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20417) );
  INV_X1 U22699 ( .A(n20417), .ZN(n19700) );
  OAI21_X1 U22700 ( .B1(n20413), .B2(n20420), .A(n19700), .ZN(n20491) );
  AOI21_X1 U22701 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20491), .ZN(n19701) );
  INV_X1 U22702 ( .A(n19701), .ZN(P2_U2815) );
  CLKBUF_X2 U22703 ( .A(n19702), .Z(n20533) );
  INV_X1 U22704 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n19705) );
  AOI21_X1 U22705 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n19703), .A(n20421), 
        .ZN(n19704) );
  OAI22_X1 U22706 ( .A1(n20533), .A2(n19705), .B1(P2_STATE_REG_0__SCAN_IN), 
        .B2(n19704), .ZN(P2_U2817) );
  OAI21_X1 U22707 ( .B1(n20421), .B2(BS16), .A(n20491), .ZN(n20489) );
  OAI21_X1 U22708 ( .B1(n20491), .B2(n20356), .A(n20489), .ZN(P2_U2818) );
  NOR2_X1 U22709 ( .A1(n19707), .A2(n19706), .ZN(n20541) );
  OAI21_X1 U22710 ( .B1(n20541), .B2(n19709), .A(n19708), .ZN(P2_U2819) );
  NOR4_X1 U22711 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19713) );
  NOR4_X1 U22712 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19712) );
  NOR4_X1 U22713 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19711) );
  NOR4_X1 U22714 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19710) );
  NAND4_X1 U22715 ( .A1(n19713), .A2(n19712), .A3(n19711), .A4(n19710), .ZN(
        n19719) );
  NOR4_X1 U22716 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19717) );
  AOI211_X1 U22717 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_28__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19716) );
  NOR4_X1 U22718 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19715) );
  NOR4_X1 U22719 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19714) );
  NAND4_X1 U22720 ( .A1(n19717), .A2(n19716), .A3(n19715), .A4(n19714), .ZN(
        n19718) );
  NOR2_X1 U22721 ( .A1(n19719), .A2(n19718), .ZN(n19729) );
  INV_X1 U22722 ( .A(n19729), .ZN(n19727) );
  NOR2_X1 U22723 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19727), .ZN(n19721) );
  INV_X1 U22724 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21654) );
  AOI22_X1 U22725 ( .A1(n19721), .A2(n19722), .B1(n21654), .B2(n19727), .ZN(
        P2_U2820) );
  OR3_X1 U22726 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19726) );
  INV_X1 U22727 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U22728 ( .A1(n19721), .A2(n19726), .B1(n19727), .B2(n19720), .ZN(
        P2_U2821) );
  INV_X1 U22729 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20490) );
  NAND2_X1 U22730 ( .A1(n19721), .A2(n20490), .ZN(n19725) );
  OAI21_X1 U22731 ( .B1(n19722), .B2(n20429), .A(n19729), .ZN(n19723) );
  OAI21_X1 U22732 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19729), .A(n19723), 
        .ZN(n19724) );
  OAI221_X1 U22733 ( .B1(n19725), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19725), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19724), .ZN(P2_U2822) );
  INV_X1 U22734 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19728) );
  OAI221_X1 U22735 ( .B1(n19729), .B2(n19728), .C1(n19727), .C2(n19726), .A(
        n19725), .ZN(P2_U2823) );
  INV_X1 U22736 ( .A(n19730), .ZN(n19732) );
  AOI22_X1 U22737 ( .A1(n19732), .A2(n19761), .B1(n19731), .B2(n19760), .ZN(
        n19744) );
  INV_X1 U22738 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19740) );
  INV_X1 U22739 ( .A(n19733), .ZN(n19735) );
  AOI21_X1 U22740 ( .B1(n15727), .B2(n19735), .A(n19734), .ZN(n19736) );
  OAI21_X1 U22741 ( .B1(n19736), .B2(n15952), .A(n15709), .ZN(n19739) );
  AOI22_X1 U22742 ( .A1(n19737), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19746), .ZN(n19738) );
  OAI211_X1 U22743 ( .C1(n19767), .C2(n19740), .A(n19739), .B(n19738), .ZN(
        n19741) );
  AOI21_X1 U22744 ( .B1(n19742), .B2(n19750), .A(n19741), .ZN(n19743) );
  NAND2_X1 U22745 ( .A1(n19744), .A2(n19743), .ZN(P2_U2835) );
  AOI21_X1 U22746 ( .B1(n19746), .B2(P2_EBX_REG_6__SCAN_IN), .A(n19745), .ZN(
        n19747) );
  OAI21_X1 U22747 ( .B1(n20438), .B2(n19748), .A(n19747), .ZN(n19749) );
  AOI21_X1 U22748 ( .B1(n19751), .B2(n19750), .A(n19749), .ZN(n19766) );
  NAND2_X1 U22749 ( .A1(n19752), .A2(n19755), .ZN(n19754) );
  MUX2_X1 U22750 ( .A(n19755), .B(n19754), .S(n19753), .Z(n19758) );
  NAND3_X1 U22751 ( .A1(n19758), .A2(n19757), .A3(n19756), .ZN(n19764) );
  AOI22_X1 U22752 ( .A1(n19762), .A2(n19761), .B1(n19760), .B2(n19759), .ZN(
        n19763) );
  AND2_X1 U22753 ( .A1(n19764), .A2(n19763), .ZN(n19765) );
  OAI211_X1 U22754 ( .C1(n16669), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U2849) );
  INV_X1 U22755 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19769) );
  OAI22_X1 U22756 ( .A1(n19771), .A2(n19770), .B1(n19769), .B2(n19768), .ZN(
        n19772) );
  INV_X1 U22757 ( .A(n19772), .ZN(n19777) );
  XNOR2_X1 U22758 ( .A(n19774), .B(n19773), .ZN(n19775) );
  NAND2_X1 U22759 ( .A1(n19775), .A2(n19790), .ZN(n19776) );
  OAI211_X1 U22760 ( .C1(n19863), .C2(n19794), .A(n19777), .B(n19776), .ZN(
        P2_U2915) );
  AOI22_X1 U22761 ( .A1(n19778), .A2(n19786), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19785), .ZN(n19784) );
  OAI21_X1 U22762 ( .B1(n19781), .B2(n19780), .A(n19779), .ZN(n19782) );
  NAND2_X1 U22763 ( .A1(n19782), .A2(n19790), .ZN(n19783) );
  OAI211_X1 U22764 ( .C1(n19859), .C2(n19794), .A(n19784), .B(n19783), .ZN(
        P2_U2916) );
  AOI22_X1 U22765 ( .A1(n19786), .A2(n20513), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19785), .ZN(n19793) );
  OAI21_X1 U22766 ( .B1(n19789), .B2(n19788), .A(n19787), .ZN(n19791) );
  NAND2_X1 U22767 ( .A1(n19791), .A2(n19790), .ZN(n19792) );
  OAI211_X1 U22768 ( .C1(n19852), .C2(n19794), .A(n19793), .B(n19792), .ZN(
        P2_U2918) );
  NOR2_X1 U22769 ( .A1(n21684), .A2(n19798), .ZN(P2_U2920) );
  AOI22_X1 U22770 ( .A1(n19795), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n20548), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19796) );
  OAI21_X1 U22771 ( .B1(n19798), .B2(n19797), .A(n19796), .ZN(P2_U2921) );
  AOI22_X1 U22772 ( .A1(n19826), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19799) );
  OAI21_X1 U22773 ( .B1(n19800), .B2(n19828), .A(n19799), .ZN(P2_U2936) );
  INV_X1 U22774 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U22775 ( .A1(n19826), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19801) );
  OAI21_X1 U22776 ( .B1(n19802), .B2(n19828), .A(n19801), .ZN(P2_U2937) );
  AOI22_X1 U22777 ( .A1(n19826), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U22778 ( .B1(n19804), .B2(n19828), .A(n19803), .ZN(P2_U2938) );
  AOI22_X1 U22779 ( .A1(n19826), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U22780 ( .B1(n19806), .B2(n19828), .A(n19805), .ZN(P2_U2939) );
  AOI22_X1 U22781 ( .A1(n19826), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U22782 ( .B1(n19808), .B2(n19828), .A(n19807), .ZN(P2_U2940) );
  AOI22_X1 U22783 ( .A1(n19826), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U22784 ( .B1(n19810), .B2(n19828), .A(n19809), .ZN(P2_U2941) );
  AOI22_X1 U22785 ( .A1(n19826), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19811) );
  OAI21_X1 U22786 ( .B1(n19812), .B2(n19828), .A(n19811), .ZN(P2_U2942) );
  AOI22_X1 U22787 ( .A1(n19826), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U22788 ( .B1(n19814), .B2(n19828), .A(n19813), .ZN(P2_U2944) );
  AOI22_X1 U22789 ( .A1(n19826), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19815) );
  OAI21_X1 U22790 ( .B1(n19816), .B2(n19828), .A(n19815), .ZN(P2_U2945) );
  INV_X1 U22791 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U22792 ( .A1(n19826), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n19817) );
  OAI21_X1 U22793 ( .B1(n19818), .B2(n19828), .A(n19817), .ZN(P2_U2946) );
  AOI22_X1 U22794 ( .A1(n19826), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19819) );
  OAI21_X1 U22795 ( .B1(n19769), .B2(n19828), .A(n19819), .ZN(P2_U2947) );
  INV_X1 U22796 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U22797 ( .A1(n19826), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19820) );
  OAI21_X1 U22798 ( .B1(n19821), .B2(n19828), .A(n19820), .ZN(P2_U2948) );
  INV_X1 U22799 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U22800 ( .A1(n19826), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19822) );
  OAI21_X1 U22801 ( .B1(n19823), .B2(n19828), .A(n19822), .ZN(P2_U2949) );
  INV_X1 U22802 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U22803 ( .A1(n19826), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19824) );
  OAI21_X1 U22804 ( .B1(n19825), .B2(n19828), .A(n19824), .ZN(P2_U2950) );
  AOI22_X1 U22805 ( .A1(n19826), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n20548), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19827) );
  OAI21_X1 U22806 ( .B1(n13532), .B2(n19828), .A(n19827), .ZN(P2_U2951) );
  AOI22_X1 U22807 ( .A1(n19836), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19835), .ZN(n19831) );
  NAND2_X1 U22808 ( .A1(n19830), .A2(n19829), .ZN(n19837) );
  NAND2_X1 U22809 ( .A1(n19831), .A2(n19837), .ZN(P2_U2966) );
  AOI21_X1 U22810 ( .B1(n19835), .B2(P2_EAX_REG_8__SCAN_IN), .A(n19832), .ZN(
        n19833) );
  OAI21_X1 U22811 ( .B1(n21715), .B2(n19834), .A(n19833), .ZN(P2_U2975) );
  AOI22_X1 U22812 ( .A1(n19836), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19835), .ZN(n19838) );
  NAND2_X1 U22813 ( .A1(n19838), .A2(n19837), .ZN(P2_U2981) );
  NAND2_X1 U22814 ( .A1(n20521), .A2(n19950), .ZN(n19888) );
  INV_X1 U22815 ( .A(n19881), .ZN(n19840) );
  AND2_X1 U22816 ( .A1(n19841), .A2(n19840), .ZN(n19843) );
  INV_X1 U22817 ( .A(n20358), .ZN(n20402) );
  OAI21_X1 U22818 ( .B1(n20402), .B2(n19881), .A(n19948), .ZN(n19842) );
  AOI22_X1 U22819 ( .A1(n19882), .A2(n20353), .B1(n20352), .B2(n19881), .ZN(
        n19850) );
  NOR2_X1 U22820 ( .A1(n20169), .A2(n20517), .ZN(n19844) );
  OAI21_X1 U22821 ( .B1(n19911), .B2(n20406), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19847) );
  AOI21_X1 U22822 ( .B1(n19847), .B2(n19846), .A(n19845), .ZN(n19848) );
  OAI21_X1 U22823 ( .B1(n19848), .B2(n19881), .A(n20361), .ZN(n19885) );
  AOI22_X1 U22824 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n20406), .B2(n20241), .ZN(n19849) );
  OAI211_X1 U22825 ( .C1(n20297), .C2(n19898), .A(n19850), .B(n19849), .ZN(
        P2_U3048) );
  INV_X1 U22826 ( .A(n19884), .ZN(n19873) );
  INV_X1 U22827 ( .A(n19883), .ZN(n19871) );
  NOR2_X2 U22828 ( .A1(n20265), .A2(n19852), .ZN(n20368) );
  NAND2_X1 U22829 ( .A1(n19880), .A2(n20549), .ZN(n20311) );
  AOI22_X1 U22830 ( .A1(n19882), .A2(n20368), .B1(n20367), .B2(n19881), .ZN(
        n19854) );
  AOI22_X1 U22831 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19883), .ZN(n20372) );
  INV_X1 U22832 ( .A(n20372), .ZN(n20273) );
  AOI22_X1 U22833 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n20406), .B2(n20273), .ZN(n19853) );
  OAI211_X1 U22834 ( .C1(n20315), .C2(n19898), .A(n19854), .B(n19853), .ZN(
        P2_U3049) );
  NOR2_X2 U22835 ( .A1(n20265), .A2(n19855), .ZN(n21751) );
  NAND2_X1 U22836 ( .A1(n19880), .A2(n19856), .ZN(n20316) );
  AOI22_X1 U22837 ( .A1(n19882), .A2(n21751), .B1(n21750), .B2(n19881), .ZN(
        n19858) );
  AOI22_X1 U22838 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19883), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19884), .ZN(n20376) );
  INV_X1 U22839 ( .A(n20376), .ZN(n21753) );
  AOI22_X1 U22840 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n20406), .B2(n21753), .ZN(n19857) );
  OAI211_X1 U22841 ( .C1(n21759), .C2(n19898), .A(n19858), .B(n19857), .ZN(
        P2_U3050) );
  AOI22_X2 U22842 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19883), .ZN(n20321) );
  NOR2_X2 U22843 ( .A1(n20265), .A2(n19859), .ZN(n20378) );
  NAND2_X1 U22844 ( .A1(n19880), .A2(n19860), .ZN(n20320) );
  AOI22_X1 U22845 ( .A1(n19882), .A2(n20378), .B1(n20377), .B2(n19881), .ZN(
        n19862) );
  AOI22_X1 U22846 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19883), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19884), .ZN(n20382) );
  INV_X1 U22847 ( .A(n20382), .ZN(n20278) );
  AOI22_X1 U22848 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n20406), .B2(n20278), .ZN(n19861) );
  OAI211_X1 U22849 ( .C1(n20321), .C2(n19898), .A(n19862), .B(n19861), .ZN(
        P2_U3051) );
  AOI22_X2 U22850 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19883), .ZN(n20329) );
  NOR2_X2 U22851 ( .A1(n20265), .A2(n19863), .ZN(n20384) );
  NAND2_X1 U22852 ( .A1(n19880), .A2(n12647), .ZN(n20325) );
  AOI22_X1 U22853 ( .A1(n19882), .A2(n20384), .B1(n20383), .B2(n19881), .ZN(
        n19865) );
  AOI22_X1 U22854 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19883), .ZN(n20388) );
  AOI22_X1 U22855 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n20406), .B2(n20281), .ZN(n19864) );
  OAI211_X1 U22856 ( .C1(n20329), .C2(n19898), .A(n19865), .B(n19864), .ZN(
        P2_U3052) );
  AOI22_X2 U22857 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19883), .ZN(n20334) );
  INV_X1 U22858 ( .A(n19866), .ZN(n19867) );
  NOR2_X2 U22859 ( .A1(n20265), .A2(n19867), .ZN(n20390) );
  NAND2_X1 U22860 ( .A1(n19880), .A2(n19868), .ZN(n20330) );
  AOI22_X1 U22861 ( .A1(n19882), .A2(n20390), .B1(n20389), .B2(n19881), .ZN(
        n19870) );
  AOI22_X1 U22862 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19883), .ZN(n20394) );
  INV_X1 U22863 ( .A(n20394), .ZN(n20250) );
  AOI22_X1 U22864 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n20406), .B2(n20250), .ZN(n19869) );
  OAI211_X1 U22865 ( .C1(n20334), .C2(n19898), .A(n19870), .B(n19869), .ZN(
        P2_U3053) );
  OAI22_X2 U22866 ( .A1(n14983), .A2(n19873), .B1(n19872), .B2(n19871), .ZN(
        n20397) );
  NOR2_X2 U22867 ( .A1(n20265), .A2(n19874), .ZN(n20396) );
  AOI22_X1 U22868 ( .A1(n19882), .A2(n20396), .B1(n20395), .B2(n19881), .ZN(
        n19877) );
  INV_X1 U22869 ( .A(n20400), .ZN(n20253) );
  AOI22_X1 U22870 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n20406), .B2(n20253), .ZN(n19876) );
  OAI211_X1 U22871 ( .C1(n20256), .C2(n19898), .A(n19877), .B(n19876), .ZN(
        P2_U3054) );
  AOI22_X2 U22872 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19884), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19883), .ZN(n20341) );
  NOR2_X2 U22873 ( .A1(n20265), .A2(n19878), .ZN(n20403) );
  NAND2_X1 U22874 ( .A1(n19880), .A2(n19879), .ZN(n20340) );
  AOI22_X1 U22875 ( .A1(n19882), .A2(n20403), .B1(n20401), .B2(n19881), .ZN(
        n19887) );
  INV_X1 U22876 ( .A(n20411), .ZN(n20257) );
  AOI22_X1 U22877 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n20406), .B2(n20257), .ZN(n19886) );
  OAI211_X1 U22878 ( .C1(n20341), .C2(n19898), .A(n19887), .B(n19886), .ZN(
        P2_U3055) );
  INV_X1 U22879 ( .A(n19950), .ZN(n19945) );
  NOR2_X1 U22880 ( .A1(n20260), .A2(n19945), .ZN(n19909) );
  NOR3_X1 U22881 ( .A1(n11059), .A2(n19909), .A3(n20552), .ZN(n19889) );
  AOI211_X2 U22882 ( .C1(n19888), .C2(n20552), .A(n20262), .B(n19889), .ZN(
        n19910) );
  AOI22_X1 U22883 ( .A1(n19910), .A2(n20353), .B1(n20352), .B2(n19909), .ZN(
        n19895) );
  INV_X1 U22884 ( .A(n19888), .ZN(n19893) );
  INV_X1 U22885 ( .A(n19909), .ZN(n19890) );
  AOI211_X1 U22886 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19890), .A(n20265), 
        .B(n19889), .ZN(n19891) );
  OAI221_X1 U22887 ( .B1(n19893), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19893), 
        .C2(n19892), .A(n19891), .ZN(n19912) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20241), .ZN(n19894) );
  OAI211_X1 U22889 ( .C1(n20297), .C2(n19943), .A(n19895), .B(n19894), .ZN(
        P2_U3056) );
  AOI22_X1 U22890 ( .A1(n19910), .A2(n20368), .B1(n20367), .B2(n19909), .ZN(
        n19897) );
  INV_X1 U22891 ( .A(n19943), .ZN(n19932) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19912), .B1(
        n19932), .B2(n20369), .ZN(n19896) );
  OAI211_X1 U22893 ( .C1(n20372), .C2(n19898), .A(n19897), .B(n19896), .ZN(
        P2_U3057) );
  AOI22_X1 U22894 ( .A1(n19910), .A2(n21751), .B1(n21750), .B2(n19909), .ZN(
        n19900) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n21753), .ZN(n19899) );
  OAI211_X1 U22896 ( .C1(n21759), .C2(n19943), .A(n19900), .B(n19899), .ZN(
        P2_U3058) );
  AOI22_X1 U22897 ( .A1(n19910), .A2(n20378), .B1(n20377), .B2(n19909), .ZN(
        n19902) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20278), .ZN(n19901) );
  OAI211_X1 U22899 ( .C1(n20321), .C2(n19943), .A(n19902), .B(n19901), .ZN(
        P2_U3059) );
  AOI22_X1 U22900 ( .A1(n19910), .A2(n20384), .B1(n20383), .B2(n19909), .ZN(
        n19904) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20281), .ZN(n19903) );
  OAI211_X1 U22902 ( .C1(n20329), .C2(n19943), .A(n19904), .B(n19903), .ZN(
        P2_U3060) );
  AOI22_X1 U22903 ( .A1(n19910), .A2(n20390), .B1(n20389), .B2(n19909), .ZN(
        n19906) );
  AOI22_X1 U22904 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20250), .ZN(n19905) );
  OAI211_X1 U22905 ( .C1(n20334), .C2(n19943), .A(n19906), .B(n19905), .ZN(
        P2_U3061) );
  AOI22_X1 U22906 ( .A1(n19910), .A2(n20396), .B1(n20395), .B2(n19909), .ZN(
        n19908) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20253), .ZN(n19907) );
  OAI211_X1 U22908 ( .C1(n20256), .C2(n19943), .A(n19908), .B(n19907), .ZN(
        P2_U3062) );
  AOI22_X1 U22909 ( .A1(n19910), .A2(n20403), .B1(n20401), .B2(n19909), .ZN(
        n19914) );
  AOI22_X1 U22910 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n20257), .ZN(n19913) );
  OAI211_X1 U22911 ( .C1(n20341), .C2(n19943), .A(n19914), .B(n19913), .ZN(
        P2_U3063) );
  NOR2_X1 U22912 ( .A1(n20295), .A2(n19945), .ZN(n19937) );
  OAI21_X1 U22913 ( .B1(n11051), .B2(n19937), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19917) );
  INV_X1 U22914 ( .A(n19915), .ZN(n20171) );
  NOR2_X1 U22915 ( .A1(n20171), .A2(n19945), .ZN(n19918) );
  INV_X1 U22916 ( .A(n19918), .ZN(n19916) );
  NAND2_X1 U22917 ( .A1(n19917), .A2(n19916), .ZN(n19938) );
  AOI22_X1 U22918 ( .A1(n19938), .A2(n20353), .B1(n20352), .B2(n19937), .ZN(
        n19923) );
  AOI21_X1 U22919 ( .B1(n19943), .B2(n19984), .A(n20356), .ZN(n19919) );
  NOR3_X1 U22920 ( .A1(n19919), .A2(n19918), .A3(n20543), .ZN(n19921) );
  AOI211_X1 U22921 ( .C1(n11051), .C2(n20501), .A(n19948), .B(n19937), .ZN(
        n19920) );
  INV_X1 U22922 ( .A(n19984), .ZN(n19939) );
  INV_X1 U22923 ( .A(n20297), .ZN(n20363) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20363), .ZN(n19922) );
  OAI211_X1 U22925 ( .C1(n20366), .C2(n19943), .A(n19923), .B(n19922), .ZN(
        P2_U3064) );
  AOI22_X1 U22926 ( .A1(n19938), .A2(n20368), .B1(n20367), .B2(n19937), .ZN(
        n19925) );
  AOI22_X1 U22927 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19940), .B1(
        n19932), .B2(n20273), .ZN(n19924) );
  OAI211_X1 U22928 ( .C1(n20315), .C2(n19984), .A(n19925), .B(n19924), .ZN(
        P2_U3065) );
  AOI22_X1 U22929 ( .A1(n19938), .A2(n21751), .B1(n21750), .B2(n19937), .ZN(
        n19927) );
  INV_X1 U22930 ( .A(n21759), .ZN(n20373) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20373), .ZN(n19926) );
  OAI211_X1 U22932 ( .C1(n20376), .C2(n19943), .A(n19927), .B(n19926), .ZN(
        P2_U3066) );
  AOI22_X1 U22933 ( .A1(n19938), .A2(n20378), .B1(n20377), .B2(n19937), .ZN(
        n19929) );
  INV_X1 U22934 ( .A(n20321), .ZN(n20379) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20379), .ZN(n19928) );
  OAI211_X1 U22936 ( .C1(n20382), .C2(n19943), .A(n19929), .B(n19928), .ZN(
        P2_U3067) );
  AOI22_X1 U22937 ( .A1(n19938), .A2(n20384), .B1(n20383), .B2(n19937), .ZN(
        n19931) );
  AOI22_X1 U22938 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19940), .B1(
        n19932), .B2(n20281), .ZN(n19930) );
  OAI211_X1 U22939 ( .C1(n20329), .C2(n19984), .A(n19931), .B(n19930), .ZN(
        P2_U3068) );
  AOI22_X1 U22940 ( .A1(n19938), .A2(n20390), .B1(n20389), .B2(n19937), .ZN(
        n19934) );
  AOI22_X1 U22941 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19940), .B1(
        n19932), .B2(n20250), .ZN(n19933) );
  OAI211_X1 U22942 ( .C1(n20334), .C2(n19984), .A(n19934), .B(n19933), .ZN(
        P2_U3069) );
  AOI22_X1 U22943 ( .A1(n19938), .A2(n20396), .B1(n20395), .B2(n19937), .ZN(
        n19936) );
  AOI22_X1 U22944 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20397), .ZN(n19935) );
  OAI211_X1 U22945 ( .C1(n20400), .C2(n19943), .A(n19936), .B(n19935), .ZN(
        P2_U3070) );
  AOI22_X1 U22946 ( .A1(n19938), .A2(n20403), .B1(n20401), .B2(n19937), .ZN(
        n19942) );
  INV_X1 U22947 ( .A(n20341), .ZN(n20405) );
  AOI22_X1 U22948 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n20405), .ZN(n19941) );
  OAI211_X1 U22949 ( .C1(n20411), .C2(n19943), .A(n19942), .B(n19941), .ZN(
        P2_U3071) );
  NOR2_X1 U22950 ( .A1(n19945), .A2(n19944), .ZN(n19974) );
  INV_X1 U22951 ( .A(n19974), .ZN(n19977) );
  OAI22_X1 U22952 ( .A1(n19984), .A2(n20366), .B1(n19977), .B2(n20296), .ZN(
        n19946) );
  INV_X1 U22953 ( .A(n19946), .ZN(n19958) );
  INV_X1 U22954 ( .A(n19947), .ZN(n19949) );
  OAI21_X1 U22955 ( .B1(n19949), .B2(n20356), .A(n19948), .ZN(n19956) );
  NAND2_X1 U22956 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19950), .ZN(
        n19955) );
  INV_X1 U22957 ( .A(n19955), .ZN(n19953) );
  INV_X1 U22958 ( .A(n11057), .ZN(n19951) );
  OAI211_X1 U22959 ( .C1(n19951), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20543), 
        .B(n19977), .ZN(n19952) );
  OAI211_X1 U22960 ( .C1(n19956), .C2(n19953), .A(n20361), .B(n19952), .ZN(
        n19981) );
  OAI21_X1 U22961 ( .B1(n11057), .B2(n19974), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19954) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19981), .B1(
        n20353), .B2(n19980), .ZN(n19957) );
  OAI211_X1 U22963 ( .C1(n20297), .C2(n19978), .A(n19958), .B(n19957), .ZN(
        P2_U3072) );
  OAI22_X1 U22964 ( .A1(n19984), .A2(n20372), .B1(n20311), .B2(n19977), .ZN(
        n19959) );
  INV_X1 U22965 ( .A(n19959), .ZN(n19961) );
  AOI22_X1 U22966 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19981), .B1(
        n20368), .B2(n19980), .ZN(n19960) );
  OAI211_X1 U22967 ( .C1(n20315), .C2(n19978), .A(n19961), .B(n19960), .ZN(
        P2_U3073) );
  OAI22_X1 U22968 ( .A1(n19984), .A2(n20376), .B1(n20316), .B2(n19977), .ZN(
        n19962) );
  INV_X1 U22969 ( .A(n19962), .ZN(n19964) );
  AOI22_X1 U22970 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19981), .B1(
        n21751), .B2(n19980), .ZN(n19963) );
  OAI211_X1 U22971 ( .C1(n21759), .C2(n19978), .A(n19964), .B(n19963), .ZN(
        P2_U3074) );
  OAI22_X1 U22972 ( .A1(n19978), .A2(n20321), .B1(n19977), .B2(n20320), .ZN(
        n19965) );
  INV_X1 U22973 ( .A(n19965), .ZN(n19967) );
  AOI22_X1 U22974 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19981), .B1(
        n20378), .B2(n19980), .ZN(n19966) );
  OAI211_X1 U22975 ( .C1(n20382), .C2(n19984), .A(n19967), .B(n19966), .ZN(
        P2_U3075) );
  OAI22_X1 U22976 ( .A1(n19984), .A2(n20388), .B1(n20325), .B2(n19977), .ZN(
        n19968) );
  INV_X1 U22977 ( .A(n19968), .ZN(n19970) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19981), .B1(
        n20384), .B2(n19980), .ZN(n19969) );
  OAI211_X1 U22979 ( .C1(n20329), .C2(n19978), .A(n19970), .B(n19969), .ZN(
        P2_U3076) );
  OAI22_X1 U22980 ( .A1(n19978), .A2(n20334), .B1(n19977), .B2(n20330), .ZN(
        n19971) );
  INV_X1 U22981 ( .A(n19971), .ZN(n19973) );
  AOI22_X1 U22982 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19981), .B1(
        n20390), .B2(n19980), .ZN(n19972) );
  OAI211_X1 U22983 ( .C1(n20394), .C2(n19984), .A(n19973), .B(n19972), .ZN(
        P2_U3077) );
  AOI22_X1 U22984 ( .A1(n20397), .A2(n20008), .B1(n19974), .B2(n20395), .ZN(
        n19976) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19981), .B1(
        n20396), .B2(n19980), .ZN(n19975) );
  OAI211_X1 U22986 ( .C1(n20400), .C2(n19984), .A(n19976), .B(n19975), .ZN(
        P2_U3078) );
  OAI22_X1 U22987 ( .A1(n19978), .A2(n20341), .B1(n19977), .B2(n20340), .ZN(
        n19979) );
  INV_X1 U22988 ( .A(n19979), .ZN(n19983) );
  AOI22_X1 U22989 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19981), .B1(
        n20403), .B2(n19980), .ZN(n19982) );
  OAI211_X1 U22990 ( .C1(n20411), .C2(n19984), .A(n19983), .B(n19982), .ZN(
        P2_U3079) );
  INV_X1 U22991 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U22992 ( .A1(n20018), .A2(n20369), .B1(n20002), .B2(n20367), .ZN(
        n19986) );
  AOI22_X1 U22993 ( .A1(n20368), .A2(n20009), .B1(n20008), .B2(n20273), .ZN(
        n19985) );
  OAI211_X1 U22994 ( .C1(n20013), .C2(n19987), .A(n19986), .B(n19985), .ZN(
        P2_U3081) );
  INV_X1 U22995 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19991) );
  OAI22_X1 U22996 ( .A1(n20040), .A2(n21759), .B1(n20006), .B2(n20316), .ZN(
        n19988) );
  INV_X1 U22997 ( .A(n19988), .ZN(n19990) );
  AOI22_X1 U22998 ( .A1(n21751), .A2(n20009), .B1(n20008), .B2(n21753), .ZN(
        n19989) );
  OAI211_X1 U22999 ( .C1(n20013), .C2(n19991), .A(n19990), .B(n19989), .ZN(
        P2_U3082) );
  OAI22_X1 U23000 ( .A1(n20040), .A2(n20321), .B1(n20006), .B2(n20320), .ZN(
        n19992) );
  INV_X1 U23001 ( .A(n19992), .ZN(n19994) );
  AOI22_X1 U23002 ( .A1(n20378), .A2(n20009), .B1(n20008), .B2(n20278), .ZN(
        n19993) );
  OAI211_X1 U23003 ( .C1(n20013), .C2(n9814), .A(n19994), .B(n19993), .ZN(
        P2_U3083) );
  INV_X1 U23004 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21683) );
  OAI22_X1 U23005 ( .A1(n20040), .A2(n20329), .B1(n20006), .B2(n20325), .ZN(
        n19995) );
  INV_X1 U23006 ( .A(n19995), .ZN(n19997) );
  AOI22_X1 U23007 ( .A1(n20384), .A2(n20009), .B1(n20008), .B2(n20281), .ZN(
        n19996) );
  OAI211_X1 U23008 ( .C1(n20013), .C2(n21683), .A(n19997), .B(n19996), .ZN(
        P2_U3084) );
  INV_X1 U23009 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n20001) );
  OAI22_X1 U23010 ( .A1(n20040), .A2(n20334), .B1(n20006), .B2(n20330), .ZN(
        n19998) );
  INV_X1 U23011 ( .A(n19998), .ZN(n20000) );
  AOI22_X1 U23012 ( .A1(n20390), .A2(n20009), .B1(n20008), .B2(n20250), .ZN(
        n19999) );
  OAI211_X1 U23013 ( .C1(n20013), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3085) );
  INV_X1 U23014 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n20005) );
  AOI22_X1 U23015 ( .A1(n20018), .A2(n20397), .B1(n20002), .B2(n20395), .ZN(
        n20004) );
  AOI22_X1 U23016 ( .A1(n20396), .A2(n20009), .B1(n20008), .B2(n20253), .ZN(
        n20003) );
  OAI211_X1 U23017 ( .C1(n20013), .C2(n20005), .A(n20004), .B(n20003), .ZN(
        P2_U3086) );
  INV_X1 U23018 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20012) );
  OAI22_X1 U23019 ( .A1(n20040), .A2(n20341), .B1(n20006), .B2(n20340), .ZN(
        n20007) );
  INV_X1 U23020 ( .A(n20007), .ZN(n20011) );
  AOI22_X1 U23021 ( .A1(n20403), .A2(n20009), .B1(n20008), .B2(n20257), .ZN(
        n20010) );
  OAI211_X1 U23022 ( .C1(n20013), .C2(n20012), .A(n20011), .B(n20010), .ZN(
        P2_U3087) );
  INV_X1 U23023 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U23024 ( .A1(n20072), .A2(n20369), .B1(n20032), .B2(n20367), .ZN(
        n20015) );
  AOI22_X1 U23025 ( .A1(n20368), .A2(n20036), .B1(n20018), .B2(n20273), .ZN(
        n20014) );
  OAI211_X1 U23026 ( .C1(n20022), .C2(n20016), .A(n20015), .B(n20014), .ZN(
        P2_U3089) );
  INV_X1 U23027 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20021) );
  OAI22_X1 U23028 ( .A1(n20041), .A2(n21759), .B1(n20043), .B2(n20316), .ZN(
        n20017) );
  INV_X1 U23029 ( .A(n20017), .ZN(n20020) );
  AOI22_X1 U23030 ( .A1(n21751), .A2(n20036), .B1(n20018), .B2(n21753), .ZN(
        n20019) );
  OAI211_X1 U23031 ( .C1(n20022), .C2(n20021), .A(n20020), .B(n20019), .ZN(
        P2_U3090) );
  OAI22_X1 U23032 ( .A1(n20040), .A2(n20382), .B1(n20043), .B2(n20320), .ZN(
        n20023) );
  INV_X1 U23033 ( .A(n20023), .ZN(n20025) );
  AOI22_X1 U23034 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20037), .B1(
        n20378), .B2(n20036), .ZN(n20024) );
  OAI211_X1 U23035 ( .C1(n20321), .C2(n20041), .A(n20025), .B(n20024), .ZN(
        P2_U3091) );
  OAI22_X1 U23036 ( .A1(n20041), .A2(n20329), .B1(n20043), .B2(n20325), .ZN(
        n20026) );
  INV_X1 U23037 ( .A(n20026), .ZN(n20028) );
  AOI22_X1 U23038 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20037), .B1(
        n20384), .B2(n20036), .ZN(n20027) );
  OAI211_X1 U23039 ( .C1(n20388), .C2(n20040), .A(n20028), .B(n20027), .ZN(
        P2_U3092) );
  OAI22_X1 U23040 ( .A1(n20040), .A2(n20394), .B1(n20043), .B2(n20330), .ZN(
        n20029) );
  INV_X1 U23041 ( .A(n20029), .ZN(n20031) );
  AOI22_X1 U23042 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20037), .B1(
        n20390), .B2(n20036), .ZN(n20030) );
  OAI211_X1 U23043 ( .C1(n20334), .C2(n20041), .A(n20031), .B(n20030), .ZN(
        P2_U3093) );
  AOI22_X1 U23044 ( .A1(n20072), .A2(n20397), .B1(n20032), .B2(n20395), .ZN(
        n20034) );
  AOI22_X1 U23045 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20037), .B1(
        n20396), .B2(n20036), .ZN(n20033) );
  OAI211_X1 U23046 ( .C1(n20400), .C2(n20040), .A(n20034), .B(n20033), .ZN(
        P2_U3094) );
  OAI22_X1 U23047 ( .A1(n20041), .A2(n20341), .B1(n20043), .B2(n20340), .ZN(
        n20035) );
  INV_X1 U23048 ( .A(n20035), .ZN(n20039) );
  AOI22_X1 U23049 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20037), .B1(
        n20403), .B2(n20036), .ZN(n20038) );
  OAI211_X1 U23050 ( .C1(n20411), .C2(n20040), .A(n20039), .B(n20038), .ZN(
        P2_U3095) );
  NAND2_X1 U23051 ( .A1(n20041), .A2(n20102), .ZN(n20042) );
  NAND2_X1 U23052 ( .A1(n20042), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20044) );
  NAND2_X1 U23053 ( .A1(n20044), .A2(n20043), .ZN(n20047) );
  INV_X1 U23054 ( .A(n11055), .ZN(n20045) );
  AOI21_X1 U23055 ( .B1(n20045), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U23056 ( .A1(n20047), .A2(n20046), .ZN(n20049) );
  NOR2_X1 U23057 ( .A1(n20295), .A2(n20079), .ZN(n20070) );
  INV_X1 U23058 ( .A(n20070), .ZN(n20048) );
  NAND2_X1 U23059 ( .A1(n20049), .A2(n20048), .ZN(n20050) );
  INV_X1 U23060 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U23061 ( .B1(n11055), .B2(n20070), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20051) );
  AOI22_X1 U23062 ( .A1(n20071), .A2(n20353), .B1(n20352), .B2(n20070), .ZN(
        n20053) );
  INV_X1 U23063 ( .A(n20102), .ZN(n20057) );
  AOI22_X1 U23064 ( .A1(n20072), .A2(n20241), .B1(n20057), .B2(n20363), .ZN(
        n20052) );
  OAI211_X1 U23065 ( .C1(n20061), .C2(n20054), .A(n20053), .B(n20052), .ZN(
        P2_U3096) );
  AOI22_X1 U23066 ( .A1(n20071), .A2(n20368), .B1(n20367), .B2(n20070), .ZN(
        n20056) );
  AOI22_X1 U23067 ( .A1(n20072), .A2(n20273), .B1(n20057), .B2(n20369), .ZN(
        n20055) );
  OAI211_X1 U23068 ( .C1(n20061), .C2(n21658), .A(n20056), .B(n20055), .ZN(
        P2_U3097) );
  AOI22_X1 U23069 ( .A1(n20071), .A2(n21751), .B1(n21750), .B2(n20070), .ZN(
        n20059) );
  AOI22_X1 U23070 ( .A1(n20072), .A2(n21753), .B1(n20057), .B2(n20373), .ZN(
        n20058) );
  OAI211_X1 U23071 ( .C1(n20061), .C2(n20060), .A(n20059), .B(n20058), .ZN(
        P2_U3098) );
  AOI22_X1 U23072 ( .A1(n20071), .A2(n20378), .B1(n20377), .B2(n20070), .ZN(
        n20063) );
  AOI22_X1 U23073 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20073), .B1(
        n20072), .B2(n20278), .ZN(n20062) );
  OAI211_X1 U23074 ( .C1(n20321), .C2(n20102), .A(n20063), .B(n20062), .ZN(
        P2_U3099) );
  AOI22_X1 U23075 ( .A1(n20071), .A2(n20384), .B1(n20383), .B2(n20070), .ZN(
        n20065) );
  AOI22_X1 U23076 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20073), .B1(
        n20072), .B2(n20281), .ZN(n20064) );
  OAI211_X1 U23077 ( .C1(n20329), .C2(n20102), .A(n20065), .B(n20064), .ZN(
        P2_U3100) );
  AOI22_X1 U23078 ( .A1(n20071), .A2(n20390), .B1(n20389), .B2(n20070), .ZN(
        n20067) );
  AOI22_X1 U23079 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20073), .B1(
        n20072), .B2(n20250), .ZN(n20066) );
  OAI211_X1 U23080 ( .C1(n20334), .C2(n20102), .A(n20067), .B(n20066), .ZN(
        P2_U3101) );
  AOI22_X1 U23081 ( .A1(n20071), .A2(n20396), .B1(n20395), .B2(n20070), .ZN(
        n20069) );
  AOI22_X1 U23082 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20073), .B1(
        n20072), .B2(n20253), .ZN(n20068) );
  OAI211_X1 U23083 ( .C1(n20256), .C2(n20102), .A(n20069), .B(n20068), .ZN(
        P2_U3102) );
  AOI22_X1 U23084 ( .A1(n20071), .A2(n20403), .B1(n20401), .B2(n20070), .ZN(
        n20075) );
  AOI22_X1 U23085 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20073), .B1(
        n20072), .B2(n20257), .ZN(n20074) );
  OAI211_X1 U23086 ( .C1(n20341), .C2(n20102), .A(n20075), .B(n20074), .ZN(
        P2_U3103) );
  NAND2_X1 U23087 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20076), .ZN(
        n20078) );
  OAI21_X1 U23088 ( .B1(n11060), .B2(n20110), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20077) );
  AOI22_X1 U23089 ( .A1(n20098), .A2(n20353), .B1(n20352), .B2(n20110), .ZN(
        n20085) );
  INV_X1 U23090 ( .A(n20492), .ZN(n20080) );
  OAI22_X1 U23091 ( .A1(n20080), .A2(n20356), .B1(n20079), .B2(n20521), .ZN(
        n20083) );
  INV_X1 U23092 ( .A(n11060), .ZN(n20081) );
  INV_X1 U23093 ( .A(n20110), .ZN(n20107) );
  OAI211_X1 U23094 ( .C1(n20081), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20543), 
        .B(n20107), .ZN(n20082) );
  NAND3_X1 U23095 ( .A1(n20083), .A2(n20361), .A3(n20082), .ZN(n20099) );
  AND2_X2 U23096 ( .A1(n20492), .A2(n20269), .ZN(n20128) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20363), .ZN(n20084) );
  OAI211_X1 U23098 ( .C1(n20366), .C2(n20102), .A(n20085), .B(n20084), .ZN(
        P2_U3104) );
  AOI22_X1 U23099 ( .A1(n20098), .A2(n20368), .B1(n20110), .B2(n20367), .ZN(
        n20087) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20369), .ZN(n20086) );
  OAI211_X1 U23101 ( .C1(n20372), .C2(n20102), .A(n20087), .B(n20086), .ZN(
        P2_U3105) );
  AOI22_X1 U23102 ( .A1(n20098), .A2(n21751), .B1(n20110), .B2(n21750), .ZN(
        n20089) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20373), .ZN(n20088) );
  OAI211_X1 U23104 ( .C1(n20376), .C2(n20102), .A(n20089), .B(n20088), .ZN(
        P2_U3106) );
  AOI22_X1 U23105 ( .A1(n20098), .A2(n20378), .B1(n20110), .B2(n20377), .ZN(
        n20091) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20379), .ZN(n20090) );
  OAI211_X1 U23107 ( .C1(n20382), .C2(n20102), .A(n20091), .B(n20090), .ZN(
        P2_U3107) );
  AOI22_X1 U23108 ( .A1(n20098), .A2(n20384), .B1(n20110), .B2(n20383), .ZN(
        n20093) );
  INV_X1 U23109 ( .A(n20329), .ZN(n20385) );
  AOI22_X1 U23110 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20385), .ZN(n20092) );
  OAI211_X1 U23111 ( .C1(n20388), .C2(n20102), .A(n20093), .B(n20092), .ZN(
        P2_U3108) );
  AOI22_X1 U23112 ( .A1(n20098), .A2(n20390), .B1(n20110), .B2(n20389), .ZN(
        n20095) );
  INV_X1 U23113 ( .A(n20334), .ZN(n20391) );
  AOI22_X1 U23114 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20391), .ZN(n20094) );
  OAI211_X1 U23115 ( .C1(n20394), .C2(n20102), .A(n20095), .B(n20094), .ZN(
        P2_U3109) );
  AOI22_X1 U23116 ( .A1(n20098), .A2(n20396), .B1(n20110), .B2(n20395), .ZN(
        n20097) );
  AOI22_X1 U23117 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20397), .ZN(n20096) );
  OAI211_X1 U23118 ( .C1(n20400), .C2(n20102), .A(n20097), .B(n20096), .ZN(
        P2_U3110) );
  AOI22_X1 U23119 ( .A1(n20098), .A2(n20403), .B1(n20110), .B2(n20401), .ZN(
        n20101) );
  AOI22_X1 U23120 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20099), .B1(
        n20128), .B2(n20405), .ZN(n20100) );
  OAI211_X1 U23121 ( .C1(n20411), .C2(n20102), .A(n20101), .B(n20100), .ZN(
        P2_U3111) );
  NAND2_X2 U23122 ( .A1(n20135), .A2(n20526), .ZN(n20162) );
  NAND2_X1 U23123 ( .A1(n20512), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20202) );
  INV_X1 U23124 ( .A(n20202), .ZN(n20198) );
  NAND2_X1 U23125 ( .A1(n20198), .A2(n20521), .ZN(n20141) );
  AOI22_X1 U23126 ( .A1(n20128), .A2(n20241), .B1(n20127), .B2(n20352), .ZN(
        n20114) );
  INV_X1 U23127 ( .A(n20128), .ZN(n20104) );
  AOI21_X1 U23128 ( .B1(n20104), .B2(n20162), .A(n20356), .ZN(n20105) );
  NOR2_X1 U23129 ( .A1(n20105), .A2(n20543), .ZN(n20109) );
  OAI21_X1 U23130 ( .B1(n11054), .B2(n20552), .A(n20501), .ZN(n20106) );
  AOI21_X1 U23131 ( .B1(n20109), .B2(n20107), .A(n20106), .ZN(n20108) );
  OAI21_X1 U23132 ( .B1(n20127), .B2(n20108), .A(n20361), .ZN(n20130) );
  OAI21_X1 U23133 ( .B1(n20110), .B2(n20127), .A(n20109), .ZN(n20112) );
  OAI21_X1 U23134 ( .B1(n11054), .B2(n20127), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20111) );
  AOI22_X1 U23135 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20130), .B1(
        n20353), .B2(n20129), .ZN(n20113) );
  OAI211_X1 U23136 ( .C1(n20297), .C2(n20162), .A(n20114), .B(n20113), .ZN(
        P2_U3112) );
  AOI22_X1 U23137 ( .A1(n20128), .A2(n20273), .B1(n20127), .B2(n20367), .ZN(
        n20116) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20368), .ZN(n20115) );
  OAI211_X1 U23139 ( .C1(n20315), .C2(n20162), .A(n20116), .B(n20115), .ZN(
        P2_U3113) );
  AOI22_X1 U23140 ( .A1(n20128), .A2(n21753), .B1(n20127), .B2(n21750), .ZN(
        n20118) );
  AOI22_X1 U23141 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n21751), .ZN(n20117) );
  OAI211_X1 U23142 ( .C1(n21759), .C2(n20162), .A(n20118), .B(n20117), .ZN(
        P2_U3114) );
  AOI22_X1 U23143 ( .A1(n20128), .A2(n20278), .B1(n20127), .B2(n20377), .ZN(
        n20120) );
  AOI22_X1 U23144 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20378), .ZN(n20119) );
  OAI211_X1 U23145 ( .C1(n20321), .C2(n20162), .A(n20120), .B(n20119), .ZN(
        P2_U3115) );
  AOI22_X1 U23146 ( .A1(n20128), .A2(n20281), .B1(n20127), .B2(n20383), .ZN(
        n20122) );
  AOI22_X1 U23147 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20384), .ZN(n20121) );
  OAI211_X1 U23148 ( .C1(n20329), .C2(n20162), .A(n20122), .B(n20121), .ZN(
        P2_U3116) );
  AOI22_X1 U23149 ( .A1(n20128), .A2(n20250), .B1(n20127), .B2(n20389), .ZN(
        n20124) );
  AOI22_X1 U23150 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20390), .ZN(n20123) );
  OAI211_X1 U23151 ( .C1(n20334), .C2(n20162), .A(n20124), .B(n20123), .ZN(
        P2_U3117) );
  AOI22_X1 U23152 ( .A1(n20128), .A2(n20253), .B1(n20127), .B2(n20395), .ZN(
        n20126) );
  AOI22_X1 U23153 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20396), .ZN(n20125) );
  OAI211_X1 U23154 ( .C1(n20256), .C2(n20162), .A(n20126), .B(n20125), .ZN(
        P2_U3118) );
  AOI22_X1 U23155 ( .A1(n20128), .A2(n20257), .B1(n20127), .B2(n20401), .ZN(
        n20132) );
  AOI22_X1 U23156 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20130), .B1(
        n20129), .B2(n20403), .ZN(n20131) );
  OAI211_X1 U23157 ( .C1(n20341), .C2(n20162), .A(n20132), .B(n20131), .ZN(
        P2_U3119) );
  NOR2_X1 U23158 ( .A1(n20260), .A2(n20202), .ZN(n20173) );
  INV_X1 U23159 ( .A(n20173), .ZN(n20161) );
  OAI22_X1 U23160 ( .A1(n20172), .A2(n20297), .B1(n20161), .B2(n20296), .ZN(
        n20133) );
  INV_X1 U23161 ( .A(n20133), .ZN(n20144) );
  INV_X1 U23162 ( .A(n20139), .ZN(n20134) );
  AOI21_X1 U23163 ( .B1(n20134), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20137) );
  AOI21_X1 U23164 ( .B1(n20135), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20543), 
        .ZN(n20138) );
  NAND2_X1 U23165 ( .A1(n20138), .A2(n20141), .ZN(n20136) );
  OAI211_X1 U23166 ( .C1(n20173), .C2(n20137), .A(n20136), .B(n20361), .ZN(
        n20165) );
  INV_X1 U23167 ( .A(n20138), .ZN(n20142) );
  OAI21_X1 U23168 ( .B1(n20139), .B2(n20173), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20140) );
  AOI22_X1 U23169 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20353), .ZN(n20143) );
  OAI211_X1 U23170 ( .C1(n20366), .C2(n20162), .A(n20144), .B(n20143), .ZN(
        P2_U3120) );
  AOI22_X1 U23171 ( .A1(n20194), .A2(n20369), .B1(n20367), .B2(n20173), .ZN(
        n20146) );
  AOI22_X1 U23172 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20368), .ZN(n20145) );
  OAI211_X1 U23173 ( .C1(n20372), .C2(n20162), .A(n20146), .B(n20145), .ZN(
        P2_U3121) );
  OAI22_X1 U23174 ( .A1(n20172), .A2(n21759), .B1(n20316), .B2(n20161), .ZN(
        n20147) );
  INV_X1 U23175 ( .A(n20147), .ZN(n20149) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n21751), .ZN(n20148) );
  OAI211_X1 U23177 ( .C1(n20376), .C2(n20162), .A(n20149), .B(n20148), .ZN(
        P2_U3122) );
  OAI22_X1 U23178 ( .A1(n20162), .A2(n20382), .B1(n20161), .B2(n20320), .ZN(
        n20150) );
  INV_X1 U23179 ( .A(n20150), .ZN(n20152) );
  AOI22_X1 U23180 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20378), .ZN(n20151) );
  OAI211_X1 U23181 ( .C1(n20321), .C2(n20172), .A(n20152), .B(n20151), .ZN(
        P2_U3123) );
  OAI22_X1 U23182 ( .A1(n20162), .A2(n20388), .B1(n20161), .B2(n20325), .ZN(
        n20153) );
  INV_X1 U23183 ( .A(n20153), .ZN(n20155) );
  AOI22_X1 U23184 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20384), .ZN(n20154) );
  OAI211_X1 U23185 ( .C1(n20329), .C2(n20172), .A(n20155), .B(n20154), .ZN(
        P2_U3124) );
  OAI22_X1 U23186 ( .A1(n20172), .A2(n20334), .B1(n20330), .B2(n20161), .ZN(
        n20156) );
  INV_X1 U23187 ( .A(n20156), .ZN(n20158) );
  AOI22_X1 U23188 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20390), .ZN(n20157) );
  OAI211_X1 U23189 ( .C1(n20394), .C2(n20162), .A(n20158), .B(n20157), .ZN(
        P2_U3125) );
  AOI22_X1 U23190 ( .A1(n20194), .A2(n20397), .B1(n20395), .B2(n20173), .ZN(
        n20160) );
  AOI22_X1 U23191 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20396), .ZN(n20159) );
  OAI211_X1 U23192 ( .C1(n20400), .C2(n20162), .A(n20160), .B(n20159), .ZN(
        P2_U3126) );
  OAI22_X1 U23193 ( .A1(n20162), .A2(n20411), .B1(n20161), .B2(n20340), .ZN(
        n20163) );
  INV_X1 U23194 ( .A(n20163), .ZN(n20167) );
  AOI22_X1 U23195 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20165), .B1(
        n20164), .B2(n20403), .ZN(n20166) );
  OAI211_X1 U23196 ( .C1(n20341), .C2(n20172), .A(n20167), .B(n20166), .ZN(
        P2_U3127) );
  NOR2_X1 U23197 ( .A1(n20295), .A2(n20202), .ZN(n20192) );
  OAI21_X1 U23198 ( .B1(n11077), .B2(n20192), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20170) );
  AOI22_X1 U23199 ( .A1(n20193), .A2(n20353), .B1(n20352), .B2(n20192), .ZN(
        n20179) );
  INV_X1 U23200 ( .A(n11077), .ZN(n20176) );
  AOI21_X1 U23201 ( .B1(n20172), .B2(n20229), .A(n20356), .ZN(n20174) );
  NOR2_X1 U23202 ( .A1(n20174), .A2(n20173), .ZN(n20175) );
  AOI211_X1 U23203 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20176), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20175), .ZN(n20177) );
  OAI21_X1 U23204 ( .B1(n20177), .B2(n20192), .A(n20361), .ZN(n20195) );
  AOI22_X1 U23205 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20241), .ZN(n20178) );
  OAI211_X1 U23206 ( .C1(n20297), .C2(n20229), .A(n20179), .B(n20178), .ZN(
        P2_U3128) );
  AOI22_X1 U23207 ( .A1(n20193), .A2(n20368), .B1(n20367), .B2(n20192), .ZN(
        n20181) );
  AOI22_X1 U23208 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20273), .ZN(n20180) );
  OAI211_X1 U23209 ( .C1(n20315), .C2(n20229), .A(n20181), .B(n20180), .ZN(
        P2_U3129) );
  AOI22_X1 U23210 ( .A1(n20193), .A2(n21751), .B1(n21750), .B2(n20192), .ZN(
        n20183) );
  AOI22_X1 U23211 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n21753), .ZN(n20182) );
  OAI211_X1 U23212 ( .C1(n21759), .C2(n20229), .A(n20183), .B(n20182), .ZN(
        P2_U3130) );
  AOI22_X1 U23213 ( .A1(n20193), .A2(n20378), .B1(n20377), .B2(n20192), .ZN(
        n20185) );
  AOI22_X1 U23214 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20278), .ZN(n20184) );
  OAI211_X1 U23215 ( .C1(n20321), .C2(n20229), .A(n20185), .B(n20184), .ZN(
        P2_U3131) );
  AOI22_X1 U23216 ( .A1(n20193), .A2(n20384), .B1(n20383), .B2(n20192), .ZN(
        n20187) );
  AOI22_X1 U23217 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20281), .ZN(n20186) );
  OAI211_X1 U23218 ( .C1(n20329), .C2(n20229), .A(n20187), .B(n20186), .ZN(
        P2_U3132) );
  AOI22_X1 U23219 ( .A1(n20193), .A2(n20390), .B1(n20389), .B2(n20192), .ZN(
        n20189) );
  AOI22_X1 U23220 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20250), .ZN(n20188) );
  OAI211_X1 U23221 ( .C1(n20334), .C2(n20229), .A(n20189), .B(n20188), .ZN(
        P2_U3133) );
  AOI22_X1 U23222 ( .A1(n20193), .A2(n20396), .B1(n20395), .B2(n20192), .ZN(
        n20191) );
  AOI22_X1 U23223 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20253), .ZN(n20190) );
  OAI211_X1 U23224 ( .C1(n20256), .C2(n20229), .A(n20191), .B(n20190), .ZN(
        P2_U3134) );
  AOI22_X1 U23225 ( .A1(n20193), .A2(n20403), .B1(n20401), .B2(n20192), .ZN(
        n20197) );
  AOI22_X1 U23226 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20195), .B1(
        n20194), .B2(n20257), .ZN(n20196) );
  OAI211_X1 U23227 ( .C1(n20341), .C2(n20229), .A(n20197), .B(n20196), .ZN(
        P2_U3135) );
  NAND2_X1 U23228 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20198), .ZN(
        n20201) );
  NAND2_X1 U23229 ( .A1(n20199), .A2(n20198), .ZN(n20205) );
  OAI21_X1 U23230 ( .B1(n20204), .B2(n20224), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20200) );
  AOI22_X1 U23231 ( .A1(n20225), .A2(n20353), .B1(n20352), .B2(n20224), .ZN(
        n20211) );
  INV_X1 U23232 ( .A(n20209), .ZN(n20203) );
  OAI22_X1 U23233 ( .A1(n20203), .A2(n20356), .B1(n20202), .B2(n20521), .ZN(
        n20208) );
  INV_X1 U23234 ( .A(n20204), .ZN(n20206) );
  OAI211_X1 U23235 ( .C1(n20206), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20543), 
        .B(n20205), .ZN(n20207) );
  NAND3_X1 U23236 ( .A1(n20208), .A2(n20361), .A3(n20207), .ZN(n20226) );
  AOI22_X1 U23237 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20363), .ZN(n20210) );
  OAI211_X1 U23238 ( .C1(n20366), .C2(n20229), .A(n20211), .B(n20210), .ZN(
        P2_U3136) );
  AOI22_X1 U23239 ( .A1(n20225), .A2(n20368), .B1(n20367), .B2(n20224), .ZN(
        n20213) );
  AOI22_X1 U23240 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20369), .ZN(n20212) );
  OAI211_X1 U23241 ( .C1(n20372), .C2(n20229), .A(n20213), .B(n20212), .ZN(
        P2_U3137) );
  AOI22_X1 U23242 ( .A1(n20225), .A2(n21751), .B1(n21750), .B2(n20224), .ZN(
        n20215) );
  AOI22_X1 U23243 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20373), .ZN(n20214) );
  OAI211_X1 U23244 ( .C1(n20376), .C2(n20229), .A(n20215), .B(n20214), .ZN(
        P2_U3138) );
  AOI22_X1 U23245 ( .A1(n20225), .A2(n20378), .B1(n20377), .B2(n20224), .ZN(
        n20217) );
  AOI22_X1 U23246 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20379), .ZN(n20216) );
  OAI211_X1 U23247 ( .C1(n20382), .C2(n20229), .A(n20217), .B(n20216), .ZN(
        P2_U3139) );
  AOI22_X1 U23248 ( .A1(n20225), .A2(n20384), .B1(n20383), .B2(n20224), .ZN(
        n20219) );
  AOI22_X1 U23249 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20385), .ZN(n20218) );
  OAI211_X1 U23250 ( .C1(n20388), .C2(n20229), .A(n20219), .B(n20218), .ZN(
        P2_U3140) );
  AOI22_X1 U23251 ( .A1(n20225), .A2(n20390), .B1(n20389), .B2(n20224), .ZN(
        n20221) );
  AOI22_X1 U23252 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20391), .ZN(n20220) );
  OAI211_X1 U23253 ( .C1(n20394), .C2(n20229), .A(n20221), .B(n20220), .ZN(
        P2_U3141) );
  AOI22_X1 U23254 ( .A1(n20225), .A2(n20396), .B1(n20395), .B2(n20224), .ZN(
        n20223) );
  AOI22_X1 U23255 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20397), .ZN(n20222) );
  OAI211_X1 U23256 ( .C1(n20400), .C2(n20229), .A(n20223), .B(n20222), .ZN(
        P2_U3142) );
  AOI22_X1 U23257 ( .A1(n20225), .A2(n20403), .B1(n20401), .B2(n20224), .ZN(
        n20228) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20226), .B1(
        n21754), .B2(n20405), .ZN(n20227) );
  OAI211_X1 U23259 ( .C1(n20411), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        P2_U3143) );
  NAND2_X1 U23260 ( .A1(n20231), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20238) );
  OR2_X1 U23261 ( .A1(n20238), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20235) );
  NAND2_X1 U23262 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20350) );
  NOR3_X2 U23263 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20350), .ZN(n21749) );
  INV_X1 U23264 ( .A(n21749), .ZN(n20232) );
  NAND2_X1 U23265 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20232), .ZN(n20233) );
  NOR2_X1 U23266 ( .A1(n20234), .A2(n20233), .ZN(n20237) );
  AOI22_X1 U23267 ( .A1(n21752), .A2(n20353), .B1(n20352), .B2(n21749), .ZN(
        n20243) );
  OAI21_X1 U23268 ( .B1(n20282), .B2(n21754), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20239) );
  OAI21_X1 U23269 ( .B1(n21749), .B2(n20501), .A(n20361), .ZN(n20236) );
  AOI211_X1 U23270 ( .C1(n20239), .C2(n20238), .A(n20237), .B(n20236), .ZN(
        n20240) );
  AOI22_X1 U23271 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n21754), .B2(n20241), .ZN(n20242) );
  OAI211_X1 U23272 ( .C1(n20297), .C2(n21758), .A(n20243), .B(n20242), .ZN(
        P2_U3144) );
  AOI22_X1 U23273 ( .A1(n21752), .A2(n20368), .B1(n20367), .B2(n21749), .ZN(
        n20245) );
  AOI22_X1 U23274 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n21754), .B2(n20273), .ZN(n20244) );
  OAI211_X1 U23275 ( .C1(n20315), .C2(n21758), .A(n20245), .B(n20244), .ZN(
        P2_U3145) );
  AOI22_X1 U23276 ( .A1(n21752), .A2(n20378), .B1(n20377), .B2(n21749), .ZN(
        n20247) );
  AOI22_X1 U23277 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n21754), .B2(n20278), .ZN(n20246) );
  OAI211_X1 U23278 ( .C1(n20321), .C2(n21758), .A(n20247), .B(n20246), .ZN(
        P2_U3147) );
  AOI22_X1 U23279 ( .A1(n21752), .A2(n20384), .B1(n20383), .B2(n21749), .ZN(
        n20249) );
  AOI22_X1 U23280 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n21754), .B2(n20281), .ZN(n20248) );
  OAI211_X1 U23281 ( .C1(n20329), .C2(n21758), .A(n20249), .B(n20248), .ZN(
        P2_U3148) );
  AOI22_X1 U23282 ( .A1(n21752), .A2(n20390), .B1(n20389), .B2(n21749), .ZN(
        n20252) );
  AOI22_X1 U23283 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n21754), .B2(n20250), .ZN(n20251) );
  OAI211_X1 U23284 ( .C1(n20334), .C2(n21758), .A(n20252), .B(n20251), .ZN(
        P2_U3149) );
  AOI22_X1 U23285 ( .A1(n21752), .A2(n20396), .B1(n20395), .B2(n21749), .ZN(
        n20255) );
  AOI22_X1 U23286 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n21754), .B2(n20253), .ZN(n20254) );
  OAI211_X1 U23287 ( .C1(n20256), .C2(n21758), .A(n20255), .B(n20254), .ZN(
        P2_U3150) );
  AOI22_X1 U23288 ( .A1(n21752), .A2(n20403), .B1(n20401), .B2(n21749), .ZN(
        n20259) );
  AOI22_X1 U23289 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n21754), .B2(n20257), .ZN(n20258) );
  OAI211_X1 U23290 ( .C1(n20341), .C2(n21758), .A(n20259), .B(n20258), .ZN(
        P2_U3151) );
  NOR2_X1 U23291 ( .A1(n20350), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20268) );
  INV_X1 U23292 ( .A(n20268), .ZN(n20263) );
  NOR2_X1 U23293 ( .A1(n20260), .A2(n20350), .ZN(n20289) );
  NOR3_X1 U23294 ( .A1(n20261), .A2(n20289), .A3(n20552), .ZN(n20264) );
  AOI211_X2 U23295 ( .C1(n20263), .C2(n20552), .A(n20262), .B(n20264), .ZN(
        n20290) );
  AOI22_X1 U23296 ( .A1(n20290), .A2(n20353), .B1(n20352), .B2(n20289), .ZN(
        n20272) );
  INV_X1 U23297 ( .A(n20289), .ZN(n20266) );
  AOI211_X1 U23298 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20266), .A(n20265), 
        .B(n20264), .ZN(n20267) );
  OAI221_X1 U23299 ( .B1(n20268), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20268), 
        .C2(n20270), .A(n20267), .ZN(n20292) );
  INV_X1 U23300 ( .A(n20347), .ZN(n20291) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20292), .B1(
        n20291), .B2(n20363), .ZN(n20271) );
  OAI211_X1 U23302 ( .C1(n20366), .C2(n21758), .A(n20272), .B(n20271), .ZN(
        P2_U3152) );
  AOI22_X1 U23303 ( .A1(n20290), .A2(n20368), .B1(n20367), .B2(n20289), .ZN(
        n20275) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20292), .B1(
        n20282), .B2(n20273), .ZN(n20274) );
  OAI211_X1 U23305 ( .C1(n20315), .C2(n20347), .A(n20275), .B(n20274), .ZN(
        P2_U3153) );
  AOI22_X1 U23306 ( .A1(n20290), .A2(n21751), .B1(n21750), .B2(n20289), .ZN(
        n20277) );
  AOI22_X1 U23307 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20292), .B1(
        n20291), .B2(n20373), .ZN(n20276) );
  OAI211_X1 U23308 ( .C1(n20376), .C2(n21758), .A(n20277), .B(n20276), .ZN(
        P2_U3154) );
  AOI22_X1 U23309 ( .A1(n20290), .A2(n20378), .B1(n20377), .B2(n20289), .ZN(
        n20280) );
  AOI22_X1 U23310 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20292), .B1(
        n20282), .B2(n20278), .ZN(n20279) );
  OAI211_X1 U23311 ( .C1(n20321), .C2(n20347), .A(n20280), .B(n20279), .ZN(
        P2_U3155) );
  AOI22_X1 U23312 ( .A1(n20290), .A2(n20384), .B1(n20383), .B2(n20289), .ZN(
        n20284) );
  AOI22_X1 U23313 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20292), .B1(
        n20282), .B2(n20281), .ZN(n20283) );
  OAI211_X1 U23314 ( .C1(n20329), .C2(n20347), .A(n20284), .B(n20283), .ZN(
        P2_U3156) );
  AOI22_X1 U23315 ( .A1(n20290), .A2(n20390), .B1(n20389), .B2(n20289), .ZN(
        n20286) );
  AOI22_X1 U23316 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20292), .B1(
        n20291), .B2(n20391), .ZN(n20285) );
  OAI211_X1 U23317 ( .C1(n20394), .C2(n21758), .A(n20286), .B(n20285), .ZN(
        P2_U3157) );
  AOI22_X1 U23318 ( .A1(n20290), .A2(n20396), .B1(n20395), .B2(n20289), .ZN(
        n20288) );
  AOI22_X1 U23319 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20292), .B1(
        n20291), .B2(n20397), .ZN(n20287) );
  OAI211_X1 U23320 ( .C1(n20400), .C2(n21758), .A(n20288), .B(n20287), .ZN(
        P2_U3158) );
  AOI22_X1 U23321 ( .A1(n20290), .A2(n20403), .B1(n20401), .B2(n20289), .ZN(
        n20294) );
  AOI22_X1 U23322 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20292), .B1(
        n20291), .B2(n20405), .ZN(n20293) );
  OAI211_X1 U23323 ( .C1(n20411), .C2(n21758), .A(n20294), .B(n20293), .ZN(
        P2_U3159) );
  NAND2_X2 U23324 ( .A1(n20354), .A2(n20526), .ZN(n20410) );
  NOR2_X1 U23325 ( .A1(n20295), .A2(n20350), .ZN(n20335) );
  INV_X1 U23326 ( .A(n20335), .ZN(n20339) );
  OAI22_X1 U23327 ( .A1(n20410), .A2(n20297), .B1(n20339), .B2(n20296), .ZN(
        n20298) );
  INV_X1 U23328 ( .A(n20298), .ZN(n20310) );
  INV_X1 U23329 ( .A(n11052), .ZN(n20299) );
  AOI21_X1 U23330 ( .B1(n20299), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20304) );
  AOI21_X1 U23331 ( .B1(n20347), .B2(n20410), .A(n20356), .ZN(n20300) );
  NOR2_X1 U23332 ( .A1(n20300), .A2(n20543), .ZN(n20305) );
  INV_X1 U23333 ( .A(n20350), .ZN(n20301) );
  NAND2_X1 U23334 ( .A1(n20302), .A2(n20301), .ZN(n20307) );
  NAND2_X1 U23335 ( .A1(n20305), .A2(n20307), .ZN(n20303) );
  OAI211_X1 U23336 ( .C1(n20335), .C2(n20304), .A(n20303), .B(n20361), .ZN(
        n20344) );
  INV_X1 U23337 ( .A(n20305), .ZN(n20308) );
  OAI21_X1 U23338 ( .B1(n11052), .B2(n20335), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20306) );
  AOI22_X1 U23339 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20344), .B1(
        n20353), .B2(n20343), .ZN(n20309) );
  OAI211_X1 U23340 ( .C1(n20366), .C2(n20347), .A(n20310), .B(n20309), .ZN(
        P2_U3160) );
  OAI22_X1 U23341 ( .A1(n20347), .A2(n20372), .B1(n20339), .B2(n20311), .ZN(
        n20312) );
  INV_X1 U23342 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U23343 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20344), .B1(
        n20368), .B2(n20343), .ZN(n20313) );
  OAI211_X1 U23344 ( .C1(n20315), .C2(n20410), .A(n20314), .B(n20313), .ZN(
        P2_U3161) );
  OAI22_X1 U23345 ( .A1(n20410), .A2(n21759), .B1(n20316), .B2(n20339), .ZN(
        n20317) );
  INV_X1 U23346 ( .A(n20317), .ZN(n20319) );
  AOI22_X1 U23347 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20344), .B1(
        n21751), .B2(n20343), .ZN(n20318) );
  OAI211_X1 U23348 ( .C1(n20376), .C2(n20347), .A(n20319), .B(n20318), .ZN(
        P2_U3162) );
  OAI22_X1 U23349 ( .A1(n20410), .A2(n20321), .B1(n20320), .B2(n20339), .ZN(
        n20322) );
  INV_X1 U23350 ( .A(n20322), .ZN(n20324) );
  AOI22_X1 U23351 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20344), .B1(
        n20378), .B2(n20343), .ZN(n20323) );
  OAI211_X1 U23352 ( .C1(n20382), .C2(n20347), .A(n20324), .B(n20323), .ZN(
        P2_U3163) );
  OAI22_X1 U23353 ( .A1(n20347), .A2(n20388), .B1(n20339), .B2(n20325), .ZN(
        n20326) );
  INV_X1 U23354 ( .A(n20326), .ZN(n20328) );
  AOI22_X1 U23355 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20344), .B1(
        n20384), .B2(n20343), .ZN(n20327) );
  OAI211_X1 U23356 ( .C1(n20329), .C2(n20410), .A(n20328), .B(n20327), .ZN(
        P2_U3164) );
  OAI22_X1 U23357 ( .A1(n20347), .A2(n20394), .B1(n20339), .B2(n20330), .ZN(
        n20331) );
  INV_X1 U23358 ( .A(n20331), .ZN(n20333) );
  AOI22_X1 U23359 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20344), .B1(
        n20390), .B2(n20343), .ZN(n20332) );
  OAI211_X1 U23360 ( .C1(n20334), .C2(n20410), .A(n20333), .B(n20332), .ZN(
        P2_U3165) );
  INV_X1 U23361 ( .A(n20410), .ZN(n20336) );
  AOI22_X1 U23362 ( .A1(n20336), .A2(n20397), .B1(n20395), .B2(n20335), .ZN(
        n20338) );
  AOI22_X1 U23363 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20344), .B1(
        n20396), .B2(n20343), .ZN(n20337) );
  OAI211_X1 U23364 ( .C1(n20400), .C2(n20347), .A(n20338), .B(n20337), .ZN(
        P2_U3166) );
  OAI22_X1 U23365 ( .A1(n20410), .A2(n20341), .B1(n20340), .B2(n20339), .ZN(
        n20342) );
  INV_X1 U23366 ( .A(n20342), .ZN(n20346) );
  AOI22_X1 U23367 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20344), .B1(
        n20403), .B2(n20343), .ZN(n20345) );
  OAI211_X1 U23368 ( .C1(n20411), .C2(n20347), .A(n20346), .B(n20345), .ZN(
        P2_U3167) );
  NAND2_X1 U23369 ( .A1(n20358), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20348) );
  OR2_X1 U23370 ( .A1(n20521), .A2(n20350), .ZN(n20355) );
  OAI21_X1 U23371 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20355), .A(n20552), 
        .ZN(n20351) );
  AOI22_X1 U23372 ( .A1(n20404), .A2(n20353), .B1(n20402), .B2(n20352), .ZN(
        n20365) );
  INV_X1 U23373 ( .A(n20354), .ZN(n20357) );
  OAI21_X1 U23374 ( .B1(n20357), .B2(n20356), .A(n20355), .ZN(n20362) );
  NAND2_X1 U23375 ( .A1(n20358), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20359) );
  NAND4_X1 U23376 ( .A1(n20362), .A2(n20361), .A3(n20360), .A4(n20359), .ZN(
        n20407) );
  AOI22_X1 U23377 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20406), .B2(n20363), .ZN(n20364) );
  OAI211_X1 U23378 ( .C1(n20366), .C2(n20410), .A(n20365), .B(n20364), .ZN(
        P2_U3168) );
  AOI22_X1 U23379 ( .A1(n20404), .A2(n20368), .B1(n20402), .B2(n20367), .ZN(
        n20371) );
  AOI22_X1 U23380 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20406), .B2(n20369), .ZN(n20370) );
  OAI211_X1 U23381 ( .C1(n20372), .C2(n20410), .A(n20371), .B(n20370), .ZN(
        P2_U3169) );
  AOI22_X1 U23382 ( .A1(n20404), .A2(n21751), .B1(n20402), .B2(n21750), .ZN(
        n20375) );
  AOI22_X1 U23383 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20406), .B2(n20373), .ZN(n20374) );
  OAI211_X1 U23384 ( .C1(n20376), .C2(n20410), .A(n20375), .B(n20374), .ZN(
        P2_U3170) );
  AOI22_X1 U23385 ( .A1(n20404), .A2(n20378), .B1(n20402), .B2(n20377), .ZN(
        n20381) );
  AOI22_X1 U23386 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20406), .B2(n20379), .ZN(n20380) );
  OAI211_X1 U23387 ( .C1(n20382), .C2(n20410), .A(n20381), .B(n20380), .ZN(
        P2_U3171) );
  AOI22_X1 U23388 ( .A1(n20404), .A2(n20384), .B1(n20402), .B2(n20383), .ZN(
        n20387) );
  AOI22_X1 U23389 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20406), .B2(n20385), .ZN(n20386) );
  OAI211_X1 U23390 ( .C1(n20388), .C2(n20410), .A(n20387), .B(n20386), .ZN(
        P2_U3172) );
  AOI22_X1 U23391 ( .A1(n20404), .A2(n20390), .B1(n20402), .B2(n20389), .ZN(
        n20393) );
  AOI22_X1 U23392 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n20406), .B2(n20391), .ZN(n20392) );
  OAI211_X1 U23393 ( .C1(n20394), .C2(n20410), .A(n20393), .B(n20392), .ZN(
        P2_U3173) );
  AOI22_X1 U23394 ( .A1(n20404), .A2(n20396), .B1(n20402), .B2(n20395), .ZN(
        n20399) );
  AOI22_X1 U23395 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n20406), .B2(n20397), .ZN(n20398) );
  OAI211_X1 U23396 ( .C1(n20400), .C2(n20410), .A(n20399), .B(n20398), .ZN(
        P2_U3174) );
  AOI22_X1 U23397 ( .A1(n20404), .A2(n20403), .B1(n20402), .B2(n20401), .ZN(
        n20409) );
  AOI22_X1 U23398 ( .A1(n20407), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n20406), .B2(n20405), .ZN(n20408) );
  OAI211_X1 U23399 ( .C1(n20411), .C2(n20410), .A(n20409), .B(n20408), .ZN(
        P2_U3175) );
  AND2_X1 U23400 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20412), .ZN(
        P2_U3179) );
  AND2_X1 U23401 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20412), .ZN(
        P2_U3180) );
  AND2_X1 U23402 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20412), .ZN(
        P2_U3181) );
  INV_X1 U23403 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21721) );
  NOR2_X1 U23404 ( .A1(n21721), .A2(n20491), .ZN(P2_U3182) );
  AND2_X1 U23405 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20412), .ZN(
        P2_U3183) );
  AND2_X1 U23406 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20412), .ZN(
        P2_U3184) );
  AND2_X1 U23407 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20412), .ZN(
        P2_U3185) );
  AND2_X1 U23408 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20412), .ZN(
        P2_U3186) );
  AND2_X1 U23409 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20412), .ZN(
        P2_U3187) );
  AND2_X1 U23410 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20412), .ZN(
        P2_U3188) );
  AND2_X1 U23411 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20412), .ZN(
        P2_U3189) );
  AND2_X1 U23412 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20412), .ZN(
        P2_U3190) );
  AND2_X1 U23413 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20412), .ZN(
        P2_U3191) );
  AND2_X1 U23414 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20412), .ZN(
        P2_U3192) );
  AND2_X1 U23415 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20412), .ZN(
        P2_U3193) );
  AND2_X1 U23416 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20412), .ZN(
        P2_U3194) );
  AND2_X1 U23417 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20412), .ZN(
        P2_U3195) );
  AND2_X1 U23418 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20412), .ZN(
        P2_U3196) );
  AND2_X1 U23419 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20412), .ZN(
        P2_U3197) );
  AND2_X1 U23420 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20412), .ZN(
        P2_U3198) );
  AND2_X1 U23421 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20412), .ZN(
        P2_U3199) );
  AND2_X1 U23422 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20412), .ZN(
        P2_U3200) );
  AND2_X1 U23423 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20412), .ZN(P2_U3201) );
  AND2_X1 U23424 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20412), .ZN(P2_U3202) );
  AND2_X1 U23425 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20412), .ZN(P2_U3203) );
  AND2_X1 U23426 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20412), .ZN(P2_U3204) );
  AND2_X1 U23427 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20412), .ZN(P2_U3205) );
  AND2_X1 U23428 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20412), .ZN(P2_U3206) );
  AND2_X1 U23429 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20412), .ZN(P2_U3207) );
  AND2_X1 U23430 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20412), .ZN(P2_U3208) );
  AND2_X1 U23431 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20553), .ZN(n20424) );
  INV_X1 U23432 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20565) );
  NOR3_X1 U23433 ( .A1(n20424), .A2(n20565), .A3(n20413), .ZN(n20416) );
  OAI211_X1 U23434 ( .C1(HOLD), .C2(n20565), .A(n20566), .B(n20414), .ZN(
        n20415) );
  NAND2_X1 U23435 ( .A1(NA), .A2(n20417), .ZN(n20422) );
  OAI211_X1 U23436 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20416), .A(n20415), 
        .B(n20422), .ZN(P2_U3209) );
  NAND2_X1 U23437 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21512), .ZN(n20423) );
  OAI21_X1 U23438 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20417), .A(n20423), 
        .ZN(n20418) );
  AOI211_X1 U23439 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20418), .A(
        n20560), .B(n20424), .ZN(n20419) );
  OAI21_X1 U23440 ( .B1(n21512), .B2(n20420), .A(n20419), .ZN(P2_U3210) );
  INV_X1 U23441 ( .A(NA), .ZN(n21517) );
  AOI22_X1 U23442 ( .A1(n20421), .A2(n20565), .B1(n20424), .B2(n21517), .ZN(
        n20427) );
  OAI21_X1 U23443 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20426) );
  OAI211_X1 U23444 ( .C1(n20424), .C2(n20423), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n20422), .ZN(n20425) );
  OAI21_X1 U23445 ( .B1(n20427), .B2(n20426), .A(n20425), .ZN(P2_U3211) );
  NAND2_X2 U23446 ( .A1(n20533), .A2(n20428), .ZN(n20484) );
  OAI222_X1 U23447 ( .A1(n20484), .A2(n20431), .B1(n20430), .B2(n20533), .C1(
        n20429), .C2(n20477), .ZN(P2_U3212) );
  OAI222_X1 U23448 ( .A1(n20484), .A2(n10136), .B1(n20432), .B2(n20533), .C1(
        n20431), .C2(n20477), .ZN(P2_U3213) );
  OAI222_X1 U23449 ( .A1(n20484), .A2(n20434), .B1(n20433), .B2(n20533), .C1(
        n10136), .C2(n20477), .ZN(P2_U3214) );
  INV_X1 U23450 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20436) );
  OAI222_X1 U23451 ( .A1(n20484), .A2(n20436), .B1(n20435), .B2(n20533), .C1(
        n20434), .C2(n20477), .ZN(P2_U3215) );
  OAI222_X1 U23452 ( .A1(n20484), .A2(n20438), .B1(n20437), .B2(n20533), .C1(
        n20436), .C2(n20477), .ZN(P2_U3216) );
  OAI222_X1 U23453 ( .A1(n20484), .A2(n20440), .B1(n20439), .B2(n20533), .C1(
        n20438), .C2(n20477), .ZN(P2_U3217) );
  OAI222_X1 U23454 ( .A1(n20484), .A2(n20442), .B1(n20441), .B2(n20533), .C1(
        n20440), .C2(n20477), .ZN(P2_U3218) );
  OAI222_X1 U23455 ( .A1(n20484), .A2(n20444), .B1(n20443), .B2(n20533), .C1(
        n20442), .C2(n20477), .ZN(P2_U3219) );
  OAI222_X1 U23456 ( .A1(n20484), .A2(n20446), .B1(n20445), .B2(n20533), .C1(
        n20444), .C2(n20477), .ZN(P2_U3220) );
  OAI222_X1 U23457 ( .A1(n20484), .A2(n20447), .B1(n21626), .B2(n20533), .C1(
        n20446), .C2(n20477), .ZN(P2_U3221) );
  OAI222_X1 U23458 ( .A1(n20484), .A2(n20449), .B1(n20448), .B2(n20533), .C1(
        n20447), .C2(n20477), .ZN(P2_U3222) );
  INV_X1 U23459 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20451) );
  OAI222_X1 U23460 ( .A1(n20484), .A2(n20451), .B1(n20450), .B2(n20533), .C1(
        n20449), .C2(n20477), .ZN(P2_U3223) );
  OAI222_X1 U23461 ( .A1(n20484), .A2(n20453), .B1(n20452), .B2(n20533), .C1(
        n20451), .C2(n20477), .ZN(P2_U3224) );
  OAI222_X1 U23462 ( .A1(n20484), .A2(n20455), .B1(n20454), .B2(n20533), .C1(
        n20453), .C2(n20477), .ZN(P2_U3225) );
  OAI222_X1 U23463 ( .A1(n20484), .A2(n20457), .B1(n20456), .B2(n20533), .C1(
        n20455), .C2(n20477), .ZN(P2_U3226) );
  OAI222_X1 U23464 ( .A1(n20484), .A2(n20459), .B1(n20458), .B2(n20533), .C1(
        n20457), .C2(n20477), .ZN(P2_U3227) );
  OAI222_X1 U23465 ( .A1(n20484), .A2(n12853), .B1(n20460), .B2(n20533), .C1(
        n20459), .C2(n20477), .ZN(P2_U3228) );
  OAI222_X1 U23466 ( .A1(n20484), .A2(n21594), .B1(n20461), .B2(n20533), .C1(
        n12853), .C2(n20477), .ZN(P2_U3229) );
  OAI222_X1 U23467 ( .A1(n20484), .A2(n12863), .B1(n20462), .B2(n20533), .C1(
        n21594), .C2(n20477), .ZN(P2_U3230) );
  OAI222_X1 U23468 ( .A1(n20484), .A2(n20464), .B1(n20463), .B2(n20533), .C1(
        n12863), .C2(n20477), .ZN(P2_U3231) );
  OAI222_X1 U23469 ( .A1(n20484), .A2(n20466), .B1(n20465), .B2(n20533), .C1(
        n20464), .C2(n20477), .ZN(P2_U3232) );
  OAI222_X1 U23470 ( .A1(n20484), .A2(n20468), .B1(n20467), .B2(n20533), .C1(
        n20466), .C2(n20477), .ZN(P2_U3233) );
  OAI222_X1 U23471 ( .A1(n20484), .A2(n16477), .B1(n20469), .B2(n20533), .C1(
        n20468), .C2(n20477), .ZN(P2_U3234) );
  OAI222_X1 U23472 ( .A1(n20484), .A2(n20471), .B1(n20470), .B2(n20533), .C1(
        n16477), .C2(n20477), .ZN(P2_U3235) );
  OAI222_X1 U23473 ( .A1(n20484), .A2(n20473), .B1(n20472), .B2(n20533), .C1(
        n20471), .C2(n20477), .ZN(P2_U3236) );
  OAI222_X1 U23474 ( .A1(n20484), .A2(n20476), .B1(n20474), .B2(n20533), .C1(
        n20473), .C2(n20477), .ZN(P2_U3237) );
  OAI222_X1 U23475 ( .A1(n20477), .A2(n20476), .B1(n20475), .B2(n20533), .C1(
        n16444), .C2(n20484), .ZN(P2_U3238) );
  OAI222_X1 U23476 ( .A1(n20484), .A2(n20479), .B1(n20478), .B2(n20533), .C1(
        n16444), .C2(n20477), .ZN(P2_U3239) );
  INV_X1 U23477 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20481) );
  OAI222_X1 U23478 ( .A1(n20484), .A2(n20481), .B1(n20480), .B2(n20533), .C1(
        n20479), .C2(n20477), .ZN(P2_U3240) );
  OAI222_X1 U23479 ( .A1(n20484), .A2(n20483), .B1(n20482), .B2(n20533), .C1(
        n20481), .C2(n20477), .ZN(P2_U3241) );
  OAI22_X1 U23480 ( .A1(n20566), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20533), .ZN(n20485) );
  INV_X1 U23481 ( .A(n20485), .ZN(P2_U3585) );
  MUX2_X1 U23482 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20566), .Z(P2_U3586) );
  OAI22_X1 U23483 ( .A1(n20566), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20533), .ZN(n20486) );
  INV_X1 U23484 ( .A(n20486), .ZN(P2_U3587) );
  OAI22_X1 U23485 ( .A1(n20566), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20533), .ZN(n20487) );
  INV_X1 U23486 ( .A(n20487), .ZN(P2_U3588) );
  OAI21_X1 U23487 ( .B1(n20491), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20489), 
        .ZN(n20488) );
  INV_X1 U23488 ( .A(n20488), .ZN(P2_U3591) );
  OAI21_X1 U23489 ( .B1(n20491), .B2(n20490), .A(n20489), .ZN(P2_U3592) );
  INV_X1 U23490 ( .A(n20530), .ZN(n20529) );
  NAND2_X1 U23491 ( .A1(n20492), .A2(n20514), .ZN(n20500) );
  INV_X1 U23492 ( .A(n20514), .ZN(n20496) );
  NAND3_X1 U23493 ( .A1(n20494), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20493), 
        .ZN(n20495) );
  NAND2_X1 U23494 ( .A1(n20495), .A2(n20515), .ZN(n20506) );
  OAI21_X1 U23495 ( .B1(n20508), .B2(n20496), .A(n20506), .ZN(n20497) );
  NAND2_X1 U23496 ( .A1(n20498), .A2(n20497), .ZN(n20499) );
  OAI211_X1 U23497 ( .C1(n20502), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        n20503) );
  INV_X1 U23498 ( .A(n20503), .ZN(n20504) );
  AOI22_X1 U23499 ( .A1(n20529), .A2(n20505), .B1(n20504), .B2(n20530), .ZN(
        P2_U3602) );
  INV_X1 U23500 ( .A(n20506), .ZN(n20507) );
  AOI222_X1 U23501 ( .A1(n20510), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n20509), 
        .B2(n20514), .C1(n20508), .C2(n20507), .ZN(n20511) );
  AOI22_X1 U23502 ( .A1(n20529), .A2(n20512), .B1(n20511), .B2(n20530), .ZN(
        P2_U3603) );
  AOI22_X1 U23503 ( .A1(n20517), .A2(n20514), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20513), .ZN(n20520) );
  INV_X1 U23504 ( .A(n20515), .ZN(n20525) );
  NOR3_X1 U23505 ( .A1(n20517), .A2(n20525), .A3(n20516), .ZN(n20518) );
  NOR2_X1 U23506 ( .A1(n20529), .A2(n20518), .ZN(n20519) );
  AOI22_X1 U23507 ( .A1(n20521), .A2(n20529), .B1(n20520), .B2(n20519), .ZN(
        P2_U3604) );
  INV_X1 U23508 ( .A(n20522), .ZN(n20523) );
  OAI22_X1 U23509 ( .A1(n20526), .A2(n20525), .B1(n20524), .B2(n20523), .ZN(
        n20527) );
  AOI21_X1 U23510 ( .B1(n20531), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20527), 
        .ZN(n20528) );
  OAI22_X1 U23511 ( .A1(n20531), .A2(n20530), .B1(n20529), .B2(n20528), .ZN(
        P2_U3605) );
  INV_X1 U23512 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20532) );
  AOI22_X1 U23513 ( .A1(n20533), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20532), 
        .B2(n20566), .ZN(P2_U3608) );
  INV_X1 U23514 ( .A(n20534), .ZN(n20535) );
  AOI22_X1 U23515 ( .A1(n20538), .A2(n20537), .B1(n20536), .B2(n20535), .ZN(
        n20539) );
  NAND2_X1 U23516 ( .A1(n20540), .A2(n20539), .ZN(n20542) );
  MUX2_X1 U23517 ( .A(P2_MORE_REG_SCAN_IN), .B(n20542), .S(n20541), .Z(
        P2_U3609) );
  OAI21_X1 U23518 ( .B1(n20544), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20543), 
        .ZN(n20546) );
  AOI211_X1 U23519 ( .C1(n20548), .C2(n20547), .A(n20546), .B(n20545), .ZN(
        n20564) );
  NAND3_X1 U23520 ( .A1(n20550), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20549), 
        .ZN(n20555) );
  OAI21_X1 U23521 ( .B1(n20553), .B2(n20552), .A(n20551), .ZN(n20554) );
  OAI21_X1 U23522 ( .B1(n20560), .B2(n20555), .A(n20554), .ZN(n20556) );
  INV_X1 U23523 ( .A(n20556), .ZN(n20563) );
  INV_X1 U23524 ( .A(n20557), .ZN(n20558) );
  AOI211_X1 U23525 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n20560), .A(n20559), 
        .B(n20558), .ZN(n20561) );
  NOR2_X1 U23526 ( .A1(n20564), .A2(n20561), .ZN(n20562) );
  AOI22_X1 U23527 ( .A1(n20565), .A2(n20564), .B1(n20563), .B2(n20562), .ZN(
        P2_U3610) );
  MUX2_X1 U23528 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n20566), .Z(P2_U3611) );
  AOI21_X1 U23529 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21520), .A(n21511), 
        .ZN(n21513) );
  INV_X1 U23530 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20567) );
  AOI21_X1 U23531 ( .B1(n21513), .B2(n20567), .A(n21579), .ZN(P1_U2802) );
  OAI21_X1 U23532 ( .B1(n20569), .B2(n20568), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20570) );
  OAI21_X1 U23533 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20571), .A(n20570), 
        .ZN(P1_U2803) );
  NOR2_X1 U23534 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20573) );
  OAI21_X1 U23535 ( .B1(n20573), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21577), .ZN(
        n20572) );
  OAI21_X1 U23536 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21577), .A(n20572), 
        .ZN(P1_U2804) );
  NOR2_X1 U23537 ( .A1(n21513), .A2(n21579), .ZN(n21569) );
  OAI21_X1 U23538 ( .B1(BS16), .B2(n20573), .A(n21569), .ZN(n21567) );
  OAI21_X1 U23539 ( .B1(n21569), .B2(n21373), .A(n21567), .ZN(P1_U2805) );
  OAI21_X1 U23540 ( .B1(n20576), .B2(n20575), .A(n20574), .ZN(P1_U2806) );
  NOR4_X1 U23541 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20580) );
  NOR4_X1 U23542 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20579) );
  NOR4_X1 U23543 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20578) );
  NOR4_X1 U23544 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20577) );
  NAND4_X1 U23545 ( .A1(n20580), .A2(n20579), .A3(n20578), .A4(n20577), .ZN(
        n20586) );
  NOR4_X1 U23546 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20584) );
  AOI211_X1 U23547 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20583) );
  NOR4_X1 U23548 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20582) );
  NOR4_X1 U23549 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20581) );
  NAND4_X1 U23550 ( .A1(n20584), .A2(n20583), .A3(n20582), .A4(n20581), .ZN(
        n20585) );
  NOR2_X1 U23551 ( .A1(n20586), .A2(n20585), .ZN(n21576) );
  INV_X1 U23552 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20588) );
  NOR3_X1 U23553 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20589) );
  OAI21_X1 U23554 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20589), .A(n21576), .ZN(
        n20587) );
  OAI21_X1 U23555 ( .B1(n21576), .B2(n20588), .A(n20587), .ZN(P1_U2807) );
  INV_X1 U23556 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21568) );
  AOI21_X1 U23557 ( .B1(n21571), .B2(n21568), .A(n20589), .ZN(n20591) );
  INV_X1 U23558 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20590) );
  INV_X1 U23559 ( .A(n21576), .ZN(n21573) );
  AOI22_X1 U23560 ( .A1(n21576), .A2(n20591), .B1(n20590), .B2(n21573), .ZN(
        P1_U2808) );
  NAND2_X1 U23561 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20601) );
  OR2_X1 U23562 ( .A1(n20593), .A2(n20592), .ZN(n20595) );
  NAND2_X1 U23563 ( .A1(n20595), .A2(n20594), .ZN(n20616) );
  AOI21_X1 U23564 ( .B1(n20596), .B2(n20601), .A(n20616), .ZN(n20617) );
  INV_X1 U23565 ( .A(n20597), .ZN(n20599) );
  INV_X1 U23566 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20598) );
  OAI22_X1 U23567 ( .A1(n20599), .A2(n20615), .B1(n20627), .B2(n20598), .ZN(
        n20600) );
  AOI211_X1 U23568 ( .C1(n20611), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20629), .B(n20600), .ZN(n20608) );
  NOR4_X1 U23569 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20631), .A3(n20601), .A4(
        n20637), .ZN(n20606) );
  OAI22_X1 U23570 ( .A1(n20604), .A2(n20603), .B1(n20602), .B2(n20649), .ZN(
        n20605) );
  NOR2_X1 U23571 ( .A1(n20606), .A2(n20605), .ZN(n20607) );
  OAI211_X1 U23572 ( .C1(n20617), .C2(n20609), .A(n20608), .B(n20607), .ZN(
        P1_U2833) );
  INV_X1 U23573 ( .A(n20610), .ZN(n20621) );
  AOI21_X1 U23574 ( .B1(n20611), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20629), .ZN(n20613) );
  NAND2_X1 U23575 ( .A1(n14862), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n20612) );
  OAI211_X1 U23576 ( .C1(n20615), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        n20619) );
  INV_X1 U23577 ( .A(n20616), .ZN(n20645) );
  NAND2_X1 U23578 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20645), .ZN(n20632) );
  AOI21_X1 U23579 ( .B1(n15267), .B2(n20632), .A(n20617), .ZN(n20618) );
  AOI211_X1 U23580 ( .C1(n20621), .C2(n20620), .A(n20619), .B(n20618), .ZN(
        n20622) );
  OAI21_X1 U23581 ( .B1(n20623), .B2(n20649), .A(n20622), .ZN(P1_U2834) );
  INV_X1 U23582 ( .A(n20624), .ZN(n20657) );
  INV_X1 U23583 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20626) );
  OAI22_X1 U23584 ( .A1(n20627), .A2(n20626), .B1(n20625), .B2(n20655), .ZN(
        n20628) );
  AOI211_X1 U23585 ( .C1(n20647), .C2(n20657), .A(n20629), .B(n20628), .ZN(
        n20635) );
  INV_X1 U23586 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20630) );
  OAI21_X1 U23587 ( .B1(n20631), .B2(n20637), .A(n20630), .ZN(n20633) );
  AOI22_X1 U23588 ( .A1(n20633), .A2(n20632), .B1(n20660), .B2(n20652), .ZN(
        n20634) );
  OAI211_X1 U23589 ( .C1(n20636), .C2(n20649), .A(n20635), .B(n20634), .ZN(
        P1_U2835) );
  NOR3_X1 U23590 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20638), .A3(n20637), .ZN(
        n20644) );
  NAND2_X1 U23591 ( .A1(n20640), .A2(n20639), .ZN(n20642) );
  NAND2_X1 U23592 ( .A1(n20642), .A2(n20641), .ZN(n20643) );
  NOR2_X1 U23593 ( .A1(n20644), .A2(n20643), .ZN(n20654) );
  INV_X1 U23594 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21523) );
  NOR2_X1 U23595 ( .A1(n20645), .A2(n21523), .ZN(n20651) );
  AOI22_X1 U23596 ( .A1(n20647), .A2(n20646), .B1(n14862), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n20648) );
  OAI21_X1 U23597 ( .B1(n20649), .B2(n20741), .A(n20648), .ZN(n20650) );
  AOI211_X1 U23598 ( .C1(n20736), .C2(n20652), .A(n20651), .B(n20650), .ZN(
        n20653) );
  OAI211_X1 U23599 ( .C1(n20656), .C2(n20655), .A(n20654), .B(n20653), .ZN(
        P1_U2836) );
  AOI22_X1 U23600 ( .A1(n20660), .A2(n20659), .B1(n20658), .B2(n20657), .ZN(
        n20661) );
  OAI21_X1 U23601 ( .B1(n20662), .B2(n20626), .A(n20661), .ZN(P1_U2867) );
  INV_X1 U23602 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n21649) );
  INV_X1 U23603 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23604 ( .A1(n20665), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20688), .ZN(n20664) );
  OAI21_X1 U23605 ( .B1(n21649), .B2(n20667), .A(n20664), .ZN(P1_U2911) );
  INV_X1 U23606 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n21624) );
  AOI22_X1 U23607 ( .A1(n20665), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20688), .ZN(n20666) );
  OAI21_X1 U23608 ( .B1(n21624), .B2(n20667), .A(n20666), .ZN(P1_U2912) );
  AOI22_X1 U23609 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20668) );
  OAI21_X1 U23610 ( .B1(n20669), .B2(n20695), .A(n20668), .ZN(P1_U2921) );
  AOI22_X1 U23611 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20670) );
  OAI21_X1 U23612 ( .B1(n15020), .B2(n20695), .A(n20670), .ZN(P1_U2922) );
  AOI22_X1 U23613 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20671) );
  OAI21_X1 U23614 ( .B1(n15022), .B2(n20695), .A(n20671), .ZN(P1_U2923) );
  AOI22_X1 U23615 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20672) );
  OAI21_X1 U23616 ( .B1(n15024), .B2(n20695), .A(n20672), .ZN(P1_U2924) );
  AOI22_X1 U23617 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20673) );
  OAI21_X1 U23618 ( .B1(n15027), .B2(n20695), .A(n20673), .ZN(P1_U2925) );
  AOI22_X1 U23619 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20674) );
  OAI21_X1 U23620 ( .B1(n15030), .B2(n20695), .A(n20674), .ZN(P1_U2926) );
  INV_X1 U23621 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U23622 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20675) );
  OAI21_X1 U23623 ( .B1(n20676), .B2(n20695), .A(n20675), .ZN(P1_U2927) );
  AOI22_X1 U23624 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20677) );
  OAI21_X1 U23625 ( .B1(n15034), .B2(n20695), .A(n20677), .ZN(P1_U2928) );
  AOI22_X1 U23626 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20678) );
  OAI21_X1 U23627 ( .B1(n20679), .B2(n20695), .A(n20678), .ZN(P1_U2929) );
  AOI22_X1 U23628 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20680) );
  OAI21_X1 U23629 ( .B1(n20681), .B2(n20695), .A(n20680), .ZN(P1_U2930) );
  AOI22_X1 U23630 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20682) );
  OAI21_X1 U23631 ( .B1(n20683), .B2(n20695), .A(n20682), .ZN(P1_U2931) );
  AOI22_X1 U23632 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20684) );
  OAI21_X1 U23633 ( .B1(n20685), .B2(n20695), .A(n20684), .ZN(P1_U2932) );
  AOI22_X1 U23634 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20686) );
  OAI21_X1 U23635 ( .B1(n20687), .B2(n20695), .A(n20686), .ZN(P1_U2933) );
  AOI22_X1 U23636 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20689) );
  OAI21_X1 U23637 ( .B1(n20690), .B2(n20695), .A(n20689), .ZN(P1_U2934) );
  AOI22_X1 U23638 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20692) );
  OAI21_X1 U23639 ( .B1(n20693), .B2(n20695), .A(n20692), .ZN(P1_U2935) );
  AOI22_X1 U23640 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20688), .B1(n20691), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20694) );
  OAI21_X1 U23641 ( .B1(n20696), .B2(n20695), .A(n20694), .ZN(P1_U2936) );
  AOI22_X1 U23642 ( .A1(n20723), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20728), .ZN(n20699) );
  INV_X1 U23643 ( .A(n20697), .ZN(n20698) );
  NAND2_X1 U23644 ( .A1(n20713), .A2(n20698), .ZN(n20715) );
  NAND2_X1 U23645 ( .A1(n20699), .A2(n20715), .ZN(P1_U2945) );
  AOI22_X1 U23646 ( .A1(n20723), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20702) );
  INV_X1 U23647 ( .A(n20700), .ZN(n20701) );
  NAND2_X1 U23648 ( .A1(n20713), .A2(n20701), .ZN(n20717) );
  NAND2_X1 U23649 ( .A1(n20702), .A2(n20717), .ZN(P1_U2946) );
  AOI22_X1 U23650 ( .A1(n20723), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20704) );
  NAND2_X1 U23651 ( .A1(n20713), .A2(n20703), .ZN(n20719) );
  NAND2_X1 U23652 ( .A1(n20704), .A2(n20719), .ZN(P1_U2947) );
  AOI22_X1 U23653 ( .A1(n20723), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20706) );
  NAND2_X1 U23654 ( .A1(n20713), .A2(n20705), .ZN(n20721) );
  NAND2_X1 U23655 ( .A1(n20706), .A2(n20721), .ZN(P1_U2948) );
  AOI22_X1 U23656 ( .A1(n20723), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20708) );
  NAND2_X1 U23657 ( .A1(n20713), .A2(n20707), .ZN(n20724) );
  NAND2_X1 U23658 ( .A1(n20708), .A2(n20724), .ZN(P1_U2949) );
  AOI22_X1 U23659 ( .A1(n20723), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20710) );
  NAND2_X1 U23660 ( .A1(n20713), .A2(n20709), .ZN(n20726) );
  NAND2_X1 U23661 ( .A1(n20710), .A2(n20726), .ZN(P1_U2950) );
  AOI22_X1 U23662 ( .A1(n20723), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20728), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20714) );
  INV_X1 U23663 ( .A(n20711), .ZN(n20712) );
  NAND2_X1 U23664 ( .A1(n20713), .A2(n20712), .ZN(n20729) );
  NAND2_X1 U23665 ( .A1(n20714), .A2(n20729), .ZN(P1_U2951) );
  AOI22_X1 U23666 ( .A1(n20723), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20716) );
  NAND2_X1 U23667 ( .A1(n20716), .A2(n20715), .ZN(P1_U2960) );
  AOI22_X1 U23668 ( .A1(n20723), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20728), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U23669 ( .A1(n20718), .A2(n20717), .ZN(P1_U2961) );
  AOI22_X1 U23670 ( .A1(n20723), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20728), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20720) );
  NAND2_X1 U23671 ( .A1(n20720), .A2(n20719), .ZN(P1_U2962) );
  AOI22_X1 U23672 ( .A1(n20723), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20728), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20722) );
  NAND2_X1 U23673 ( .A1(n20722), .A2(n20721), .ZN(P1_U2963) );
  AOI22_X1 U23674 ( .A1(n20723), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20728), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20725) );
  NAND2_X1 U23675 ( .A1(n20725), .A2(n20724), .ZN(P1_U2964) );
  AOI22_X1 U23676 ( .A1(n20723), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20728), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20727) );
  NAND2_X1 U23677 ( .A1(n20727), .A2(n20726), .ZN(P1_U2965) );
  AOI22_X1 U23678 ( .A1(n20723), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20728), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20730) );
  NAND2_X1 U23679 ( .A1(n20730), .A2(n20729), .ZN(P1_U2966) );
  AOI22_X1 U23680 ( .A1(n20732), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20731), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20740) );
  AOI21_X1 U23681 ( .B1(n20735), .B2(n20734), .A(n20733), .ZN(n20750) );
  AOI22_X1 U23682 ( .A1(n20750), .A2(n20738), .B1(n20737), .B2(n20736), .ZN(
        n20739) );
  OAI211_X1 U23683 ( .C1(n20742), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        P1_U2995) );
  NOR2_X1 U23684 ( .A1(n20744), .A2(n20743), .ZN(n20775) );
  NOR2_X1 U23685 ( .A1(n20775), .A2(n20768), .ZN(n20765) );
  INV_X1 U23686 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20752) );
  INV_X1 U23687 ( .A(n20745), .ZN(n20746) );
  AOI211_X1 U23688 ( .C1(n20764), .C2(n20752), .A(n20746), .B(n20758), .ZN(
        n20749) );
  OAI22_X1 U23689 ( .A1(n20788), .A2(n20747), .B1(n21523), .B2(n20786), .ZN(
        n20748) );
  AOI211_X1 U23690 ( .C1(n20750), .C2(n20760), .A(n20749), .B(n20748), .ZN(
        n20751) );
  OAI21_X1 U23691 ( .B1(n20765), .B2(n20752), .A(n20751), .ZN(P1_U3027) );
  INV_X1 U23692 ( .A(n20753), .ZN(n20754) );
  AOI21_X1 U23693 ( .B1(n20756), .B2(n20755), .A(n20754), .ZN(n20763) );
  INV_X1 U23694 ( .A(n20757), .ZN(n20761) );
  INV_X1 U23695 ( .A(n20758), .ZN(n20759) );
  AOI22_X1 U23696 ( .A1(n20761), .A2(n20760), .B1(n20759), .B2(n20764), .ZN(
        n20762) );
  OAI211_X1 U23697 ( .C1(n20765), .C2(n20764), .A(n20763), .B(n20762), .ZN(
        P1_U3028) );
  OR2_X1 U23698 ( .A1(n20793), .A2(n20766), .ZN(n20781) );
  INV_X1 U23699 ( .A(n20767), .ZN(n20769) );
  AOI21_X1 U23700 ( .B1(n20770), .B2(n20769), .A(n20768), .ZN(n20779) );
  NOR2_X1 U23701 ( .A1(n20771), .A2(n20784), .ZN(n20777) );
  INV_X1 U23702 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20772) );
  OAI22_X1 U23703 ( .A1(n20788), .A2(n20773), .B1(n20772), .B2(n20786), .ZN(
        n20774) );
  AOI211_X1 U23704 ( .C1(n20777), .C2(n20776), .A(n20775), .B(n20774), .ZN(
        n20778) );
  OAI221_X1 U23705 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20781), .C1(
        n20780), .C2(n20779), .A(n20778), .ZN(P1_U3029) );
  NAND2_X1 U23706 ( .A1(n20783), .A2(n20782), .ZN(n20794) );
  NOR2_X1 U23707 ( .A1(n20785), .A2(n20784), .ZN(n20790) );
  OAI22_X1 U23708 ( .A1(n20788), .A2(n20787), .B1(n21571), .B2(n20786), .ZN(
        n20789) );
  AOI21_X1 U23709 ( .B1(n20790), .B2(n13824), .A(n20789), .ZN(n20791) );
  OAI221_X1 U23710 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20794), .C1(
        n20793), .C2(n20792), .A(n20791), .ZN(P1_U3030) );
  NOR2_X1 U23711 ( .A1(n21623), .A2(n20795), .ZN(P1_U3032) );
  AOI22_X2 U23712 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9584), .B1(DATAI_16_), 
        .B2(n9613), .ZN(n21445) );
  AOI22_X1 U23713 ( .A1(DATAI_24_), .A2(n20844), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n9584), .ZN(n21385) );
  NOR3_X1 U23714 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20864) );
  NAND2_X1 U23715 ( .A1(n21327), .A2(n20864), .ZN(n20847) );
  OAI22_X1 U23716 ( .A1(n21498), .A2(n21385), .B1(n21429), .B2(n20847), .ZN(
        n20801) );
  INV_X1 U23717 ( .A(n20801), .ZN(n20814) );
  INV_X1 U23718 ( .A(n21198), .ZN(n20802) );
  NOR2_X1 U23719 ( .A1(n20802), .A2(n21120), .ZN(n20968) );
  NAND2_X1 U23720 ( .A1(n20809), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21286) );
  NAND2_X1 U23721 ( .A1(n20880), .A2(n21498), .ZN(n20804) );
  AOI21_X1 U23722 ( .B1(n20804), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21433), 
        .ZN(n20808) );
  OR2_X1 U23723 ( .A1(n21118), .A2(n20805), .ZN(n20856) );
  NAND2_X1 U23724 ( .A1(n20932), .A2(n14245), .ZN(n20811) );
  AOI22_X1 U23725 ( .A1(n20808), .A2(n20811), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20847), .ZN(n20806) );
  INV_X1 U23726 ( .A(n20808), .ZN(n20812) );
  NOR2_X1 U23727 ( .A1(n20809), .A2(n21503), .ZN(n21121) );
  INV_X1 U23728 ( .A(n21121), .ZN(n21202) );
  INV_X1 U23729 ( .A(n20968), .ZN(n20810) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20851), .B1(
        n21289), .B2(n20850), .ZN(n20813) );
  OAI211_X1 U23731 ( .C1(n21445), .C2(n20880), .A(n20814), .B(n20813), .ZN(
        P1_U3033) );
  AOI22_X2 U23732 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9584), .B1(DATAI_17_), 
        .B2(n9613), .ZN(n21452) );
  AOI22_X1 U23733 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9584), .B1(DATAI_25_), 
        .B2(n20844), .ZN(n21390) );
  OAI22_X1 U23734 ( .A1(n21498), .A2(n21390), .B1(n21446), .B2(n20847), .ZN(
        n20815) );
  INV_X1 U23735 ( .A(n20815), .ZN(n20818) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20851), .B1(
        n21293), .B2(n20850), .ZN(n20817) );
  OAI211_X1 U23737 ( .C1(n21452), .C2(n20880), .A(n20818), .B(n20817), .ZN(
        P1_U3034) );
  AOI22_X2 U23738 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9584), .B1(DATAI_18_), 
        .B2(n9613), .ZN(n21459) );
  AOI22_X1 U23739 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9584), .B1(DATAI_26_), 
        .B2(n20844), .ZN(n21395) );
  OAI22_X1 U23740 ( .A1(n21498), .A2(n21395), .B1(n21453), .B2(n20847), .ZN(
        n20820) );
  INV_X1 U23741 ( .A(n20820), .ZN(n20823) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20851), .B1(
        n21297), .B2(n20850), .ZN(n20822) );
  OAI211_X1 U23743 ( .C1(n21459), .C2(n20880), .A(n20823), .B(n20822), .ZN(
        P1_U3035) );
  AOI22_X1 U23744 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n9584), .B1(DATAI_19_), 
        .B2(n9613), .ZN(n21466) );
  OAI22_X1 U23745 ( .A1(n21498), .A2(n21399), .B1(n21460), .B2(n20847), .ZN(
        n20825) );
  INV_X1 U23746 ( .A(n20825), .ZN(n20828) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20851), .B1(
        n21301), .B2(n20850), .ZN(n20827) );
  OAI211_X1 U23748 ( .C1(n9779), .C2(n20880), .A(n20828), .B(n20827), .ZN(
        P1_U3036) );
  AOI22_X2 U23749 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9584), .B1(DATAI_20_), 
        .B2(n9613), .ZN(n21473) );
  AOI22_X1 U23750 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9584), .B1(DATAI_28_), 
        .B2(n20844), .ZN(n21404) );
  OAI22_X1 U23751 ( .A1(n21498), .A2(n21404), .B1(n21467), .B2(n20847), .ZN(
        n20830) );
  INV_X1 U23752 ( .A(n20830), .ZN(n20833) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20851), .B1(
        n21305), .B2(n20850), .ZN(n20832) );
  OAI211_X1 U23754 ( .C1(n21473), .C2(n20880), .A(n20833), .B(n20832), .ZN(
        P1_U3037) );
  AOI22_X2 U23755 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9584), .B1(DATAI_21_), 
        .B2(n9613), .ZN(n21480) );
  AOI22_X1 U23756 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9584), .B1(DATAI_29_), 
        .B2(n20844), .ZN(n21409) );
  OAI22_X1 U23757 ( .A1(n21498), .A2(n21409), .B1(n21474), .B2(n20847), .ZN(
        n20835) );
  INV_X1 U23758 ( .A(n20835), .ZN(n20838) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20851), .B1(
        n21309), .B2(n20850), .ZN(n20837) );
  OAI211_X1 U23760 ( .C1(n21480), .C2(n20880), .A(n20838), .B(n20837), .ZN(
        P1_U3038) );
  AOI22_X2 U23761 ( .A1(DATAI_22_), .A2(n9613), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9584), .ZN(n21487) );
  AOI22_X1 U23762 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9584), .B1(DATAI_30_), 
        .B2(n20844), .ZN(n21414) );
  OAI22_X1 U23763 ( .A1(n21498), .A2(n21414), .B1(n21481), .B2(n20847), .ZN(
        n20840) );
  INV_X1 U23764 ( .A(n20840), .ZN(n20843) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20851), .B1(
        n21313), .B2(n20850), .ZN(n20842) );
  OAI211_X1 U23766 ( .C1(n21487), .C2(n20880), .A(n20843), .B(n20842), .ZN(
        P1_U3039) );
  AOI22_X2 U23767 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9584), .B1(DATAI_23_), 
        .B2(n9613), .ZN(n21499) );
  AOI22_X1 U23768 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n9584), .B1(DATAI_31_), 
        .B2(n20844), .ZN(n21423) );
  OAI22_X1 U23769 ( .A1(n21498), .A2(n21423), .B1(n21488), .B2(n20847), .ZN(
        n20848) );
  INV_X1 U23770 ( .A(n20848), .ZN(n20853) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20851), .B1(
        n21319), .B2(n20850), .ZN(n20852) );
  OAI211_X1 U23772 ( .C1(n21499), .C2(n20880), .A(n20853), .B(n20852), .ZN(
        P1_U3040) );
  INV_X1 U23773 ( .A(n20864), .ZN(n20855) );
  OAI21_X1 U23774 ( .B1(n20856), .B2(n20854), .A(n20887), .ZN(n20860) );
  NAND2_X1 U23775 ( .A1(n20860), .A2(n9585), .ZN(n20858) );
  NAND2_X1 U23776 ( .A1(n20864), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20857) );
  OAI22_X1 U23777 ( .A1(n21430), .A2(n20888), .B1(n21429), .B2(n20887), .ZN(
        n20859) );
  INV_X1 U23778 ( .A(n20859), .ZN(n20866) );
  INV_X1 U23779 ( .A(n20933), .ZN(n20862) );
  INV_X1 U23780 ( .A(n20860), .ZN(n20861) );
  OAI211_X1 U23781 ( .C1(n20862), .C2(n21373), .A(n9585), .B(n20861), .ZN(
        n20863) );
  OAI211_X1 U23782 ( .C1(n9585), .C2(n20864), .A(n21439), .B(n20863), .ZN(
        n20891) );
  INV_X1 U23783 ( .A(n20880), .ZN(n20890) );
  INV_X1 U23784 ( .A(n21385), .ZN(n21442) );
  AOI22_X1 U23785 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20891), .B1(
        n20890), .B2(n21442), .ZN(n20865) );
  OAI211_X1 U23786 ( .C1(n21445), .C2(n20927), .A(n20866), .B(n20865), .ZN(
        P1_U3041) );
  OAI22_X1 U23787 ( .A1(n21447), .A2(n20888), .B1(n21446), .B2(n20887), .ZN(
        n20867) );
  INV_X1 U23788 ( .A(n20867), .ZN(n20869) );
  INV_X1 U23789 ( .A(n20927), .ZN(n20877) );
  INV_X1 U23790 ( .A(n21452), .ZN(n21387) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20891), .B1(
        n20877), .B2(n21387), .ZN(n20868) );
  OAI211_X1 U23792 ( .C1(n21390), .C2(n20880), .A(n20869), .B(n20868), .ZN(
        P1_U3042) );
  OAI22_X1 U23793 ( .A1(n21454), .A2(n20888), .B1(n21453), .B2(n20887), .ZN(
        n20870) );
  INV_X1 U23794 ( .A(n20870), .ZN(n20872) );
  INV_X1 U23795 ( .A(n21395), .ZN(n21456) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20891), .B1(
        n20890), .B2(n21456), .ZN(n20871) );
  OAI211_X1 U23797 ( .C1(n21459), .C2(n20927), .A(n20872), .B(n20871), .ZN(
        P1_U3043) );
  OAI22_X1 U23798 ( .A1(n21461), .A2(n20888), .B1(n21460), .B2(n20887), .ZN(
        n20873) );
  INV_X1 U23799 ( .A(n20873), .ZN(n20875) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20891), .B1(
        n20877), .B2(n9778), .ZN(n20874) );
  OAI211_X1 U23801 ( .C1(n21399), .C2(n20880), .A(n20875), .B(n20874), .ZN(
        P1_U3044) );
  OAI22_X1 U23802 ( .A1(n21468), .A2(n20888), .B1(n21467), .B2(n20887), .ZN(
        n20876) );
  INV_X1 U23803 ( .A(n20876), .ZN(n20879) );
  INV_X1 U23804 ( .A(n21473), .ZN(n21401) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20891), .B1(
        n20877), .B2(n21401), .ZN(n20878) );
  OAI211_X1 U23806 ( .C1(n21404), .C2(n20880), .A(n20879), .B(n20878), .ZN(
        P1_U3045) );
  OAI22_X1 U23807 ( .A1(n21475), .A2(n20888), .B1(n21474), .B2(n20887), .ZN(
        n20881) );
  INV_X1 U23808 ( .A(n20881), .ZN(n20883) );
  INV_X1 U23809 ( .A(n21409), .ZN(n21477) );
  AOI22_X1 U23810 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20891), .B1(
        n20890), .B2(n21477), .ZN(n20882) );
  OAI211_X1 U23811 ( .C1(n21480), .C2(n20927), .A(n20883), .B(n20882), .ZN(
        P1_U3046) );
  OAI22_X1 U23812 ( .A1(n21482), .A2(n20888), .B1(n21481), .B2(n20887), .ZN(
        n20884) );
  INV_X1 U23813 ( .A(n20884), .ZN(n20886) );
  INV_X1 U23814 ( .A(n21414), .ZN(n21484) );
  AOI22_X1 U23815 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20891), .B1(
        n20890), .B2(n21484), .ZN(n20885) );
  OAI211_X1 U23816 ( .C1(n21487), .C2(n20927), .A(n20886), .B(n20885), .ZN(
        P1_U3047) );
  OAI22_X1 U23817 ( .A1(n21491), .A2(n20888), .B1(n21488), .B2(n20887), .ZN(
        n20889) );
  INV_X1 U23818 ( .A(n20889), .ZN(n20893) );
  INV_X1 U23819 ( .A(n21423), .ZN(n21493) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20891), .B1(
        n20890), .B2(n21493), .ZN(n20892) );
  OAI211_X1 U23821 ( .C1(n21499), .C2(n20927), .A(n20893), .B(n20892), .ZN(
        P1_U3048) );
  NAND3_X1 U23822 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21275), .A3(
        n21276), .ZN(n20937) );
  OR2_X1 U23823 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20937), .ZN(
        n20921) );
  OAI22_X1 U23824 ( .A1(n20966), .A2(n21445), .B1(n21429), .B2(n20921), .ZN(
        n20895) );
  INV_X1 U23825 ( .A(n20895), .ZN(n20902) );
  NAND2_X1 U23826 ( .A1(n20966), .A2(n20927), .ZN(n20896) );
  AOI21_X1 U23827 ( .B1(n20896), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21433), 
        .ZN(n20898) );
  NAND2_X1 U23828 ( .A1(n20932), .A2(n21375), .ZN(n20899) );
  AOI22_X1 U23829 ( .A1(n20898), .A2(n20899), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20921), .ZN(n20897) );
  OR2_X1 U23830 ( .A1(n21198), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21051) );
  NAND2_X1 U23831 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21051), .ZN(n21048) );
  NAND3_X1 U23832 ( .A1(n21200), .A2(n20897), .A3(n21048), .ZN(n20924) );
  INV_X1 U23833 ( .A(n20898), .ZN(n20900) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20924), .B1(
        n21289), .B2(n20923), .ZN(n20901) );
  OAI211_X1 U23835 ( .C1(n21385), .C2(n20927), .A(n20902), .B(n20901), .ZN(
        P1_U3049) );
  OAI22_X1 U23836 ( .A1(n20927), .A2(n21390), .B1(n21446), .B2(n20921), .ZN(
        n20903) );
  INV_X1 U23837 ( .A(n20903), .ZN(n20905) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20924), .B1(
        n21293), .B2(n20923), .ZN(n20904) );
  OAI211_X1 U23839 ( .C1(n21452), .C2(n20966), .A(n20905), .B(n20904), .ZN(
        P1_U3050) );
  OAI22_X1 U23840 ( .A1(n20966), .A2(n21459), .B1(n21453), .B2(n20921), .ZN(
        n20906) );
  INV_X1 U23841 ( .A(n20906), .ZN(n20908) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20924), .B1(
        n21297), .B2(n20923), .ZN(n20907) );
  OAI211_X1 U23843 ( .C1(n21395), .C2(n20927), .A(n20908), .B(n20907), .ZN(
        P1_U3051) );
  OAI22_X1 U23844 ( .A1(n20927), .A2(n21399), .B1(n21460), .B2(n20921), .ZN(
        n20909) );
  INV_X1 U23845 ( .A(n20909), .ZN(n20911) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20924), .B1(
        n21301), .B2(n20923), .ZN(n20910) );
  OAI211_X1 U23847 ( .C1(n9779), .C2(n20966), .A(n20911), .B(n20910), .ZN(
        P1_U3052) );
  OAI22_X1 U23848 ( .A1(n20966), .A2(n21473), .B1(n21467), .B2(n20921), .ZN(
        n20912) );
  INV_X1 U23849 ( .A(n20912), .ZN(n20914) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20924), .B1(
        n21305), .B2(n20923), .ZN(n20913) );
  OAI211_X1 U23851 ( .C1(n21404), .C2(n20927), .A(n20914), .B(n20913), .ZN(
        P1_U3053) );
  OAI22_X1 U23852 ( .A1(n20927), .A2(n21409), .B1(n21474), .B2(n20921), .ZN(
        n20915) );
  INV_X1 U23853 ( .A(n20915), .ZN(n20917) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20924), .B1(
        n21309), .B2(n20923), .ZN(n20916) );
  OAI211_X1 U23855 ( .C1(n21480), .C2(n20966), .A(n20917), .B(n20916), .ZN(
        P1_U3054) );
  OAI22_X1 U23856 ( .A1(n20966), .A2(n21487), .B1(n21481), .B2(n20921), .ZN(
        n20918) );
  INV_X1 U23857 ( .A(n20918), .ZN(n20920) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20924), .B1(
        n21313), .B2(n20923), .ZN(n20919) );
  OAI211_X1 U23859 ( .C1(n21414), .C2(n20927), .A(n20920), .B(n20919), .ZN(
        P1_U3055) );
  OAI22_X1 U23860 ( .A1(n20966), .A2(n21499), .B1(n21488), .B2(n20921), .ZN(
        n20922) );
  INV_X1 U23861 ( .A(n20922), .ZN(n20926) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20924), .B1(
        n21319), .B2(n20923), .ZN(n20925) );
  OAI211_X1 U23863 ( .C1(n21423), .C2(n20927), .A(n20926), .B(n20925), .ZN(
        P1_U3056) );
  INV_X1 U23864 ( .A(n20928), .ZN(n21234) );
  NAND2_X1 U23865 ( .A1(n21234), .A2(n21275), .ZN(n20960) );
  OAI22_X1 U23866 ( .A1(n20978), .A2(n21445), .B1(n21429), .B2(n20960), .ZN(
        n20929) );
  INV_X1 U23867 ( .A(n20929), .ZN(n20941) );
  INV_X1 U23868 ( .A(n20960), .ZN(n20931) );
  AOI21_X1 U23869 ( .B1(n20932), .B2(n21424), .A(n20931), .ZN(n20939) );
  OR2_X1 U23870 ( .A1(n20933), .A2(n21433), .ZN(n20934) );
  INV_X1 U23871 ( .A(n20938), .ZN(n20935) );
  AOI22_X1 U23872 ( .A1(n20939), .A2(n20935), .B1(n21433), .B2(n20937), .ZN(
        n20936) );
  NAND2_X1 U23873 ( .A1(n21439), .A2(n20936), .ZN(n20963) );
  AOI22_X1 U23874 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20963), .B1(
        n21289), .B2(n20962), .ZN(n20940) );
  OAI211_X1 U23875 ( .C1(n21385), .C2(n20966), .A(n20941), .B(n20940), .ZN(
        P1_U3057) );
  OAI22_X1 U23876 ( .A1(n20978), .A2(n21452), .B1(n21446), .B2(n20960), .ZN(
        n20942) );
  INV_X1 U23877 ( .A(n20942), .ZN(n20944) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20963), .B1(
        n21293), .B2(n20962), .ZN(n20943) );
  OAI211_X1 U23879 ( .C1(n21390), .C2(n20966), .A(n20944), .B(n20943), .ZN(
        P1_U3058) );
  OAI22_X1 U23880 ( .A1(n20966), .A2(n21395), .B1(n21453), .B2(n20960), .ZN(
        n20945) );
  INV_X1 U23881 ( .A(n20945), .ZN(n20947) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20963), .B1(
        n21297), .B2(n20962), .ZN(n20946) );
  OAI211_X1 U23883 ( .C1(n21459), .C2(n20978), .A(n20947), .B(n20946), .ZN(
        P1_U3059) );
  OAI22_X1 U23884 ( .A1(n20978), .A2(n9779), .B1(n21460), .B2(n20960), .ZN(
        n20948) );
  INV_X1 U23885 ( .A(n20948), .ZN(n20950) );
  AOI22_X1 U23886 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20963), .B1(
        n21301), .B2(n20962), .ZN(n20949) );
  OAI211_X1 U23887 ( .C1(n21399), .C2(n20966), .A(n20950), .B(n20949), .ZN(
        P1_U3060) );
  OAI22_X1 U23888 ( .A1(n20966), .A2(n21404), .B1(n21467), .B2(n20960), .ZN(
        n20951) );
  INV_X1 U23889 ( .A(n20951), .ZN(n20953) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20963), .B1(
        n21305), .B2(n20962), .ZN(n20952) );
  OAI211_X1 U23891 ( .C1(n21473), .C2(n20978), .A(n20953), .B(n20952), .ZN(
        P1_U3061) );
  OAI22_X1 U23892 ( .A1(n20966), .A2(n21409), .B1(n21474), .B2(n20960), .ZN(
        n20954) );
  INV_X1 U23893 ( .A(n20954), .ZN(n20956) );
  AOI22_X1 U23894 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20963), .B1(
        n21309), .B2(n20962), .ZN(n20955) );
  OAI211_X1 U23895 ( .C1(n21480), .C2(n20978), .A(n20956), .B(n20955), .ZN(
        P1_U3062) );
  OAI22_X1 U23896 ( .A1(n20978), .A2(n21487), .B1(n21481), .B2(n20960), .ZN(
        n20957) );
  INV_X1 U23897 ( .A(n20957), .ZN(n20959) );
  AOI22_X1 U23898 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20963), .B1(
        n21313), .B2(n20962), .ZN(n20958) );
  OAI211_X1 U23899 ( .C1(n21414), .C2(n20966), .A(n20959), .B(n20958), .ZN(
        P1_U3063) );
  OAI22_X1 U23900 ( .A1(n20978), .A2(n21499), .B1(n21488), .B2(n20960), .ZN(
        n20961) );
  INV_X1 U23901 ( .A(n20961), .ZN(n20965) );
  AOI22_X1 U23902 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20963), .B1(
        n21319), .B2(n20962), .ZN(n20964) );
  OAI211_X1 U23903 ( .C1(n21423), .C2(n20966), .A(n20965), .B(n20964), .ZN(
        P1_U3064) );
  INV_X1 U23904 ( .A(n21117), .ZN(n21274) );
  OR2_X1 U23905 ( .A1(n21279), .A2(n20967), .ZN(n20972) );
  NOR2_X1 U23906 ( .A1(n20972), .A2(n21433), .ZN(n21081) );
  NAND2_X1 U23907 ( .A1(n21081), .A2(n14245), .ZN(n20970) );
  INV_X1 U23908 ( .A(n21286), .ZN(n21366) );
  NAND2_X1 U23909 ( .A1(n20968), .A2(n21366), .ZN(n20969) );
  NOR3_X1 U23910 ( .A1(n21276), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21014) );
  INV_X1 U23911 ( .A(n21014), .ZN(n21007) );
  NOR2_X1 U23912 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21007), .ZN(
        n20977) );
  INV_X1 U23913 ( .A(n20977), .ZN(n20999) );
  OAI22_X1 U23914 ( .A1(n21430), .A2(n21000), .B1(n21429), .B2(n20999), .ZN(
        n20971) );
  INV_X1 U23915 ( .A(n20971), .ZN(n20980) );
  INV_X1 U23916 ( .A(n20972), .ZN(n21047) );
  AOI21_X1 U23917 ( .B1(n20978), .B2(n21044), .A(n21373), .ZN(n20973) );
  AOI21_X1 U23918 ( .B1(n21047), .B2(n14245), .A(n20973), .ZN(n20974) );
  NOR2_X1 U23919 ( .A1(n20974), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U23920 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21442), .ZN(n20979) );
  OAI211_X1 U23921 ( .C1(n21445), .C2(n21044), .A(n20980), .B(n20979), .ZN(
        P1_U3065) );
  OAI22_X1 U23922 ( .A1(n21447), .A2(n21000), .B1(n21446), .B2(n20999), .ZN(
        n20981) );
  INV_X1 U23923 ( .A(n20981), .ZN(n20983) );
  INV_X1 U23924 ( .A(n21390), .ZN(n21449) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21449), .ZN(n20982) );
  OAI211_X1 U23926 ( .C1(n21452), .C2(n21044), .A(n20983), .B(n20982), .ZN(
        P1_U3066) );
  OAI22_X1 U23927 ( .A1(n21454), .A2(n21000), .B1(n21453), .B2(n20999), .ZN(
        n20984) );
  INV_X1 U23928 ( .A(n20984), .ZN(n20986) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21456), .ZN(n20985) );
  OAI211_X1 U23930 ( .C1(n21459), .C2(n21044), .A(n20986), .B(n20985), .ZN(
        P1_U3067) );
  OAI22_X1 U23931 ( .A1(n21461), .A2(n21000), .B1(n21460), .B2(n20999), .ZN(
        n20987) );
  INV_X1 U23932 ( .A(n20987), .ZN(n20989) );
  INV_X1 U23933 ( .A(n21399), .ZN(n21463) );
  AOI22_X1 U23934 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21463), .ZN(n20988) );
  OAI211_X1 U23935 ( .C1(n9779), .C2(n21044), .A(n20989), .B(n20988), .ZN(
        P1_U3068) );
  OAI22_X1 U23936 ( .A1(n21468), .A2(n21000), .B1(n21467), .B2(n20999), .ZN(
        n20990) );
  INV_X1 U23937 ( .A(n20990), .ZN(n20992) );
  INV_X1 U23938 ( .A(n21404), .ZN(n21470) );
  AOI22_X1 U23939 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21470), .ZN(n20991) );
  OAI211_X1 U23940 ( .C1(n21473), .C2(n21044), .A(n20992), .B(n20991), .ZN(
        P1_U3069) );
  OAI22_X1 U23941 ( .A1(n21475), .A2(n21000), .B1(n21474), .B2(n20999), .ZN(
        n20993) );
  INV_X1 U23942 ( .A(n20993), .ZN(n20995) );
  AOI22_X1 U23943 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21477), .ZN(n20994) );
  OAI211_X1 U23944 ( .C1(n21480), .C2(n21044), .A(n20995), .B(n20994), .ZN(
        P1_U3070) );
  OAI22_X1 U23945 ( .A1(n21482), .A2(n21000), .B1(n21481), .B2(n20999), .ZN(
        n20996) );
  INV_X1 U23946 ( .A(n20996), .ZN(n20998) );
  AOI22_X1 U23947 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21484), .ZN(n20997) );
  OAI211_X1 U23948 ( .C1(n21487), .C2(n21044), .A(n20998), .B(n20997), .ZN(
        P1_U3071) );
  OAI22_X1 U23949 ( .A1(n21491), .A2(n21000), .B1(n21488), .B2(n20999), .ZN(
        n21001) );
  INV_X1 U23950 ( .A(n21001), .ZN(n21005) );
  AOI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21003), .B1(
        n21002), .B2(n21493), .ZN(n21004) );
  OAI211_X1 U23952 ( .C1(n21499), .C2(n21044), .A(n21005), .B(n21004), .ZN(
        P1_U3072) );
  INV_X1 U23953 ( .A(n21324), .ZN(n21006) );
  INV_X1 U23954 ( .A(n20854), .ZN(n21325) );
  NAND2_X1 U23955 ( .A1(n21081), .A2(n21325), .ZN(n21009) );
  NOR2_X1 U23956 ( .A1(n21327), .A2(n21007), .ZN(n21010) );
  AOI22_X1 U23957 ( .A1(n9585), .A2(n21010), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21014), .ZN(n21008) );
  INV_X1 U23958 ( .A(n21010), .ZN(n21037) );
  OAI22_X1 U23959 ( .A1(n21430), .A2(n21038), .B1(n21429), .B2(n21037), .ZN(
        n21011) );
  INV_X1 U23960 ( .A(n21011), .ZN(n21017) );
  NOR3_X1 U23961 ( .A1(n21013), .A2(n21012), .A3(n21432), .ZN(n21015) );
  INV_X1 U23962 ( .A(n21044), .ZN(n21034) );
  AOI22_X1 U23963 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21041), .B1(
        n21034), .B2(n21442), .ZN(n21016) );
  OAI211_X1 U23964 ( .C1(n21445), .C2(n21075), .A(n21017), .B(n21016), .ZN(
        P1_U3073) );
  OAI22_X1 U23965 ( .A1(n21447), .A2(n21038), .B1(n21446), .B2(n21037), .ZN(
        n21018) );
  INV_X1 U23966 ( .A(n21018), .ZN(n21020) );
  AOI22_X1 U23967 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21041), .B1(
        n21034), .B2(n21449), .ZN(n21019) );
  OAI211_X1 U23968 ( .C1(n21452), .C2(n21075), .A(n21020), .B(n21019), .ZN(
        P1_U3074) );
  OAI22_X1 U23969 ( .A1(n21454), .A2(n21038), .B1(n21453), .B2(n21037), .ZN(
        n21021) );
  INV_X1 U23970 ( .A(n21021), .ZN(n21023) );
  INV_X1 U23971 ( .A(n21459), .ZN(n21392) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21041), .B1(
        n21040), .B2(n21392), .ZN(n21022) );
  OAI211_X1 U23973 ( .C1(n21395), .C2(n21044), .A(n21023), .B(n21022), .ZN(
        P1_U3075) );
  OAI22_X1 U23974 ( .A1(n21461), .A2(n21038), .B1(n21460), .B2(n21037), .ZN(
        n21024) );
  INV_X1 U23975 ( .A(n21024), .ZN(n21026) );
  AOI22_X1 U23976 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21041), .B1(
        n21040), .B2(n9778), .ZN(n21025) );
  OAI211_X1 U23977 ( .C1(n21399), .C2(n21044), .A(n21026), .B(n21025), .ZN(
        P1_U3076) );
  OAI22_X1 U23978 ( .A1(n21468), .A2(n21038), .B1(n21467), .B2(n21037), .ZN(
        n21027) );
  INV_X1 U23979 ( .A(n21027), .ZN(n21029) );
  AOI22_X1 U23980 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21041), .B1(
        n21040), .B2(n21401), .ZN(n21028) );
  OAI211_X1 U23981 ( .C1(n21404), .C2(n21044), .A(n21029), .B(n21028), .ZN(
        P1_U3077) );
  OAI22_X1 U23982 ( .A1(n21475), .A2(n21038), .B1(n21474), .B2(n21037), .ZN(
        n21030) );
  INV_X1 U23983 ( .A(n21030), .ZN(n21032) );
  INV_X1 U23984 ( .A(n21480), .ZN(n21406) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21041), .B1(
        n21040), .B2(n21406), .ZN(n21031) );
  OAI211_X1 U23986 ( .C1(n21409), .C2(n21044), .A(n21032), .B(n21031), .ZN(
        P1_U3078) );
  OAI22_X1 U23987 ( .A1(n21482), .A2(n21038), .B1(n21481), .B2(n21037), .ZN(
        n21033) );
  INV_X1 U23988 ( .A(n21033), .ZN(n21036) );
  AOI22_X1 U23989 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21041), .B1(
        n21034), .B2(n21484), .ZN(n21035) );
  OAI211_X1 U23990 ( .C1(n21487), .C2(n21075), .A(n21036), .B(n21035), .ZN(
        P1_U3079) );
  OAI22_X1 U23991 ( .A1(n21491), .A2(n21038), .B1(n21488), .B2(n21037), .ZN(
        n21039) );
  INV_X1 U23992 ( .A(n21039), .ZN(n21043) );
  INV_X1 U23993 ( .A(n21499), .ZN(n21418) );
  AOI22_X1 U23994 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21041), .B1(
        n21040), .B2(n21418), .ZN(n21042) );
  OAI211_X1 U23995 ( .C1(n21423), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        P1_U3080) );
  INV_X1 U23996 ( .A(n21194), .ZN(n21371) );
  NAND2_X1 U23997 ( .A1(n21327), .A2(n10565), .ZN(n21074) );
  OAI22_X1 U23998 ( .A1(n21075), .A2(n21385), .B1(n21074), .B2(n21429), .ZN(
        n21045) );
  INV_X1 U23999 ( .A(n21045), .ZN(n21055) );
  AOI21_X1 U24000 ( .B1(n21109), .B2(n21075), .A(n21373), .ZN(n21046) );
  NOR2_X1 U24001 ( .A1(n21046), .A2(n21433), .ZN(n21050) );
  NAND2_X1 U24002 ( .A1(n21047), .A2(n21375), .ZN(n21052) );
  AOI22_X1 U24003 ( .A1(n21050), .A2(n21052), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21074), .ZN(n21049) );
  NAND3_X1 U24004 ( .A1(n21378), .A2(n21049), .A3(n21048), .ZN(n21078) );
  INV_X1 U24005 ( .A(n21050), .ZN(n21053) );
  AOI22_X1 U24006 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21078), .B1(
        n21289), .B2(n21077), .ZN(n21054) );
  OAI211_X1 U24007 ( .C1(n21445), .C2(n21109), .A(n21055), .B(n21054), .ZN(
        P1_U3081) );
  OAI22_X1 U24008 ( .A1(n21075), .A2(n21390), .B1(n21074), .B2(n21446), .ZN(
        n21056) );
  INV_X1 U24009 ( .A(n21056), .ZN(n21058) );
  AOI22_X1 U24010 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21078), .B1(
        n21293), .B2(n21077), .ZN(n21057) );
  OAI211_X1 U24011 ( .C1(n21452), .C2(n21109), .A(n21058), .B(n21057), .ZN(
        P1_U3082) );
  OAI22_X1 U24012 ( .A1(n21109), .A2(n21459), .B1(n21074), .B2(n21453), .ZN(
        n21059) );
  INV_X1 U24013 ( .A(n21059), .ZN(n21061) );
  AOI22_X1 U24014 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21078), .B1(
        n21297), .B2(n21077), .ZN(n21060) );
  OAI211_X1 U24015 ( .C1(n21395), .C2(n21075), .A(n21061), .B(n21060), .ZN(
        P1_U3083) );
  OAI22_X1 U24016 ( .A1(n21109), .A2(n9779), .B1(n21074), .B2(n21460), .ZN(
        n21062) );
  INV_X1 U24017 ( .A(n21062), .ZN(n21064) );
  AOI22_X1 U24018 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21078), .B1(
        n21301), .B2(n21077), .ZN(n21063) );
  OAI211_X1 U24019 ( .C1(n21399), .C2(n21075), .A(n21064), .B(n21063), .ZN(
        P1_U3084) );
  OAI22_X1 U24020 ( .A1(n21109), .A2(n21473), .B1(n21074), .B2(n21467), .ZN(
        n21065) );
  INV_X1 U24021 ( .A(n21065), .ZN(n21067) );
  AOI22_X1 U24022 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21078), .B1(
        n21305), .B2(n21077), .ZN(n21066) );
  OAI211_X1 U24023 ( .C1(n21404), .C2(n21075), .A(n21067), .B(n21066), .ZN(
        P1_U3085) );
  OAI22_X1 U24024 ( .A1(n21075), .A2(n21409), .B1(n21074), .B2(n21474), .ZN(
        n21068) );
  INV_X1 U24025 ( .A(n21068), .ZN(n21070) );
  AOI22_X1 U24026 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21078), .B1(
        n21309), .B2(n21077), .ZN(n21069) );
  OAI211_X1 U24027 ( .C1(n21480), .C2(n21109), .A(n21070), .B(n21069), .ZN(
        P1_U3086) );
  OAI22_X1 U24028 ( .A1(n21075), .A2(n21414), .B1(n21074), .B2(n21481), .ZN(
        n21071) );
  INV_X1 U24029 ( .A(n21071), .ZN(n21073) );
  AOI22_X1 U24030 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21078), .B1(
        n21313), .B2(n21077), .ZN(n21072) );
  OAI211_X1 U24031 ( .C1(n21487), .C2(n21109), .A(n21073), .B(n21072), .ZN(
        P1_U3087) );
  OAI22_X1 U24032 ( .A1(n21075), .A2(n21423), .B1(n21488), .B2(n21074), .ZN(
        n21076) );
  INV_X1 U24033 ( .A(n21076), .ZN(n21080) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21078), .B1(
        n21319), .B2(n21077), .ZN(n21079) );
  OAI211_X1 U24035 ( .C1(n21499), .C2(n21109), .A(n21080), .B(n21079), .ZN(
        P1_U3088) );
  NAND2_X1 U24036 ( .A1(n21081), .A2(n21424), .ZN(n21084) );
  INV_X1 U24037 ( .A(n21110), .ZN(n21082) );
  AOI22_X1 U24038 ( .A1(n9585), .A2(n21082), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n10565), .ZN(n21083) );
  OAI22_X1 U24039 ( .A1(n21430), .A2(n21111), .B1(n21110), .B2(n21429), .ZN(
        n21085) );
  INV_X1 U24040 ( .A(n21085), .ZN(n21090) );
  NOR2_X1 U24041 ( .A1(n21088), .A2(n21241), .ZN(n21086) );
  INV_X1 U24042 ( .A(n21445), .ZN(n21382) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21114), .B1(
        n21153), .B2(n21382), .ZN(n21089) );
  OAI211_X1 U24044 ( .C1(n21385), .C2(n21109), .A(n21090), .B(n21089), .ZN(
        P1_U3089) );
  OAI22_X1 U24045 ( .A1(n21447), .A2(n21111), .B1(n21110), .B2(n21446), .ZN(
        n21091) );
  INV_X1 U24046 ( .A(n21091), .ZN(n21093) );
  AOI22_X1 U24047 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21114), .B1(
        n21153), .B2(n21387), .ZN(n21092) );
  OAI211_X1 U24048 ( .C1(n21390), .C2(n21109), .A(n21093), .B(n21092), .ZN(
        P1_U3090) );
  OAI22_X1 U24049 ( .A1(n21454), .A2(n21111), .B1(n21110), .B2(n21453), .ZN(
        n21094) );
  INV_X1 U24050 ( .A(n21094), .ZN(n21096) );
  INV_X1 U24051 ( .A(n21109), .ZN(n21113) );
  AOI22_X1 U24052 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21456), .ZN(n21095) );
  OAI211_X1 U24053 ( .C1(n21459), .C2(n21125), .A(n21096), .B(n21095), .ZN(
        P1_U3091) );
  OAI22_X1 U24054 ( .A1(n21461), .A2(n21111), .B1(n21110), .B2(n21460), .ZN(
        n21097) );
  INV_X1 U24055 ( .A(n21097), .ZN(n21099) );
  AOI22_X1 U24056 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21463), .ZN(n21098) );
  OAI211_X1 U24057 ( .C1(n9779), .C2(n21125), .A(n21099), .B(n21098), .ZN(
        P1_U3092) );
  OAI22_X1 U24058 ( .A1(n21468), .A2(n21111), .B1(n21110), .B2(n21467), .ZN(
        n21100) );
  INV_X1 U24059 ( .A(n21100), .ZN(n21102) );
  AOI22_X1 U24060 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21470), .ZN(n21101) );
  OAI211_X1 U24061 ( .C1(n21473), .C2(n21125), .A(n21102), .B(n21101), .ZN(
        P1_U3093) );
  OAI22_X1 U24062 ( .A1(n21475), .A2(n21111), .B1(n21110), .B2(n21474), .ZN(
        n21103) );
  INV_X1 U24063 ( .A(n21103), .ZN(n21105) );
  AOI22_X1 U24064 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21477), .ZN(n21104) );
  OAI211_X1 U24065 ( .C1(n21480), .C2(n21125), .A(n21105), .B(n21104), .ZN(
        P1_U3094) );
  OAI22_X1 U24066 ( .A1(n21482), .A2(n21111), .B1(n21110), .B2(n21481), .ZN(
        n21106) );
  INV_X1 U24067 ( .A(n21106), .ZN(n21108) );
  INV_X1 U24068 ( .A(n21487), .ZN(n21411) );
  AOI22_X1 U24069 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21114), .B1(
        n21153), .B2(n21411), .ZN(n21107) );
  OAI211_X1 U24070 ( .C1(n21414), .C2(n21109), .A(n21108), .B(n21107), .ZN(
        P1_U3095) );
  OAI22_X1 U24071 ( .A1(n21491), .A2(n21111), .B1(n21110), .B2(n21488), .ZN(
        n21112) );
  INV_X1 U24072 ( .A(n21112), .ZN(n21116) );
  AOI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21114), .B1(
        n21113), .B2(n21493), .ZN(n21115) );
  OAI211_X1 U24074 ( .C1(n21499), .C2(n21125), .A(n21116), .B(n21115), .ZN(
        P1_U3096) );
  NAND2_X1 U24075 ( .A1(n21118), .A2(n21279), .ZN(n21236) );
  OR2_X1 U24076 ( .A1(n21236), .A2(n21375), .ZN(n21119) );
  NOR3_X1 U24077 ( .A1(n21275), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21165) );
  INV_X1 U24078 ( .A(n21165), .ZN(n21157) );
  NOR2_X1 U24079 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21157), .ZN(
        n21129) );
  INV_X1 U24080 ( .A(n21129), .ZN(n21150) );
  NAND2_X1 U24081 ( .A1(n21119), .A2(n21150), .ZN(n21126) );
  NAND2_X1 U24082 ( .A1(n21126), .A2(n9585), .ZN(n21123) );
  AND2_X1 U24083 ( .A1(n21120), .A2(n21198), .ZN(n21280) );
  NAND2_X1 U24084 ( .A1(n21121), .A2(n21280), .ZN(n21122) );
  OAI22_X1 U24085 ( .A1(n21430), .A2(n21151), .B1(n21429), .B2(n21150), .ZN(
        n21124) );
  INV_X1 U24086 ( .A(n21124), .ZN(n21131) );
  AOI21_X1 U24087 ( .B1(n21193), .B2(n21125), .A(n21373), .ZN(n21127) );
  OR2_X1 U24088 ( .A1(n21127), .A2(n21126), .ZN(n21128) );
  AOI22_X1 U24089 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21442), .ZN(n21130) );
  OAI211_X1 U24090 ( .C1(n21445), .C2(n21193), .A(n21131), .B(n21130), .ZN(
        P1_U3097) );
  OAI22_X1 U24091 ( .A1(n21447), .A2(n21151), .B1(n21446), .B2(n21150), .ZN(
        n21132) );
  INV_X1 U24092 ( .A(n21132), .ZN(n21134) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21449), .ZN(n21133) );
  OAI211_X1 U24094 ( .C1(n21452), .C2(n21193), .A(n21134), .B(n21133), .ZN(
        P1_U3098) );
  OAI22_X1 U24095 ( .A1(n21454), .A2(n21151), .B1(n21453), .B2(n21150), .ZN(
        n21135) );
  INV_X1 U24096 ( .A(n21135), .ZN(n21137) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21456), .ZN(n21136) );
  OAI211_X1 U24098 ( .C1(n21459), .C2(n21193), .A(n21137), .B(n21136), .ZN(
        P1_U3099) );
  OAI22_X1 U24099 ( .A1(n21461), .A2(n21151), .B1(n21460), .B2(n21150), .ZN(
        n21138) );
  INV_X1 U24100 ( .A(n21138), .ZN(n21140) );
  AOI22_X1 U24101 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21463), .ZN(n21139) );
  OAI211_X1 U24102 ( .C1(n9779), .C2(n21193), .A(n21140), .B(n21139), .ZN(
        P1_U3100) );
  OAI22_X1 U24103 ( .A1(n21468), .A2(n21151), .B1(n21467), .B2(n21150), .ZN(
        n21141) );
  INV_X1 U24104 ( .A(n21141), .ZN(n21143) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21470), .ZN(n21142) );
  OAI211_X1 U24106 ( .C1(n21473), .C2(n21193), .A(n21143), .B(n21142), .ZN(
        P1_U3101) );
  OAI22_X1 U24107 ( .A1(n21475), .A2(n21151), .B1(n21474), .B2(n21150), .ZN(
        n21144) );
  INV_X1 U24108 ( .A(n21144), .ZN(n21146) );
  AOI22_X1 U24109 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21477), .ZN(n21145) );
  OAI211_X1 U24110 ( .C1(n21480), .C2(n21193), .A(n21146), .B(n21145), .ZN(
        P1_U3102) );
  OAI22_X1 U24111 ( .A1(n21482), .A2(n21151), .B1(n21481), .B2(n21150), .ZN(
        n21147) );
  INV_X1 U24112 ( .A(n21147), .ZN(n21149) );
  AOI22_X1 U24113 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21484), .ZN(n21148) );
  OAI211_X1 U24114 ( .C1(n21487), .C2(n21193), .A(n21149), .B(n21148), .ZN(
        P1_U3103) );
  OAI22_X1 U24115 ( .A1(n21491), .A2(n21151), .B1(n21488), .B2(n21150), .ZN(
        n21152) );
  INV_X1 U24116 ( .A(n21152), .ZN(n21156) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21154), .B1(
        n21153), .B2(n21493), .ZN(n21155) );
  OAI211_X1 U24118 ( .C1(n21499), .C2(n21193), .A(n21156), .B(n21155), .ZN(
        P1_U3104) );
  OR2_X1 U24119 ( .A1(n21236), .A2(n20854), .ZN(n21158) );
  OR2_X1 U24120 ( .A1(n21327), .A2(n21157), .ZN(n21186) );
  NAND2_X1 U24121 ( .A1(n21158), .A2(n21186), .ZN(n21162) );
  NAND2_X1 U24122 ( .A1(n21162), .A2(n9585), .ZN(n21160) );
  NAND2_X1 U24123 ( .A1(n21165), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21159) );
  OAI22_X1 U24124 ( .A1(n21430), .A2(n21187), .B1(n21429), .B2(n21186), .ZN(
        n21161) );
  INV_X1 U24125 ( .A(n21161), .ZN(n21167) );
  INV_X1 U24126 ( .A(n21233), .ZN(n21242) );
  AOI21_X1 U24127 ( .B1(n9585), .B2(n21373), .A(n21242), .ZN(n21163) );
  OR2_X1 U24128 ( .A1(n21163), .A2(n21162), .ZN(n21164) );
  OAI211_X1 U24129 ( .C1(n9585), .C2(n21165), .A(n21439), .B(n21164), .ZN(
        n21190) );
  AOI22_X1 U24130 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21382), .ZN(n21166) );
  OAI211_X1 U24131 ( .C1(n21385), .C2(n21193), .A(n21167), .B(n21166), .ZN(
        P1_U3105) );
  OAI22_X1 U24132 ( .A1(n21447), .A2(n21187), .B1(n21446), .B2(n21186), .ZN(
        n21168) );
  INV_X1 U24133 ( .A(n21168), .ZN(n21170) );
  AOI22_X1 U24134 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21387), .ZN(n21169) );
  OAI211_X1 U24135 ( .C1(n21390), .C2(n21193), .A(n21170), .B(n21169), .ZN(
        P1_U3106) );
  OAI22_X1 U24136 ( .A1(n21454), .A2(n21187), .B1(n21453), .B2(n21186), .ZN(
        n21171) );
  INV_X1 U24137 ( .A(n21171), .ZN(n21173) );
  AOI22_X1 U24138 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21392), .ZN(n21172) );
  OAI211_X1 U24139 ( .C1(n21395), .C2(n21193), .A(n21173), .B(n21172), .ZN(
        P1_U3107) );
  OAI22_X1 U24140 ( .A1(n21461), .A2(n21187), .B1(n21460), .B2(n21186), .ZN(
        n21174) );
  INV_X1 U24141 ( .A(n21174), .ZN(n21176) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n9778), .ZN(n21175) );
  OAI211_X1 U24143 ( .C1(n21399), .C2(n21193), .A(n21176), .B(n21175), .ZN(
        P1_U3108) );
  OAI22_X1 U24144 ( .A1(n21468), .A2(n21187), .B1(n21467), .B2(n21186), .ZN(
        n21177) );
  INV_X1 U24145 ( .A(n21177), .ZN(n21179) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21401), .ZN(n21178) );
  OAI211_X1 U24147 ( .C1(n21404), .C2(n21193), .A(n21179), .B(n21178), .ZN(
        P1_U3109) );
  OAI22_X1 U24148 ( .A1(n21475), .A2(n21187), .B1(n21474), .B2(n21186), .ZN(
        n21180) );
  INV_X1 U24149 ( .A(n21180), .ZN(n21182) );
  AOI22_X1 U24150 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21406), .ZN(n21181) );
  OAI211_X1 U24151 ( .C1(n21409), .C2(n21193), .A(n21182), .B(n21181), .ZN(
        P1_U3110) );
  OAI22_X1 U24152 ( .A1(n21482), .A2(n21187), .B1(n21481), .B2(n21186), .ZN(
        n21183) );
  INV_X1 U24153 ( .A(n21183), .ZN(n21185) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21411), .ZN(n21184) );
  OAI211_X1 U24155 ( .C1(n21414), .C2(n21193), .A(n21185), .B(n21184), .ZN(
        P1_U3111) );
  OAI22_X1 U24156 ( .A1(n21491), .A2(n21187), .B1(n21488), .B2(n21186), .ZN(
        n21188) );
  INV_X1 U24157 ( .A(n21188), .ZN(n21192) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21190), .B1(
        n21189), .B2(n21418), .ZN(n21191) );
  OAI211_X1 U24159 ( .C1(n21423), .C2(n21193), .A(n21192), .B(n21191), .ZN(
        P1_U3112) );
  NOR3_X1 U24160 ( .A1(n21275), .A2(n21195), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21243) );
  NAND2_X1 U24161 ( .A1(n21327), .A2(n21243), .ZN(n21225) );
  OAI22_X1 U24162 ( .A1(n21231), .A2(n21385), .B1(n21225), .B2(n21429), .ZN(
        n21196) );
  INV_X1 U24163 ( .A(n21196), .ZN(n21206) );
  AOI21_X1 U24164 ( .B1(n21273), .B2(n21231), .A(n21373), .ZN(n21197) );
  NOR2_X1 U24165 ( .A1(n21197), .A2(n21433), .ZN(n21201) );
  OR2_X1 U24166 ( .A1(n21236), .A2(n14245), .ZN(n21203) );
  AOI22_X1 U24167 ( .A1(n21201), .A2(n21203), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21225), .ZN(n21199) );
  OR2_X1 U24168 ( .A1(n21198), .A2(n21275), .ZN(n21364) );
  NAND2_X1 U24169 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21364), .ZN(n21377) );
  NAND3_X1 U24170 ( .A1(n21200), .A2(n21199), .A3(n21377), .ZN(n21228) );
  INV_X1 U24171 ( .A(n21201), .ZN(n21204) );
  AOI22_X1 U24172 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21228), .B1(
        n21289), .B2(n21227), .ZN(n21205) );
  OAI211_X1 U24173 ( .C1(n21445), .C2(n21273), .A(n21206), .B(n21205), .ZN(
        P1_U3113) );
  OAI22_X1 U24174 ( .A1(n21273), .A2(n21452), .B1(n21446), .B2(n21225), .ZN(
        n21207) );
  INV_X1 U24175 ( .A(n21207), .ZN(n21209) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21228), .B1(
        n21293), .B2(n21227), .ZN(n21208) );
  OAI211_X1 U24177 ( .C1(n21390), .C2(n21231), .A(n21209), .B(n21208), .ZN(
        P1_U3114) );
  OAI22_X1 U24178 ( .A1(n21231), .A2(n21395), .B1(n21225), .B2(n21453), .ZN(
        n21210) );
  INV_X1 U24179 ( .A(n21210), .ZN(n21212) );
  AOI22_X1 U24180 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21228), .B1(
        n21297), .B2(n21227), .ZN(n21211) );
  OAI211_X1 U24181 ( .C1(n21459), .C2(n21273), .A(n21212), .B(n21211), .ZN(
        P1_U3115) );
  OAI22_X1 U24182 ( .A1(n21231), .A2(n21399), .B1(n21225), .B2(n21460), .ZN(
        n21213) );
  INV_X1 U24183 ( .A(n21213), .ZN(n21215) );
  AOI22_X1 U24184 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21228), .B1(
        n21301), .B2(n21227), .ZN(n21214) );
  OAI211_X1 U24185 ( .C1(n9779), .C2(n21273), .A(n21215), .B(n21214), .ZN(
        P1_U3116) );
  OAI22_X1 U24186 ( .A1(n21273), .A2(n21473), .B1(n21225), .B2(n21467), .ZN(
        n21216) );
  INV_X1 U24187 ( .A(n21216), .ZN(n21218) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21228), .B1(
        n21305), .B2(n21227), .ZN(n21217) );
  OAI211_X1 U24189 ( .C1(n21404), .C2(n21231), .A(n21218), .B(n21217), .ZN(
        P1_U3117) );
  OAI22_X1 U24190 ( .A1(n21231), .A2(n21409), .B1(n21225), .B2(n21474), .ZN(
        n21219) );
  INV_X1 U24191 ( .A(n21219), .ZN(n21221) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21228), .B1(
        n21309), .B2(n21227), .ZN(n21220) );
  OAI211_X1 U24193 ( .C1(n21480), .C2(n21273), .A(n21221), .B(n21220), .ZN(
        P1_U3118) );
  OAI22_X1 U24194 ( .A1(n21231), .A2(n21414), .B1(n21225), .B2(n21481), .ZN(
        n21222) );
  INV_X1 U24195 ( .A(n21222), .ZN(n21224) );
  AOI22_X1 U24196 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21228), .B1(
        n21313), .B2(n21227), .ZN(n21223) );
  OAI211_X1 U24197 ( .C1(n21487), .C2(n21273), .A(n21224), .B(n21223), .ZN(
        P1_U3119) );
  OAI22_X1 U24198 ( .A1(n21273), .A2(n21499), .B1(n21225), .B2(n21488), .ZN(
        n21226) );
  INV_X1 U24199 ( .A(n21226), .ZN(n21230) );
  AOI22_X1 U24200 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21228), .B1(
        n21319), .B2(n21227), .ZN(n21229) );
  OAI211_X1 U24201 ( .C1(n21423), .C2(n21231), .A(n21230), .B(n21229), .ZN(
        P1_U3120) );
  NAND2_X1 U24202 ( .A1(n21234), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21266) );
  OAI21_X1 U24203 ( .B1(n21236), .B2(n21235), .A(n21266), .ZN(n21237) );
  NAND2_X1 U24204 ( .A1(n21237), .A2(n9585), .ZN(n21239) );
  NAND2_X1 U24205 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21243), .ZN(n21238) );
  OAI22_X1 U24206 ( .A1(n21430), .A2(n21267), .B1(n21429), .B2(n21266), .ZN(
        n21240) );
  INV_X1 U24207 ( .A(n21240), .ZN(n21246) );
  NOR2_X1 U24208 ( .A1(n21242), .A2(n21241), .ZN(n21244) );
  INV_X1 U24209 ( .A(n21273), .ZN(n21263) );
  AOI22_X1 U24210 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n21263), .B2(n21442), .ZN(n21245) );
  OAI211_X1 U24211 ( .C1(n21445), .C2(n21323), .A(n21246), .B(n21245), .ZN(
        P1_U3121) );
  OAI22_X1 U24212 ( .A1(n21447), .A2(n21267), .B1(n21446), .B2(n21266), .ZN(
        n21247) );
  INV_X1 U24213 ( .A(n21247), .ZN(n21249) );
  AOI22_X1 U24214 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n21263), .B2(n21449), .ZN(n21248) );
  OAI211_X1 U24215 ( .C1(n21452), .C2(n21323), .A(n21249), .B(n21248), .ZN(
        P1_U3122) );
  OAI22_X1 U24216 ( .A1(n21454), .A2(n21267), .B1(n21453), .B2(n21266), .ZN(
        n21250) );
  INV_X1 U24217 ( .A(n21250), .ZN(n21252) );
  INV_X1 U24218 ( .A(n21323), .ZN(n21269) );
  AOI22_X1 U24219 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n21269), .B2(n21392), .ZN(n21251) );
  OAI211_X1 U24220 ( .C1(n21395), .C2(n21273), .A(n21252), .B(n21251), .ZN(
        P1_U3123) );
  OAI22_X1 U24221 ( .A1(n21461), .A2(n21267), .B1(n21460), .B2(n21266), .ZN(
        n21253) );
  INV_X1 U24222 ( .A(n21253), .ZN(n21255) );
  AOI22_X1 U24223 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n21269), .B2(n9778), .ZN(n21254) );
  OAI211_X1 U24224 ( .C1(n21399), .C2(n21273), .A(n21255), .B(n21254), .ZN(
        P1_U3124) );
  OAI22_X1 U24225 ( .A1(n21468), .A2(n21267), .B1(n21467), .B2(n21266), .ZN(
        n21256) );
  INV_X1 U24226 ( .A(n21256), .ZN(n21258) );
  AOI22_X1 U24227 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n21263), .B2(n21470), .ZN(n21257) );
  OAI211_X1 U24228 ( .C1(n21473), .C2(n21323), .A(n21258), .B(n21257), .ZN(
        P1_U3125) );
  OAI22_X1 U24229 ( .A1(n21475), .A2(n21267), .B1(n21474), .B2(n21266), .ZN(
        n21259) );
  INV_X1 U24230 ( .A(n21259), .ZN(n21261) );
  AOI22_X1 U24231 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n21269), .B2(n21406), .ZN(n21260) );
  OAI211_X1 U24232 ( .C1(n21409), .C2(n21273), .A(n21261), .B(n21260), .ZN(
        P1_U3126) );
  OAI22_X1 U24233 ( .A1(n21482), .A2(n21267), .B1(n21481), .B2(n21266), .ZN(
        n21262) );
  INV_X1 U24234 ( .A(n21262), .ZN(n21265) );
  AOI22_X1 U24235 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n21263), .B2(n21484), .ZN(n21264) );
  OAI211_X1 U24236 ( .C1(n21487), .C2(n21323), .A(n21265), .B(n21264), .ZN(
        P1_U3127) );
  OAI22_X1 U24237 ( .A1(n21491), .A2(n21267), .B1(n21488), .B2(n21266), .ZN(
        n21268) );
  INV_X1 U24238 ( .A(n21268), .ZN(n21272) );
  AOI22_X1 U24239 ( .A1(n21270), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n21269), .B2(n21418), .ZN(n21271) );
  OAI211_X1 U24240 ( .C1(n21423), .C2(n21273), .A(n21272), .B(n21271), .ZN(
        P1_U3128) );
  NOR3_X1 U24241 ( .A1(n21276), .A2(n21275), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21335) );
  INV_X1 U24242 ( .A(n21335), .ZN(n21326) );
  NOR2_X1 U24243 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21326), .ZN(
        n21283) );
  OAI22_X1 U24244 ( .A1(n21336), .A2(n21445), .B1(n21429), .B2(n21316), .ZN(
        n21277) );
  INV_X1 U24245 ( .A(n21277), .ZN(n21291) );
  AOI21_X1 U24246 ( .B1(n21323), .B2(n21336), .A(n21373), .ZN(n21278) );
  NOR2_X1 U24247 ( .A1(n21278), .A2(n21433), .ZN(n21284) );
  NAND2_X1 U24248 ( .A1(n21425), .A2(n14245), .ZN(n21287) );
  INV_X1 U24249 ( .A(n21280), .ZN(n21285) );
  AOI22_X1 U24250 ( .A1(n21284), .A2(n21287), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21285), .ZN(n21281) );
  OAI211_X1 U24251 ( .C1(n21283), .C2(n21282), .A(n21378), .B(n21281), .ZN(
        n21320) );
  INV_X1 U24252 ( .A(n21284), .ZN(n21288) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21320), .B1(
        n21289), .B2(n21318), .ZN(n21290) );
  OAI211_X1 U24254 ( .C1(n21385), .C2(n21323), .A(n21291), .B(n21290), .ZN(
        P1_U3129) );
  OAI22_X1 U24255 ( .A1(n21336), .A2(n21452), .B1(n21446), .B2(n21316), .ZN(
        n21292) );
  INV_X1 U24256 ( .A(n21292), .ZN(n21295) );
  AOI22_X1 U24257 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21320), .B1(
        n21293), .B2(n21318), .ZN(n21294) );
  OAI211_X1 U24258 ( .C1(n21390), .C2(n21323), .A(n21295), .B(n21294), .ZN(
        P1_U3130) );
  OAI22_X1 U24259 ( .A1(n21336), .A2(n21459), .B1(n21453), .B2(n21316), .ZN(
        n21296) );
  INV_X1 U24260 ( .A(n21296), .ZN(n21299) );
  AOI22_X1 U24261 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21320), .B1(
        n21297), .B2(n21318), .ZN(n21298) );
  OAI211_X1 U24262 ( .C1(n21395), .C2(n21323), .A(n21299), .B(n21298), .ZN(
        P1_U3131) );
  OAI22_X1 U24263 ( .A1(n21336), .A2(n9779), .B1(n21460), .B2(n21316), .ZN(
        n21300) );
  INV_X1 U24264 ( .A(n21300), .ZN(n21303) );
  AOI22_X1 U24265 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21320), .B1(
        n21301), .B2(n21318), .ZN(n21302) );
  OAI211_X1 U24266 ( .C1(n21399), .C2(n21323), .A(n21303), .B(n21302), .ZN(
        P1_U3132) );
  OAI22_X1 U24267 ( .A1(n21336), .A2(n21473), .B1(n21467), .B2(n21316), .ZN(
        n21304) );
  INV_X1 U24268 ( .A(n21304), .ZN(n21307) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21320), .B1(
        n21305), .B2(n21318), .ZN(n21306) );
  OAI211_X1 U24270 ( .C1(n21404), .C2(n21323), .A(n21307), .B(n21306), .ZN(
        P1_U3133) );
  OAI22_X1 U24271 ( .A1(n21336), .A2(n21480), .B1(n21474), .B2(n21316), .ZN(
        n21308) );
  INV_X1 U24272 ( .A(n21308), .ZN(n21311) );
  AOI22_X1 U24273 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21320), .B1(
        n21309), .B2(n21318), .ZN(n21310) );
  OAI211_X1 U24274 ( .C1(n21409), .C2(n21323), .A(n21311), .B(n21310), .ZN(
        P1_U3134) );
  OAI22_X1 U24275 ( .A1(n21336), .A2(n21487), .B1(n21481), .B2(n21316), .ZN(
        n21312) );
  INV_X1 U24276 ( .A(n21312), .ZN(n21315) );
  AOI22_X1 U24277 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21320), .B1(
        n21313), .B2(n21318), .ZN(n21314) );
  OAI211_X1 U24278 ( .C1(n21414), .C2(n21323), .A(n21315), .B(n21314), .ZN(
        P1_U3135) );
  OAI22_X1 U24279 ( .A1(n21336), .A2(n21499), .B1(n21488), .B2(n21316), .ZN(
        n21317) );
  INV_X1 U24280 ( .A(n21317), .ZN(n21322) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21320), .B1(
        n21319), .B2(n21318), .ZN(n21321) );
  OAI211_X1 U24282 ( .C1(n21423), .C2(n21323), .A(n21322), .B(n21321), .ZN(
        P1_U3136) );
  NAND2_X1 U24283 ( .A1(n21425), .A2(n21325), .ZN(n21328) );
  OR2_X1 U24284 ( .A1(n21327), .A2(n21326), .ZN(n21357) );
  NAND2_X1 U24285 ( .A1(n21328), .A2(n21357), .ZN(n21332) );
  NAND2_X1 U24286 ( .A1(n21332), .A2(n9585), .ZN(n21330) );
  NAND2_X1 U24287 ( .A1(n21335), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21329) );
  OAI22_X1 U24288 ( .A1(n21430), .A2(n21358), .B1(n21429), .B2(n21357), .ZN(
        n21331) );
  INV_X1 U24289 ( .A(n21331), .ZN(n21338) );
  INV_X1 U24290 ( .A(n21332), .ZN(n21333) );
  OAI211_X1 U24291 ( .C1(n21372), .C2(n21373), .A(n9585), .B(n21333), .ZN(
        n21334) );
  OAI211_X1 U24292 ( .C1(n9585), .C2(n21335), .A(n21439), .B(n21334), .ZN(
        n21361) );
  AOI22_X1 U24293 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21442), .ZN(n21337) );
  OAI211_X1 U24294 ( .C1(n21445), .C2(n21422), .A(n21338), .B(n21337), .ZN(
        P1_U3137) );
  OAI22_X1 U24295 ( .A1(n21447), .A2(n21358), .B1(n21446), .B2(n21357), .ZN(
        n21339) );
  INV_X1 U24296 ( .A(n21339), .ZN(n21341) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21449), .ZN(n21340) );
  OAI211_X1 U24298 ( .C1(n21452), .C2(n21422), .A(n21341), .B(n21340), .ZN(
        P1_U3138) );
  OAI22_X1 U24299 ( .A1(n21454), .A2(n21358), .B1(n21453), .B2(n21357), .ZN(
        n21342) );
  INV_X1 U24300 ( .A(n21342), .ZN(n21344) );
  AOI22_X1 U24301 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21456), .ZN(n21343) );
  OAI211_X1 U24302 ( .C1(n21459), .C2(n21422), .A(n21344), .B(n21343), .ZN(
        P1_U3139) );
  OAI22_X1 U24303 ( .A1(n21461), .A2(n21358), .B1(n21460), .B2(n21357), .ZN(
        n21345) );
  INV_X1 U24304 ( .A(n21345), .ZN(n21347) );
  AOI22_X1 U24305 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21463), .ZN(n21346) );
  OAI211_X1 U24306 ( .C1(n9779), .C2(n21422), .A(n21347), .B(n21346), .ZN(
        P1_U3140) );
  OAI22_X1 U24307 ( .A1(n21468), .A2(n21358), .B1(n21467), .B2(n21357), .ZN(
        n21348) );
  INV_X1 U24308 ( .A(n21348), .ZN(n21350) );
  AOI22_X1 U24309 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21470), .ZN(n21349) );
  OAI211_X1 U24310 ( .C1(n21473), .C2(n21422), .A(n21350), .B(n21349), .ZN(
        P1_U3141) );
  OAI22_X1 U24311 ( .A1(n21475), .A2(n21358), .B1(n21474), .B2(n21357), .ZN(
        n21351) );
  INV_X1 U24312 ( .A(n21351), .ZN(n21353) );
  AOI22_X1 U24313 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21477), .ZN(n21352) );
  OAI211_X1 U24314 ( .C1(n21480), .C2(n21422), .A(n21353), .B(n21352), .ZN(
        P1_U3142) );
  OAI22_X1 U24315 ( .A1(n21482), .A2(n21358), .B1(n21481), .B2(n21357), .ZN(
        n21354) );
  INV_X1 U24316 ( .A(n21354), .ZN(n21356) );
  AOI22_X1 U24317 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21484), .ZN(n21355) );
  OAI211_X1 U24318 ( .C1(n21487), .C2(n21422), .A(n21356), .B(n21355), .ZN(
        P1_U3143) );
  OAI22_X1 U24319 ( .A1(n21491), .A2(n21358), .B1(n21488), .B2(n21357), .ZN(
        n21359) );
  INV_X1 U24320 ( .A(n21359), .ZN(n21363) );
  AOI22_X1 U24321 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21361), .B1(
        n21360), .B2(n21493), .ZN(n21362) );
  OAI211_X1 U24322 ( .C1(n21499), .C2(n21422), .A(n21363), .B(n21362), .ZN(
        P1_U3144) );
  NAND3_X1 U24323 ( .A1(n21425), .A2(n21375), .A3(n9585), .ZN(n21368) );
  INV_X1 U24324 ( .A(n21364), .ZN(n21365) );
  NAND2_X1 U24325 ( .A1(n21366), .A2(n21365), .ZN(n21367) );
  INV_X1 U24326 ( .A(n21441), .ZN(n21369) );
  NOR2_X1 U24327 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21369), .ZN(
        n21380) );
  INV_X1 U24328 ( .A(n21380), .ZN(n21415) );
  OAI22_X1 U24329 ( .A1(n21430), .A2(n21416), .B1(n21429), .B2(n21415), .ZN(
        n21370) );
  INV_X1 U24330 ( .A(n21370), .ZN(n21384) );
  AOI21_X1 U24331 ( .B1(n21422), .B2(n21381), .A(n21373), .ZN(n21374) );
  AOI21_X1 U24332 ( .B1(n21425), .B2(n21375), .A(n21374), .ZN(n21376) );
  NOR2_X1 U24333 ( .A1(n21376), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21379) );
  AOI22_X1 U24334 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21382), .ZN(n21383) );
  OAI211_X1 U24335 ( .C1(n21385), .C2(n21422), .A(n21384), .B(n21383), .ZN(
        P1_U3145) );
  OAI22_X1 U24336 ( .A1(n21447), .A2(n21416), .B1(n21446), .B2(n21415), .ZN(
        n21386) );
  INV_X1 U24337 ( .A(n21386), .ZN(n21389) );
  AOI22_X1 U24338 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21387), .ZN(n21388) );
  OAI211_X1 U24339 ( .C1(n21390), .C2(n21422), .A(n21389), .B(n21388), .ZN(
        P1_U3146) );
  OAI22_X1 U24340 ( .A1(n21454), .A2(n21416), .B1(n21453), .B2(n21415), .ZN(
        n21391) );
  INV_X1 U24341 ( .A(n21391), .ZN(n21394) );
  AOI22_X1 U24342 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21392), .ZN(n21393) );
  OAI211_X1 U24343 ( .C1(n21395), .C2(n21422), .A(n21394), .B(n21393), .ZN(
        P1_U3147) );
  OAI22_X1 U24344 ( .A1(n21461), .A2(n21416), .B1(n21460), .B2(n21415), .ZN(
        n21396) );
  INV_X1 U24345 ( .A(n21396), .ZN(n21398) );
  AOI22_X1 U24346 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n9778), .ZN(n21397) );
  OAI211_X1 U24347 ( .C1(n21399), .C2(n21422), .A(n21398), .B(n21397), .ZN(
        P1_U3148) );
  OAI22_X1 U24348 ( .A1(n21468), .A2(n21416), .B1(n21467), .B2(n21415), .ZN(
        n21400) );
  INV_X1 U24349 ( .A(n21400), .ZN(n21403) );
  AOI22_X1 U24350 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21401), .ZN(n21402) );
  OAI211_X1 U24351 ( .C1(n21404), .C2(n21422), .A(n21403), .B(n21402), .ZN(
        P1_U3149) );
  OAI22_X1 U24352 ( .A1(n21475), .A2(n21416), .B1(n21474), .B2(n21415), .ZN(
        n21405) );
  INV_X1 U24353 ( .A(n21405), .ZN(n21408) );
  AOI22_X1 U24354 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21406), .ZN(n21407) );
  OAI211_X1 U24355 ( .C1(n21409), .C2(n21422), .A(n21408), .B(n21407), .ZN(
        P1_U3150) );
  OAI22_X1 U24356 ( .A1(n21482), .A2(n21416), .B1(n21481), .B2(n21415), .ZN(
        n21410) );
  INV_X1 U24357 ( .A(n21410), .ZN(n21413) );
  AOI22_X1 U24358 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21411), .ZN(n21412) );
  OAI211_X1 U24359 ( .C1(n21414), .C2(n21422), .A(n21413), .B(n21412), .ZN(
        P1_U3151) );
  OAI22_X1 U24360 ( .A1(n21491), .A2(n21416), .B1(n21488), .B2(n21415), .ZN(
        n21417) );
  INV_X1 U24361 ( .A(n21417), .ZN(n21421) );
  AOI22_X1 U24362 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21419), .B1(
        n21494), .B2(n21418), .ZN(n21420) );
  OAI211_X1 U24363 ( .C1(n21423), .C2(n21422), .A(n21421), .B(n21420), .ZN(
        P1_U3152) );
  NAND2_X1 U24364 ( .A1(n21425), .A2(n21424), .ZN(n21426) );
  NAND2_X1 U24365 ( .A1(n21426), .A2(n21489), .ZN(n21435) );
  NAND2_X1 U24366 ( .A1(n21435), .A2(n9585), .ZN(n21428) );
  NAND2_X1 U24367 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21441), .ZN(n21427) );
  OAI22_X1 U24368 ( .A1(n21430), .A2(n21490), .B1(n21489), .B2(n21429), .ZN(
        n21431) );
  INV_X1 U24369 ( .A(n21431), .ZN(n21444) );
  OAI21_X1 U24370 ( .B1(n21434), .B2(n21433), .A(n21432), .ZN(n21437) );
  INV_X1 U24371 ( .A(n21435), .ZN(n21436) );
  NAND2_X1 U24372 ( .A1(n21437), .A2(n21436), .ZN(n21438) );
  OAI211_X1 U24373 ( .C1(n21441), .C2(n9585), .A(n21439), .B(n21438), .ZN(
        n21495) );
  AOI22_X1 U24374 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21442), .ZN(n21443) );
  OAI211_X1 U24375 ( .C1(n21445), .C2(n21498), .A(n21444), .B(n21443), .ZN(
        P1_U3153) );
  OAI22_X1 U24376 ( .A1(n21447), .A2(n21490), .B1(n21489), .B2(n21446), .ZN(
        n21448) );
  INV_X1 U24377 ( .A(n21448), .ZN(n21451) );
  AOI22_X1 U24378 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21449), .ZN(n21450) );
  OAI211_X1 U24379 ( .C1(n21452), .C2(n21498), .A(n21451), .B(n21450), .ZN(
        P1_U3154) );
  OAI22_X1 U24380 ( .A1(n21454), .A2(n21490), .B1(n21489), .B2(n21453), .ZN(
        n21455) );
  INV_X1 U24381 ( .A(n21455), .ZN(n21458) );
  AOI22_X1 U24382 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21456), .ZN(n21457) );
  OAI211_X1 U24383 ( .C1(n21459), .C2(n21498), .A(n21458), .B(n21457), .ZN(
        P1_U3155) );
  OAI22_X1 U24384 ( .A1(n21461), .A2(n21490), .B1(n21489), .B2(n21460), .ZN(
        n21462) );
  INV_X1 U24385 ( .A(n21462), .ZN(n21465) );
  AOI22_X1 U24386 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21463), .ZN(n21464) );
  OAI211_X1 U24387 ( .C1(n9779), .C2(n21498), .A(n21465), .B(n21464), .ZN(
        P1_U3156) );
  OAI22_X1 U24388 ( .A1(n21468), .A2(n21490), .B1(n21489), .B2(n21467), .ZN(
        n21469) );
  INV_X1 U24389 ( .A(n21469), .ZN(n21472) );
  AOI22_X1 U24390 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21470), .ZN(n21471) );
  OAI211_X1 U24391 ( .C1(n21473), .C2(n21498), .A(n21472), .B(n21471), .ZN(
        P1_U3157) );
  OAI22_X1 U24392 ( .A1(n21475), .A2(n21490), .B1(n21489), .B2(n21474), .ZN(
        n21476) );
  INV_X1 U24393 ( .A(n21476), .ZN(n21479) );
  AOI22_X1 U24394 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21477), .ZN(n21478) );
  OAI211_X1 U24395 ( .C1(n21480), .C2(n21498), .A(n21479), .B(n21478), .ZN(
        P1_U3158) );
  OAI22_X1 U24396 ( .A1(n21482), .A2(n21490), .B1(n21489), .B2(n21481), .ZN(
        n21483) );
  INV_X1 U24397 ( .A(n21483), .ZN(n21486) );
  AOI22_X1 U24398 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21484), .ZN(n21485) );
  OAI211_X1 U24399 ( .C1(n21487), .C2(n21498), .A(n21486), .B(n21485), .ZN(
        P1_U3159) );
  OAI22_X1 U24400 ( .A1(n21491), .A2(n21490), .B1(n21489), .B2(n21488), .ZN(
        n21492) );
  INV_X1 U24401 ( .A(n21492), .ZN(n21497) );
  AOI22_X1 U24402 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21493), .ZN(n21496) );
  OAI211_X1 U24403 ( .C1(n21499), .C2(n21498), .A(n21497), .B(n21496), .ZN(
        P1_U3160) );
  NOR2_X1 U24404 ( .A1(n21501), .A2(n21500), .ZN(n21504) );
  OAI21_X1 U24405 ( .B1(n21504), .B2(n21503), .A(n21502), .ZN(P1_U3163) );
  AND2_X1 U24406 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21505), .ZN(
        P1_U3164) );
  AND2_X1 U24407 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21505), .ZN(
        P1_U3165) );
  AND2_X1 U24408 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21505), .ZN(
        P1_U3166) );
  AND2_X1 U24409 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21505), .ZN(
        P1_U3167) );
  AND2_X1 U24410 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21505), .ZN(
        P1_U3168) );
  AND2_X1 U24411 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21505), .ZN(
        P1_U3169) );
  AND2_X1 U24412 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21505), .ZN(
        P1_U3170) );
  AND2_X1 U24413 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21505), .ZN(
        P1_U3171) );
  AND2_X1 U24414 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21505), .ZN(
        P1_U3172) );
  AND2_X1 U24415 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21505), .ZN(
        P1_U3173) );
  AND2_X1 U24416 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21505), .ZN(
        P1_U3174) );
  AND2_X1 U24417 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21505), .ZN(
        P1_U3175) );
  AND2_X1 U24418 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21505), .ZN(
        P1_U3176) );
  AND2_X1 U24419 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21505), .ZN(
        P1_U3177) );
  AND2_X1 U24420 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21505), .ZN(
        P1_U3178) );
  AND2_X1 U24421 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21505), .ZN(
        P1_U3179) );
  AND2_X1 U24422 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21505), .ZN(
        P1_U3180) );
  AND2_X1 U24423 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21505), .ZN(
        P1_U3181) );
  AND2_X1 U24424 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21505), .ZN(
        P1_U3182) );
  AND2_X1 U24425 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21505), .ZN(
        P1_U3183) );
  AND2_X1 U24426 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21505), .ZN(
        P1_U3184) );
  AND2_X1 U24427 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21505), .ZN(
        P1_U3185) );
  AND2_X1 U24428 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21505), .ZN(P1_U3186) );
  AND2_X1 U24429 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21505), .ZN(P1_U3187) );
  AND2_X1 U24430 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21505), .ZN(P1_U3188) );
  AND2_X1 U24431 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21505), .ZN(P1_U3189) );
  AND2_X1 U24432 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21505), .ZN(P1_U3190) );
  AND2_X1 U24433 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21505), .ZN(P1_U3191) );
  AND2_X1 U24434 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21505), .ZN(P1_U3192) );
  AND2_X1 U24435 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21505), .ZN(P1_U3193) );
  NAND2_X1 U24436 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21510), .ZN(n21516) );
  INV_X1 U24437 ( .A(n21516), .ZN(n21509) );
  NOR2_X1 U24438 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21506) );
  OAI21_X1 U24439 ( .B1(n21506), .B2(n21512), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21507) );
  AOI21_X1 U24440 ( .B1(NA), .B2(n21511), .A(n21507), .ZN(n21508) );
  OAI22_X1 U24441 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21509), .B1(n21579), 
        .B2(n21508), .ZN(P1_U3194) );
  NOR3_X1 U24442 ( .A1(NA), .A2(n21511), .A3(n21510), .ZN(n21515) );
  AOI21_X1 U24443 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n21520), .A(n21512), .ZN(n21514) );
  AOI222_X1 U24444 ( .A1(n21515), .A2(n21514), .B1(n21515), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n21514), .C2(n21513), .ZN(n21519)
         );
  OAI211_X1 U24445 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21517), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21516), .ZN(n21518) );
  NAND2_X1 U24446 ( .A1(n21519), .A2(n21518), .ZN(P1_U3196) );
  OR2_X1 U24447 ( .A1(n21577), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21546) );
  INV_X1 U24448 ( .A(n21546), .ZN(n21559) );
  INV_X1 U24449 ( .A(n21543), .ZN(n21560) );
  AOI222_X1 U24450 ( .A1(n21559), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21560), .ZN(n21521) );
  INV_X1 U24451 ( .A(n21521), .ZN(P1_U3197) );
  AOI222_X1 U24452 ( .A1(n21560), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21559), .ZN(n21522) );
  INV_X1 U24453 ( .A(n21522), .ZN(P1_U3198) );
  INV_X1 U24454 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21525) );
  OAI222_X1 U24455 ( .A1(n21543), .A2(n21525), .B1(n21524), .B2(n21579), .C1(
        n21523), .C2(n21546), .ZN(P1_U3199) );
  AOI222_X1 U24456 ( .A1(n21559), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21560), .ZN(n21526) );
  INV_X1 U24457 ( .A(n21526), .ZN(P1_U3200) );
  AOI222_X1 U24458 ( .A1(n21560), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21559), .ZN(n21527) );
  INV_X1 U24459 ( .A(n21527), .ZN(P1_U3201) );
  AOI222_X1 U24460 ( .A1(n21560), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21559), .ZN(n21528) );
  INV_X1 U24461 ( .A(n21528), .ZN(P1_U3202) );
  AOI222_X1 U24462 ( .A1(n21560), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21559), .ZN(n21529) );
  INV_X1 U24463 ( .A(n21529), .ZN(P1_U3203) );
  AOI222_X1 U24464 ( .A1(n21560), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n21559), .ZN(n21530) );
  INV_X1 U24465 ( .A(n21530), .ZN(P1_U3204) );
  AOI222_X1 U24466 ( .A1(n21560), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21559), .ZN(n21531) );
  INV_X1 U24467 ( .A(n21531), .ZN(P1_U3205) );
  AOI222_X1 U24468 ( .A1(n21559), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21560), .ZN(n21532) );
  INV_X1 U24469 ( .A(n21532), .ZN(P1_U3206) );
  AOI22_X1 U24470 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21559), .ZN(n21533) );
  OAI21_X1 U24471 ( .B1(n21534), .B2(n21543), .A(n21533), .ZN(P1_U3207) );
  AOI22_X1 U24472 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21560), .ZN(n21535) );
  OAI21_X1 U24473 ( .B1(n21537), .B2(n21546), .A(n21535), .ZN(P1_U3208) );
  AOI22_X1 U24474 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21559), .ZN(n21536) );
  OAI21_X1 U24475 ( .B1(n21537), .B2(n21543), .A(n21536), .ZN(P1_U3209) );
  AOI22_X1 U24476 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21560), .ZN(n21538) );
  OAI21_X1 U24477 ( .B1(n21540), .B2(n21546), .A(n21538), .ZN(P1_U3210) );
  AOI22_X1 U24478 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21559), .ZN(n21539) );
  OAI21_X1 U24479 ( .B1(n21540), .B2(n21543), .A(n21539), .ZN(P1_U3211) );
  AOI22_X1 U24480 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21560), .ZN(n21541) );
  OAI21_X1 U24481 ( .B1(n21544), .B2(n21546), .A(n21541), .ZN(P1_U3212) );
  AOI22_X1 U24482 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21559), .ZN(n21542) );
  OAI21_X1 U24483 ( .B1(n21544), .B2(n21543), .A(n21542), .ZN(P1_U3213) );
  AOI22_X1 U24484 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21577), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21560), .ZN(n21545) );
  OAI21_X1 U24485 ( .B1(n21547), .B2(n21546), .A(n21545), .ZN(P1_U3214) );
  AOI222_X1 U24486 ( .A1(n21559), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21560), .ZN(n21548) );
  INV_X1 U24487 ( .A(n21548), .ZN(P1_U3215) );
  AOI222_X1 U24488 ( .A1(n21560), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21559), .ZN(n21549) );
  INV_X1 U24489 ( .A(n21549), .ZN(P1_U3216) );
  AOI222_X1 U24490 ( .A1(n21560), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21559), .ZN(n21550) );
  INV_X1 U24491 ( .A(n21550), .ZN(P1_U3217) );
  AOI222_X1 U24492 ( .A1(n21560), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21559), .ZN(n21551) );
  INV_X1 U24493 ( .A(n21551), .ZN(P1_U3218) );
  AOI222_X1 U24494 ( .A1(n21560), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n21559), .ZN(n21552) );
  INV_X1 U24495 ( .A(n21552), .ZN(P1_U3219) );
  AOI222_X1 U24496 ( .A1(n21560), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21559), .ZN(n21553) );
  INV_X1 U24497 ( .A(n21553), .ZN(P1_U3220) );
  AOI222_X1 U24498 ( .A1(n21560), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21559), .ZN(n21554) );
  INV_X1 U24499 ( .A(n21554), .ZN(P1_U3221) );
  AOI222_X1 U24500 ( .A1(n21560), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21559), .ZN(n21555) );
  INV_X1 U24501 ( .A(n21555), .ZN(P1_U3222) );
  AOI222_X1 U24502 ( .A1(n21560), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21559), .ZN(n21556) );
  INV_X1 U24503 ( .A(n21556), .ZN(P1_U3223) );
  AOI222_X1 U24504 ( .A1(n21560), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21559), .ZN(n21557) );
  INV_X1 U24505 ( .A(n21557), .ZN(P1_U3224) );
  AOI222_X1 U24506 ( .A1(n21559), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21560), .ZN(n21558) );
  INV_X1 U24507 ( .A(n21558), .ZN(P1_U3225) );
  AOI222_X1 U24508 ( .A1(n21560), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21577), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21559), .ZN(n21561) );
  INV_X1 U24509 ( .A(n21561), .ZN(P1_U3226) );
  OAI22_X1 U24510 ( .A1(n21577), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21579), .ZN(n21562) );
  INV_X1 U24511 ( .A(n21562), .ZN(P1_U3458) );
  OAI22_X1 U24512 ( .A1(n21577), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21579), .ZN(n21563) );
  INV_X1 U24513 ( .A(n21563), .ZN(P1_U3459) );
  OAI22_X1 U24514 ( .A1(n21577), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21579), .ZN(n21564) );
  INV_X1 U24515 ( .A(n21564), .ZN(P1_U3460) );
  OAI22_X1 U24516 ( .A1(n21577), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21579), .ZN(n21565) );
  INV_X1 U24517 ( .A(n21565), .ZN(P1_U3461) );
  OAI21_X1 U24518 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21569), .A(n21567), 
        .ZN(n21566) );
  INV_X1 U24519 ( .A(n21566), .ZN(P1_U3464) );
  OAI21_X1 U24520 ( .B1(n21569), .B2(n21568), .A(n21567), .ZN(P1_U3465) );
  AOI21_X1 U24521 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21570) );
  OAI22_X1 U24522 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n21571), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21570), .ZN(n21572) );
  INV_X1 U24523 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21699) );
  AOI22_X1 U24524 ( .A1(n21576), .A2(n21572), .B1(n21699), .B2(n21573), .ZN(
        P1_U3481) );
  NOR2_X1 U24525 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21575) );
  INV_X1 U24526 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21574) );
  AOI22_X1 U24527 ( .A1(n21576), .A2(n21575), .B1(n21574), .B2(n21573), .ZN(
        P1_U3482) );
  AOI22_X1 U24528 ( .A1(n21579), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21578), 
        .B2(n21577), .ZN(P1_U3483) );
  OAI21_X1 U24529 ( .B1(n21581), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21580), 
        .ZN(n21582) );
  OAI21_X1 U24530 ( .B1(n21584), .B2(n21583), .A(n21582), .ZN(n21585) );
  NAND3_X1 U24531 ( .A1(n21585), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21590), 
        .ZN(n21586) );
  OAI21_X1 U24532 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21587), .A(n21586), 
        .ZN(n21593) );
  AOI211_X1 U24533 ( .C1(n20688), .C2(n21590), .A(n21589), .B(n21588), .ZN(
        n21592) );
  NAND2_X1 U24534 ( .A1(n21592), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21591) );
  OAI21_X1 U24535 ( .B1(n21593), .B2(n21592), .A(n21591), .ZN(P1_U3485) );
  MUX2_X1 U24536 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21577), .Z(P1_U3486) );
  NAND4_X1 U24537 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A4(n21594), .ZN(n21598) );
  INV_X1 U24538 ( .A(DATAI_3_), .ZN(n21698) );
  NAND4_X1 U24539 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(n21699), .A4(n21698), .ZN(n21597)
         );
  NAND4_X1 U24540 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_22__SCAN_IN), .A3(P2_DATAO_REG_31__SCAN_IN), .A4(
        n21686), .ZN(n21596) );
  INV_X1 U24541 ( .A(DATAI_27_), .ZN(n21689) );
  NAND4_X1 U24542 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n21689), .A3(n21691), .A4(
        n21692), .ZN(n21595) );
  NOR4_X1 U24543 ( .A1(n21598), .A2(n21597), .A3(n21596), .A4(n21595), .ZN(
        n21748) );
  NOR4_X1 U24544 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__5__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__7__SCAN_IN), 
        .A4(n21626), .ZN(n21604) );
  NOR4_X1 U24545 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P1_DATAO_REG_24__SCAN_IN), .A4(n21618), .ZN(n21603) );
  NOR4_X1 U24546 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_14__5__SCAN_IN), .A4(n21639), .ZN(n21599) );
  NAND2_X1 U24547 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21599), .ZN(
        n21600) );
  NOR4_X1 U24548 ( .A1(n21601), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .A4(n21600), .ZN(n21602) );
  NAND3_X1 U24549 ( .A1(n21604), .A2(n21603), .A3(n21602), .ZN(n21616) );
  NAND4_X1 U24550 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_BYTEENABLE_REG_1__SCAN_IN), .A3(n21648), .A4(n21655), .ZN(n21615)
         );
  NOR3_X1 U24551 ( .A1(DATAI_26_), .A2(P1_DATAO_REG_25__SCAN_IN), .A3(n21605), 
        .ZN(n21608) );
  NOR4_X1 U24552 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        P1_REIP_REG_21__SCAN_IN), .A3(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A4(
        P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21607) );
  NOR4_X1 U24553 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n21667), .A3(n21670), .A4(
        n21668), .ZN(n21606) );
  NAND4_X1 U24554 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n21608), .A3(n21607), 
        .A4(n21606), .ZN(n21614) );
  INV_X1 U24555 ( .A(DATAI_21_), .ZN(n21733) );
  NOR4_X1 U24556 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_1__6__SCAN_IN), .A3(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(n21733), .ZN(n21612) );
  NOR4_X1 U24557 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .A3(P2_DATAO_REG_19__SCAN_IN), .A4(
        n21729), .ZN(n21611) );
  NOR4_X1 U24558 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_EBX_REG_15__SCAN_IN), .A3(P2_LWORD_REG_8__SCAN_IN), .A4(n17916), 
        .ZN(n21610) );
  NOR4_X1 U24559 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n21722), .A4(n21718), .ZN(
        n21609) );
  NAND4_X1 U24560 ( .A1(n21612), .A2(n21611), .A3(n21610), .A4(n21609), .ZN(
        n21613) );
  NOR4_X1 U24561 ( .A1(n21616), .A2(n21615), .A3(n21614), .A4(n21613), .ZN(
        n21747) );
  AOI22_X1 U24562 ( .A1(n21619), .A2(keyinput24), .B1(n21618), .B2(keyinput40), 
        .ZN(n21617) );
  OAI221_X1 U24563 ( .B1(n21619), .B2(keyinput24), .C1(n21618), .C2(keyinput40), .A(n21617), .ZN(n21631) );
  AOI22_X1 U24564 ( .A1(n14083), .A2(keyinput58), .B1(keyinput26), .B2(n21621), 
        .ZN(n21620) );
  OAI221_X1 U24565 ( .B1(n14083), .B2(keyinput58), .C1(n21621), .C2(keyinput26), .A(n21620), .ZN(n21630) );
  AOI22_X1 U24566 ( .A1(n21624), .A2(keyinput52), .B1(n21623), .B2(keyinput34), 
        .ZN(n21622) );
  OAI221_X1 U24567 ( .B1(n21624), .B2(keyinput52), .C1(n21623), .C2(keyinput34), .A(n21622), .ZN(n21629) );
  AOI22_X1 U24568 ( .A1(n21627), .A2(keyinput16), .B1(n21626), .B2(keyinput19), 
        .ZN(n21625) );
  OAI221_X1 U24569 ( .B1(n21627), .B2(keyinput16), .C1(n21626), .C2(keyinput19), .A(n21625), .ZN(n21628) );
  NOR4_X1 U24570 ( .A1(n21631), .A2(n21630), .A3(n21629), .A4(n21628), .ZN(
        n21681) );
  INV_X1 U24571 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21634) );
  AOI22_X1 U24572 ( .A1(n21634), .A2(keyinput55), .B1(keyinput28), .B2(n21633), 
        .ZN(n21632) );
  OAI221_X1 U24573 ( .B1(n21634), .B2(keyinput55), .C1(n21633), .C2(keyinput28), .A(n21632), .ZN(n21646) );
  INV_X1 U24574 ( .A(DATAI_26_), .ZN(n21637) );
  AOI22_X1 U24575 ( .A1(n21637), .A2(keyinput9), .B1(keyinput23), .B2(n21636), 
        .ZN(n21635) );
  OAI221_X1 U24576 ( .B1(n21637), .B2(keyinput9), .C1(n21636), .C2(keyinput23), 
        .A(n21635), .ZN(n21645) );
  INV_X1 U24577 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21640) );
  AOI22_X1 U24578 ( .A1(n21640), .A2(keyinput31), .B1(keyinput61), .B2(n21639), 
        .ZN(n21638) );
  OAI221_X1 U24579 ( .B1(n21640), .B2(keyinput31), .C1(n21639), .C2(keyinput61), .A(n21638), .ZN(n21644) );
  XNOR2_X1 U24580 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput60), .ZN(
        n21642) );
  XNOR2_X1 U24581 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput39), .ZN(n21641)
         );
  NAND2_X1 U24582 ( .A1(n21642), .A2(n21641), .ZN(n21643) );
  NOR4_X1 U24583 ( .A1(n21646), .A2(n21645), .A3(n21644), .A4(n21643), .ZN(
        n21680) );
  AOI22_X1 U24584 ( .A1(n21649), .A2(keyinput3), .B1(n21648), .B2(keyinput4), 
        .ZN(n21647) );
  OAI221_X1 U24585 ( .B1(n21649), .B2(keyinput3), .C1(n21648), .C2(keyinput4), 
        .A(n21647), .ZN(n21662) );
  AOI22_X1 U24586 ( .A1(n21652), .A2(keyinput7), .B1(keyinput32), .B2(n21651), 
        .ZN(n21650) );
  OAI221_X1 U24587 ( .B1(n21652), .B2(keyinput7), .C1(n21651), .C2(keyinput32), 
        .A(n21650), .ZN(n21661) );
  AOI22_X1 U24588 ( .A1(n21655), .A2(keyinput6), .B1(keyinput30), .B2(n21654), 
        .ZN(n21653) );
  OAI221_X1 U24589 ( .B1(n21655), .B2(keyinput6), .C1(n21654), .C2(keyinput30), 
        .A(n21653), .ZN(n21660) );
  AOI22_X1 U24590 ( .A1(n21658), .A2(keyinput59), .B1(keyinput14), .B2(n21657), 
        .ZN(n21656) );
  OAI221_X1 U24591 ( .B1(n21658), .B2(keyinput59), .C1(n21657), .C2(keyinput14), .A(n21656), .ZN(n21659) );
  NOR4_X1 U24592 ( .A1(n21662), .A2(n21661), .A3(n21660), .A4(n21659), .ZN(
        n21679) );
  AOI22_X1 U24593 ( .A1(n21665), .A2(keyinput53), .B1(n21664), .B2(keyinput22), 
        .ZN(n21663) );
  OAI221_X1 U24594 ( .B1(n21665), .B2(keyinput53), .C1(n21664), .C2(keyinput22), .A(n21663), .ZN(n21677) );
  AOI22_X1 U24595 ( .A1(n21668), .A2(keyinput29), .B1(n21667), .B2(keyinput1), 
        .ZN(n21666) );
  OAI221_X1 U24596 ( .B1(n21668), .B2(keyinput29), .C1(n21667), .C2(keyinput1), 
        .A(n21666), .ZN(n21676) );
  INV_X1 U24597 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21671) );
  AOI22_X1 U24598 ( .A1(n21671), .A2(keyinput47), .B1(keyinput5), .B2(n21670), 
        .ZN(n21669) );
  OAI221_X1 U24599 ( .B1(n21671), .B2(keyinput47), .C1(n21670), .C2(keyinput5), 
        .A(n21669), .ZN(n21675) );
  XOR2_X1 U24600 ( .A(n15119), .B(keyinput50), .Z(n21673) );
  XNOR2_X1 U24601 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput49), .ZN(
        n21672) );
  NAND2_X1 U24602 ( .A1(n21673), .A2(n21672), .ZN(n21674) );
  NOR4_X1 U24603 ( .A1(n21677), .A2(n21676), .A3(n21675), .A4(n21674), .ZN(
        n21678) );
  NAND4_X1 U24604 ( .A1(n21681), .A2(n21680), .A3(n21679), .A4(n21678), .ZN(
        n21746) );
  AOI22_X1 U24605 ( .A1(n21684), .A2(keyinput18), .B1(n21683), .B2(keyinput46), 
        .ZN(n21682) );
  OAI221_X1 U24606 ( .B1(n21684), .B2(keyinput18), .C1(n21683), .C2(keyinput46), .A(n21682), .ZN(n21696) );
  AOI22_X1 U24607 ( .A1(n21687), .A2(keyinput2), .B1(n21686), .B2(keyinput0), 
        .ZN(n21685) );
  OAI221_X1 U24608 ( .B1(n21687), .B2(keyinput2), .C1(n21686), .C2(keyinput0), 
        .A(n21685), .ZN(n21695) );
  AOI22_X1 U24609 ( .A1(n11155), .A2(keyinput62), .B1(keyinput57), .B2(n21689), 
        .ZN(n21688) );
  OAI221_X1 U24610 ( .B1(n11155), .B2(keyinput62), .C1(n21689), .C2(keyinput57), .A(n21688), .ZN(n21694) );
  AOI22_X1 U24611 ( .A1(n21692), .A2(keyinput11), .B1(n21691), .B2(keyinput27), 
        .ZN(n21690) );
  OAI221_X1 U24612 ( .B1(n21692), .B2(keyinput11), .C1(n21691), .C2(keyinput27), .A(n21690), .ZN(n21693) );
  NOR4_X1 U24613 ( .A1(n21696), .A2(n21695), .A3(n21694), .A4(n21693), .ZN(
        n21744) );
  AOI22_X1 U24614 ( .A1(n21699), .A2(keyinput43), .B1(n21698), .B2(keyinput35), 
        .ZN(n21697) );
  OAI221_X1 U24615 ( .B1(n21699), .B2(keyinput43), .C1(n21698), .C2(keyinput35), .A(n21697), .ZN(n21711) );
  AOI22_X1 U24616 ( .A1(n21702), .A2(keyinput37), .B1(n21701), .B2(keyinput8), 
        .ZN(n21700) );
  OAI221_X1 U24617 ( .B1(n21702), .B2(keyinput37), .C1(n21701), .C2(keyinput8), 
        .A(n21700), .ZN(n21710) );
  AOI22_X1 U24618 ( .A1(n21705), .A2(keyinput56), .B1(n21704), .B2(keyinput48), 
        .ZN(n21703) );
  OAI221_X1 U24619 ( .B1(n21705), .B2(keyinput56), .C1(n21704), .C2(keyinput48), .A(n21703), .ZN(n21709) );
  XNOR2_X1 U24620 ( .A(P2_REIP_REG_19__SCAN_IN), .B(keyinput63), .ZN(n21707)
         );
  XNOR2_X1 U24621 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B(keyinput21), .ZN(
        n21706) );
  NAND2_X1 U24622 ( .A1(n21707), .A2(n21706), .ZN(n21708) );
  NOR4_X1 U24623 ( .A1(n21711), .A2(n21710), .A3(n21709), .A4(n21708), .ZN(
        n21743) );
  AOI22_X1 U24624 ( .A1(n21713), .A2(keyinput45), .B1(n17916), .B2(keyinput20), 
        .ZN(n21712) );
  OAI221_X1 U24625 ( .B1(n21713), .B2(keyinput45), .C1(n17916), .C2(keyinput20), .A(n21712), .ZN(n21726) );
  AOI22_X1 U24626 ( .A1(n21716), .A2(keyinput36), .B1(keyinput17), .B2(n21715), 
        .ZN(n21714) );
  OAI221_X1 U24627 ( .B1(n21716), .B2(keyinput36), .C1(n21715), .C2(keyinput17), .A(n21714), .ZN(n21725) );
  AOI22_X1 U24628 ( .A1(n21719), .A2(keyinput54), .B1(keyinput44), .B2(n21718), 
        .ZN(n21717) );
  OAI221_X1 U24629 ( .B1(n21719), .B2(keyinput54), .C1(n21718), .C2(keyinput44), .A(n21717), .ZN(n21724) );
  AOI22_X1 U24630 ( .A1(n21722), .A2(keyinput13), .B1(keyinput33), .B2(n21721), 
        .ZN(n21720) );
  OAI221_X1 U24631 ( .B1(n21722), .B2(keyinput13), .C1(n21721), .C2(keyinput33), .A(n21720), .ZN(n21723) );
  NOR4_X1 U24632 ( .A1(n21726), .A2(n21725), .A3(n21724), .A4(n21723), .ZN(
        n21742) );
  AOI22_X1 U24633 ( .A1(n21729), .A2(keyinput38), .B1(keyinput12), .B2(n21728), 
        .ZN(n21727) );
  OAI221_X1 U24634 ( .B1(n21729), .B2(keyinput38), .C1(n21728), .C2(keyinput12), .A(n21727), .ZN(n21740) );
  INV_X1 U24635 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21731) );
  AOI22_X1 U24636 ( .A1(n13532), .A2(keyinput25), .B1(keyinput15), .B2(n21731), 
        .ZN(n21730) );
  OAI221_X1 U24637 ( .B1(n13532), .B2(keyinput25), .C1(n21731), .C2(keyinput15), .A(n21730), .ZN(n21739) );
  AOI22_X1 U24638 ( .A1(n21734), .A2(keyinput51), .B1(n21733), .B2(keyinput10), 
        .ZN(n21732) );
  OAI221_X1 U24639 ( .B1(n21734), .B2(keyinput51), .C1(n21733), .C2(keyinput10), .A(n21732), .ZN(n21738) );
  XNOR2_X1 U24640 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B(keyinput41), .ZN(
        n21736) );
  XNOR2_X1 U24641 ( .A(keyinput42), .B(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n21735) );
  NAND2_X1 U24642 ( .A1(n21736), .A2(n21735), .ZN(n21737) );
  NOR4_X1 U24643 ( .A1(n21740), .A2(n21739), .A3(n21738), .A4(n21737), .ZN(
        n21741) );
  NAND4_X1 U24644 ( .A1(n21744), .A2(n21743), .A3(n21742), .A4(n21741), .ZN(
        n21745) );
  AOI211_X1 U24645 ( .C1(n21748), .C2(n21747), .A(n21746), .B(n21745), .ZN(
        n21761) );
  AOI22_X1 U24646 ( .A1(n21752), .A2(n21751), .B1(n21750), .B2(n21749), .ZN(
        n21757) );
  AOI22_X1 U24647 ( .A1(n21755), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n21754), .B2(n21753), .ZN(n21756) );
  OAI211_X1 U24648 ( .C1(n21759), .C2(n21758), .A(n21757), .B(n21756), .ZN(
        n21760) );
  XOR2_X1 U24649 ( .A(n21761), .B(n21760), .Z(P2_U3146) );
  CLKBUF_X1 U11067 ( .A(n12538), .Z(n12604) );
  CLKBUF_X1 U11068 ( .A(n12015), .Z(n14530) );
  CLKBUF_X1 U11071 ( .A(n11058), .Z(n20204) );
  CLKBUF_X1 U11110 ( .A(n11878), .Z(n13777) );
  CLKBUF_X1 U11503 ( .A(n20894), .Z(n9587) );
  CLKBUF_X1 U11841 ( .A(n11158), .Z(n12932) );
  CLKBUF_X1 U12000 ( .A(n10590), .Z(n17748) );
endmodule

