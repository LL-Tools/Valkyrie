

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6415, n6416, n6417, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888;

  NAND3_X1 U7163 ( .A1(n7365), .A2(n9835), .A3(n13401), .ZN(n13051) );
  NAND2_X1 U7164 ( .A1(n9870), .A2(n9871), .ZN(n9835) );
  CLKBUF_X2 U7165 ( .A(n10416), .Z(n10191) );
  INV_X2 U7166 ( .A(n9708), .ZN(n10423) );
  INV_X1 U7167 ( .A(n8470), .ZN(n10097) );
  NAND2_X2 U7168 ( .A1(n14563), .A2(n12912), .ZN(n12539) );
  INV_X1 U7169 ( .A(n6892), .ZN(n8470) );
  AND4_X1 U7170 ( .A1(n9084), .A2(n8903), .A3(n8836), .A4(n8864), .ZN(n8839)
         );
  NOR2_X1 U7171 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8865) );
  BUF_X1 U7172 ( .A(n12737), .Z(n12803) );
  AOI21_X1 U7173 ( .B1(n7527), .B2(n7529), .A(n7526), .ZN(n7525) );
  INV_X2 U7174 ( .A(n6617), .ZN(n12381) );
  AND2_X1 U7175 ( .A1(n8850), .A2(n8046), .ZN(n9143) );
  INV_X1 U7176 ( .A(n8645), .ZN(n8775) );
  NAND2_X1 U7177 ( .A1(n7128), .A2(n10614), .ZN(n7205) );
  AND2_X1 U7179 ( .A1(n14363), .A2(n7889), .ZN(n14304) );
  CLKBUF_X2 U7180 ( .A(n8239), .Z(n6415) );
  INV_X1 U7181 ( .A(n8239), .ZN(n8644) );
  NAND2_X1 U7182 ( .A1(n11716), .A2(n10312), .ZN(n12162) );
  NAND2_X1 U7183 ( .A1(n9844), .A2(n9874), .ZN(n9867) );
  OAI211_X1 U7184 ( .C1(n9708), .C2(SI_2_), .A(n9486), .B(n9485), .ZN(n15790)
         );
  XNOR2_X1 U7185 ( .A(n14252), .B(n14253), .ZN(n14254) );
  AND2_X1 U7186 ( .A1(n8189), .A2(n12670), .ZN(n10397) );
  AND2_X1 U7187 ( .A1(n8235), .A2(n10769), .ZN(n8355) );
  INV_X2 U7188 ( .A(n8644), .ZN(n8732) );
  CLKBUF_X2 U7189 ( .A(n9533), .Z(n10424) );
  NAND2_X1 U7190 ( .A1(n10482), .A2(n10483), .ZN(n11503) );
  NAND2_X1 U7191 ( .A1(n9068), .A2(n9067), .ZN(n14504) );
  INV_X1 U7192 ( .A(n15064), .ZN(n15200) );
  CLKBUF_X3 U7193 ( .A(n8227), .Z(n8296) );
  INV_X2 U7194 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n11181) );
  XNOR2_X1 U7195 ( .A(n6856), .B(n8424), .ZN(n10833) );
  AND2_X1 U7196 ( .A1(n7765), .A2(n6593), .ZN(n12948) );
  NAND4_X2 U7197 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n15797)
         );
  NAND4_X1 U7198 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n8949), .ZN(n14021)
         );
  INV_X2 U7199 ( .A(n14352), .ZN(n14396) );
  INV_X1 U7200 ( .A(n12534), .ZN(n8895) );
  INV_X1 U7201 ( .A(n8170), .ZN(n12929) );
  XNOR2_X1 U7202 ( .A(n15379), .B(n15380), .ZN(n15878) );
  INV_X1 U7203 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9411) );
  INV_X1 U7204 ( .A(n8301), .ZN(n6420) );
  NOR2_X2 U7205 ( .A1(n9404), .A2(n9475), .ZN(n7586) );
  NAND2_X2 U7206 ( .A1(n15370), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15369) );
  INV_X2 U7207 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n15370) );
  NAND2_X2 U7208 ( .A1(n15008), .A2(n7964), .ZN(n14966) );
  NAND2_X2 U7209 ( .A1(n10330), .A2(n10329), .ZN(n15008) );
  NAND2_X1 U7210 ( .A1(n7254), .A2(n7252), .ZN(n8274) );
  NOR2_X2 U7211 ( .A1(n12890), .A2(n13004), .ZN(n13008) );
  XNOR2_X2 U7212 ( .A(n8694), .B(n8692), .ZN(n12228) );
  INV_X1 U7213 ( .A(n6893), .ZN(n13827) );
  NAND2_X2 U7214 ( .A1(n7859), .A2(n15377), .ZN(n15380) );
  NAND2_X1 U7215 ( .A1(n11216), .A2(n11441), .ZN(n11295) );
  NAND4_X4 U7216 ( .A1(n8272), .A2(n8271), .A3(n8270), .A4(n8269), .ZN(n14745)
         );
  NAND3_X2 U7217 ( .A1(n8886), .A2(n8885), .A3(n6769), .ZN(n10044) );
  OAI21_X2 U7218 ( .B1(n14373), .B2(n6483), .A(n7161), .ZN(n14313) );
  NAND2_X2 U7219 ( .A1(n7841), .A2(n8250), .ZN(n14746) );
  AND2_X1 U7220 ( .A1(n10597), .A2(n12816), .ZN(n8239) );
  XNOR2_X2 U7221 ( .A(n7564), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10676) );
  XNOR2_X2 U7222 ( .A(n8089), .B(SI_9_), .ZN(n8401) );
  OAI21_X2 U7223 ( .B1(n8694), .B2(n7514), .A(n7512), .ZN(n8737) );
  OAI211_X2 U7224 ( .C1(n9218), .C2(n8001), .A(n6621), .B(n7119), .ZN(n8694)
         );
  AOI211_X2 U7225 ( .C1(n13410), .C2(n10160), .A(n13385), .B(n13384), .ZN(
        n13386) );
  OAI21_X2 U7226 ( .B1(n7111), .B2(n8401), .A(n6854), .ZN(n6856) );
  AND2_X2 U7227 ( .A1(n8859), .A2(n8858), .ZN(n14386) );
  NAND2_X4 U7228 ( .A1(n14337), .A2(n8861), .ZN(n8899) );
  BUF_X2 U7229 ( .A(n8115), .Z(n6416) );
  INV_X1 U7230 ( .A(n14023), .ZN(n11578) );
  NAND2_X1 U7231 ( .A1(n7275), .A2(n7274), .ZN(n13974) );
  NAND2_X1 U7232 ( .A1(n14929), .A2(n14928), .ZN(n10337) );
  NAND2_X1 U7233 ( .A1(n8578), .A2(n8577), .ZN(n15188) );
  AND2_X1 U7234 ( .A1(n12735), .A2(n12733), .ZN(n15099) );
  AND2_X1 U7235 ( .A1(n9157), .A2(n9156), .ZN(n14546) );
  AND2_X1 U7236 ( .A1(n12267), .A2(n10315), .ZN(n12181) );
  XNOR2_X1 U7237 ( .A(n6703), .B(n8548), .ZN(n11305) );
  NAND2_X2 U7238 ( .A1(n10494), .A2(n10496), .ZN(n11602) );
  NAND2_X1 U7239 ( .A1(n14743), .A2(n15580), .ZN(n10306) );
  NAND2_X2 U7240 ( .A1(n10472), .A2(n10475), .ZN(n10442) );
  INV_X1 U7241 ( .A(n13122), .ZN(n12042) );
  INV_X1 U7242 ( .A(n13126), .ZN(n15784) );
  INV_X4 U7243 ( .A(n10564), .ZN(n6417) );
  OAI21_X1 U7244 ( .B1(n7993), .B2(n7528), .A(n7525), .ZN(n7264) );
  NAND4_X1 U7245 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(n14743)
         );
  INV_X1 U7246 ( .A(n14022), .ZN(n11330) );
  NAND4_X1 U7247 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n14023)
         );
  NAND4_X1 U7248 ( .A1(n8908), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n14025)
         );
  BUF_X2 U7249 ( .A(n9009), .Z(n9302) );
  CLKBUF_X3 U7250 ( .A(n6420), .Z(n6422) );
  BUF_X2 U7251 ( .A(n8355), .Z(n10091) );
  NAND2_X1 U7252 ( .A1(n12929), .A2(n8171), .ZN(n8227) );
  NAND2_X1 U7253 ( .A1(n8801), .A2(n15526), .ZN(n12670) );
  INV_X1 U7254 ( .A(n8863), .ZN(n8857) );
  NAND2_X1 U7255 ( .A1(n7878), .A2(n7876), .ZN(n15366) );
  AND3_X1 U7256 ( .A1(n8842), .A2(n8841), .A3(n8840), .ZN(n8872) );
  INV_X1 U7257 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9476) );
  NOR2_X1 U7258 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8837) );
  NOR2_X1 U7259 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8838) );
  MUX2_X1 U7260 ( .A(n10398), .B(n10402), .S(n15618), .Z(n10401) );
  AND2_X1 U7261 ( .A1(n6669), .A2(n6668), .ZN(n10402) );
  NOR2_X1 U7262 ( .A1(n6874), .A2(n7881), .ZN(n7880) );
  AND2_X1 U7263 ( .A1(n6932), .A2(n7757), .ZN(n12972) );
  OAI21_X1 U7264 ( .B1(n6558), .B2(n15558), .A(n7171), .ZN(n14856) );
  NAND2_X1 U7265 ( .A1(n13974), .A2(n7750), .ZN(n9366) );
  XNOR2_X1 U7266 ( .A(n14832), .B(n14852), .ZN(n15134) );
  AND2_X1 U7267 ( .A1(n6887), .A2(n6885), .ZN(n15252) );
  OR2_X1 U7268 ( .A1(n15143), .A2(n15558), .ZN(n6887) );
  XNOR2_X1 U7269 ( .A(n15444), .B(n15443), .ZN(n7879) );
  AND2_X1 U7270 ( .A1(n7952), .A2(n6601), .ZN(n14832) );
  AND2_X1 U7271 ( .A1(n7160), .A2(n10281), .ZN(n12935) );
  AOI21_X1 U7272 ( .B1(n6704), .B2(n6452), .A(n6426), .ZN(n6981) );
  NAND2_X1 U7273 ( .A1(n13885), .A2(n9288), .ZN(n13976) );
  AND2_X1 U7274 ( .A1(n8045), .A2(n6683), .ZN(n14417) );
  AOI21_X1 U7275 ( .B1(n10279), .B2(n10270), .A(n14302), .ZN(n7154) );
  NAND2_X1 U7276 ( .A1(n10337), .A2(n6449), .ZN(n7402) );
  OAI21_X1 U7277 ( .B1(n14929), .B2(n6889), .A(n6554), .ZN(n14895) );
  AOI21_X1 U7278 ( .B1(n6685), .B2(n6684), .A(n7362), .ZN(n6683) );
  NAND2_X1 U7279 ( .A1(n6843), .A2(n10151), .ZN(n13388) );
  NAND2_X1 U7280 ( .A1(n13887), .A2(n13886), .ZN(n13885) );
  NAND2_X1 U7281 ( .A1(n7560), .A2(n13298), .ZN(n7559) );
  AND2_X1 U7282 ( .A1(n6848), .A2(n6847), .ZN(n13347) );
  OR2_X1 U7283 ( .A1(n9272), .A2(n9271), .ZN(n13887) );
  NOR2_X1 U7284 ( .A1(n14837), .A2(n14838), .ZN(n15128) );
  OAI21_X1 U7285 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(n12873) );
  AOI211_X1 U7286 ( .C1(n15750), .C2(n14440), .A(n14439), .B(n14438), .ZN(
        n14441) );
  OAI21_X1 U7287 ( .B1(n12507), .B2(n6542), .A(n6758), .ZN(n12509) );
  NAND2_X1 U7288 ( .A1(n6780), .A2(n6778), .ZN(n13920) );
  NAND2_X1 U7289 ( .A1(n13400), .A2(n10563), .ZN(n6843) );
  AOI21_X1 U7290 ( .B1(n7348), .B2(n14379), .A(n7346), .ZN(n14427) );
  NAND2_X1 U7291 ( .A1(n13280), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13279) );
  OAI21_X1 U7292 ( .B1(n14263), .B2(n7808), .A(n7806), .ZN(n14225) );
  NAND2_X1 U7293 ( .A1(n14208), .A2(n9977), .ZN(n14195) );
  OAI21_X1 U7294 ( .B1(n9973), .B2(n7387), .A(n7384), .ZN(n14210) );
  NAND2_X1 U7295 ( .A1(n12973), .A2(n9778), .ZN(n12975) );
  OAI211_X1 U7296 ( .C1(n7383), .C2(n14261), .A(n6682), .B(n14209), .ZN(n14208) );
  NAND2_X1 U7297 ( .A1(n13966), .A2(n9190), .ZN(n13871) );
  NOR2_X1 U7298 ( .A1(n14180), .A2(n10041), .ZN(n8025) );
  INV_X1 U7299 ( .A(n12854), .ZN(n10393) );
  NAND2_X1 U7300 ( .A1(n10344), .A2(n14831), .ZN(n12854) );
  NAND2_X1 U7301 ( .A1(n7062), .A2(n7064), .ZN(n14335) );
  NAND2_X1 U7302 ( .A1(n7458), .A2(n10175), .ZN(n13549) );
  AOI22_X1 U7303 ( .A1(n15404), .A2(n15340), .B1(P3_ADDR_REG_13__SCAN_IN), 
        .B2(n15341), .ZN(n15406) );
  NAND2_X1 U7304 ( .A1(n9322), .A2(n9321), .ZN(n12934) );
  INV_X1 U7305 ( .A(n14880), .ZN(n6419) );
  NAND2_X1 U7306 ( .A1(n8010), .A2(n8008), .ZN(n14476) );
  NOR2_X1 U7307 ( .A1(n13205), .A2(n12214), .ZN(n13222) );
  NAND2_X1 U7308 ( .A1(n15338), .A2(n7373), .ZN(n15404) );
  NAND2_X1 U7309 ( .A1(n12346), .A2(n12345), .ZN(n12344) );
  NAND2_X1 U7310 ( .A1(n6783), .A2(n6779), .ZN(n6778) );
  AOI21_X1 U7311 ( .B1(n7395), .B2(n9966), .A(n7394), .ZN(n7393) );
  NAND2_X1 U7312 ( .A1(n15354), .A2(n15355), .ZN(n15338) );
  NAND2_X1 U7313 ( .A1(n15336), .A2(n6954), .ZN(n15354) );
  OAI21_X1 U7314 ( .B1(n8014), .B2(n7054), .A(n7052), .ZN(n10022) );
  OR2_X1 U7315 ( .A1(n14381), .A2(n14477), .ZN(n14382) );
  AND2_X1 U7316 ( .A1(n6953), .A2(n6952), .ZN(n15399) );
  NAND2_X1 U7317 ( .A1(n7284), .A2(n6850), .ZN(n12210) );
  NAND2_X1 U7318 ( .A1(n6679), .A2(n9247), .ZN(n14440) );
  NAND2_X1 U7319 ( .A1(n12168), .A2(n6444), .ZN(n15091) );
  INV_X1 U7320 ( .A(n7078), .ZN(n10155) );
  AND2_X1 U7321 ( .A1(n10372), .A2(n12747), .ZN(n15070) );
  NAND2_X1 U7322 ( .A1(n9220), .A2(n9219), .ZN(n14277) );
  NAND2_X1 U7323 ( .A1(n10361), .A2(n10360), .ZN(n11719) );
  AOI21_X1 U7324 ( .B1(n11530), .B2(n6499), .A(n8033), .ZN(n12021) );
  OAI21_X1 U7325 ( .B1(n7081), .B2(n7080), .A(n7079), .ZN(n7078) );
  NAND2_X1 U7326 ( .A1(n11384), .A2(n11385), .ZN(n11383) );
  NAND2_X1 U7327 ( .A1(n9147), .A2(n9146), .ZN(n14477) );
  NAND2_X1 U7328 ( .A1(n11531), .A2(n11534), .ZN(n11530) );
  NAND2_X1 U7329 ( .A1(n7263), .A2(n8484), .ZN(n15212) );
  OAI21_X1 U7330 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15332), .A(n15331), .ZN(
        n15396) );
  NOR2_X1 U7331 ( .A1(n15419), .A2(n15386), .ZN(n15388) );
  OR2_X1 U7332 ( .A1(n15234), .A2(n10314), .ZN(n12267) );
  NAND2_X1 U7333 ( .A1(n15329), .A2(n15330), .ZN(n15361) );
  NOR2_X1 U7334 ( .A1(n11738), .A2(n14509), .ZN(n11762) );
  OR2_X1 U7335 ( .A1(n11533), .A2(n12428), .ZN(n11738) );
  AND4_X1 U7336 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n13389)
         );
  NAND2_X1 U7337 ( .A1(n8994), .A2(n8993), .ZN(n12428) );
  NOR2_X1 U7338 ( .A1(n10167), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10177) );
  AND2_X1 U7339 ( .A1(n9935), .A2(n9934), .ZN(n12595) );
  INV_X1 U7340 ( .A(n14688), .ZN(n12700) );
  INV_X1 U7341 ( .A(n11749), .ZN(n13123) );
  NAND2_X1 U7342 ( .A1(n7131), .A2(n6536), .ZN(n13154) );
  NAND2_X1 U7343 ( .A1(n6837), .A2(n10121), .ZN(n10472) );
  AND2_X1 U7344 ( .A1(n11572), .A2(n11039), .ZN(n11643) );
  AND2_X1 U7345 ( .A1(n8357), .A2(n8356), .ZN(n14688) );
  NAND2_X1 U7346 ( .A1(n9605), .A2(n6514), .ZN(n13121) );
  NAND2_X1 U7347 ( .A1(n8982), .A2(n8981), .ZN(n12420) );
  NAND2_X1 U7348 ( .A1(n11340), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U7349 ( .A1(n6488), .A2(n9480), .ZN(n13126) );
  INV_X1 U7350 ( .A(n7264), .ZN(n6799) );
  NAND2_X1 U7351 ( .A1(n6939), .A2(n6532), .ZN(n11365) );
  NAND4_X1 U7352 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n13125)
         );
  NAND2_X1 U7353 ( .A1(n10597), .A2(n12670), .ZN(n8645) );
  INV_X1 U7354 ( .A(n10045), .ZN(n15742) );
  OAI211_X1 U7355 ( .C1(n8301), .C2(n10780), .A(n8310), .B(n8309), .ZN(n15569)
         );
  INV_X1 U7356 ( .A(n11204), .ZN(n10303) );
  INV_X2 U7357 ( .A(n10397), .ZN(n8755) );
  AND2_X1 U7358 ( .A1(n7071), .A2(n6511), .ZN(n10045) );
  AOI21_X1 U7359 ( .B1(n8114), .B2(n8523), .A(n8525), .ZN(n8115) );
  NAND2_X1 U7360 ( .A1(n7245), .A2(n8790), .ZN(n10597) );
  CLKBUF_X2 U7361 ( .A(n9598), .Z(n9744) );
  CLKBUF_X1 U7362 ( .A(n9422), .Z(n10622) );
  NAND4_X1 U7363 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(n14022)
         );
  AND2_X1 U7364 ( .A1(n9413), .A2(n13827), .ZN(n9598) );
  AND2_X2 U7365 ( .A1(n12371), .A2(n13827), .ZN(n10416) );
  NAND2_X1 U7366 ( .A1(n12371), .A2(n6893), .ZN(n9506) );
  INV_X2 U7367 ( .A(n9422), .ZN(n9484) );
  INV_X2 U7368 ( .A(n9561), .ZN(n10180) );
  NAND2_X1 U7369 ( .A1(n9434), .A2(n9436), .ZN(n12237) );
  AND2_X1 U7370 ( .A1(n9439), .A2(n9438), .ZN(n9908) );
  AND2_X1 U7371 ( .A1(n12534), .A2(n12626), .ZN(n12582) );
  INV_X1 U7372 ( .A(n8926), .ZN(n9009) );
  NAND2_X2 U7373 ( .A1(n9413), .A2(n6893), .ZN(n9561) );
  NOR2_X1 U7374 ( .A1(n9590), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U7375 ( .A1(n8849), .A2(n9343), .ZN(n12625) );
  MUX2_X1 U7376 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9437), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9439) );
  INV_X2 U7377 ( .A(n8235), .ZN(n8594) );
  MUX2_X1 U7378 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9431), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9434) );
  AND2_X1 U7379 ( .A1(n8100), .A2(n8099), .ZN(n8191) );
  XNOR2_X1 U7380 ( .A(n6853), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9413) );
  INV_X1 U7381 ( .A(n7999), .ZN(n7998) );
  AND2_X2 U7382 ( .A1(n8894), .A2(n8891), .ZN(n9374) );
  AND2_X2 U7383 ( .A1(n12912), .A2(n8894), .ZN(n6474) );
  INV_X2 U7384 ( .A(n12539), .ZN(n9991) );
  NAND2_X1 U7385 ( .A1(n9447), .A2(n9893), .ZN(n11660) );
  NAND2_X1 U7386 ( .A1(n7317), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7316) );
  NAND3_X1 U7387 ( .A1(n14386), .A2(n10278), .A3(n12626), .ZN(n12373) );
  NAND2_X4 U7388 ( .A1(n11054), .A2(n12942), .ZN(n8940) );
  XNOR2_X1 U7389 ( .A(n8187), .B(P1_IR_REG_19__SCAN_IN), .ZN(n12652) );
  MUX2_X1 U7390 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8843), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7754) );
  NOR2_X1 U7391 ( .A1(n8423), .A2(SI_10_), .ZN(n8000) );
  XNOR2_X1 U7392 ( .A(n8086), .B(SI_8_), .ZN(n8383) );
  AND2_X1 U7393 ( .A1(n9501), .A2(n9520), .ZN(n9553) );
  NAND2_X1 U7394 ( .A1(n8857), .A2(n13610), .ZN(n8844) );
  MUX2_X1 U7395 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8142), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8143) );
  OR2_X1 U7396 ( .A1(n9446), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U7397 ( .A1(n7847), .A2(n7842), .ZN(n8171) );
  NOR2_X1 U7398 ( .A1(n15886), .A2(n15372), .ZN(n15416) );
  INV_X1 U7399 ( .A(n8408), .ZN(n6673) );
  XNOR2_X1 U7400 ( .A(n8162), .B(n8161), .ZN(n15526) );
  AND2_X1 U7401 ( .A1(n7753), .A2(n7752), .ZN(n9417) );
  INV_X1 U7402 ( .A(n9519), .ZN(n9501) );
  CLKBUF_X1 U7403 ( .A(n6664), .Z(n8167) );
  OR2_X1 U7404 ( .A1(n8160), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n8178) );
  OAI21_X1 U7405 ( .B1(n8080), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n8066), .ZN(
        n8251) );
  NAND2_X2 U7406 ( .A1(n10769), .A2(P1_U3086), .ZN(n15305) );
  NAND2_X1 U7407 ( .A1(n7151), .A2(n9519), .ZN(n10788) );
  XNOR2_X1 U7408 ( .A(n7132), .B(n9476), .ZN(n11033) );
  NAND3_X1 U7409 ( .A1(n7239), .A2(n7238), .A3(n7237), .ZN(n10999) );
  AND2_X2 U7410 ( .A1(n7002), .A2(n7001), .ZN(n8080) );
  AND3_X1 U7411 ( .A1(n8869), .A2(n8868), .A3(n8867), .ZN(n8873) );
  AND2_X1 U7412 ( .A1(n8140), .A2(n8139), .ZN(n8146) );
  NOR2_X1 U7413 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8840) );
  INV_X1 U7414 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9593) );
  INV_X1 U7415 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9609) );
  NOR2_X1 U7416 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n8140) );
  NOR2_X1 U7417 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n8139) );
  NOR2_X1 U7418 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8842) );
  INV_X1 U7419 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8148) );
  INV_X4 U7420 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7421 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8841) );
  NOR2_X1 U7422 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9396) );
  INV_X4 U7423 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7424 ( .A(P2_RD_REG_SCAN_IN), .ZN(n13609) );
  NOR2_X1 U7425 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9401) );
  NOR2_X1 U7426 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8868) );
  NOR2_X1 U7427 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n8869) );
  NOR2_X1 U7428 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8130) );
  INV_X1 U7429 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8331) );
  INV_X1 U7430 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8133) );
  INV_X4 U7431 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7432 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9554) );
  INV_X1 U7433 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9552) );
  INV_X1 U7435 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8929) );
  INV_X1 U7436 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9084) );
  INV_X1 U7437 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8864) );
  NOR2_X2 U7438 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7778) );
  NAND2_X1 U7439 ( .A1(n8138), .A2(n8183), .ZN(n8160) );
  NAND2_X2 U7440 ( .A1(n8470), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8228) );
  NAND2_X2 U7441 ( .A1(n8879), .A2(n8878), .ZN(n12942) );
  OAI21_X2 U7442 ( .B1(n8863), .B2(n8862), .A(n8875), .ZN(n8879) );
  NAND2_X2 U7443 ( .A1(n7967), .A2(n7966), .ZN(n11716) );
  INV_X2 U7444 ( .A(n7244), .ZN(n15549) );
  OAI21_X2 U7445 ( .B1(n14871), .B2(n14870), .A(n15604), .ZN(n14873) );
  CLKBUF_X2 U7446 ( .A(n14400), .Z(n6421) );
  OAI211_X1 U7447 ( .C1(n10778), .C2(n8926), .A(n8915), .B(n8914), .ZN(n14400)
         );
  AND2_X4 U7448 ( .A1(n6951), .A2(n12534), .ZN(n6617) );
  INV_X1 U7449 ( .A(n12373), .ZN(n6951) );
  NAND2_X1 U7450 ( .A1(n7070), .A2(n7068), .ZN(n7193) );
  AND2_X1 U7451 ( .A1(n7069), .A2(n10038), .ZN(n7068) );
  NAND2_X1 U7452 ( .A1(n6423), .A2(n6456), .ZN(n7675) );
  AOI21_X1 U7453 ( .B1(n7998), .B2(n7995), .A(n7994), .ZN(n7993) );
  INV_X1 U7454 ( .A(n8096), .ZN(n7994) );
  AND2_X1 U7455 ( .A1(n8000), .A2(n7997), .ZN(n7995) );
  NAND2_X1 U7456 ( .A1(n6870), .A2(n15319), .ZN(n15320) );
  NAND2_X1 U7457 ( .A1(n15375), .A2(n15374), .ZN(n6870) );
  INV_X1 U7458 ( .A(n7288), .ZN(n6847) );
  OAI21_X1 U7459 ( .B1(n13400), .B2(n6846), .A(n6844), .ZN(n6848) );
  OAI21_X1 U7460 ( .B1(n7290), .B2(n7289), .A(n6570), .ZN(n7288) );
  OR2_X1 U7461 ( .A1(n12988), .A2(n13418), .ZN(n10558) );
  NOR2_X1 U7462 ( .A1(n9410), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7752) );
  AND2_X1 U7463 ( .A1(n7462), .A2(n7102), .ZN(n6819) );
  NAND2_X1 U7464 ( .A1(n9534), .A2(n9537), .ZN(n7102) );
  NOR2_X1 U7465 ( .A1(n12934), .A2(n14420), .ZN(n7895) );
  AOI21_X1 U7466 ( .B1(n6436), .B2(n7792), .A(n6548), .ZN(n7788) );
  NAND2_X1 U7467 ( .A1(n6436), .A2(n14195), .ZN(n6690) );
  INV_X1 U7468 ( .A(n9979), .ZN(n7792) );
  NOR2_X1 U7469 ( .A1(n10030), .A2(n8049), .ZN(n10036) );
  NOR2_X1 U7470 ( .A1(n14902), .A2(n7850), .ZN(n7849) );
  NOR2_X1 U7471 ( .A1(n12851), .A2(n14910), .ZN(n8062) );
  INV_X1 U7472 ( .A(n7962), .ZN(n7961) );
  NAND2_X1 U7473 ( .A1(n14746), .A2(n11204), .ZN(n12668) );
  NAND2_X1 U7474 ( .A1(n8355), .A2(n8219), .ZN(n7242) );
  OAI21_X1 U7475 ( .B1(n8759), .B2(n7533), .A(n7531), .ZN(n10088) );
  INV_X1 U7476 ( .A(n7534), .ZN(n7533) );
  AOI21_X1 U7477 ( .B1(n7534), .B2(n7536), .A(n7532), .ZN(n7531) );
  INV_X1 U7478 ( .A(n10068), .ZN(n7532) );
  INV_X1 U7479 ( .A(n7123), .ZN(n7122) );
  AOI21_X1 U7480 ( .B1(n7123), .B2(n7121), .A(n6563), .ZN(n7120) );
  AOI21_X1 U7481 ( .B1(n6416), .B2(n8003), .A(n6573), .ZN(n7123) );
  INV_X1 U7482 ( .A(n9561), .ZN(n7746) );
  OR2_X1 U7483 ( .A1(n10160), .A2(n13389), .ZN(n10573) );
  NAND2_X1 U7484 ( .A1(n10022), .A2(n8011), .ZN(n8010) );
  NOR2_X1 U7485 ( .A1(n12333), .A2(n8012), .ZN(n8011) );
  INV_X1 U7486 ( .A(n12239), .ZN(n8012) );
  CLKBUF_X3 U7487 ( .A(n8470), .Z(n12657) );
  NAND2_X1 U7488 ( .A1(n6665), .A2(n10392), .ZN(n10394) );
  AND2_X1 U7489 ( .A1(n14868), .A2(n10391), .ZN(n7126) );
  XNOR2_X1 U7490 ( .A(n14721), .B(n6419), .ZN(n14868) );
  NOR2_X1 U7491 ( .A1(n14987), .A2(n7965), .ZN(n7964) );
  INV_X1 U7492 ( .A(n10331), .ZN(n7965) );
  AOI21_X1 U7493 ( .B1(n8168), .B2(n6513), .A(n7843), .ZN(n7842) );
  OR2_X1 U7494 ( .A1(n8168), .A2(n7848), .ZN(n7847) );
  NAND2_X1 U7495 ( .A1(n12417), .A2(n12416), .ZN(n12415) );
  NAND2_X1 U7496 ( .A1(n12409), .A2(n12408), .ZN(n12414) );
  OAI21_X1 U7497 ( .B1(n6960), .B2(n12702), .A(n12701), .ZN(n6959) );
  NAND2_X1 U7498 ( .A1(n12492), .A2(n12493), .ZN(n6744) );
  NAND2_X1 U7499 ( .A1(n12494), .A2(n6746), .ZN(n6745) );
  NAND2_X1 U7500 ( .A1(n6747), .A2(n6749), .ZN(n6746) );
  AND2_X1 U7501 ( .A1(n7819), .A2(n12505), .ZN(n7817) );
  NAND2_X1 U7502 ( .A1(n7664), .A2(n6490), .ZN(n7663) );
  NAND2_X1 U7503 ( .A1(n7665), .A2(n7667), .ZN(n7664) );
  XNOR2_X1 U7504 ( .A(n12652), .B(n12651), .ZN(n12655) );
  OR2_X1 U7505 ( .A1(n6982), .A2(n12801), .ZN(n6979) );
  INV_X1 U7506 ( .A(n12800), .ZN(n6982) );
  NAND2_X1 U7507 ( .A1(n13051), .A2(n9835), .ZN(n9844) );
  XNOR2_X1 U7508 ( .A(n13411), .B(n12895), .ZN(n9874) );
  INV_X1 U7509 ( .A(n7314), .ZN(n7676) );
  INV_X1 U7510 ( .A(n11155), .ZN(n7688) );
  INV_X1 U7511 ( .A(n11154), .ZN(n7685) );
  NAND2_X1 U7512 ( .A1(n13191), .A2(n10609), .ZN(n10610) );
  INV_X1 U7513 ( .A(n10619), .ZN(n7552) );
  OAI21_X1 U7514 ( .B1(n13259), .B2(n10700), .A(n7137), .ZN(n10707) );
  AND2_X1 U7515 ( .A1(n7138), .A2(n13287), .ZN(n7137) );
  OR2_X1 U7516 ( .A1(n13260), .A2(n10700), .ZN(n7138) );
  OR2_X1 U7517 ( .A1(n13340), .A2(n10200), .ZN(n10577) );
  NAND2_X1 U7518 ( .A1(n7369), .A2(n13350), .ZN(n10572) );
  OR2_X1 U7519 ( .A1(n13814), .A2(n13117), .ZN(n10516) );
  NOR2_X1 U7520 ( .A1(n6443), .A2(n7345), .ZN(n7344) );
  INV_X1 U7521 ( .A(n10137), .ZN(n7345) );
  AND2_X1 U7522 ( .A1(n10232), .A2(n7503), .ZN(n7502) );
  NAND2_X1 U7523 ( .A1(n11440), .A2(n11509), .ZN(n10482) );
  AOI21_X1 U7524 ( .B1(n7090), .B2(n7933), .A(n9766), .ZN(n7088) );
  AND2_X1 U7525 ( .A1(n7461), .A2(n7930), .ZN(n7460) );
  NAND2_X1 U7526 ( .A1(n7462), .A2(n7464), .ZN(n7461) );
  NAND2_X1 U7527 ( .A1(n9517), .A2(n9516), .ZN(n6817) );
  NAND2_X1 U7528 ( .A1(n6428), .A2(n6507), .ZN(n6743) );
  INV_X1 U7529 ( .A(n6739), .ZN(n6738) );
  OAI21_X1 U7530 ( .B1(n7838), .B2(n6742), .A(n12529), .ZN(n6739) );
  INV_X1 U7531 ( .A(n14563), .ZN(n8894) );
  NAND2_X1 U7532 ( .A1(n7197), .A2(n10038), .ZN(n7196) );
  INV_X1 U7533 ( .A(n10037), .ZN(n7197) );
  AND2_X1 U7534 ( .A1(n6689), .A2(n7806), .ZN(n7805) );
  INV_X1 U7535 ( .A(n14298), .ZN(n10029) );
  NAND2_X1 U7536 ( .A1(n7067), .A2(n10024), .ZN(n7066) );
  INV_X1 U7537 ( .A(n10023), .ZN(n7067) );
  NOR2_X1 U7538 ( .A1(n14504), .A2(n12460), .ZN(n7886) );
  INV_X1 U7539 ( .A(n11588), .ZN(n7802) );
  INV_X1 U7540 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8867) );
  NOR2_X1 U7541 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n8871) );
  OAI21_X1 U7542 ( .B1(n7263), .B2(n8645), .A(n6556), .ZN(n6805) );
  NAND2_X1 U7543 ( .A1(n7262), .A2(n8775), .ZN(n6804) );
  NAND2_X1 U7544 ( .A1(n11371), .A2(n7236), .ZN(n7979) );
  AND2_X1 U7545 ( .A1(n7984), .A2(n11373), .ZN(n7236) );
  AND2_X1 U7546 ( .A1(n7988), .A2(n7229), .ZN(n6793) );
  INV_X1 U7547 ( .A(n7989), .ZN(n7988) );
  INV_X1 U7548 ( .A(n8403), .ZN(n8465) );
  AND2_X1 U7549 ( .A1(n10324), .A2(n15033), .ZN(n10325) );
  NAND2_X1 U7550 ( .A1(n7263), .A2(n7261), .ZN(n12733) );
  NOR2_X1 U7551 ( .A1(n10323), .A2(n7262), .ZN(n7261) );
  NOR2_X1 U7552 ( .A1(n14887), .A2(n14880), .ZN(n10065) );
  NAND2_X1 U7553 ( .A1(n8188), .A2(n15526), .ZN(n12814) );
  NAND2_X1 U7554 ( .A1(n8739), .A2(n8738), .ZN(n8759) );
  OAI21_X1 U7555 ( .B1(n8737), .B2(n13837), .A(n8736), .ZN(n8739) );
  NAND2_X1 U7556 ( .A1(n8122), .A2(n11193), .ZN(n8125) );
  NAND2_X1 U7557 ( .A1(n6799), .A2(n6797), .ZN(n6691) );
  AND2_X1 U7558 ( .A1(n6796), .A2(n6795), .ZN(n8500) );
  NAND2_X1 U7559 ( .A1(n7264), .A2(n10972), .ZN(n6796) );
  OR2_X1 U7560 ( .A1(n8466), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U7561 ( .A1(n8191), .A2(n8192), .ZN(n8194) );
  NAND2_X1 U7562 ( .A1(n8384), .A2(n6786), .ZN(n7111) );
  INV_X1 U7563 ( .A(n8383), .ZN(n6786) );
  INV_X1 U7564 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7865) );
  INV_X1 U7565 ( .A(n13127), .ZN(n6837) );
  XNOR2_X1 U7566 ( .A(n9531), .B(n13125), .ZN(n11363) );
  NAND2_X1 U7567 ( .A1(n13016), .A2(n13017), .ZN(n9731) );
  NAND2_X1 U7568 ( .A1(n9513), .A2(n9514), .ZN(n7321) );
  NAND2_X1 U7569 ( .A1(n9731), .A2(n7761), .ZN(n7760) );
  NOR2_X1 U7570 ( .A1(n13025), .A2(n7762), .ZN(n7761) );
  INV_X1 U7571 ( .A(n13018), .ZN(n7762) );
  NOR2_X1 U7572 ( .A1(n10405), .A2(n10404), .ZN(n10435) );
  NAND2_X1 U7573 ( .A1(n10416), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9462) );
  AND2_X1 U7574 ( .A1(n10681), .A2(n11154), .ZN(n11018) );
  NAND2_X1 U7575 ( .A1(n7685), .A2(n7688), .ZN(n7684) );
  NAND2_X1 U7576 ( .A1(n11018), .A2(n6481), .ZN(n7686) );
  OR2_X1 U7577 ( .A1(n13190), .A2(n10660), .ZN(n7588) );
  OAI21_X1 U7578 ( .B1(n13222), .B2(n13220), .A(n13221), .ZN(n13219) );
  NAND2_X1 U7579 ( .A1(n7691), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U7580 ( .A1(n7552), .A2(n7562), .ZN(n7560) );
  INV_X1 U7581 ( .A(n10153), .ZN(n7292) );
  AND2_X1 U7582 ( .A1(n10573), .A2(n10571), .ZN(n13379) );
  BUF_X1 U7583 ( .A(n10423), .Z(n6931) );
  AOI21_X1 U7584 ( .B1(n7920), .B2(n7922), .A(n10560), .ZN(n7918) );
  NAND2_X1 U7585 ( .A1(n13451), .A2(n7920), .ZN(n7919) );
  OR2_X1 U7586 ( .A1(n13587), .A2(n13480), .ZN(n13452) );
  NOR2_X1 U7587 ( .A1(n7710), .A2(n6530), .ZN(n7379) );
  AND2_X1 U7588 ( .A1(n13477), .A2(n7711), .ZN(n7710) );
  INV_X1 U7589 ( .A(n10145), .ZN(n7711) );
  NAND2_X1 U7590 ( .A1(n9922), .A2(n6417), .ZN(n15783) );
  INV_X1 U7591 ( .A(n15799), .ZN(n15785) );
  AND2_X2 U7592 ( .A1(n9422), .A2(n10769), .ZN(n9533) );
  NAND2_X2 U7593 ( .A1(n9422), .A2(n10071), .ZN(n9708) );
  NAND2_X1 U7594 ( .A1(n10410), .A2(n10409), .ZN(n10422) );
  NAND2_X1 U7595 ( .A1(n9417), .A2(n9418), .ZN(n7317) );
  NAND2_X1 U7596 ( .A1(n10173), .A2(n10172), .ZN(n10186) );
  NOR2_X1 U7597 ( .A1(n10171), .A2(n7470), .ZN(n7469) );
  NAND2_X1 U7598 ( .A1(n9818), .A2(n6620), .ZN(n9837) );
  OR2_X1 U7599 ( .A1(n9736), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n9755) );
  OAI21_X1 U7600 ( .B1(n9705), .B2(n9717), .A(n7455), .ZN(n9734) );
  NAND2_X1 U7601 ( .A1(n7459), .A2(n7462), .ZN(n9588) );
  OR2_X1 U7602 ( .A1(n9557), .A2(n7464), .ZN(n7459) );
  INV_X1 U7603 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7152) );
  AND2_X1 U7604 ( .A1(n7150), .A2(n7778), .ZN(n7153) );
  NAND2_X1 U7605 ( .A1(n7736), .A2(n9131), .ZN(n7735) );
  INV_X1 U7606 ( .A(n9170), .ZN(n7736) );
  INV_X1 U7607 ( .A(n6474), .ZN(n9379) );
  INV_X1 U7608 ( .A(n9374), .ZN(n9326) );
  AND2_X1 U7609 ( .A1(n14563), .A2(n8891), .ZN(n9001) );
  OAI21_X1 U7610 ( .B1(n8023), .B2(n8022), .A(n8024), .ZN(n10269) );
  AOI21_X1 U7611 ( .B1(n8025), .B2(n6442), .A(n6550), .ZN(n8024) );
  INV_X1 U7612 ( .A(n8025), .ZN(n8022) );
  NAND2_X1 U7613 ( .A1(n9275), .A2(n6471), .ZN(n9323) );
  AOI21_X1 U7614 ( .B1(n14187), .B2(n12934), .A(n14380), .ZN(n10282) );
  NAND2_X1 U7615 ( .A1(n14195), .A2(n9978), .ZN(n7789) );
  AND2_X1 U7616 ( .A1(n7883), .A2(n6860), .ZN(n6859) );
  INV_X1 U7617 ( .A(n14425), .ZN(n6860) );
  INV_X1 U7618 ( .A(n7162), .ZN(n7161) );
  OAI21_X1 U7619 ( .B1(n6483), .B2(n14389), .A(n9964), .ZN(n7162) );
  NAND2_X1 U7620 ( .A1(n10027), .A2(n10026), .ZN(n14333) );
  INV_X1 U7621 ( .A(n14335), .ZN(n10027) );
  INV_X1 U7622 ( .A(n7053), .ZN(n7052) );
  INV_X1 U7623 ( .A(n10021), .ZN(n7054) );
  INV_X1 U7624 ( .A(n8020), .ZN(n8019) );
  AOI21_X1 U7625 ( .B1(n8020), .B2(n8018), .A(n6519), .ZN(n8017) );
  INV_X1 U7626 ( .A(n10019), .ZN(n8018) );
  NAND2_X1 U7627 ( .A1(n7181), .A2(n8027), .ZN(n11531) );
  AOI21_X1 U7628 ( .B1(n8030), .B2(n8028), .A(n8029), .ZN(n8027) );
  NAND2_X1 U7629 ( .A1(n11626), .A2(n8031), .ZN(n7181) );
  NOR2_X1 U7630 ( .A1(n14019), .A2(n12420), .ZN(n8029) );
  NOR2_X1 U7631 ( .A1(n11663), .A2(n10044), .ZN(n11572) );
  XNOR2_X1 U7632 ( .A(n12625), .B(n12582), .ZN(n8860) );
  INV_X1 U7633 ( .A(n15721), .ZN(n10289) );
  NAND2_X1 U7634 ( .A1(n7542), .A2(n12551), .ZN(n12552) );
  NAND2_X1 U7635 ( .A1(n14557), .A2(n9302), .ZN(n7542) );
  INV_X1 U7636 ( .A(n8940), .ZN(n11049) );
  AND3_X1 U7637 ( .A1(n12640), .A2(n12625), .A3(n8895), .ZN(n15750) );
  AND2_X1 U7638 ( .A1(n9358), .A2(n9357), .ZN(n15716) );
  XNOR2_X1 U7639 ( .A(n8890), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U7640 ( .A1(n8889), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8890) );
  INV_X1 U7641 ( .A(n8889), .ZN(n7168) );
  NOR2_X1 U7642 ( .A1(n14603), .A2(n7233), .ZN(n7232) );
  INV_X1 U7643 ( .A(n8591), .ZN(n7233) );
  NAND2_X1 U7644 ( .A1(n6670), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8600) );
  INV_X1 U7645 ( .A(n8598), .ZN(n6670) );
  NAND2_X1 U7646 ( .A1(n14696), .A2(n7973), .ZN(n7972) );
  AND2_X1 U7647 ( .A1(n8222), .A2(n8221), .ZN(n8225) );
  XNOR2_X1 U7648 ( .A(n7350), .B(n10397), .ZN(n7219) );
  NAND2_X1 U7649 ( .A1(n7244), .A2(n7243), .ZN(n8223) );
  NAND2_X1 U7650 ( .A1(n11371), .A2(n11373), .ZN(n8322) );
  INV_X1 U7651 ( .A(n14725), .ZN(n14666) );
  INV_X1 U7652 ( .A(n8296), .ZN(n12656) );
  AND2_X1 U7653 ( .A1(n10964), .A2(n6508), .ZN(n7417) );
  NAND2_X1 U7654 ( .A1(n12075), .A2(n7410), .ZN(n7409) );
  OR2_X1 U7655 ( .A1(n12076), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7410) );
  XNOR2_X1 U7656 ( .A(n14834), .B(n14720), .ZN(n14852) );
  INV_X1 U7657 ( .A(n15131), .ZN(n14834) );
  NOR2_X2 U7658 ( .A1(n12804), .A2(n14876), .ZN(n14833) );
  OR2_X1 U7659 ( .A1(n10394), .A2(n10393), .ZN(n14850) );
  OR2_X1 U7660 ( .A1(n8722), .A2(n8721), .ZN(n8746) );
  NAND2_X1 U7661 ( .A1(n7402), .A2(n7403), .ZN(n14869) );
  OR2_X1 U7662 ( .A1(n6591), .A2(n8062), .ZN(n7850) );
  NAND2_X1 U7663 ( .A1(n14953), .A2(n10388), .ZN(n14935) );
  OR2_X1 U7664 ( .A1(n14994), .A2(n14611), .ZN(n14968) );
  NAND2_X1 U7665 ( .A1(n15000), .A2(n15006), .ZN(n10385) );
  NAND2_X1 U7666 ( .A1(n12306), .A2(n7008), .ZN(n12350) );
  AOI21_X1 U7667 ( .B1(n10317), .B2(n7010), .A(n7008), .ZN(n7007) );
  OR2_X1 U7668 ( .A1(n12651), .A2(n8801), .ZN(n15524) );
  NOR2_X1 U7669 ( .A1(n15128), .A2(n15132), .ZN(n7495) );
  NAND2_X1 U7670 ( .A1(n8621), .A2(n8620), .ZN(n14974) );
  INV_X1 U7671 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8166) );
  XNOR2_X1 U7672 ( .A(n7381), .B(n8442), .ZN(n10865) );
  OAI21_X1 U7673 ( .B1(n8091), .B2(n8000), .A(n7998), .ZN(n7381) );
  NAND2_X1 U7674 ( .A1(n7877), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7876) );
  INV_X1 U7675 ( .A(n13105), .ZN(n13402) );
  AOI21_X1 U7676 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n10167), .A(n10177), .ZN(
        n13370) );
  NOR2_X1 U7677 ( .A1(n7388), .A2(n10270), .ZN(n6684) );
  XNOR2_X1 U7678 ( .A(n7057), .B(n9989), .ZN(n14418) );
  NAND2_X1 U7679 ( .A1(n10273), .A2(n10042), .ZN(n7057) );
  NOR2_X1 U7680 ( .A1(n12284), .A2(n12229), .ZN(n7245) );
  AND2_X1 U7681 ( .A1(n14880), .A2(n15598), .ZN(n15135) );
  NAND2_X1 U7682 ( .A1(n8596), .A2(n8595), .ZN(n15012) );
  NAND2_X1 U7683 ( .A1(n7198), .A2(n8691), .ZN(n14618) );
  NAND2_X1 U7684 ( .A1(n7124), .A2(n8699), .ZN(n14903) );
  NAND2_X1 U7685 ( .A1(n12282), .A2(n10091), .ZN(n7124) );
  MUX2_X1 U7686 ( .A(n11181), .B(n15310), .S(n8235), .Z(n15525) );
  OR2_X1 U7687 ( .A1(n8235), .A2(n8254), .ZN(n8255) );
  NAND2_X1 U7688 ( .A1(n8752), .A2(n8751), .ZN(n14721) );
  NOR2_X1 U7689 ( .A1(n10843), .A2(n10844), .ZN(n10894) );
  NOR2_X1 U7690 ( .A1(n14816), .A2(n14805), .ZN(n6710) );
  NAND2_X1 U7691 ( .A1(n7862), .A2(n7864), .ZN(n7861) );
  INV_X1 U7692 ( .A(n15451), .ZN(n7863) );
  INV_X1 U7693 ( .A(n12679), .ZN(n12683) );
  AND2_X1 U7694 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  AND2_X1 U7695 ( .A1(n12694), .A2(n15488), .ZN(n12695) );
  OR2_X1 U7696 ( .A1(n12693), .A2(n12692), .ZN(n12694) );
  NAND2_X1 U7697 ( .A1(n12394), .A2(n12393), .ZN(n6752) );
  OR2_X1 U7698 ( .A1(n12703), .A2(n12705), .ZN(n6957) );
  NAND2_X1 U7699 ( .A1(n12707), .A2(n6986), .ZN(n6985) );
  OR2_X1 U7700 ( .A1(n6732), .A2(n6731), .ZN(n6950) );
  AOI21_X1 U7701 ( .B1(n6733), .B2(n12457), .A(n12456), .ZN(n6731) );
  AND2_X1 U7702 ( .A1(n12475), .A2(n12476), .ZN(n7830) );
  OAI21_X1 U7703 ( .B1(n12477), .B2(n7830), .A(n6935), .ZN(n12484) );
  AND2_X1 U7704 ( .A1(n7827), .A2(n6936), .ZN(n6935) );
  INV_X1 U7705 ( .A(n12483), .ZN(n6936) );
  NAND2_X1 U7706 ( .A1(n12489), .A2(n12488), .ZN(n7834) );
  INV_X1 U7707 ( .A(n12489), .ZN(n7836) );
  AOI21_X1 U7708 ( .B1(n7644), .B2(n7643), .A(n6447), .ZN(n10485) );
  INV_X1 U7709 ( .A(n10500), .ZN(n10501) );
  AND2_X1 U7710 ( .A1(n12774), .A2(n12773), .ZN(n7442) );
  NAND2_X1 U7711 ( .A1(n6462), .A2(n7905), .ZN(n7439) );
  AOI21_X1 U7712 ( .B1(n6701), .B2(n15001), .A(n12771), .ZN(n12772) );
  INV_X1 U7713 ( .A(n7666), .ZN(n7665) );
  OAI21_X1 U7714 ( .B1(n7667), .B2(n7669), .A(n10539), .ZN(n7666) );
  NOR2_X1 U7715 ( .A1(n10534), .A2(n7670), .ZN(n7669) );
  NAND2_X1 U7716 ( .A1(n7812), .A2(n7811), .ZN(n7810) );
  NAND2_X1 U7717 ( .A1(n12504), .A2(n7819), .ZN(n7811) );
  INV_X1 U7718 ( .A(n7814), .ZN(n7813) );
  OAI21_X1 U7719 ( .B1(n7818), .B2(n7816), .A(n7815), .ZN(n7814) );
  AOI21_X1 U7720 ( .B1(n6480), .B2(n7819), .A(n12505), .ZN(n7818) );
  NAND2_X1 U7721 ( .A1(n6697), .A2(n6696), .ZN(n12783) );
  INV_X1 U7722 ( .A(n12779), .ZN(n6696) );
  NAND2_X1 U7723 ( .A1(n6698), .A2(n12778), .ZN(n12782) );
  NAND2_X1 U7724 ( .A1(n12782), .A2(n12783), .ZN(n6974) );
  OR2_X1 U7725 ( .A1(n6974), .A2(n12785), .ZN(n12791) );
  OAI21_X1 U7726 ( .B1(n10553), .B2(n7655), .A(n7654), .ZN(n7653) );
  NAND2_X1 U7727 ( .A1(n7657), .A2(n7656), .ZN(n7655) );
  NOR2_X1 U7728 ( .A1(n13430), .A2(n10556), .ZN(n7654) );
  NOR2_X1 U7729 ( .A1(n13421), .A2(n10561), .ZN(n7652) );
  NAND2_X1 U7730 ( .A1(n10572), .A2(n10564), .ZN(n7314) );
  NAND2_X1 U7731 ( .A1(n13158), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7576) );
  NOR2_X1 U7732 ( .A1(n6430), .A2(n13175), .ZN(n7141) );
  INV_X1 U7733 ( .A(n10138), .ZN(n7748) );
  INV_X1 U7734 ( .A(n11400), .ZN(n10126) );
  AND3_X1 U7735 ( .A1(n9409), .A2(n13720), .A3(n9432), .ZN(n8038) );
  INV_X1 U7736 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U7737 ( .A1(n12526), .A2(n7839), .ZN(n7838) );
  OAI21_X1 U7738 ( .B1(n12518), .B2(n6756), .A(n6754), .ZN(n12525) );
  NAND2_X1 U7739 ( .A1(n6484), .A2(n6757), .ZN(n6756) );
  AOI21_X1 U7740 ( .B1(n6484), .B2(n6755), .A(n6448), .ZN(n6754) );
  INV_X1 U7741 ( .A(n8715), .ZN(n7513) );
  OR2_X1 U7742 ( .A1(n8002), .A2(n8652), .ZN(n8001) );
  NAND2_X1 U7743 ( .A1(n8105), .A2(n8523), .ZN(n8003) );
  INV_X1 U7744 ( .A(n8104), .ZN(n7526) );
  AND2_X1 U7745 ( .A1(n7998), .A2(n7997), .ZN(n7996) );
  INV_X1 U7746 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8063) );
  NAND2_X1 U7747 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n15367), .ZN(n7328) );
  NAND2_X1 U7748 ( .A1(n9870), .A2(n9869), .ZN(n12883) );
  NOR2_X1 U7749 ( .A1(n11216), .A2(n11441), .ZN(n9493) );
  INV_X1 U7750 ( .A(n9621), .ZN(n6921) );
  AND2_X1 U7751 ( .A1(n9695), .A2(n9656), .ZN(n6918) );
  OR2_X1 U7752 ( .A1(n9561), .A2(n13341), .ZN(n10195) );
  NAND2_X1 U7753 ( .A1(n7608), .A2(n7601), .ZN(n10627) );
  AND2_X1 U7754 ( .A1(n7603), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U7755 ( .A1(n10989), .A2(n10604), .ZN(n7549) );
  NAND2_X1 U7756 ( .A1(n7595), .A2(n6479), .ZN(n7597) );
  INV_X1 U7757 ( .A(n11026), .ZN(n7596) );
  NAND2_X1 U7758 ( .A1(n7681), .A2(n7679), .ZN(n7682) );
  INV_X1 U7759 ( .A(n7680), .ZN(n7679) );
  OR2_X1 U7760 ( .A1(n7685), .A2(n7687), .ZN(n7681) );
  OAI21_X1 U7761 ( .B1(n7688), .B2(n7687), .A(n10791), .ZN(n7680) );
  INV_X1 U7762 ( .A(n11162), .ZN(n7600) );
  NAND2_X1 U7763 ( .A1(n7597), .A2(n10640), .ZN(n7593) );
  NAND2_X1 U7764 ( .A1(n6577), .A2(n13142), .ZN(n7131) );
  AOI21_X1 U7765 ( .B1(n10606), .B2(n10684), .A(n10607), .ZN(n11233) );
  NAND2_X1 U7766 ( .A1(n7131), .A2(n7130), .ZN(n10606) );
  INV_X1 U7767 ( .A(n13154), .ZN(n10607) );
  NAND2_X1 U7768 ( .A1(n7571), .A2(n7570), .ZN(n7569) );
  NOR2_X1 U7769 ( .A1(n13155), .A2(n10688), .ZN(n7570) );
  INV_X1 U7770 ( .A(n13156), .ZN(n7571) );
  NAND2_X1 U7771 ( .A1(n7574), .A2(n11490), .ZN(n7568) );
  INV_X1 U7772 ( .A(n7699), .ZN(n7698) );
  OAI21_X1 U7773 ( .B1(n7703), .B2(n7700), .A(n6560), .ZN(n7699) );
  OR2_X1 U7774 ( .A1(n10688), .A2(n7706), .ZN(n7700) );
  NAND2_X1 U7775 ( .A1(n11858), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7701) );
  AND2_X1 U7776 ( .A1(n11869), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U7777 ( .A1(n7578), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7577) );
  INV_X1 U7778 ( .A(n10655), .ZN(n7622) );
  NOR2_X1 U7779 ( .A1(n7614), .A2(n7612), .ZN(n7611) );
  INV_X1 U7780 ( .A(n13162), .ZN(n7612) );
  INV_X1 U7781 ( .A(n7615), .ZN(n7614) );
  AND2_X1 U7782 ( .A1(n7616), .A2(n7619), .ZN(n7615) );
  INV_X1 U7783 ( .A(n11856), .ZN(n7616) );
  OR2_X1 U7784 ( .A1(n10613), .A2(n7129), .ZN(n7128) );
  NAND2_X1 U7785 ( .A1(n10695), .A2(n6997), .ZN(n7693) );
  INV_X1 U7786 ( .A(n10618), .ZN(n7562) );
  OR2_X1 U7787 ( .A1(n7547), .A2(n10615), .ZN(n7204) );
  NAND2_X1 U7788 ( .A1(n9802), .A2(n12986), .ZN(n9827) );
  NOR2_X1 U7789 ( .A1(n13442), .A2(n7924), .ZN(n7923) );
  AND2_X1 U7790 ( .A1(n9724), .A2(n9741), .ZN(n7312) );
  NOR2_X1 U7791 ( .A1(n10144), .A2(n7716), .ZN(n7715) );
  INV_X1 U7792 ( .A(n10142), .ZN(n7716) );
  NAND2_X1 U7793 ( .A1(n13118), .A2(n7110), .ZN(n10524) );
  NAND2_X1 U7794 ( .A1(n12211), .A2(n12201), .ZN(n10522) );
  AND2_X1 U7795 ( .A1(n10507), .A2(n6895), .ZN(n10231) );
  OR2_X1 U7796 ( .A1(n9708), .A2(n10775), .ZN(n9424) );
  INV_X1 U7797 ( .A(n11702), .ZN(n10243) );
  NAND2_X1 U7798 ( .A1(n9797), .A2(n9799), .ZN(n7082) );
  AOI21_X1 U7799 ( .B1(n9799), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n9815), .ZN(
        n7083) );
  NOR2_X1 U7800 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n9397) );
  NAND2_X1 U7801 ( .A1(n9784), .A2(n9783), .ZN(n9798) );
  INV_X1 U7802 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9768) );
  AOI21_X1 U7803 ( .B1(n7935), .B2(n7937), .A(n6630), .ZN(n7933) );
  INV_X1 U7804 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U7805 ( .B1(n9704), .B2(n9717), .A(n9719), .ZN(n7456) );
  INV_X1 U7806 ( .A(n7931), .ZN(n7930) );
  OAI21_X1 U7807 ( .B1(n9587), .B2(n7932), .A(n9607), .ZN(n7931) );
  INV_X1 U7808 ( .A(n9589), .ZN(n7932) );
  AOI21_X1 U7809 ( .B1(n7466), .B2(n7463), .A(n6568), .ZN(n7462) );
  INV_X1 U7810 ( .A(n9558), .ZN(n7463) );
  INV_X1 U7811 ( .A(n7742), .ZN(n7741) );
  OAI21_X1 U7812 ( .B1(n13869), .B2(n7743), .A(n13934), .ZN(n7742) );
  AOI21_X1 U7813 ( .B1(n13869), .B2(n7743), .A(n7741), .ZN(n7740) );
  AND2_X1 U7814 ( .A1(n7838), .A2(n6742), .ZN(n6740) );
  NAND2_X1 U7815 ( .A1(n12624), .A2(n7544), .ZN(n12574) );
  INV_X1 U7816 ( .A(n7545), .ZN(n7544) );
  OAI21_X1 U7817 ( .B1(n12570), .B2(n12571), .A(n7546), .ZN(n7545) );
  INV_X1 U7818 ( .A(n11065), .ZN(n6713) );
  NAND2_X1 U7819 ( .A1(n14095), .A2(n11791), .ZN(n11792) );
  OR2_X1 U7820 ( .A1(n6861), .A2(n14420), .ZN(n14187) );
  INV_X1 U7821 ( .A(n9276), .ZN(n9275) );
  AND2_X1 U7822 ( .A1(n6445), .A2(n14527), .ZN(n7883) );
  NOR2_X1 U7823 ( .A1(n10035), .A2(n6689), .ZN(n7069) );
  NOR2_X1 U7824 ( .A1(n14440), .A2(n14277), .ZN(n7884) );
  AND2_X1 U7825 ( .A1(n9950), .A2(n12605), .ZN(n11926) );
  NAND2_X1 U7826 ( .A1(n8028), .A2(n9940), .ZN(n6761) );
  AND2_X1 U7827 ( .A1(n7781), .A2(n9961), .ZN(n7165) );
  NOR2_X1 U7828 ( .A1(n8844), .A2(n8848), .ZN(n9334) );
  OR2_X1 U7829 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n8848) );
  INV_X1 U7830 ( .A(n7978), .ZN(n7977) );
  OAI21_X1 U7831 ( .B1(n14582), .B2(n8498), .A(n8542), .ZN(n7978) );
  INV_X1 U7832 ( .A(n14656), .ZN(n7987) );
  NOR2_X1 U7833 ( .A1(n7213), .A2(n6551), .ZN(n7212) );
  NOR2_X1 U7834 ( .A1(n8533), .A2(n8532), .ZN(n6672) );
  AOI21_X1 U7835 ( .B1(n6980), .B2(n6979), .A(n6695), .ZN(n6694) );
  INV_X1 U7836 ( .A(n7446), .ZN(n7445) );
  OAI21_X1 U7837 ( .B1(n6981), .B2(n6978), .A(n6975), .ZN(n7446) );
  AOI21_X1 U7838 ( .B1(n6977), .B2(n6976), .A(n7447), .ZN(n6975) );
  INV_X1 U7839 ( .A(n6494), .ZN(n6976) );
  INV_X1 U7840 ( .A(n12811), .ZN(n7444) );
  NAND2_X1 U7841 ( .A1(n7487), .A2(n6948), .ZN(n6666) );
  NAND2_X1 U7842 ( .A1(n14935), .A2(n10390), .ZN(n6948) );
  NAND2_X1 U7843 ( .A1(n7487), .A2(n7260), .ZN(n6667) );
  INV_X1 U7844 ( .A(n10389), .ZN(n7260) );
  OR2_X1 U7845 ( .A1(n7968), .A2(n7406), .ZN(n7405) );
  AND2_X1 U7846 ( .A1(n14902), .A2(n10339), .ZN(n7968) );
  INV_X1 U7847 ( .A(n6924), .ZN(n8701) );
  AND2_X1 U7848 ( .A1(n12851), .A2(n10336), .ZN(n7180) );
  NOR2_X1 U7849 ( .A1(n14940), .A2(n14921), .ZN(n7642) );
  AOI21_X1 U7850 ( .B1(n7480), .B2(n15001), .A(n6582), .ZN(n7267) );
  INV_X1 U7851 ( .A(n10386), .ZN(n7857) );
  INV_X1 U7852 ( .A(n7480), .ZN(n7268) );
  AND2_X1 U7853 ( .A1(n14987), .A2(n10384), .ZN(n7480) );
  NOR2_X1 U7854 ( .A1(n7635), .A2(n15188), .ZN(n7634) );
  NAND2_X1 U7855 ( .A1(n15182), .A2(n7636), .ZN(n7635) );
  INV_X1 U7856 ( .A(n6672), .ZN(n8555) );
  OR2_X1 U7857 ( .A1(n14715), .A2(n14586), .ZN(n10372) );
  OR2_X1 U7858 ( .A1(n12738), .A2(n14584), .ZN(n10322) );
  NAND2_X1 U7859 ( .A1(n12181), .A2(n7963), .ZN(n7962) );
  INV_X1 U7860 ( .A(n8059), .ZN(n7963) );
  INV_X1 U7861 ( .A(n7960), .ZN(n7959) );
  OAI21_X1 U7862 ( .B1(n7962), .B2(n7011), .A(n12267), .ZN(n7960) );
  NOR2_X1 U7863 ( .A1(n15234), .A2(n15291), .ZN(n7637) );
  NOR2_X1 U7864 ( .A1(n15597), .A2(n12706), .ZN(n7628) );
  NAND2_X1 U7865 ( .A1(n14936), .A2(n7638), .ZN(n14887) );
  NOR2_X1 U7866 ( .A1(n14890), .A2(n7640), .ZN(n7638) );
  AND2_X1 U7867 ( .A1(n14977), .A2(n15263), .ZN(n14936) );
  NOR2_X2 U7868 ( .A1(n6473), .A2(n14974), .ZN(n14977) );
  INV_X1 U7869 ( .A(n8593), .ZN(n7524) );
  INV_X1 U7870 ( .A(n8592), .ZN(n7523) );
  AND2_X1 U7871 ( .A1(n8546), .A2(n8547), .ZN(n8568) );
  NAND2_X1 U7872 ( .A1(n8119), .A2(SI_17_), .ZN(n8570) );
  NAND2_X1 U7873 ( .A1(n8383), .A2(n8087), .ZN(n6687) );
  AND2_X1 U7874 ( .A1(n8507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U7875 ( .A1(n8075), .A2(SI_4_), .ZN(n7000) );
  INV_X1 U7876 ( .A(n8075), .ZN(n8305) );
  INV_X1 U7877 ( .A(n7327), .ZN(n7325) );
  AND2_X1 U7878 ( .A1(n7328), .A2(n15317), .ZN(n6873) );
  NAND2_X1 U7879 ( .A1(n15316), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U7880 ( .A1(n15321), .A2(n15322), .ZN(n15323) );
  XNOR2_X1 U7881 ( .A(n15323), .B(n7363), .ZN(n15362) );
  NAND2_X1 U7882 ( .A1(n15326), .A2(n15327), .ZN(n15328) );
  INV_X1 U7883 ( .A(n15357), .ZN(n6952) );
  OR2_X1 U7884 ( .A1(n15356), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n6953) );
  INV_X1 U7885 ( .A(n13121), .ZN(n6903) );
  AND2_X1 U7886 ( .A1(n9606), .A2(n9584), .ZN(n7770) );
  NAND3_X1 U7887 ( .A1(n9477), .A2(n6572), .A3(n6454), .ZN(n11299) );
  NAND2_X1 U7888 ( .A1(n13084), .A2(n12894), .ZN(n7766) );
  AND2_X1 U7889 ( .A1(n7320), .A2(n6505), .ZN(n6933) );
  NAND2_X1 U7890 ( .A1(n13817), .A2(n9450), .ZN(n9455) );
  INV_X1 U7891 ( .A(n6918), .ZN(n6915) );
  AND2_X1 U7892 ( .A1(n15798), .A2(n11358), .ZN(n10473) );
  NOR2_X1 U7893 ( .A1(n7759), .A2(n8043), .ZN(n7758) );
  INV_X1 U7894 ( .A(n13072), .ZN(n7759) );
  AND2_X1 U7895 ( .A1(n9532), .A2(n11524), .ZN(n7774) );
  NAND2_X1 U7896 ( .A1(n7319), .A2(n6644), .ZN(n11361) );
  NOR2_X1 U7897 ( .A1(n7768), .A2(n13093), .ZN(n7767) );
  INV_X1 U7898 ( .A(n9698), .ZN(n7768) );
  INV_X1 U7899 ( .A(n10575), .ZN(n7472) );
  AOI21_X1 U7900 ( .B1(n7674), .B2(n7673), .A(n6559), .ZN(n7671) );
  NAND2_X1 U7901 ( .A1(n10586), .A2(n7359), .ZN(n7358) );
  INV_X1 U7902 ( .A(n10428), .ZN(n7359) );
  AND4_X1 U7903 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10457) );
  AND4_X1 U7904 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n11749)
         );
  NAND2_X1 U7905 ( .A1(n10416), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9508) );
  OR2_X1 U7906 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  NAND2_X1 U7907 ( .A1(n9744), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U7908 ( .A1(n10990), .A2(n10991), .ZN(n10989) );
  NAND2_X1 U7909 ( .A1(n10626), .A2(n10676), .ZN(n10986) );
  INV_X1 U7910 ( .A(n10627), .ZN(n10626) );
  XNOR2_X1 U7911 ( .A(n7549), .B(n7206), .ZN(n11019) );
  NAND2_X1 U7912 ( .A1(n11018), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U7913 ( .A1(n7549), .A2(n11033), .ZN(n11149) );
  AOI21_X1 U7914 ( .B1(n11151), .B2(n11149), .A(n11150), .ZN(n11153) );
  AND2_X1 U7915 ( .A1(n6605), .A2(n7686), .ZN(n10682) );
  NAND2_X1 U7916 ( .A1(n7625), .A2(n10687), .ZN(n7624) );
  INV_X1 U7917 ( .A(n10653), .ZN(n7625) );
  NAND2_X1 U7918 ( .A1(n6658), .A2(n7620), .ZN(n7619) );
  INV_X1 U7919 ( .A(n11484), .ZN(n7620) );
  NAND2_X1 U7920 ( .A1(n13163), .A2(n13162), .ZN(n13161) );
  NOR2_X1 U7921 ( .A1(n7577), .A2(n13194), .ZN(n13193) );
  NAND2_X1 U7922 ( .A1(n10610), .A2(n10893), .ZN(n10611) );
  NAND2_X1 U7923 ( .A1(n7583), .A2(n13215), .ZN(n7582) );
  INV_X1 U7924 ( .A(n7588), .ZN(n6991) );
  INV_X1 U7925 ( .A(n7128), .ZN(n13254) );
  NAND2_X1 U7926 ( .A1(n13219), .A2(n7692), .ZN(n7691) );
  XNOR2_X1 U7927 ( .A(n10668), .B(n6997), .ZN(n13247) );
  NOR2_X1 U7928 ( .A1(n13247), .A2(n13246), .ZN(n13245) );
  AOI21_X1 U7929 ( .B1(n10614), .B2(n13738), .A(n7548), .ZN(n7547) );
  INV_X1 U7930 ( .A(n13272), .ZN(n7548) );
  NAND2_X1 U7931 ( .A1(n13254), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U7932 ( .A1(n7690), .A2(n7693), .ZN(n13259) );
  NAND2_X1 U7933 ( .A1(n13259), .A2(n13260), .ZN(n13258) );
  OAI211_X1 U7934 ( .C1(n7205), .C2(n10615), .A(n7204), .B(n13287), .ZN(n10619) );
  NAND2_X1 U7935 ( .A1(n10192), .A2(n13665), .ZN(n12921) );
  INV_X1 U7936 ( .A(n7941), .ZN(n7940) );
  AND2_X1 U7937 ( .A1(n13348), .A2(n13330), .ZN(n13333) );
  NAND2_X1 U7938 ( .A1(n13347), .A2(n13358), .ZN(n13348) );
  NAND2_X1 U7939 ( .A1(n13349), .A2(n15796), .ZN(n13352) );
  INV_X1 U7940 ( .A(n10571), .ZN(n6813) );
  AND2_X1 U7941 ( .A1(n10574), .A2(n10572), .ZN(n13368) );
  AOI21_X1 U7942 ( .B1(n7291), .B2(n10152), .A(n6566), .ZN(n7290) );
  NAND2_X1 U7943 ( .A1(n7303), .A2(n7302), .ZN(n9923) );
  INV_X1 U7944 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U7945 ( .A1(n6904), .A2(n7504), .ZN(n13376) );
  AOI21_X1 U7946 ( .B1(n7506), .B2(n10563), .A(n7505), .ZN(n7504) );
  NAND2_X1 U7947 ( .A1(n10237), .A2(n7506), .ZN(n6904) );
  INV_X1 U7948 ( .A(n10567), .ZN(n7505) );
  AND2_X1 U7949 ( .A1(n10565), .A2(n6828), .ZN(n7508) );
  NAND2_X1 U7950 ( .A1(n13420), .A2(n10467), .ZN(n10237) );
  OAI21_X1 U7951 ( .B1(n13455), .B2(n10450), .A(n10449), .ZN(n13443) );
  NAND2_X1 U7952 ( .A1(n13443), .A2(n13442), .ZN(n13441) );
  OAI21_X1 U7953 ( .B1(n13494), .B2(n13477), .A(n6567), .ZN(n13451) );
  NAND2_X1 U7954 ( .A1(n13482), .A2(n10538), .ZN(n6902) );
  NAND2_X1 U7955 ( .A1(n7296), .A2(n7294), .ZN(n13464) );
  NOR2_X1 U7956 ( .A1(n7295), .A2(n13467), .ZN(n7294) );
  INV_X1 U7957 ( .A(n7379), .ZN(n7295) );
  AND2_X1 U7958 ( .A1(n9749), .A2(n9748), .ZN(n13469) );
  AND2_X1 U7959 ( .A1(n9765), .A2(n9764), .ZN(n13480) );
  NAND2_X1 U7960 ( .A1(n13494), .A2(n10535), .ZN(n13483) );
  NAND2_X1 U7961 ( .A1(n13483), .A2(n13482), .ZN(n13481) );
  NAND2_X1 U7962 ( .A1(n7713), .A2(n13522), .ZN(n7712) );
  AND2_X1 U7963 ( .A1(n10533), .A2(n10535), .ZN(n13495) );
  AND2_X1 U7964 ( .A1(n10532), .A2(n10536), .ZN(n13508) );
  INV_X1 U7965 ( .A(n6900), .ZN(n6899) );
  OAI21_X1 U7966 ( .B1(n13517), .B2(n6901), .A(n13508), .ZN(n6900) );
  INV_X1 U7967 ( .A(n10530), .ZN(n6901) );
  NAND2_X1 U7968 ( .A1(n12210), .A2(n12205), .ZN(n6849) );
  NAND2_X1 U7969 ( .A1(n7106), .A2(n6533), .ZN(n7105) );
  INV_X1 U7970 ( .A(n10233), .ZN(n7497) );
  AND3_X1 U7971 ( .A1(n9678), .A2(n9677), .A3(n9676), .ZN(n13045) );
  NAND2_X1 U7972 ( .A1(n7286), .A2(n7344), .ZN(n10139) );
  INV_X1 U7973 ( .A(n10235), .ZN(n12001) );
  AND2_X1 U7974 ( .A1(n10524), .A2(n10522), .ZN(n10235) );
  AND2_X1 U7975 ( .A1(n10235), .A2(n10525), .ZN(n7939) );
  NAND2_X1 U7976 ( .A1(n7502), .A2(n10233), .ZN(n7500) );
  NAND2_X1 U7977 ( .A1(n11878), .A2(n7502), .ZN(n7501) );
  OR2_X1 U7978 ( .A1(n12092), .A2(n12091), .ZN(n12094) );
  NAND2_X1 U7979 ( .A1(n11612), .A2(n10228), .ZN(n10229) );
  AND2_X1 U7980 ( .A1(n9560), .A2(n9559), .ZN(n11607) );
  OR2_X1 U7981 ( .A1(n13125), .A2(n11547), .ZN(n11611) );
  AND3_X1 U7982 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(n10130) );
  NAND2_X1 U7983 ( .A1(n9525), .A2(n9524), .ZN(n9544) );
  NAND2_X1 U7984 ( .A1(n10440), .A2(n6836), .ZN(n6833) );
  INV_X1 U7985 ( .A(n11365), .ZN(n11440) );
  BUF_X1 U7986 ( .A(n10440), .Z(n15781) );
  AND2_X1 U7987 ( .A1(n9466), .A2(n9465), .ZN(n15795) );
  AND2_X1 U7988 ( .A1(n9910), .A2(n6417), .ZN(n15799) );
  OAI211_X1 U7989 ( .C1(n11315), .C2(n11314), .A(n11313), .B(n11312), .ZN(
        n11318) );
  NAND2_X1 U7990 ( .A1(n9801), .A2(n9800), .ZN(n12988) );
  NAND2_X1 U7991 ( .A1(n9786), .A2(n9785), .ZN(n13037) );
  NAND2_X1 U7992 ( .A1(n9758), .A2(n9757), .ZN(n13587) );
  NAND2_X1 U7993 ( .A1(n15805), .A2(n15841), .ZN(n15851) );
  INV_X1 U7994 ( .A(n15783), .ZN(n15796) );
  CLKBUF_X1 U7995 ( .A(n9878), .Z(n10800) );
  OR2_X1 U7996 ( .A1(n13819), .A2(n9411), .ZN(n6853) );
  NAND2_X1 U7997 ( .A1(n7945), .A2(n7946), .ZN(n10408) );
  AOI21_X1 U7998 ( .B1(n7947), .B2(n10185), .A(n6650), .ZN(n7946) );
  NAND2_X1 U7999 ( .A1(n7468), .A2(n7944), .ZN(n7471) );
  AND2_X1 U8000 ( .A1(n10156), .A2(n6655), .ZN(n7468) );
  XNOR2_X1 U8001 ( .A(n10155), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n10154) );
  NOR2_X1 U8002 ( .A1(n9841), .A2(n7452), .ZN(n6827) );
  INV_X1 U8003 ( .A(n7083), .ZN(n7081) );
  NAND2_X1 U8004 ( .A1(n7082), .A2(n9836), .ZN(n7077) );
  NOR2_X1 U8005 ( .A1(n9893), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U8006 ( .A1(n7082), .A2(n7083), .ZN(n9818) );
  OR2_X1 U8007 ( .A1(n9426), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n9446) );
  INV_X1 U8008 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9448) );
  XNOR2_X1 U8009 ( .A(n9798), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9797) );
  INV_X1 U8010 ( .A(n7933), .ZN(n7089) );
  INV_X1 U8011 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U8012 ( .A1(n6820), .A2(n6824), .ZN(n9705) );
  INV_X1 U8013 ( .A(n6825), .ZN(n6824) );
  NAND2_X1 U8014 ( .A1(n7449), .A2(n6821), .ZN(n6820) );
  OAI21_X1 U8015 ( .B1(n9658), .B2(n6618), .A(n9700), .ZN(n6825) );
  OR2_X1 U8016 ( .A1(n6476), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U8017 ( .A1(n9627), .A2(n9626), .ZN(n9642) );
  XNOR2_X1 U8018 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .ZN(n9607) );
  AND2_X1 U8019 ( .A1(n10747), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9556) );
  XNOR2_X1 U8020 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .ZN(n9572) );
  NAND2_X1 U8021 ( .A1(n7101), .A2(n9537), .ZN(n9557) );
  NAND2_X1 U8022 ( .A1(n9536), .A2(n9535), .ZN(n7101) );
  AND2_X1 U8023 ( .A1(n7777), .A2(n9476), .ZN(n7150) );
  NAND2_X1 U8024 ( .A1(n7778), .A2(n7777), .ZN(n9475) );
  NAND2_X1 U8025 ( .A1(n7777), .A2(n7241), .ZN(n7240) );
  INV_X1 U8026 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7241) );
  OR2_X1 U8027 ( .A1(n14571), .A2(n9342), .ZN(n10596) );
  NOR2_X1 U8028 ( .A1(n11427), .A2(n7273), .ZN(n7272) );
  INV_X1 U8029 ( .A(n8978), .ZN(n7273) );
  XNOR2_X1 U8030 ( .A(n13920), .B(n13919), .ZN(n13856) );
  NAND2_X1 U8031 ( .A1(n11694), .A2(n6434), .ZN(n7270) );
  NAND2_X1 U8032 ( .A1(n11383), .A2(n7271), .ZN(n6773) );
  AND2_X1 U8033 ( .A1(n7272), .A2(n11694), .ZN(n7271) );
  NAND2_X1 U8034 ( .A1(n6773), .A2(n6771), .ZN(n11844) );
  NOR2_X1 U8035 ( .A1(n6432), .A2(n6772), .ZN(n6771) );
  INV_X1 U8036 ( .A(n11845), .ZN(n6772) );
  INV_X1 U8037 ( .A(n8897), .ZN(n7725) );
  NAND2_X1 U8038 ( .A1(n8898), .A2(n8897), .ZN(n7727) );
  INV_X1 U8039 ( .A(n13842), .ZN(n9128) );
  NAND2_X1 U8040 ( .A1(n7793), .A2(n12912), .ZN(n7797) );
  NAND2_X1 U8041 ( .A1(n7795), .A2(n7794), .ZN(n7793) );
  NAND2_X1 U8042 ( .A1(n14563), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U8043 ( .A1(n8894), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U8044 ( .A1(n7278), .A2(n7276), .ZN(n12288) );
  NAND2_X1 U8045 ( .A1(n13959), .A2(n13961), .ZN(n13960) );
  NAND2_X1 U8046 ( .A1(n9138), .A2(n6465), .ZN(n9180) );
  NOR2_X1 U8047 ( .A1(n7734), .A2(n9169), .ZN(n7733) );
  NOR2_X1 U8048 ( .A1(n7735), .A2(n9127), .ZN(n7734) );
  INV_X1 U8049 ( .A(n9174), .ZN(n7731) );
  INV_X1 U8050 ( .A(n7735), .ZN(n7732) );
  NOR2_X1 U8051 ( .A1(n12625), .A2(n8895), .ZN(n11051) );
  NOR2_X1 U8052 ( .A1(n6719), .A2(n11064), .ZN(n6717) );
  NAND2_X1 U8053 ( .A1(n15682), .A2(n15680), .ZN(n11787) );
  INV_X1 U8054 ( .A(n14131), .ZN(n6722) );
  NOR2_X1 U8055 ( .A1(n6442), .A2(n7195), .ZN(n7192) );
  INV_X1 U8056 ( .A(n14203), .ZN(n7349) );
  NAND2_X1 U8057 ( .A1(n7382), .A2(n7804), .ZN(n6682) );
  AND2_X1 U8058 ( .A1(n7385), .A2(n7387), .ZN(n7382) );
  NAND2_X1 U8059 ( .A1(n7070), .A2(n7069), .ZN(n14234) );
  AND2_X1 U8060 ( .A1(n9976), .A2(n6681), .ZN(n7806) );
  INV_X1 U8061 ( .A(n9974), .ZN(n7807) );
  OR2_X1 U8062 ( .A1(n14277), .A2(n14255), .ZN(n9974) );
  OR2_X1 U8063 ( .A1(n9209), .A2(n9208), .ZN(n9231) );
  NOR2_X1 U8064 ( .A1(n14300), .A2(n7396), .ZN(n7395) );
  INV_X1 U8065 ( .A(n9967), .ZN(n7396) );
  OR2_X1 U8066 ( .A1(n14313), .A2(n9966), .ZN(n7397) );
  AOI21_X1 U8067 ( .B1(n7061), .B2(n7060), .A(n8006), .ZN(n7059) );
  INV_X1 U8068 ( .A(n10024), .ZN(n7060) );
  NAND2_X1 U8069 ( .A1(n7063), .A2(n10024), .ZN(n7062) );
  INV_X1 U8070 ( .A(n14476), .ZN(n7063) );
  NAND2_X1 U8071 ( .A1(n6858), .A2(n13902), .ZN(n8013) );
  INV_X1 U8072 ( .A(n9960), .ZN(n7785) );
  AOI21_X1 U8073 ( .B1(n8017), .B2(n8019), .A(n6543), .ZN(n8016) );
  NAND2_X1 U8074 ( .A1(n9088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U8075 ( .A1(n11930), .A2(n9957), .ZN(n12151) );
  NAND2_X1 U8076 ( .A1(n12151), .A2(n12150), .ZN(n12149) );
  NOR2_X1 U8077 ( .A1(n12608), .A2(n10018), .ZN(n8020) );
  OR2_X1 U8078 ( .A1(n6501), .A2(n8058), .ZN(n8033) );
  NAND2_X1 U8079 ( .A1(n11530), .A2(n6482), .ZN(n11731) );
  INV_X1 U8080 ( .A(n7800), .ZN(n7799) );
  OAI21_X1 U8081 ( .B1(n7802), .B2(n12598), .A(n12596), .ZN(n7800) );
  NAND2_X1 U8082 ( .A1(n9009), .A2(n10740), .ZN(n7071) );
  NAND2_X1 U8083 ( .A1(n7189), .A2(n12942), .ZN(n7188) );
  NAND2_X1 U8084 ( .A1(n11576), .A2(n9933), .ZN(n11035) );
  AND2_X1 U8085 ( .A1(n11051), .A2(n11074), .ZN(n14376) );
  INV_X1 U8086 ( .A(n14376), .ZN(n14329) );
  INV_X1 U8087 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8903) );
  OAI21_X1 U8088 ( .B1(n10280), .B2(n7158), .A(n7155), .ZN(n7159) );
  AOI21_X1 U8089 ( .B1(n10279), .B2(n7157), .A(n7156), .ZN(n7155) );
  NOR2_X1 U8090 ( .A1(n7158), .A2(n12620), .ZN(n7157) );
  NOR2_X1 U8091 ( .A1(n14379), .A2(n7158), .ZN(n7156) );
  NAND2_X1 U8092 ( .A1(n7072), .A2(n15764), .ZN(n10283) );
  NAND2_X1 U8093 ( .A1(n9177), .A2(n9176), .ZN(n14466) );
  NAND2_X1 U8094 ( .A1(n9013), .A2(n9012), .ZN(n14509) );
  NAND2_X1 U8095 ( .A1(n11663), .A2(n10044), .ZN(n11570) );
  AND2_X1 U8096 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n8875) );
  INV_X1 U8097 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9133) );
  AND2_X1 U8098 ( .A1(n7215), .A2(n7216), .ZN(n14581) );
  NAND2_X1 U8099 ( .A1(n14581), .A2(n14582), .ZN(n14580) );
  NOR2_X1 U8100 ( .A1(n7974), .A2(n7971), .ZN(n7970) );
  INV_X1 U8101 ( .A(n14619), .ZN(n7971) );
  NAND2_X1 U8102 ( .A1(n14609), .A2(n7990), .ZN(n7989) );
  INV_X1 U8103 ( .A(n7991), .ZN(n7990) );
  NOR2_X1 U8104 ( .A1(n11707), .A2(n7982), .ZN(n7981) );
  AND2_X1 U8105 ( .A1(n12218), .A2(n7212), .ZN(n7208) );
  NAND2_X1 U8106 ( .A1(n14637), .A2(n14638), .ZN(n14636) );
  AOI21_X1 U8107 ( .B1(n7232), .B2(n7230), .A(n8613), .ZN(n7229) );
  INV_X1 U8108 ( .A(n14673), .ZN(n7230) );
  INV_X1 U8109 ( .A(n7232), .ZN(n7231) );
  INV_X1 U8110 ( .A(n6678), .ZN(n8656) );
  INV_X1 U8111 ( .A(n11125), .ZN(n8246) );
  INV_X1 U8112 ( .A(n7378), .ZN(n7980) );
  NOR2_X1 U8113 ( .A1(n12878), .A2(n8814), .ZN(n11826) );
  NAND2_X1 U8114 ( .A1(n8485), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8533) );
  AND2_X1 U8115 ( .A1(n8605), .A2(n8604), .ZN(n14677) );
  NAND2_X1 U8116 ( .A1(n8226), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8215) );
  INV_X1 U8117 ( .A(n6890), .ZN(n7179) );
  NAND2_X1 U8118 ( .A1(n10725), .A2(n6518), .ZN(n10838) );
  OR2_X1 U8119 ( .A1(n7021), .A2(n14756), .ZN(n7029) );
  OR2_X1 U8120 ( .A1(n14752), .A2(n7031), .ZN(n7021) );
  NAND2_X1 U8121 ( .A1(n7023), .A2(n14773), .ZN(n7028) );
  INV_X1 U8122 ( .A(n10850), .ZN(n7023) );
  NAND2_X1 U8123 ( .A1(n7020), .A2(n6439), .ZN(n7025) );
  INV_X1 U8124 ( .A(n7029), .ZN(n7020) );
  OAI21_X1 U8125 ( .B1(n14772), .B2(n7022), .A(n6439), .ZN(n7026) );
  INV_X1 U8126 ( .A(n7028), .ZN(n7022) );
  NAND2_X1 U8127 ( .A1(n10931), .A2(n7424), .ZN(n7421) );
  INV_X1 U8128 ( .A(n6486), .ZN(n7420) );
  OR2_X1 U8129 ( .A1(n8443), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8445) );
  NOR2_X1 U8130 ( .A1(n11143), .A2(n11142), .ZN(n11284) );
  OR2_X1 U8131 ( .A1(n8385), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8507) );
  INV_X1 U8132 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8065) );
  AND2_X1 U8133 ( .A1(n8746), .A2(n8723), .ZN(n14885) );
  NAND2_X1 U8134 ( .A1(n14914), .A2(n10339), .ZN(n14896) );
  NAND2_X1 U8135 ( .A1(n14936), .A2(n7642), .ZN(n14919) );
  INV_X1 U8136 ( .A(n8062), .ZN(n7851) );
  NAND2_X1 U8137 ( .A1(n14970), .A2(n6503), .ZN(n14947) );
  NAND2_X1 U8138 ( .A1(n10385), .A2(n7480), .ZN(n14986) );
  AND2_X1 U8139 ( .A1(n8177), .A2(n8176), .ZN(n14611) );
  AOI21_X1 U8140 ( .B1(n10325), .B2(n6700), .A(n6699), .ZN(n10329) );
  INV_X1 U8141 ( .A(n15004), .ZN(n6700) );
  NOR2_X1 U8142 ( .A1(n10380), .A2(n7258), .ZN(n7257) );
  NAND2_X1 U8143 ( .A1(n6565), .A2(n12350), .ZN(n6787) );
  AND2_X1 U8144 ( .A1(n10373), .A2(n10369), .ZN(n7485) );
  NOR2_X1 U8145 ( .A1(n15070), .A2(n15069), .ZN(n10373) );
  NAND2_X1 U8146 ( .A1(n7854), .A2(n7476), .ZN(n12306) );
  AOI21_X1 U8147 ( .B1(n6435), .B2(n7856), .A(n6541), .ZN(n7854) );
  OAI211_X1 U8148 ( .C1(n11719), .C2(n7479), .A(n7478), .B(n6435), .ZN(n7476)
         );
  OAI21_X1 U8149 ( .B1(n7959), .B2(n7010), .A(n10317), .ZN(n7005) );
  OR2_X1 U8150 ( .A1(n7958), .A2(n7010), .ZN(n7006) );
  AOI21_X1 U8151 ( .B1(n10306), .B2(n7950), .A(n6545), .ZN(n7949) );
  INV_X1 U8152 ( .A(n10305), .ZN(n7950) );
  NAND2_X1 U8153 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8323) );
  NAND2_X1 U8154 ( .A1(n7840), .A2(n11204), .ZN(n7474) );
  NAND2_X1 U8155 ( .A1(n6574), .A2(n11824), .ZN(n7475) );
  NAND2_X1 U8156 ( .A1(n12668), .A2(n12667), .ZN(n11824) );
  NAND2_X1 U8157 ( .A1(n12676), .A2(n7957), .ZN(n7956) );
  INV_X1 U8158 ( .A(n14675), .ZN(n15111) );
  NAND2_X1 U8159 ( .A1(n10077), .A2(n10076), .ZN(n14826) );
  OR2_X1 U8160 ( .A1(n11828), .A2(n12814), .ZN(n15588) );
  AND2_X1 U8161 ( .A1(n8797), .A2(n8812), .ZN(n15598) );
  NAND2_X1 U8162 ( .A1(n6632), .A2(n6464), .ZN(n7543) );
  AND2_X1 U8163 ( .A1(n8151), .A2(n8150), .ZN(n8790) );
  OAI211_X1 U8164 ( .C1(n7119), .C2(n8692), .A(n7117), .B(n7114), .ZN(n8717)
         );
  AOI21_X1 U8165 ( .B1(n8693), .B2(n7118), .A(n6627), .ZN(n7117) );
  OR2_X1 U8166 ( .A1(n9218), .A2(n7115), .ZN(n7114) );
  NOR2_X1 U8167 ( .A1(n8160), .A2(n8147), .ZN(n7352) );
  XNOR2_X1 U8168 ( .A(n6680), .B(n8653), .ZN(n12098) );
  OAI21_X1 U8169 ( .B1(n9218), .B2(n8652), .A(n8651), .ZN(n6680) );
  NAND2_X1 U8170 ( .A1(n7907), .A2(n7906), .ZN(n8793) );
  AND2_X1 U8171 ( .A1(n8161), .A2(n8179), .ZN(n7906) );
  INV_X1 U8172 ( .A(n8160), .ZN(n7907) );
  INV_X1 U8173 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U8174 ( .A1(n7516), .A2(n7518), .ZN(n8632) );
  NAND2_X1 U8175 ( .A1(n8593), .A2(n7521), .ZN(n7516) );
  XNOR2_X1 U8176 ( .A(n6947), .B(n8504), .ZN(n11257) );
  OAI21_X1 U8177 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n6947) );
  AND2_X1 U8178 ( .A1(n8482), .A2(n8467), .ZN(n11684) );
  OR2_X1 U8179 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  AOI21_X1 U8180 ( .B1(n8088), .B2(n6688), .A(n6855), .ZN(n6854) );
  NAND2_X1 U8181 ( .A1(n7111), .A2(n8087), .ZN(n8402) );
  NAND2_X1 U8182 ( .A1(n8901), .A2(n8234), .ZN(n8216) );
  XNOR2_X1 U8183 ( .A(n15363), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n15365) );
  NAND2_X1 U8184 ( .A1(n6878), .A2(n7860), .ZN(n6877) );
  INV_X1 U8185 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7860) );
  INV_X1 U8186 ( .A(n15431), .ZN(n6879) );
  NAND2_X1 U8187 ( .A1(n7875), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7874) );
  INV_X1 U8188 ( .A(n15460), .ZN(n7875) );
  OAI21_X1 U8189 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15343), .A(n15342), .ZN(
        n15352) );
  AOI21_X1 U8190 ( .B1(n7870), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7871), .ZN(
        n7869) );
  NAND2_X1 U8191 ( .A1(n7871), .A2(n7867), .ZN(n7866) );
  INV_X1 U8192 ( .A(n7874), .ZN(n7867) );
  NAND2_X1 U8193 ( .A1(n7873), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7868) );
  OAI21_X1 U8194 ( .B1(n7874), .B2(n6491), .A(n15463), .ZN(n7873) );
  AND2_X1 U8195 ( .A1(n7340), .A2(n15465), .ZN(n15412) );
  OAI21_X1 U8196 ( .B1(n15466), .B2(n15467), .A(n7342), .ZN(n7340) );
  INV_X1 U8197 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U8198 ( .A1(n9672), .A2(n9671), .ZN(n13523) );
  AND2_X1 U8199 ( .A1(n9793), .A2(n9792), .ZN(n13457) );
  NAND2_X1 U8200 ( .A1(n9723), .A2(n9722), .ZN(n13497) );
  NAND2_X1 U8201 ( .A1(n9740), .A2(n9739), .ZN(n13484) );
  AOI21_X1 U8202 ( .B1(n6910), .B2(n9867), .A(n6909), .ZN(n6906) );
  NOR2_X1 U8203 ( .A1(n13007), .A2(n13106), .ZN(n6910) );
  AND2_X1 U8204 ( .A1(n6912), .A2(n9873), .ZN(n6909) );
  AOI21_X1 U8205 ( .B1(n9868), .B2(n6912), .A(n13100), .ZN(n6908) );
  NOR2_X1 U8206 ( .A1(n7756), .A2(n9873), .ZN(n6911) );
  AND3_X1 U8207 ( .A1(n9504), .A2(n9503), .A3(n9502), .ZN(n11509) );
  OR2_X1 U8208 ( .A1(n9708), .A2(SI_4_), .ZN(n9504) );
  NAND2_X1 U8209 ( .A1(n9826), .A2(n9825), .ZN(n13057) );
  AND2_X1 U8210 ( .A1(n13086), .A2(n15799), .ZN(n13076) );
  AOI21_X1 U8211 ( .B1(n10180), .B2(n13458), .A(n9776), .ZN(n13470) );
  INV_X1 U8212 ( .A(n13088), .ZN(n13094) );
  NAND2_X1 U8213 ( .A1(n11361), .A2(n7774), .ZN(n11523) );
  INV_X1 U8214 ( .A(n13084), .ZN(n6956) );
  NAND2_X1 U8215 ( .A1(n13833), .A2(n10424), .ZN(n10165) );
  INV_X1 U8216 ( .A(n13083), .ZN(n13098) );
  OAI21_X1 U8217 ( .B1(n13370), .B2(n9561), .A(n7297), .ZN(n13350) );
  NOR2_X1 U8218 ( .A1(n6623), .A2(n7298), .ZN(n7297) );
  NAND2_X1 U8219 ( .A1(n10169), .A2(n10168), .ZN(n7298) );
  NAND4_X1 U8220 ( .A1(n9581), .A2(n9580), .A3(n9579), .A4(n9578), .ZN(n13122)
         );
  OR2_X1 U8221 ( .A1(n9506), .A2(n15861), .ZN(n6839) );
  AND3_X1 U8222 ( .A1(n9416), .A2(n9414), .A3(n9415), .ZN(n6838) );
  NAND2_X1 U8223 ( .A1(n7145), .A2(n10658), .ZN(n7144) );
  NAND2_X1 U8224 ( .A1(n13199), .A2(n13198), .ZN(n13197) );
  NAND2_X1 U8225 ( .A1(n7200), .A2(n6470), .ZN(n7127) );
  NOR2_X1 U8226 ( .A1(n10716), .A2(n10715), .ZN(n6998) );
  OAI21_X1 U8227 ( .B1(n7559), .B2(n7556), .A(n7555), .ZN(n7554) );
  NAND2_X1 U8228 ( .A1(n7293), .A2(n7291), .ZN(n13382) );
  NAND2_X1 U8229 ( .A1(n7293), .A2(n10153), .ZN(n13380) );
  NAND2_X1 U8230 ( .A1(n9843), .A2(n9842), .ZN(n13411) );
  NAND2_X1 U8231 ( .A1(n11782), .A2(n10424), .ZN(n9843) );
  NAND2_X1 U8232 ( .A1(n9770), .A2(n9769), .ZN(n13794) );
  OR2_X1 U8233 ( .A1(n9417), .A2(n9411), .ZN(n6913) );
  NAND2_X1 U8234 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  NAND2_X1 U8235 ( .A1(n13974), .A2(n9301), .ZN(n10056) );
  NAND2_X1 U8236 ( .A1(n12360), .A2(n9115), .ZN(n13842) );
  NAND2_X1 U8237 ( .A1(n9120), .A2(n9119), .ZN(n14490) );
  AND2_X1 U8238 ( .A1(n9257), .A2(n9256), .ZN(n14256) );
  NOR2_X1 U8239 ( .A1(n10055), .A2(n7751), .ZN(n7750) );
  INV_X1 U8240 ( .A(n9301), .ZN(n7751) );
  INV_X1 U8241 ( .A(n14285), .ZN(n14255) );
  AND2_X1 U8242 ( .A1(n9282), .A2(n9281), .ZN(n13980) );
  OR2_X1 U8243 ( .A1(n14218), .A2(n9326), .ZN(n9282) );
  AND2_X1 U8244 ( .A1(n9238), .A2(n9237), .ZN(n14303) );
  INV_X1 U8245 ( .A(n6776), .ZN(n6775) );
  OR2_X1 U8246 ( .A1(n7278), .A2(n6495), .ZN(n6774) );
  OAI21_X1 U8247 ( .B1(n7276), .B2(n6495), .A(n12321), .ZN(n6776) );
  OR2_X1 U8248 ( .A1(n9383), .A2(n12640), .ZN(n13952) );
  AND2_X1 U8249 ( .A1(n9314), .A2(n9313), .ZN(n13979) );
  NAND2_X1 U8250 ( .A1(n9290), .A2(n9289), .ZN(n14425) );
  NAND2_X1 U8251 ( .A1(n9373), .A2(n14385), .ZN(n13998) );
  NAND2_X1 U8252 ( .A1(n9331), .A2(n9330), .ZN(n14005) );
  OR2_X1 U8253 ( .A1(n12932), .A2(n9326), .ZN(n9331) );
  INV_X1 U8254 ( .A(n13979), .ZN(n14196) );
  OR2_X1 U8255 ( .A1(n14201), .A2(n9326), .ZN(n9298) );
  INV_X1 U8256 ( .A(n13980), .ZN(n14226) );
  NAND2_X1 U8257 ( .A1(n9186), .A2(n9185), .ZN(n14360) );
  OR2_X1 U8258 ( .A1(n9126), .A2(n9125), .ZN(n14010) );
  NAND4_X1 U8259 ( .A1(n8986), .A2(n8985), .A3(n8984), .A4(n8983), .ZN(n14019)
         );
  NAND4_X1 U8260 ( .A1(n8972), .A2(n8971), .A3(n8970), .A4(n8969), .ZN(n14020)
         );
  NAND2_X1 U8261 ( .A1(n6711), .A2(n11061), .ZN(n14061) );
  NAND2_X1 U8262 ( .A1(n15655), .A2(n14047), .ZN(n6711) );
  NAND2_X1 U8263 ( .A1(n6945), .A2(n6944), .ZN(n14159) );
  INV_X1 U8264 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6944) );
  INV_X1 U8265 ( .A(n14139), .ZN(n6945) );
  NOR2_X1 U8266 ( .A1(n8857), .A2(n8048), .ZN(n8858) );
  NAND2_X1 U8267 ( .A1(n9154), .A2(n8852), .ZN(n8859) );
  NAND2_X1 U8268 ( .A1(n14476), .A2(n10023), .ZN(n14354) );
  INV_X1 U8269 ( .A(n12552), .ZN(n14516) );
  AND2_X1 U8270 ( .A1(n14407), .A2(n14410), .ZN(n14513) );
  OAI211_X1 U8271 ( .C1(n14418), .C2(n15748), .A(n14416), .B(n14417), .ZN(
        n14521) );
  NAND2_X1 U8272 ( .A1(n9365), .A2(n9364), .ZN(n15721) );
  NAND3_X1 U8273 ( .A1(n7896), .A2(n7897), .A3(n6540), .ZN(n8889) );
  INV_X1 U8274 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8888) );
  INV_X1 U8275 ( .A(n14386), .ZN(n12630) );
  NOR2_X1 U8276 ( .A1(n7223), .A2(n14717), .ZN(n7221) );
  NOR2_X1 U8277 ( .A1(n7226), .A2(n7224), .ZN(n7223) );
  INV_X1 U8278 ( .A(n7227), .ZN(n7224) );
  NAND2_X1 U8279 ( .A1(n7227), .A2(n7228), .ZN(n7225) );
  NOR2_X1 U8280 ( .A1(n14657), .A2(n14656), .ZN(n14655) );
  AND2_X1 U8281 ( .A1(n8820), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14698) );
  NAND2_X1 U8282 ( .A1(n7975), .A2(n8714), .ZN(n7353) );
  NAND2_X1 U8283 ( .A1(n8663), .A2(n8662), .ZN(n14725) );
  OR2_X1 U8284 ( .A1(n14594), .A2(n8267), .ZN(n8663) );
  INV_X1 U8285 ( .A(n14707), .ZN(n14731) );
  NAND2_X1 U8286 ( .A1(n14758), .A2(n14759), .ZN(n14757) );
  XNOR2_X1 U8287 ( .A(n7425), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U8288 ( .A1(n8281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U8289 ( .A1(n11186), .A2(n6526), .ZN(n10843) );
  NAND2_X1 U8290 ( .A1(n10945), .A2(n6705), .ZN(n10963) );
  NAND2_X1 U8291 ( .A1(n6706), .A2(n10921), .ZN(n6705) );
  OR2_X1 U8292 ( .A1(n10963), .A2(n7416), .ZN(n7413) );
  INV_X1 U8293 ( .A(n7417), .ZN(n7416) );
  AOI21_X1 U8294 ( .B1(n7417), .B2(n7415), .A(n6576), .ZN(n7414) );
  INV_X1 U8295 ( .A(n10962), .ZN(n7415) );
  AND2_X1 U8296 ( .A1(n7413), .A2(n7411), .ZN(n11282) );
  NOR2_X1 U8297 ( .A1(n7412), .A2(n11138), .ZN(n7411) );
  INV_X1 U8298 ( .A(n7414), .ZN(n7412) );
  NOR2_X1 U8299 ( .A1(n11284), .A2(n7018), .ZN(n11286) );
  NOR2_X1 U8300 ( .A1(n7019), .A2(n12276), .ZN(n7018) );
  NAND2_X1 U8301 ( .A1(n11286), .A2(n11287), .ZN(n11466) );
  AOI21_X1 U8302 ( .B1(n15474), .B2(n15473), .A(n6527), .ZN(n12080) );
  NAND2_X1 U8303 ( .A1(n12080), .A2(n12079), .ZN(n14779) );
  OAI21_X1 U8304 ( .B1(n14818), .B2(n14817), .A(n14765), .ZN(n7035) );
  XNOR2_X1 U8305 ( .A(n6707), .B(n14808), .ZN(n14818) );
  NAND2_X1 U8306 ( .A1(n7427), .A2(n6708), .ZN(n6707) );
  INV_X1 U8307 ( .A(n14807), .ZN(n6708) );
  XNOR2_X1 U8308 ( .A(n14815), .B(n7036), .ZN(n14816) );
  OR2_X1 U8309 ( .A1(n15483), .A2(n8065), .ZN(n7431) );
  NAND2_X1 U8310 ( .A1(n14850), .A2(n6785), .ZN(n14853) );
  NAND2_X1 U8311 ( .A1(n12804), .A2(n14839), .ZN(n6785) );
  INV_X1 U8312 ( .A(n14836), .ZN(n14837) );
  INV_X1 U8313 ( .A(n7174), .ZN(n7173) );
  NAND2_X1 U8314 ( .A1(n7858), .A2(n10391), .ZN(n14865) );
  OAI21_X1 U8315 ( .B1(n7853), .B2(n7489), .A(n7487), .ZN(n7858) );
  NAND2_X2 U8316 ( .A1(n8743), .A2(n8742), .ZN(n14880) );
  NAND2_X1 U8317 ( .A1(n14895), .A2(n10340), .ZN(n14884) );
  NAND2_X1 U8318 ( .A1(n14899), .A2(n10390), .ZN(n14892) );
  NAND2_X1 U8319 ( .A1(n7012), .A2(n14898), .ZN(n15147) );
  NAND2_X1 U8320 ( .A1(n7013), .A2(n15604), .ZN(n7012) );
  NAND2_X1 U8321 ( .A1(n7014), .A2(n14895), .ZN(n7013) );
  NAND2_X1 U8322 ( .A1(n14896), .A2(n14897), .ZN(n7014) );
  NAND2_X1 U8323 ( .A1(n7853), .A2(n7852), .ZN(n14901) );
  INV_X1 U8324 ( .A(n7850), .ZN(n7852) );
  INV_X1 U8325 ( .A(n15531), .ZN(n15511) );
  OAI21_X1 U8326 ( .B1(n8575), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8187) );
  NOR2_X1 U8327 ( .A1(n7492), .A2(n8137), .ZN(n7491) );
  AND2_X1 U8328 ( .A1(n8131), .A2(n8463), .ZN(n6881) );
  NAND2_X1 U8329 ( .A1(n8141), .A2(n8166), .ZN(n7492) );
  XNOR2_X1 U8330 ( .A(n15367), .B(P1_ADDR_REG_2__SCAN_IN), .ZN(n7341) );
  INV_X1 U8331 ( .A(n15392), .ZN(n6942) );
  NAND2_X1 U8332 ( .A1(n7336), .A2(n7329), .ZN(n15425) );
  AND2_X1 U8333 ( .A1(n7330), .A2(n15426), .ZN(n7329) );
  NAND2_X1 U8334 ( .A1(n15430), .A2(n15431), .ZN(n15429) );
  OR2_X1 U8335 ( .A1(n15455), .A2(n15405), .ZN(n6862) );
  NOR2_X1 U8336 ( .A1(n6491), .A2(n15463), .ZN(n7871) );
  INV_X1 U8337 ( .A(n6491), .ZN(n7870) );
  NAND2_X1 U8338 ( .A1(n15459), .A2(n7874), .ZN(n7872) );
  NAND2_X1 U8339 ( .A1(n15412), .A2(n15411), .ZN(n15436) );
  XNOR2_X1 U8340 ( .A(n15437), .B(n6876), .ZN(n15442) );
  NAND2_X1 U8341 ( .A1(n12675), .A2(n12674), .ZN(n12678) );
  NAND2_X1 U8342 ( .A1(n6968), .A2(n6969), .ZN(n6965) );
  NAND2_X1 U8343 ( .A1(n12691), .A2(n12668), .ZN(n6969) );
  OR2_X1 U8344 ( .A1(n12669), .A2(n12691), .ZN(n6968) );
  NAND2_X1 U8345 ( .A1(n10044), .A2(n12556), .ZN(n12382) );
  NAND2_X1 U8346 ( .A1(n12547), .A2(n12396), .ZN(n7831) );
  AOI21_X1 U8347 ( .B1(n14020), .B2(n12381), .A(n12403), .ZN(n12417) );
  INV_X1 U8348 ( .A(n12698), .ZN(n6962) );
  NAND2_X1 U8349 ( .A1(n6964), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U8350 ( .A1(n6963), .A2(n6962), .ZN(n6961) );
  NAND2_X1 U8351 ( .A1(n12696), .A2(n12695), .ZN(n6964) );
  INV_X1 U8352 ( .A(n12697), .ZN(n6963) );
  NOR2_X1 U8353 ( .A1(n12407), .A2(n6751), .ZN(n6750) );
  NAND2_X1 U8354 ( .A1(n6960), .A2(n12702), .ZN(n6958) );
  NAND2_X1 U8355 ( .A1(n12463), .A2(n6515), .ZN(n7832) );
  NAND2_X1 U8356 ( .A1(n6984), .A2(n6983), .ZN(n12714) );
  AOI21_X1 U8357 ( .B1(n6440), .B2(n6987), .A(n6557), .ZN(n6983) );
  NOR2_X1 U8358 ( .A1(n6986), .A2(n12707), .ZN(n6987) );
  NAND2_X1 U8359 ( .A1(n7826), .A2(n12483), .ZN(n7825) );
  NAND2_X1 U8360 ( .A1(n7830), .A2(n7827), .ZN(n7826) );
  NAND2_X1 U8361 ( .A1(n7829), .A2(n7828), .ZN(n7827) );
  INV_X1 U8362 ( .A(n12475), .ZN(n7828) );
  INV_X1 U8363 ( .A(n12476), .ZN(n7829) );
  OAI22_X1 U8364 ( .A1(n12721), .A2(n7903), .B1(n12722), .B2(n7902), .ZN(
        n12727) );
  INV_X1 U8365 ( .A(n12720), .ZN(n7902) );
  NOR2_X1 U8366 ( .A1(n12720), .A2(n12723), .ZN(n7903) );
  NAND2_X1 U8367 ( .A1(n7647), .A2(n6417), .ZN(n7646) );
  NAND2_X1 U8368 ( .A1(n10480), .A2(n6417), .ZN(n7643) );
  INV_X1 U8369 ( .A(n12493), .ZN(n6747) );
  NAND2_X1 U8370 ( .A1(n7836), .A2(n7837), .ZN(n7835) );
  INV_X1 U8371 ( .A(n10531), .ZN(n7670) );
  NAND2_X1 U8372 ( .A1(n10491), .A2(n11770), .ZN(n10505) );
  NAND2_X1 U8373 ( .A1(n7668), .A2(n10535), .ZN(n7667) );
  NAND2_X1 U8374 ( .A1(n7658), .A2(n13504), .ZN(n7668) );
  INV_X1 U8375 ( .A(n10534), .ZN(n7658) );
  OAI21_X1 U8376 ( .B1(n12498), .B2(n12497), .A(n12496), .ZN(n6748) );
  INV_X1 U8377 ( .A(n7817), .ZN(n7812) );
  NAND2_X1 U8378 ( .A1(n12503), .A2(n12502), .ZN(n7819) );
  INV_X1 U8379 ( .A(n12503), .ZN(n7820) );
  NAND2_X1 U8380 ( .A1(n7817), .A2(n6480), .ZN(n7815) );
  NAND2_X1 U8381 ( .A1(n12775), .A2(n12777), .ZN(n7899) );
  NOR2_X1 U8382 ( .A1(n7900), .A2(n7442), .ZN(n7441) );
  OAI21_X1 U8383 ( .B1(n7660), .B2(n7662), .A(n7659), .ZN(n10548) );
  AOI21_X1 U8384 ( .B1(n7661), .B2(n7663), .A(n6555), .ZN(n7659) );
  INV_X1 U8385 ( .A(n13442), .ZN(n7656) );
  INV_X1 U8386 ( .A(n10552), .ZN(n7657) );
  NAND2_X1 U8387 ( .A1(n12506), .A2(n12508), .ZN(n6758) );
  INV_X1 U8388 ( .A(n12784), .ZN(n6973) );
  NAND2_X1 U8389 ( .A1(n7433), .A2(n12784), .ZN(n6972) );
  NAND2_X1 U8390 ( .A1(n12655), .A2(n12821), .ZN(n6988) );
  OR2_X1 U8391 ( .A1(n12655), .A2(n8801), .ZN(n6989) );
  INV_X1 U8392 ( .A(n7343), .ZN(n7607) );
  NOR2_X1 U8393 ( .A1(n12515), .A2(n12516), .ZN(n6755) );
  NAND2_X1 U8394 ( .A1(n12515), .A2(n12516), .ZN(n6757) );
  NAND2_X1 U8395 ( .A1(n6971), .A2(n12784), .ZN(n12788) );
  NAND2_X1 U8396 ( .A1(n6974), .A2(n12785), .ZN(n6971) );
  NAND2_X1 U8397 ( .A1(n7438), .A2(n12796), .ZN(n7435) );
  INV_X1 U8398 ( .A(n8572), .ZN(n8121) );
  NOR2_X1 U8399 ( .A1(n8121), .A2(SI_18_), .ZN(n8120) );
  INV_X1 U8400 ( .A(n8100), .ZN(n7529) );
  INV_X1 U8401 ( .A(n8442), .ZN(n7997) );
  NAND2_X1 U8402 ( .A1(n7651), .A2(n7650), .ZN(n7649) );
  NOR2_X1 U8403 ( .A1(n10563), .A2(n10562), .ZN(n7650) );
  NAND2_X1 U8404 ( .A1(n7653), .A2(n7652), .ZN(n7651) );
  OR2_X1 U8405 ( .A1(n13106), .A2(n10564), .ZN(n7648) );
  NAND2_X1 U8406 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n7605), .ZN(n7604) );
  INV_X1 U8407 ( .A(n8037), .ZN(n7605) );
  NOR2_X1 U8408 ( .A1(n7607), .A2(n15815), .ZN(n7606) );
  NAND2_X1 U8409 ( .A1(n7607), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U8410 ( .A1(n11163), .A2(n10633), .ZN(n7594) );
  INV_X1 U8411 ( .A(n10170), .ZN(n7289) );
  AND2_X1 U8412 ( .A1(n6592), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U8413 ( .A1(n13399), .A2(n10151), .ZN(n6845) );
  INV_X1 U8414 ( .A(n10151), .ZN(n6846) );
  NAND2_X1 U8415 ( .A1(n6903), .A2(n12107), .ZN(n11972) );
  OR2_X1 U8416 ( .A1(n12107), .A2(n13121), .ZN(n10517) );
  NAND2_X1 U8417 ( .A1(n13126), .A2(n11299), .ZN(n10481) );
  INV_X1 U8418 ( .A(n9735), .ZN(n7937) );
  INV_X1 U8419 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9400) );
  INV_X1 U8420 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9403) );
  NOR2_X1 U8421 ( .A1(n7103), .A2(n6816), .ZN(n6815) );
  INV_X1 U8422 ( .A(n9518), .ZN(n6816) );
  INV_X1 U8423 ( .A(n9537), .ZN(n7103) );
  AND2_X1 U8424 ( .A1(n7467), .A2(n9572), .ZN(n7466) );
  NAND2_X1 U8425 ( .A1(n9556), .A2(n9558), .ZN(n7467) );
  NAND2_X1 U8426 ( .A1(n12569), .A2(n12568), .ZN(n7546) );
  NAND2_X1 U8427 ( .A1(n7791), .A2(n9979), .ZN(n7790) );
  INV_X1 U8428 ( .A(n9978), .ZN(n7791) );
  INV_X1 U8429 ( .A(n12590), .ZN(n8007) );
  NOR2_X1 U8430 ( .A1(n12614), .A2(n7784), .ZN(n7783) );
  AND2_X1 U8431 ( .A1(n7786), .A2(n9960), .ZN(n7784) );
  NAND2_X1 U8432 ( .A1(n7783), .A2(n7785), .ZN(n7781) );
  NAND2_X1 U8433 ( .A1(n12810), .A2(n12809), .ZN(n7448) );
  OAI21_X1 U8434 ( .B1(n12655), .B2(n12822), .A(n7901), .ZN(n12737) );
  NAND2_X1 U8435 ( .A1(n12655), .A2(n15526), .ZN(n7901) );
  INV_X1 U8436 ( .A(n10340), .ZN(n7408) );
  NOR2_X1 U8437 ( .A1(n8677), .A2(n8676), .ZN(n6924) );
  INV_X1 U8438 ( .A(n8616), .ZN(n8618) );
  INV_X1 U8439 ( .A(n6416), .ZN(n7121) );
  OAI21_X1 U8440 ( .B1(n10769), .B2(n10747), .A(n6930), .ZN(n8081) );
  NAND2_X1 U8441 ( .A1(n10769), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6930) );
  AND2_X1 U8442 ( .A1(n8302), .A2(n7000), .ZN(n8074) );
  INV_X1 U8443 ( .A(n8251), .ZN(n8073) );
  XNOR2_X1 U8444 ( .A(n11109), .B(n11509), .ZN(n9511) );
  XNOR2_X1 U8445 ( .A(n11519), .B(n11109), .ZN(n9531) );
  AOI21_X1 U8446 ( .B1(n13368), .B2(n10571), .A(n7314), .ZN(n7313) );
  NAND2_X1 U8447 ( .A1(n6437), .A2(n13141), .ZN(n7130) );
  NAND2_X1 U8448 ( .A1(n7143), .A2(n7142), .ZN(n7678) );
  AOI21_X1 U8449 ( .B1(n7145), .B2(n7141), .A(n7140), .ZN(n7139) );
  NAND2_X1 U8450 ( .A1(n7678), .A2(n10893), .ZN(n10694) );
  AOI21_X1 U8451 ( .B1(n6813), .B2(n10573), .A(n6812), .ZN(n6811) );
  INV_X1 U8452 ( .A(n10574), .ZN(n6812) );
  INV_X1 U8453 ( .A(n10572), .ZN(n6808) );
  NOR2_X1 U8454 ( .A1(n9845), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7303) );
  AND2_X1 U8455 ( .A1(n6586), .A2(n7508), .ZN(n7506) );
  INV_X1 U8456 ( .A(n7303), .ZN(n9856) );
  OR2_X1 U8457 ( .A1(n9827), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9845) );
  INV_X1 U8458 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7311) );
  INV_X1 U8459 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9741) );
  NOR2_X1 U8460 ( .A1(n9712), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9725) );
  INV_X1 U8461 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7306) );
  AND2_X1 U8462 ( .A1(n11488), .A2(n7308), .ZN(n7307) );
  INV_X1 U8463 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7308) );
  CLKBUF_X1 U8464 ( .A(n11882), .Z(n11884) );
  INV_X1 U8465 ( .A(n11616), .ZN(n10129) );
  INV_X1 U8466 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7301) );
  AND2_X1 U8467 ( .A1(n10470), .A2(n11436), .ZN(n10476) );
  NAND2_X1 U8468 ( .A1(n11448), .A2(n15784), .ZN(n10470) );
  NOR2_X1 U8469 ( .A1(n10124), .A2(n6831), .ZN(n6830) );
  AND2_X1 U8470 ( .A1(n10127), .A2(n11399), .ZN(n6834) );
  INV_X1 U8471 ( .A(n10187), .ZN(n7948) );
  AOI21_X1 U8472 ( .B1(n9438), .B2(P3_IR_REG_31__SCAN_IN), .A(n9419), .ZN(
        n9420) );
  INV_X1 U8473 ( .A(n10162), .ZN(n7470) );
  INV_X1 U8474 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9432) );
  NAND4_X1 U8475 ( .A1(n9448), .A2(n9407), .A3(n9408), .A4(n9406), .ZN(n9427)
         );
  INV_X1 U8476 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9407) );
  INV_X1 U8477 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U8478 ( .A1(n7451), .A2(n9852), .ZN(n7079) );
  NOR2_X1 U8479 ( .A1(n6618), .A2(n6822), .ZN(n6821) );
  INV_X1 U8480 ( .A(n9643), .ZN(n6822) );
  NAND2_X1 U8481 ( .A1(n6927), .A2(n9554), .ZN(n9590) );
  INV_X1 U8482 ( .A(n9574), .ZN(n6927) );
  INV_X1 U8483 ( .A(n7466), .ZN(n7464) );
  AND2_X1 U8484 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8995) );
  NAND2_X1 U8485 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  INV_X1 U8486 ( .A(n9139), .ZN(n9138) );
  NOR2_X1 U8487 ( .A1(n7074), .A2(n14122), .ZN(n7073) );
  AND2_X1 U8488 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8965) );
  AND2_X1 U8489 ( .A1(n12581), .A2(n12553), .ZN(n12624) );
  NOR2_X1 U8490 ( .A1(n13978), .A2(n13888), .ZN(n7076) );
  AOI21_X1 U8491 ( .B1(n7805), .B2(n7808), .A(n6547), .ZN(n7804) );
  NAND2_X1 U8492 ( .A1(n7805), .A2(n7386), .ZN(n7385) );
  NOR2_X1 U8493 ( .A1(n13951), .A2(n9230), .ZN(n7075) );
  INV_X1 U8494 ( .A(n9231), .ZN(n9221) );
  INV_X1 U8495 ( .A(n9969), .ZN(n7394) );
  INV_X1 U8496 ( .A(n9962), .ZN(n7163) );
  NAND2_X1 U8497 ( .A1(n9138), .A2(n7073), .ZN(n9158) );
  NAND2_X1 U8498 ( .A1(n9138), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9148) );
  INV_X1 U8499 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n13603) );
  OR2_X1 U8500 ( .A1(n9121), .A2(n13603), .ZN(n9139) );
  INV_X1 U8501 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9069) );
  OR2_X1 U8502 ( .A1(n9070), .A2(n9069), .ZN(n9090) );
  NAND2_X1 U8503 ( .A1(n9053), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9070) );
  INV_X1 U8504 ( .A(n9054), .ZN(n9053) );
  INV_X1 U8505 ( .A(n10014), .ZN(n8034) );
  NAND3_X1 U8506 ( .A1(n8996), .A2(P2_REG3_REG_9__SCAN_IN), .A3(n6431), .ZN(
        n9054) );
  NAND2_X1 U8507 ( .A1(n8996), .A2(n6431), .ZN(n9038) );
  NOR2_X1 U8508 ( .A1(n12599), .A2(n8032), .ZN(n8031) );
  INV_X1 U8509 ( .A(n10011), .ZN(n8032) );
  AND2_X1 U8510 ( .A1(n6493), .A2(n10011), .ZN(n8030) );
  INV_X1 U8511 ( .A(n9935), .ZN(n7803) );
  AND2_X1 U8512 ( .A1(n11054), .A2(n11086), .ZN(n7189) );
  NAND2_X1 U8513 ( .A1(n8940), .A2(n7190), .ZN(n7191) );
  AND2_X1 U8514 ( .A1(n10769), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7190) );
  AND2_X1 U8515 ( .A1(n6424), .A2(n14308), .ZN(n7889) );
  INV_X1 U8516 ( .A(n14546), .ZN(n14364) );
  NAND2_X1 U8517 ( .A1(n12153), .A2(n12248), .ZN(n12337) );
  OR2_X1 U8518 ( .A1(n9010), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9028) );
  INV_X1 U8519 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n13592) );
  AND2_X1 U8520 ( .A1(n8912), .A2(n8929), .ZN(n8943) );
  NOR2_X1 U8521 ( .A1(n8473), .A2(n8472), .ZN(n8471) );
  INV_X1 U8522 ( .A(n8714), .ZN(n7973) );
  INV_X1 U8523 ( .A(n14682), .ZN(n7982) );
  NAND2_X1 U8524 ( .A1(n7378), .A2(n7984), .ZN(n7377) );
  NOR2_X1 U8525 ( .A1(n8636), .A2(n6649), .ZN(n6678) );
  NAND2_X1 U8526 ( .A1(n11372), .A2(n6648), .ZN(n7378) );
  AND2_X1 U8527 ( .A1(n8471), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8485) );
  OAI22_X1 U8528 ( .A1(n8213), .A2(n8227), .B1(n6892), .B2(n6891), .ZN(n6890)
         );
  NAND2_X1 U8529 ( .A1(n6924), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U8530 ( .A1(n6678), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U8531 ( .A1(n15001), .A2(n15005), .ZN(n6699) );
  INV_X1 U8532 ( .A(n10381), .ZN(n7258) );
  NAND2_X1 U8533 ( .A1(n12835), .A2(n10362), .ZN(n7478) );
  INV_X1 U8534 ( .A(n10362), .ZN(n7479) );
  NAND2_X1 U8535 ( .A1(n10363), .A2(n7011), .ZN(n7855) );
  INV_X1 U8536 ( .A(n10363), .ZN(n7856) );
  INV_X1 U8537 ( .A(n8323), .ZN(n6674) );
  INV_X1 U8538 ( .A(n10306), .ZN(n7951) );
  NOR2_X1 U8539 ( .A1(n15495), .A2(n12700), .ZN(n7630) );
  NAND2_X1 U8540 ( .A1(n11960), .A2(n11961), .ZN(n10304) );
  NAND2_X1 U8541 ( .A1(n11205), .A2(n10091), .ZN(n7263) );
  NAND2_X1 U8542 ( .A1(n13695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7848) );
  INV_X1 U8543 ( .A(n7844), .ZN(n7843) );
  OAI21_X1 U8544 ( .B1(n7846), .B2(P1_IR_REG_30__SCAN_IN), .A(n7845), .ZN(
        n7844) );
  NAND2_X1 U8545 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7845) );
  NOR2_X1 U8546 ( .A1(n8169), .A2(n15296), .ZN(n7846) );
  INV_X1 U8547 ( .A(n8761), .ZN(n7538) );
  AOI21_X1 U8548 ( .B1(n7537), .B2(n8758), .A(n7535), .ZN(n7534) );
  INV_X1 U8549 ( .A(n9981), .ZN(n7535) );
  INV_X1 U8550 ( .A(n7515), .ZN(n7514) );
  AOI21_X1 U8551 ( .B1(n8692), .B2(n7515), .A(n7513), .ZN(n7512) );
  NOR2_X1 U8552 ( .A1(n8716), .A2(n6627), .ZN(n7515) );
  NAND2_X1 U8553 ( .A1(n8693), .A2(n7116), .ZN(n7115) );
  INV_X1 U8554 ( .A(n8001), .ZN(n7116) );
  INV_X1 U8555 ( .A(n6621), .ZN(n7118) );
  NAND2_X1 U8556 ( .A1(n6692), .A2(n8672), .ZN(n7119) );
  INV_X1 U8557 ( .A(n8651), .ZN(n6692) );
  NAND2_X1 U8558 ( .A1(n6686), .A2(n8634), .ZN(n8650) );
  OAI21_X1 U8559 ( .B1(n8593), .B2(n7519), .A(n7517), .ZN(n6686) );
  AOI21_X1 U8560 ( .B1(n7518), .B2(n7520), .A(n8631), .ZN(n7517) );
  NOR2_X1 U8561 ( .A1(n8110), .A2(n8503), .ZN(n8521) );
  NOR2_X1 U8562 ( .A1(n8501), .A2(SI_14_), .ZN(n8522) );
  NAND2_X1 U8563 ( .A1(n8106), .A2(n13693), .ZN(n8523) );
  NAND2_X1 U8564 ( .A1(n6798), .A2(n8500), .ZN(n8502) );
  OAI21_X1 U8565 ( .B1(n8090), .B2(n8000), .A(n8092), .ZN(n7999) );
  INV_X1 U8566 ( .A(n8090), .ZN(n6855) );
  INV_X1 U8567 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U8568 ( .A1(n7380), .A2(n8085), .ZN(n8384) );
  OR2_X1 U8569 ( .A1(n8351), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U8570 ( .A(n8081), .B(SI_6_), .ZN(n8353) );
  NAND2_X1 U8571 ( .A1(n15390), .A2(n15389), .ZN(n15329) );
  NAND2_X1 U8572 ( .A1(n7372), .A2(n7370), .ZN(n15334) );
  NAND2_X1 U8573 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n7371), .ZN(n7370) );
  NAND2_X1 U8574 ( .A1(n15396), .A2(n15395), .ZN(n7372) );
  INV_X1 U8575 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7371) );
  INV_X1 U8576 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U8577 ( .A1(n15348), .A2(n15347), .ZN(n15349) );
  OR2_X1 U8578 ( .A1(n9682), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9712) );
  INV_X1 U8579 ( .A(n9551), .ZN(n7773) );
  AND2_X1 U8580 ( .A1(n9813), .A2(n9796), .ZN(n7775) );
  INV_X1 U8581 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12986) );
  OR2_X1 U8582 ( .A1(n9877), .A2(n9876), .ZN(n12885) );
  INV_X1 U8583 ( .A(n15795), .ZN(n11110) );
  AND2_X1 U8584 ( .A1(n9787), .A2(n13036), .ZN(n9802) );
  AND2_X1 U8585 ( .A1(n9725), .A2(n7309), .ZN(n9787) );
  AND2_X1 U8586 ( .A1(n6622), .A2(n7310), .ZN(n7309) );
  INV_X1 U8587 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7310) );
  INV_X1 U8588 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U8589 ( .A1(n9680), .A2(n9679), .ZN(n9682) );
  AND2_X1 U8590 ( .A1(n9600), .A2(n7304), .ZN(n9680) );
  AND2_X1 U8591 ( .A1(n6492), .A2(n7305), .ZN(n7304) );
  INV_X1 U8592 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U8593 ( .A1(n6922), .A2(n9637), .ZN(n13061) );
  NAND2_X1 U8594 ( .A1(n12996), .A2(n6918), .ZN(n7769) );
  OR2_X1 U8595 ( .A1(n9561), .A2(n12921), .ZN(n10420) );
  AND4_X1 U8596 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10200) );
  NAND2_X1 U8597 ( .A1(n10416), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U8598 ( .A1(n10986), .A2(n10628), .ZN(n11009) );
  NAND2_X1 U8599 ( .A1(n6996), .A2(n6995), .ZN(n11006) );
  INV_X1 U8600 ( .A(n11009), .ZN(n6995) );
  INV_X1 U8601 ( .A(n11008), .ZN(n6996) );
  NAND2_X1 U8602 ( .A1(n7599), .A2(n11026), .ZN(n11164) );
  OR2_X1 U8603 ( .A1(n11028), .A2(n11027), .ZN(n7599) );
  NAND2_X1 U8604 ( .A1(n11028), .A2(n6641), .ZN(n7598) );
  AND2_X1 U8605 ( .A1(n7592), .A2(n7591), .ZN(n13130) );
  NAND2_X1 U8606 ( .A1(n7593), .A2(n11343), .ZN(n7592) );
  NAND2_X1 U8607 ( .A1(n7573), .A2(n7567), .ZN(n7566) );
  AND2_X1 U8608 ( .A1(n13155), .A2(n10688), .ZN(n7567) );
  NOR2_X1 U8609 ( .A1(n7707), .A2(n11859), .ZN(n11493) );
  NAND2_X1 U8610 ( .A1(n7697), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7705) );
  INV_X1 U8611 ( .A(n7707), .ZN(n7697) );
  INV_X1 U8612 ( .A(n11859), .ZN(n7704) );
  NAND2_X1 U8613 ( .A1(n7696), .A2(n7694), .ZN(n10691) );
  INV_X1 U8614 ( .A(n7695), .ZN(n7694) );
  OAI21_X1 U8615 ( .B1(n10689), .B2(n7701), .A(n7698), .ZN(n7695) );
  AOI21_X1 U8616 ( .B1(n7615), .B2(n7621), .A(n6575), .ZN(n7613) );
  OAI21_X1 U8617 ( .B1(n7678), .B2(n10893), .A(n10694), .ZN(n13205) );
  AND2_X1 U8618 ( .A1(n13232), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7581) );
  INV_X1 U8619 ( .A(n10611), .ZN(n13231) );
  NOR2_X1 U8620 ( .A1(n13245), .A2(n6528), .ZN(n13263) );
  OR2_X1 U8621 ( .A1(n13263), .A2(n13262), .ZN(n7590) );
  AND2_X1 U8622 ( .A1(n7135), .A2(n10707), .ZN(n13280) );
  AND2_X1 U8623 ( .A1(n10701), .A2(n10976), .ZN(n7136) );
  AND2_X1 U8624 ( .A1(n7590), .A2(n7589), .ZN(n13284) );
  NAND2_X1 U8625 ( .A1(n10669), .A2(n13266), .ZN(n7589) );
  NOR2_X1 U8626 ( .A1(n13284), .A2(n13283), .ZN(n13281) );
  INV_X1 U8627 ( .A(n7559), .ZN(n7558) );
  OAI21_X1 U8628 ( .B1(n7552), .B2(n13299), .A(n7550), .ZN(n7555) );
  AND2_X1 U8629 ( .A1(n13307), .A2(n7551), .ZN(n7550) );
  OR2_X1 U8630 ( .A1(n7562), .A2(n13299), .ZN(n7551) );
  NOR2_X1 U8631 ( .A1(n6470), .A2(n7561), .ZN(n7556) );
  NAND2_X1 U8632 ( .A1(n10615), .A2(n10976), .ZN(n7202) );
  AND2_X1 U8633 ( .A1(n12921), .A2(n10194), .ZN(n13341) );
  OAI21_X1 U8634 ( .B1(n13376), .B2(n6810), .A(n6807), .ZN(n13357) );
  AOI21_X1 U8635 ( .B1(n6811), .B2(n6809), .A(n6808), .ZN(n6807) );
  INV_X1 U8636 ( .A(n6811), .ZN(n6810) );
  INV_X1 U8637 ( .A(n10573), .ZN(n6809) );
  NAND2_X1 U8638 ( .A1(n6923), .A2(n6423), .ZN(n13355) );
  INV_X1 U8639 ( .A(n13357), .ZN(n6923) );
  NOR2_X1 U8640 ( .A1(n9923), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n10166) );
  AND2_X1 U8641 ( .A1(n9809), .A2(n9808), .ZN(n13418) );
  AOI21_X1 U8642 ( .B1(n7923), .B2(n7921), .A(n6549), .ZN(n7920) );
  INV_X1 U8643 ( .A(n10540), .ZN(n7921) );
  INV_X1 U8644 ( .A(n7923), .ZN(n7922) );
  NAND2_X1 U8645 ( .A1(n13464), .A2(n10146), .ZN(n13455) );
  NAND2_X1 U8646 ( .A1(n9725), .A2(n7312), .ZN(n9759) );
  NAND2_X1 U8647 ( .A1(n9725), .A2(n6622), .ZN(n9771) );
  AOI21_X1 U8648 ( .B1(n6899), .B2(n6901), .A(n10537), .ZN(n6897) );
  NAND2_X1 U8649 ( .A1(n13518), .A2(n13519), .ZN(n10143) );
  AOI21_X1 U8650 ( .B1(n7939), .B2(n12091), .A(n7938), .ZN(n7108) );
  INV_X1 U8651 ( .A(n10522), .ZN(n7938) );
  INV_X1 U8652 ( .A(n6851), .ZN(n6850) );
  OAI21_X1 U8653 ( .B1(n7344), .B2(n7285), .A(n10140), .ZN(n6851) );
  NAND2_X1 U8654 ( .A1(n9600), .A2(n6492), .ZN(n9647) );
  NAND2_X1 U8655 ( .A1(n9600), .A2(n7307), .ZN(n9631) );
  OR2_X1 U8656 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  NAND2_X1 U8657 ( .A1(n6894), .A2(n11770), .ZN(n10233) );
  INV_X1 U8658 ( .A(n10231), .ZN(n6894) );
  AND2_X1 U8659 ( .A1(n9599), .A2(n11747), .ZN(n9600) );
  INV_X1 U8660 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U8661 ( .A1(n9600), .A2(n11488), .ZN(n9614) );
  AND3_X1 U8662 ( .A1(n7301), .A2(n9525), .A3(n7299), .ZN(n9599) );
  AND2_X1 U8663 ( .A1(n9524), .A2(n7300), .ZN(n7299) );
  INV_X1 U8664 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U8665 ( .A1(n7914), .A2(n10496), .ZN(n11878) );
  NOR2_X1 U8666 ( .A1(n11602), .A2(n7916), .ZN(n7915) );
  INV_X1 U8667 ( .A(n10493), .ZN(n7916) );
  AND2_X1 U8668 ( .A1(n10227), .A2(n10493), .ZN(n11616) );
  CLKBUF_X1 U8669 ( .A(n11615), .Z(n7366) );
  NOR2_X1 U8670 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9525) );
  NAND2_X1 U8671 ( .A1(n11611), .A2(n10488), .ZN(n11399) );
  AND2_X1 U8672 ( .A1(n10263), .A2(n15836), .ZN(n11316) );
  INV_X1 U8673 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n13720) );
  OR2_X1 U8674 ( .A1(n11314), .A2(n10247), .ZN(n11311) );
  AND2_X1 U8675 ( .A1(n10253), .A2(n10252), .ZN(n11312) );
  INV_X1 U8676 ( .A(n15851), .ZN(n13745) );
  NAND2_X1 U8677 ( .A1(n11977), .A2(n6624), .ZN(n11978) );
  INV_X1 U8678 ( .A(n15806), .ZN(n15836) );
  AND2_X1 U8679 ( .A1(n13816), .A2(n10599), .ZN(n10263) );
  OR2_X1 U8680 ( .A1(n10253), .A2(n9900), .ZN(n10260) );
  NAND2_X1 U8681 ( .A1(n10243), .A2(n11660), .ZN(n15806) );
  NAND2_X1 U8682 ( .A1(n9880), .A2(n9879), .ZN(n11315) );
  AND2_X1 U8683 ( .A1(n7752), .A2(n7926), .ZN(n6852) );
  AND2_X1 U8684 ( .A1(n9418), .A2(n9412), .ZN(n7926) );
  INV_X1 U8685 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9418) );
  INV_X1 U8686 ( .A(n9417), .ZN(n7343) );
  OR2_X1 U8687 ( .A1(n9420), .A2(n8037), .ZN(n7609) );
  OR2_X1 U8688 ( .A1(n10155), .A2(n12231), .ZN(n10156) );
  AOI21_X1 U8689 ( .B1(n7088), .B2(n7089), .A(n6631), .ZN(n7085) );
  INV_X1 U8690 ( .A(n7088), .ZN(n7086) );
  INV_X1 U8691 ( .A(n6823), .ZN(n9701) );
  AOI21_X1 U8692 ( .B1(n9659), .B2(n9658), .A(n6618), .ZN(n6823) );
  NAND2_X1 U8693 ( .A1(n7449), .A2(n9643), .ZN(n9659) );
  XNOR2_X1 U8694 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .ZN(n9641) );
  AOI21_X1 U8695 ( .B1(n7930), .B2(n7932), .A(n6569), .ZN(n7928) );
  XNOR2_X1 U8696 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .ZN(n9624) );
  NAND2_X1 U8697 ( .A1(n6817), .A2(n9518), .ZN(n9536) );
  INV_X1 U8698 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9520) );
  OAI21_X1 U8699 ( .B1(n7913), .B2(n7912), .A(n7910), .ZN(n9517) );
  AOI21_X1 U8700 ( .B1(n7911), .B2(n9498), .A(n6564), .ZN(n7910) );
  INV_X1 U8701 ( .A(n9474), .ZN(n7911) );
  XNOR2_X1 U8702 ( .A(n13590), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n9481) );
  XNOR2_X1 U8703 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n9469) );
  NAND2_X1 U8704 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7564) );
  AND2_X1 U8705 ( .A1(n9421), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U8706 ( .A1(n8996), .A2(n8995), .ZN(n9016) );
  NAND2_X1 U8707 ( .A1(n9128), .A2(n9127), .ZN(n13840) );
  OR2_X1 U8708 ( .A1(n9250), .A2(n13927), .ZN(n9276) );
  NAND2_X1 U8709 ( .A1(n7741), .A2(n7743), .ZN(n7737) );
  INV_X1 U8710 ( .A(n7740), .ZN(n7739) );
  NOR2_X1 U8711 ( .A1(n12290), .A2(n7277), .ZN(n7276) );
  INV_X1 U8712 ( .A(n9064), .ZN(n7277) );
  INV_X1 U8713 ( .A(n9081), .ZN(n6777) );
  NAND2_X1 U8714 ( .A1(n11893), .A2(n6521), .ZN(n7278) );
  INV_X1 U8715 ( .A(n9049), .ZN(n7279) );
  NAND2_X1 U8716 ( .A1(n8965), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8999) );
  INV_X1 U8717 ( .A(n13977), .ZN(n7274) );
  INV_X1 U8718 ( .A(n13976), .ZN(n7275) );
  NAND2_X1 U8719 ( .A1(n13840), .A2(n9131), .ZN(n13897) );
  NAND2_X1 U8720 ( .A1(n12523), .A2(n6457), .ZN(n6736) );
  NOR2_X1 U8721 ( .A1(n12579), .A2(n7822), .ZN(n7821) );
  AND2_X1 U8722 ( .A1(n12580), .A2(n6602), .ZN(n7822) );
  NAND2_X1 U8723 ( .A1(n9991), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U8724 ( .A1(n9991), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U8725 ( .A1(n6717), .A2(n11067), .ZN(n6716) );
  NAND2_X1 U8726 ( .A1(n6718), .A2(n11067), .ZN(n6715) );
  OR2_X1 U8727 ( .A1(n11266), .A2(n11265), .ZN(n11263) );
  OR2_X1 U8728 ( .A1(n14101), .A2(n14100), .ZN(n14103) );
  XNOR2_X1 U8729 ( .A(n11792), .B(n11806), .ZN(n14108) );
  NOR2_X1 U8730 ( .A1(n14169), .A2(n7893), .ZN(n7891) );
  OR2_X1 U8731 ( .A1(n12621), .A2(n14302), .ZN(n7388) );
  NAND2_X1 U8732 ( .A1(n8057), .A2(n9999), .ZN(n7362) );
  NOR2_X1 U8733 ( .A1(n9323), .A2(n9389), .ZN(n10049) );
  AND2_X1 U8734 ( .A1(n9308), .A2(n9323), .ZN(n14188) );
  NAND2_X1 U8735 ( .A1(n7193), .A2(n7194), .ZN(n14202) );
  NAND2_X1 U8736 ( .A1(n9275), .A2(n7076), .ZN(n9307) );
  NAND2_X1 U8737 ( .A1(n14288), .A2(n7883), .ZN(n14214) );
  INV_X1 U8738 ( .A(n14261), .ZN(n9973) );
  INV_X1 U8739 ( .A(n7805), .ZN(n7387) );
  AND2_X1 U8740 ( .A1(n14288), .A2(n6445), .ZN(n14229) );
  INV_X1 U8741 ( .A(n9975), .ZN(n7808) );
  NAND2_X1 U8742 ( .A1(n14288), .A2(n14533), .ZN(n14272) );
  NAND2_X1 U8743 ( .A1(n9221), .A2(n7075), .ZN(n9239) );
  OR2_X1 U8744 ( .A1(n14267), .A2(n14266), .ZN(n14269) );
  NAND2_X1 U8745 ( .A1(n9178), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9209) );
  INV_X1 U8746 ( .A(n9180), .ZN(n9178) );
  AND2_X1 U8747 ( .A1(n9216), .A2(n9215), .ZN(n14315) );
  NAND2_X1 U8748 ( .A1(n14363), .A2(n6424), .ZN(n14319) );
  NAND2_X1 U8749 ( .A1(n14363), .A2(n14347), .ZN(n14341) );
  AND2_X1 U8750 ( .A1(n12593), .A2(n12592), .ZN(n14353) );
  NAND2_X1 U8751 ( .A1(n7164), .A2(n9962), .ZN(n14356) );
  NAND2_X1 U8752 ( .A1(n14373), .A2(n14389), .ZN(n7164) );
  OR2_X1 U8753 ( .A1(n9104), .A2(n14097), .ZN(n9121) );
  NAND2_X1 U8754 ( .A1(n9955), .A2(n9954), .ZN(n11930) );
  AND2_X1 U8755 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  NAND2_X1 U8756 ( .A1(n11926), .A2(n7400), .ZN(n9952) );
  NAND2_X1 U8757 ( .A1(n11763), .A2(n7886), .ZN(n12125) );
  NAND2_X1 U8758 ( .A1(n11763), .A2(n12120), .ZN(n12127) );
  NAND2_X1 U8759 ( .A1(n6763), .A2(n9942), .ZN(n11733) );
  OAI21_X1 U8760 ( .B1(n11475), .B2(n6762), .A(n6562), .ZN(n6763) );
  INV_X1 U8761 ( .A(n9940), .ZN(n6762) );
  NAND2_X1 U8762 ( .A1(n11643), .A2(n6425), .ZN(n11627) );
  NAND2_X1 U8763 ( .A1(n6759), .A2(n9937), .ZN(n11631) );
  NAND2_X1 U8764 ( .A1(n10045), .A2(n14022), .ZN(n9936) );
  NAND2_X1 U8765 ( .A1(n11034), .A2(n9935), .ZN(n11647) );
  INV_X1 U8766 ( .A(n14273), .ZN(n14380) );
  NAND2_X1 U8767 ( .A1(n11643), .A2(n10045), .ZN(n11644) );
  AND2_X1 U8768 ( .A1(n14422), .A2(n14421), .ZN(n7185) );
  NAND2_X1 U8769 ( .A1(n6760), .A2(n9940), .ZN(n11535) );
  NAND2_X1 U8770 ( .A1(n11475), .A2(n12599), .ZN(n6760) );
  AND2_X1 U8771 ( .A1(n10596), .A2(n11050), .ZN(n9386) );
  AND2_X1 U8772 ( .A1(n9341), .A2(n9340), .ZN(n9363) );
  INV_X1 U8773 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n13610) );
  INV_X1 U8774 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9132) );
  INV_X1 U8775 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8836) );
  OR2_X1 U8776 ( .A1(n9028), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9030) );
  OR2_X1 U8777 ( .A1(n8960), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U8778 ( .A1(n8080), .A2(n8070), .ZN(n8901) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U8780 ( .A1(n6673), .A2(n6539), .ZN(n8450) );
  OR2_X1 U8781 ( .A1(n8450), .A2(n13649), .ZN(n8473) );
  INV_X1 U8782 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13649) );
  NAND2_X1 U8783 ( .A1(n7976), .A2(n6806), .ZN(n14637) );
  AOI21_X1 U8784 ( .B1(n7977), .B2(n8498), .A(n6580), .ZN(n7976) );
  NAND2_X1 U8785 ( .A1(n8313), .A2(n8318), .ZN(n11371) );
  OR2_X1 U8786 ( .A1(n8391), .A2(n8390), .ZN(n8408) );
  OR2_X1 U8787 ( .A1(n8600), .A2(n8164), .ZN(n8636) );
  NAND2_X1 U8788 ( .A1(n6792), .A2(n6791), .ZN(n14662) );
  AOI21_X1 U8789 ( .B1(n6793), .B2(n7231), .A(n7986), .ZN(n6791) );
  NAND2_X1 U8790 ( .A1(n14672), .A2(n6793), .ZN(n6792) );
  OR2_X1 U8791 ( .A1(n8441), .A2(n7213), .ZN(n7211) );
  NAND2_X1 U8792 ( .A1(n8553), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U8793 ( .A1(n14672), .A2(n14673), .ZN(n14671) );
  NAND2_X1 U8794 ( .A1(n14580), .A2(n8499), .ZN(n14627) );
  AND2_X1 U8795 ( .A1(n6693), .A2(n6609), .ZN(n12875) );
  NAND2_X1 U8796 ( .A1(n12813), .A2(n12812), .ZN(n7443) );
  NOR4_X1 U8797 ( .A1(n12855), .A2(n14868), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  AND2_X1 U8798 ( .A1(n8810), .A2(n8809), .ZN(n12653) );
  AND3_X1 U8799 ( .A1(n8539), .A2(n8538), .A3(n8537), .ZN(n14707) );
  AND4_X1 U8800 ( .A1(n8516), .A2(n8515), .A3(n8514), .A4(n8513), .ZN(n14586)
         );
  AND4_X1 U8801 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n10323)
         );
  AND4_X1 U8802 ( .A1(n8478), .A2(n8477), .A3(n8476), .A4(n8475), .ZN(n14584)
         );
  AND4_X1 U8803 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n12699)
         );
  NAND2_X1 U8804 ( .A1(n11181), .A2(n8253), .ZN(n8281) );
  NAND2_X1 U8805 ( .A1(n11187), .A2(n11188), .ZN(n11186) );
  NAND2_X1 U8806 ( .A1(n7049), .A2(n10900), .ZN(n10917) );
  OR2_X1 U8807 ( .A1(n10935), .A2(n10901), .ZN(n7049) );
  NAND2_X1 U8808 ( .A1(n10923), .A2(n10922), .ZN(n10945) );
  NAND2_X1 U8809 ( .A1(n7048), .A2(n7050), .ZN(n7047) );
  NAND2_X1 U8810 ( .A1(n7040), .A2(n10916), .ZN(n7048) );
  NAND2_X1 U8811 ( .A1(n10900), .A2(n10901), .ZN(n7040) );
  NAND2_X1 U8812 ( .A1(n10963), .A2(n10962), .ZN(n7418) );
  NAND2_X1 U8813 ( .A1(n10950), .A2(n10959), .ZN(n7044) );
  AND2_X1 U8814 ( .A1(n7050), .A2(n10900), .ZN(n7046) );
  OR2_X1 U8815 ( .A1(n14789), .A2(n7039), .ZN(n7038) );
  NOR2_X1 U8816 ( .A1(n12078), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7039) );
  NAND2_X1 U8817 ( .A1(n7430), .A2(n7429), .ZN(n7428) );
  NAND2_X1 U8818 ( .A1(n7428), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7427) );
  AND2_X1 U8819 ( .A1(n14798), .A2(n14809), .ZN(n14807) );
  NAND2_X1 U8820 ( .A1(n14795), .A2(n6645), .ZN(n14810) );
  AND2_X1 U8821 ( .A1(n10067), .A2(n10066), .ZN(n15131) );
  XNOR2_X1 U8822 ( .A(n14844), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14858) );
  NAND2_X1 U8823 ( .A1(n7175), .A2(n15604), .ZN(n7174) );
  NOR2_X1 U8824 ( .A1(n10393), .A2(n10345), .ZN(n7175) );
  NOR2_X1 U8825 ( .A1(n7954), .A2(n7404), .ZN(n7401) );
  NAND2_X1 U8826 ( .A1(n10393), .A2(n7955), .ZN(n7954) );
  NAND2_X1 U8827 ( .A1(n10393), .A2(n10345), .ZN(n7953) );
  OAI21_X1 U8828 ( .B1(n7174), .B2(n7955), .A(n10348), .ZN(n7172) );
  NAND2_X1 U8829 ( .A1(n8744), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n14844) );
  INV_X1 U8830 ( .A(n8746), .ZN(n8744) );
  INV_X1 U8831 ( .A(n7488), .ZN(n7487) );
  INV_X1 U8832 ( .A(n14706), .ZN(n14697) );
  INV_X1 U8833 ( .A(n7180), .ZN(n6889) );
  NAND2_X1 U8834 ( .A1(n7180), .A2(n14934), .ZN(n6888) );
  NAND2_X1 U8835 ( .A1(n7853), .A2(n7849), .ZN(n14899) );
  NAND2_X1 U8836 ( .A1(n8675), .A2(n8674), .ZN(n14921) );
  NAND2_X1 U8837 ( .A1(n14936), .A2(n14944), .ZN(n14937) );
  NAND2_X1 U8838 ( .A1(n14970), .A2(n10334), .ZN(n14949) );
  AOI21_X1 U8839 ( .B1(n7267), .B2(n7268), .A(n6546), .ZN(n7265) );
  NAND2_X1 U8840 ( .A1(n7634), .A2(n15271), .ZN(n7633) );
  INV_X1 U8841 ( .A(n7634), .ZN(n7632) );
  NOR3_X1 U8842 ( .A1(n15058), .A2(n15188), .A3(n15045), .ZN(n15027) );
  INV_X1 U8843 ( .A(n10325), .ZN(n15003) );
  NOR2_X1 U8844 ( .A1(n15058), .A2(n15045), .ZN(n15044) );
  INV_X1 U8845 ( .A(n15002), .ZN(n15074) );
  INV_X1 U8846 ( .A(n10369), .ZN(n10370) );
  INV_X1 U8847 ( .A(n7486), .ZN(n7484) );
  NAND2_X1 U8848 ( .A1(n15085), .A2(n15099), .ZN(n15089) );
  NAND2_X1 U8849 ( .A1(n12344), .A2(n10322), .ZN(n15085) );
  INV_X1 U8850 ( .A(n12181), .ZN(n12839) );
  AND2_X1 U8851 ( .A1(n12168), .A2(n7637), .ZN(n12314) );
  NAND2_X1 U8852 ( .A1(n12168), .A2(n10064), .ZN(n12272) );
  NAND2_X1 U8853 ( .A1(n6673), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U8854 ( .A1(n12173), .A2(n12837), .ZN(n12178) );
  NAND2_X1 U8855 ( .A1(n7477), .A2(n10362), .ZN(n12173) );
  NAND2_X1 U8856 ( .A1(n11719), .A2(n11718), .ZN(n7477) );
  AND2_X1 U8857 ( .A1(n7627), .A2(n7630), .ZN(n11939) );
  NOR2_X1 U8858 ( .A1(n15498), .A2(n15597), .ZN(n7627) );
  INV_X1 U8859 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8368) );
  OR2_X1 U8860 ( .A1(n8369), .A2(n8368), .ZN(n8391) );
  NAND2_X1 U8861 ( .A1(n6675), .A2(n6674), .ZN(n8369) );
  NOR2_X1 U8862 ( .A1(n6677), .A2(n6676), .ZN(n6675) );
  NAND2_X1 U8863 ( .A1(n6674), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8345) );
  XNOR2_X1 U8864 ( .A(n14743), .B(n15495), .ZN(n15488) );
  NAND2_X1 U8865 ( .A1(n7629), .A2(n15580), .ZN(n15499) );
  NAND2_X1 U8866 ( .A1(n15506), .A2(n12831), .ZN(n7473) );
  NAND2_X1 U8867 ( .A1(n10304), .A2(n12828), .ZN(n7178) );
  NOR2_X1 U8868 ( .A1(n15518), .A2(n15564), .ZN(n15516) );
  NAND2_X1 U8869 ( .A1(n15549), .A2(n15525), .ZN(n15107) );
  NAND2_X1 U8870 ( .A1(n7626), .A2(n11204), .ZN(n15518) );
  INV_X1 U8871 ( .A(n15107), .ZN(n7626) );
  INV_X1 U8872 ( .A(n11824), .ZN(n12829) );
  OR2_X1 U8873 ( .A1(n12815), .A2(n10881), .ZN(n14706) );
  NOR2_X1 U8874 ( .A1(n12163), .A2(n8059), .ZN(n12180) );
  AND3_X1 U8875 ( .A1(n10110), .A2(n10109), .A3(n10108), .ZN(n10115) );
  INV_X1 U8876 ( .A(n15572), .ZN(n15601) );
  INV_X1 U8877 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8794) );
  OAI21_X1 U8878 ( .B1(n8793), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8795) );
  INV_X1 U8879 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8136) );
  INV_X1 U8880 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8135) );
  XNOR2_X1 U8881 ( .A(n10075), .B(n10074), .ZN(n12910) );
  XNOR2_X1 U8882 ( .A(n10069), .B(n10068), .ZN(n12928) );
  NAND2_X1 U8883 ( .A1(n7530), .A2(n7534), .ZN(n10069) );
  NAND2_X1 U8884 ( .A1(n8759), .A2(n7537), .ZN(n7530) );
  XNOR2_X1 U8885 ( .A(n9983), .B(n9982), .ZN(n12945) );
  OAI21_X1 U8886 ( .B1(n8759), .B2(n8758), .A(n8761), .ZN(n9983) );
  XNOR2_X1 U8887 ( .A(n8759), .B(n8741), .ZN(n12941) );
  NAND2_X1 U8888 ( .A1(n7522), .A2(n8125), .ZN(n8617) );
  NAND2_X1 U8889 ( .A1(n7524), .A2(n7523), .ZN(n7522) );
  NAND2_X1 U8890 ( .A1(n8186), .A2(n8185), .ZN(n8575) );
  INV_X1 U8891 ( .A(n8549), .ZN(n8186) );
  XNOR2_X1 U8892 ( .A(n8574), .B(n8573), .ZN(n11309) );
  AND2_X1 U8893 ( .A1(n8571), .A2(n8570), .ZN(n8574) );
  NAND2_X1 U8894 ( .A1(n8569), .A2(n8546), .ZN(n6703) );
  XNOR2_X1 U8895 ( .A(n8483), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12076) );
  AND2_X1 U8896 ( .A1(n8405), .A2(n8425), .ZN(n10949) );
  NAND2_X1 U8897 ( .A1(n7000), .A2(n8334), .ZN(n8336) );
  NAND2_X1 U8898 ( .A1(n7112), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U8899 ( .A1(n7113), .A2(n8065), .ZN(n8004) );
  NAND3_X1 U8900 ( .A1(n6871), .A2(n6872), .A3(n6534), .ZN(n15375) );
  INV_X1 U8901 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15374) );
  XNOR2_X1 U8902 ( .A(n15362), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n15378) );
  NOR2_X1 U8903 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n6867) );
  NAND2_X1 U8904 ( .A1(n15325), .A2(n15324), .ZN(n15385) );
  XNOR2_X1 U8905 ( .A(n15328), .B(n7375), .ZN(n15390) );
  INV_X1 U8906 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n7375) );
  AND2_X1 U8907 ( .A1(n15335), .A2(n15334), .ZN(n15356) );
  NOR2_X1 U8908 ( .A1(n15335), .A2(n15334), .ZN(n15357) );
  NAND2_X1 U8909 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n6955), .ZN(n6954) );
  INV_X1 U8910 ( .A(n15455), .ZN(n6864) );
  NAND2_X1 U8911 ( .A1(n13829), .A2(n10424), .ZN(n7458) );
  NAND2_X1 U8912 ( .A1(n7756), .A2(n9867), .ZN(n12967) );
  NAND2_X1 U8913 ( .A1(n10190), .A2(n10189), .ZN(n13340) );
  INV_X1 U8914 ( .A(n7766), .ZN(n7764) );
  NAND2_X1 U8915 ( .A1(n10472), .A2(n11109), .ZN(n7367) );
  NAND2_X1 U8916 ( .A1(n10442), .A2(n12896), .ZN(n7368) );
  NAND2_X1 U8917 ( .A1(n7776), .A2(n9796), .ZN(n12984) );
  AOI21_X1 U8918 ( .B1(n7767), .B2(n6915), .A(n6517), .ZN(n6914) );
  INV_X1 U8919 ( .A(n7767), .ZN(n6916) );
  NAND2_X1 U8920 ( .A1(n9731), .A2(n13018), .ZN(n13026) );
  INV_X1 U8921 ( .A(n7318), .ZN(n7755) );
  INV_X1 U8922 ( .A(n7321), .ZN(n11247) );
  NAND2_X1 U8923 ( .A1(n7365), .A2(n9835), .ZN(n13053) );
  AND2_X1 U8924 ( .A1(n7760), .A2(n7763), .ZN(n13073) );
  AND2_X1 U8925 ( .A1(n11361), .A2(n9532), .ZN(n11525) );
  NAND2_X1 U8926 ( .A1(n7769), .A2(n9698), .ZN(n13092) );
  AOI21_X1 U8927 ( .B1(n10587), .B2(n10586), .A(n10585), .ZN(n10588) );
  NAND2_X1 U8928 ( .A1(n10590), .A2(n10592), .ZN(n7094) );
  OAI21_X1 U8929 ( .B1(n10435), .B2(n7358), .A(n6525), .ZN(n10466) );
  INV_X1 U8930 ( .A(n10457), .ZN(n13322) );
  NAND2_X1 U8931 ( .A1(n9863), .A2(n9862), .ZN(n13105) );
  INV_X1 U8932 ( .A(n13418), .ZN(n13108) );
  INV_X1 U8933 ( .A(n13457), .ZN(n13109) );
  INV_X1 U8934 ( .A(n13480), .ZN(n13111) );
  INV_X1 U8935 ( .A(n13469), .ZN(n13112) );
  INV_X1 U8936 ( .A(n13045), .ZN(n13116) );
  NAND2_X1 U8937 ( .A1(n10416), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9527) );
  NOR2_X1 U8938 ( .A1(n6453), .A2(n6561), .ZN(n6939) );
  OR2_X1 U8939 ( .A1(n9506), .A2(n9487), .ZN(n9488) );
  NAND2_X1 U8940 ( .A1(n10180), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9491) );
  NAND4_X1 U8941 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9461), .ZN(n15798)
         );
  AND2_X1 U8942 ( .A1(n6994), .A2(n6993), .ZN(n11028) );
  INV_X1 U8943 ( .A(n10985), .ZN(n6993) );
  NAND2_X1 U8944 ( .A1(n11006), .A2(n10986), .ZN(n6994) );
  NAND2_X1 U8945 ( .A1(n7686), .A2(n7684), .ZN(n11158) );
  AND2_X1 U8946 ( .A1(n6661), .A2(n7146), .ZN(n11348) );
  AOI21_X1 U8947 ( .B1(n13142), .B2(n7563), .A(n13141), .ZN(n13144) );
  AOI21_X1 U8948 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(n13132) );
  NAND2_X1 U8949 ( .A1(n13156), .A2(n13154), .ZN(n7572) );
  AND2_X1 U8950 ( .A1(n11493), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U8951 ( .A1(n13161), .A2(n7624), .ZN(n11486) );
  NAND2_X1 U8952 ( .A1(n7617), .A2(n7619), .ZN(n11857) );
  NAND2_X1 U8953 ( .A1(n13161), .A2(n7618), .ZN(n7617) );
  NAND2_X1 U8954 ( .A1(n7235), .A2(n7578), .ZN(n13176) );
  OAI21_X1 U8955 ( .B1(n13185), .B2(n6619), .A(n13184), .ZN(n13183) );
  NOR2_X1 U8956 ( .A1(n13204), .A2(n13748), .ZN(n13233) );
  NAND2_X1 U8957 ( .A1(n7582), .A2(n10611), .ZN(n13204) );
  NAND2_X1 U8958 ( .A1(n13197), .A2(n7588), .ZN(n13210) );
  NAND2_X1 U8959 ( .A1(n6992), .A2(n6990), .ZN(n13236) );
  AND2_X1 U8960 ( .A1(n13237), .A2(n6446), .ZN(n6990) );
  AND2_X1 U8961 ( .A1(n6992), .A2(n6446), .ZN(n13238) );
  NAND2_X1 U8962 ( .A1(n7689), .A2(n7693), .ZN(n13243) );
  AND2_X1 U8963 ( .A1(n7693), .A2(n7691), .ZN(n13244) );
  INV_X1 U8964 ( .A(n7690), .ZN(n7689) );
  NAND2_X1 U8965 ( .A1(n13253), .A2(n10614), .ZN(n13271) );
  AOI21_X1 U8966 ( .B1(n12369), .B2(n10424), .A(n8055), .ZN(n13327) );
  XNOR2_X1 U8967 ( .A(n6829), .B(n13329), .ZN(n13546) );
  NAND2_X1 U8968 ( .A1(n13355), .A2(n13328), .ZN(n6829) );
  NAND2_X1 U8969 ( .A1(n13339), .A2(n13338), .ZN(n13545) );
  INV_X1 U8970 ( .A(n13337), .ZN(n13338) );
  AOI21_X1 U8971 ( .B1(n13354), .B2(n15801), .A(n13353), .ZN(n13551) );
  NAND2_X1 U8972 ( .A1(n13352), .A2(n13351), .ZN(n13353) );
  NAND2_X1 U8973 ( .A1(n13348), .A2(n8044), .ZN(n13354) );
  OAI21_X1 U8974 ( .B1(n13376), .B2(n6813), .A(n10573), .ZN(n13369) );
  NAND2_X1 U8975 ( .A1(n7287), .A2(n7290), .ZN(n13365) );
  NAND2_X1 U8976 ( .A1(n13388), .A2(n7291), .ZN(n7287) );
  OR2_X1 U8977 ( .A1(n10237), .A2(n10563), .ZN(n7507) );
  NAND2_X1 U8978 ( .A1(n9855), .A2(n9854), .ZN(n10238) );
  NAND2_X1 U8979 ( .A1(n10237), .A2(n10468), .ZN(n13398) );
  NAND2_X1 U8980 ( .A1(n7925), .A2(n10550), .ZN(n13440) );
  NAND2_X1 U8981 ( .A1(n13451), .A2(n10540), .ZN(n7925) );
  NAND2_X1 U8982 ( .A1(n7296), .A2(n7379), .ZN(n13466) );
  NAND2_X1 U8983 ( .A1(n13481), .A2(n10541), .ZN(n13463) );
  NAND2_X1 U8984 ( .A1(n7708), .A2(n6441), .ZN(n7709) );
  NAND2_X1 U8985 ( .A1(n7708), .A2(n7712), .ZN(n13490) );
  OAI21_X1 U8986 ( .B1(n13516), .B2(n6901), .A(n6899), .ZN(n13507) );
  NAND2_X1 U8987 ( .A1(n6898), .A2(n10530), .ZN(n13509) );
  NAND2_X1 U8988 ( .A1(n13516), .A2(n13517), .ZN(n6898) );
  NAND2_X1 U8989 ( .A1(n10139), .A2(n10138), .ZN(n12002) );
  NAND2_X1 U8990 ( .A1(n12094), .A2(n7939), .ZN(n12000) );
  AND2_X1 U8991 ( .A1(n15813), .A2(n11514), .ZN(n13537) );
  NAND2_X1 U8992 ( .A1(n10229), .A2(n10493), .ZN(n7917) );
  NOR2_X1 U8993 ( .A1(n11318), .A2(n15809), .ZN(n11777) );
  NAND2_X1 U8994 ( .A1(n10123), .A2(n10122), .ZN(n15780) );
  INV_X2 U8995 ( .A(n15813), .ZN(n15816) );
  AND2_X2 U8996 ( .A1(n11316), .A2(n15809), .ZN(n15812) );
  NAND2_X1 U8997 ( .A1(n11777), .A2(n15836), .ZN(n13534) );
  INV_X1 U8998 ( .A(n10221), .ZN(n7510) );
  AND2_X1 U8999 ( .A1(n15873), .A2(n15836), .ZN(n13754) );
  INV_X1 U9000 ( .A(n13754), .ZN(n13750) );
  INV_X1 U9001 ( .A(n10458), .ZN(n13758) );
  INV_X1 U9002 ( .A(n13327), .ZN(n13760) );
  NAND2_X1 U9003 ( .A1(n10206), .A2(n10205), .ZN(n12920) );
  AOI21_X1 U9004 ( .B1(n13546), .B2(n15851), .A(n13545), .ZN(n13766) );
  NAND2_X1 U9005 ( .A1(n9693), .A2(n9692), .ZN(n13814) );
  INV_X1 U9006 ( .A(n11547), .ZN(n11519) );
  INV_X1 U9007 ( .A(n9466), .ZN(n11358) );
  AND2_X1 U9008 ( .A1(n10621), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13816) );
  INV_X1 U9009 ( .A(n9413), .ZN(n12371) );
  XNOR2_X1 U9010 ( .A(n7091), .B(n10163), .ZN(n13833) );
  NAND2_X1 U9011 ( .A1(n7471), .A2(n10162), .ZN(n7091) );
  NAND2_X1 U9012 ( .A1(n6826), .A2(n9853), .ZN(n11782) );
  OAI21_X1 U9013 ( .B1(n7081), .B2(n7077), .A(n7450), .ZN(n9853) );
  NAND2_X1 U9014 ( .A1(n9837), .A2(n6827), .ZN(n6826) );
  NOR2_X1 U9015 ( .A1(n9894), .A2(n9902), .ZN(n11702) );
  INV_X1 U9016 ( .A(n9892), .ZN(n9894) );
  NAND2_X1 U9017 ( .A1(n9818), .A2(n9817), .ZN(n9823) );
  OAI21_X1 U9018 ( .B1(n9797), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n9799), .ZN(
        n9816) );
  XNOR2_X1 U9019 ( .A(n9449), .B(n9448), .ZN(n11454) );
  INV_X1 U9020 ( .A(SI_19_), .ZN(n11193) );
  INV_X1 U9021 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9452) );
  OAI21_X1 U9022 ( .B1(n9755), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9453) );
  INV_X1 U9023 ( .A(n7087), .ZN(n9767) );
  AOI21_X1 U9024 ( .B1(n7453), .B2(n7454), .A(n7089), .ZN(n7087) );
  NAND2_X1 U9025 ( .A1(n7934), .A2(n9735), .ZN(n9754) );
  NAND2_X1 U9026 ( .A1(n9734), .A2(n9733), .ZN(n7934) );
  INV_X1 U9027 ( .A(SI_16_), .ZN(n10957) );
  INV_X1 U9028 ( .A(SI_15_), .ZN(n13693) );
  XNOR2_X1 U9029 ( .A(n9669), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13230) );
  INV_X1 U9030 ( .A(SI_12_), .ZN(n10860) );
  NAND2_X1 U9031 ( .A1(n9664), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9644) );
  INV_X1 U9032 ( .A(SI_11_), .ZN(n10863) );
  NAND2_X1 U9033 ( .A1(n7929), .A2(n9589), .ZN(n9608) );
  NAND2_X1 U9034 ( .A1(n9588), .A2(n9587), .ZN(n7929) );
  NAND2_X1 U9035 ( .A1(n7465), .A2(n9558), .ZN(n9573) );
  OR2_X1 U9036 ( .A1(n9557), .A2(n9556), .ZN(n7465) );
  NAND2_X1 U9037 ( .A1(n7149), .A2(n7148), .ZN(n7151) );
  XNOR2_X1 U9038 ( .A(P3_IR_REG_31__SCAN_IN), .B(P3_IR_REG_4__SCAN_IN), .ZN(
        n7148) );
  NAND2_X1 U9039 ( .A1(n9475), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U9040 ( .A1(n7913), .A2(n9474), .ZN(n9499) );
  NAND2_X1 U9041 ( .A1(n9411), .A2(n9483), .ZN(n7238) );
  AOI21_X1 U9042 ( .B1(n11383), .B2(n7272), .A(n6434), .ZN(n7269) );
  NAND2_X1 U9043 ( .A1(n12098), .A2(n9302), .ZN(n6679) );
  NAND2_X1 U9044 ( .A1(n9052), .A2(n9051), .ZN(n12460) );
  NAND2_X1 U9045 ( .A1(n13960), .A2(n8925), .ZN(n13862) );
  NOR2_X1 U9046 ( .A1(n6770), .A2(n6432), .ZN(n11846) );
  INV_X1 U9047 ( .A(n6773), .ZN(n6770) );
  INV_X1 U9048 ( .A(n7723), .ZN(n7722) );
  NAND2_X1 U9049 ( .A1(n7724), .A2(n7727), .ZN(n11421) );
  OR2_X1 U9050 ( .A1(n13878), .A2(n13879), .ZN(n13944) );
  NAND2_X1 U9051 ( .A1(n12288), .A2(n9081), .ZN(n12324) );
  OAI21_X1 U9052 ( .B1(n9128), .B2(n7735), .A(n7733), .ZN(n13911) );
  AND2_X1 U9053 ( .A1(n8939), .A2(n8925), .ZN(n7720) );
  NOR2_X1 U9054 ( .A1(n7796), .A2(n7170), .ZN(n12380) );
  AND2_X1 U9055 ( .A1(n9374), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U9056 ( .A1(n9204), .A2(n13869), .ZN(n13937) );
  NAND2_X1 U9057 ( .A1(n7278), .A2(n9064), .ZN(n12291) );
  AND2_X1 U9058 ( .A1(n9165), .A2(n9164), .ZN(n14330) );
  NAND2_X1 U9059 ( .A1(n6487), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U9060 ( .A1(n13968), .A2(n13967), .ZN(n13966) );
  NAND2_X1 U9061 ( .A1(n11383), .A2(n8978), .ZN(n11428) );
  AND2_X1 U9062 ( .A1(n11392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13873) );
  NAND2_X1 U9063 ( .A1(n9137), .A2(n9136), .ZN(n13999) );
  NAND2_X1 U9064 ( .A1(n9246), .A2(n9245), .ZN(n14227) );
  OR2_X1 U9065 ( .A1(n14257), .A2(n9326), .ZN(n9246) );
  INV_X1 U9066 ( .A(n14303), .ZN(n14008) );
  OR2_X1 U9067 ( .A1(n9094), .A2(n9093), .ZN(n14012) );
  INV_X1 U9068 ( .A(n12380), .ZN(n14024) );
  NAND2_X1 U9069 ( .A1(n15642), .A2(n15643), .ZN(n15641) );
  NAND2_X1 U9070 ( .A1(n15656), .A2(n15657), .ZN(n15655) );
  NAND2_X1 U9071 ( .A1(n14061), .A2(n14060), .ZN(n11063) );
  NAND2_X1 U9072 ( .A1(n11065), .A2(n11064), .ZN(n14087) );
  OAI211_X1 U9073 ( .C1(n11065), .C2(n6719), .A(n6714), .B(n11066), .ZN(n14089) );
  INV_X1 U9074 ( .A(n6717), .ZN(n6714) );
  NAND2_X1 U9075 ( .A1(n11263), .A2(n6723), .ZN(n15682) );
  NOR2_X1 U9076 ( .A1(n6725), .A2(n6724), .ZN(n6723) );
  INV_X1 U9077 ( .A(n11071), .ZN(n6724) );
  INV_X1 U9078 ( .A(n11072), .ZN(n6725) );
  AND2_X1 U9079 ( .A1(n11263), .A2(n11071), .ZN(n11073) );
  NAND2_X1 U9080 ( .A1(n15684), .A2(n6625), .ZN(n14095) );
  INV_X1 U9081 ( .A(n14093), .ZN(n6726) );
  NAND2_X1 U9082 ( .A1(n15684), .A2(n11789), .ZN(n14094) );
  NAND2_X1 U9083 ( .A1(n11797), .A2(n11796), .ZN(n14132) );
  AND2_X1 U9084 ( .A1(n11813), .A2(n11812), .ZN(n14142) );
  OAI21_X1 U9085 ( .B1(n11797), .B2(n6722), .A(n6720), .ZN(n15711) );
  INV_X1 U9086 ( .A(n6721), .ZN(n6720) );
  OAI21_X1 U9087 ( .B1(n11796), .B2(n6722), .A(n14133), .ZN(n6721) );
  NAND2_X1 U9088 ( .A1(n15711), .A2(n15710), .ZN(n15709) );
  XNOR2_X1 U9089 ( .A(n6727), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14162) );
  INV_X1 U9090 ( .A(n14161), .ZN(n15708) );
  NAND2_X1 U9091 ( .A1(n10280), .A2(n7154), .ZN(n7160) );
  NAND2_X1 U9092 ( .A1(n7789), .A2(n9979), .ZN(n14181) );
  AND2_X1 U9093 ( .A1(n8026), .A2(n10040), .ZN(n14186) );
  NAND2_X1 U9094 ( .A1(n8026), .A2(n8025), .ZN(n14419) );
  INV_X1 U9095 ( .A(n7347), .ZN(n7346) );
  XNOR2_X1 U9096 ( .A(n14195), .B(n7349), .ZN(n7348) );
  NAND2_X1 U9097 ( .A1(n14234), .A2(n10037), .ZN(n14207) );
  AND2_X1 U9098 ( .A1(n7070), .A2(n10034), .ZN(n14235) );
  NAND2_X1 U9099 ( .A1(n14263), .A2(n9974), .ZN(n14252) );
  NAND2_X1 U9100 ( .A1(n7397), .A2(n9967), .ZN(n14299) );
  NAND2_X1 U9101 ( .A1(n14333), .A2(n10028), .ZN(n14311) );
  NOR2_X1 U9102 ( .A1(n14389), .A2(n8009), .ZN(n8008) );
  INV_X1 U9103 ( .A(n8013), .ZN(n8009) );
  NAND2_X1 U9104 ( .A1(n8010), .A2(n8013), .ZN(n14390) );
  NAND2_X1 U9105 ( .A1(n10022), .A2(n12239), .ZN(n12332) );
  INV_X1 U9106 ( .A(n7782), .ZN(n12334) );
  AOI21_X1 U9107 ( .B1(n12241), .B2(n9959), .A(n7785), .ZN(n7782) );
  NAND2_X1 U9108 ( .A1(n7051), .A2(n10021), .ZN(n12238) );
  NAND2_X1 U9109 ( .A1(n8014), .A2(n8016), .ZN(n7051) );
  NAND2_X1 U9110 ( .A1(n8015), .A2(n8017), .ZN(n12148) );
  OR2_X1 U9111 ( .A1(n12118), .A2(n8019), .ZN(n8015) );
  NAND2_X1 U9112 ( .A1(n8021), .A2(n8020), .ZN(n11920) );
  AND2_X1 U9113 ( .A1(n8021), .A2(n10017), .ZN(n11921) );
  NAND2_X1 U9114 ( .A1(n12118), .A2(n10019), .ZN(n8021) );
  NAND2_X1 U9115 ( .A1(n11731), .A2(n10014), .ZN(n11754) );
  NOR2_X1 U9116 ( .A1(n8036), .A2(n8035), .ZN(n11732) );
  INV_X1 U9117 ( .A(n10012), .ZN(n8035) );
  INV_X1 U9118 ( .A(n11530), .ZN(n8036) );
  OAI21_X1 U9119 ( .B1(n11626), .B2(n6493), .A(n10011), .ZN(n11473) );
  INV_X1 U9120 ( .A(n10044), .ZN(n11574) );
  NAND2_X1 U9121 ( .A1(n7186), .A2(n7184), .ZN(n14522) );
  NAND2_X1 U9122 ( .A1(n6498), .A2(n7187), .ZN(n7186) );
  AND2_X1 U9123 ( .A1(n14423), .A2(n7185), .ZN(n7184) );
  AND2_X1 U9124 ( .A1(n14419), .A2(n15764), .ZN(n7187) );
  AND2_X1 U9125 ( .A1(n9274), .A2(n9273), .ZN(n14527) );
  AND2_X1 U9126 ( .A1(n9229), .A2(n9228), .ZN(n14537) );
  INV_X1 U9127 ( .A(n12460), .ZN(n12120) );
  NAND2_X1 U9128 ( .A1(n9036), .A2(n9035), .ZN(n12455) );
  NOR2_X1 U9129 ( .A1(n15733), .A2(n6784), .ZN(n15734) );
  AND2_X1 U9130 ( .A1(n15750), .A2(n10044), .ZN(n6784) );
  AND2_X1 U9131 ( .A1(n9386), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15722) );
  INV_X1 U9132 ( .A(n8891), .ZN(n12912) );
  NAND2_X1 U9133 ( .A1(n7169), .A2(n7166), .ZN(n14563) );
  NOR2_X1 U9134 ( .A1(n7168), .A2(n7167), .ZN(n7166) );
  NOR2_X1 U9135 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7167) );
  XNOR2_X1 U9136 ( .A(n9336), .B(n9335), .ZN(n14571) );
  INV_X1 U9137 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9335) );
  OAI21_X1 U9138 ( .B1(n9340), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9336) );
  INV_X1 U9139 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12285) );
  MUX2_X1 U9140 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8847), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8849) );
  INV_X1 U9141 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11541) );
  INV_X1 U9142 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11408) );
  INV_X1 U9143 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11360) );
  INV_X1 U9144 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11323) );
  INV_X1 U9145 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11132) );
  INV_X1 U9146 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11308) );
  INV_X1 U9147 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n13593) );
  INV_X1 U9148 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10912) );
  INV_X1 U9149 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10867) );
  INV_X1 U9150 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10753) );
  MUX2_X1 U9151 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8911), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8913) );
  NAND2_X1 U9152 ( .A1(n8910), .A2(n6728), .ZN(n15619) );
  INV_X1 U9153 ( .A(n6729), .ZN(n6728) );
  OAI21_X1 U9154 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_1__SCAN_IN), .A(
        n6730), .ZN(n6729) );
  NAND2_X1 U9155 ( .A1(n7983), .A2(n14682), .ZN(n11708) );
  NAND3_X1 U9156 ( .A1(n11196), .A2(n8266), .A3(n11210), .ZN(n8317) );
  AND2_X1 U9157 ( .A1(n11196), .A2(n8266), .ZN(n11209) );
  AND2_X1 U9158 ( .A1(n14671), .A2(n7232), .ZN(n14601) );
  NAND2_X1 U9159 ( .A1(n14671), .A2(n8591), .ZN(n14602) );
  AOI21_X1 U9160 ( .B1(n7970), .B2(n6801), .A(n6571), .ZN(n6800) );
  INV_X1 U9161 ( .A(n7970), .ZN(n6802) );
  INV_X1 U9162 ( .A(n8225), .ZN(n7360) );
  OR2_X1 U9163 ( .A1(n11171), .A2(n8755), .ZN(n8244) );
  NAND2_X1 U9164 ( .A1(n11172), .A2(n11171), .ZN(n8245) );
  OR2_X1 U9165 ( .A1(n14655), .A2(n7989), .ZN(n14607) );
  NOR2_X1 U9166 ( .A1(n14655), .A2(n7991), .ZN(n14608) );
  OAI211_X1 U9167 ( .C1(n8441), .C2(n7209), .A(n7214), .B(n7207), .ZN(n12253)
         );
  AND2_X1 U9168 ( .A1(n12254), .A2(n12251), .ZN(n7214) );
  NAND2_X1 U9169 ( .A1(n7199), .A2(n8670), .ZN(n14646) );
  OR2_X1 U9170 ( .A1(n14672), .A2(n7231), .ZN(n6794) );
  NAND2_X1 U9171 ( .A1(n7985), .A2(n11411), .ZN(n14684) );
  OR2_X1 U9172 ( .A1(n8817), .A2(P1_U3086), .ZN(n12878) );
  OR3_X1 U9173 ( .A1(n10100), .A2(n10099), .A3(n10098), .ZN(n14719) );
  INV_X1 U9174 ( .A(n12653), .ZN(n14720) );
  NAND2_X1 U9175 ( .A1(n8728), .A2(n8727), .ZN(n14722) );
  NAND2_X1 U9176 ( .A1(n8684), .A2(n8683), .ZN(n14724) );
  AND2_X1 U9177 ( .A1(n8642), .A2(n8641), .ZN(n14612) );
  NAND2_X1 U9178 ( .A1(n8226), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8299) );
  INV_X1 U9179 ( .A(n7493), .ZN(n7841) );
  OAI211_X1 U9180 ( .C1(n8267), .C2(n14749), .A(n8249), .B(n7494), .ZN(n7493)
         );
  CLKBUF_X1 U9181 ( .A(n10302), .Z(n14747) );
  NAND2_X1 U9182 ( .A1(n7032), .A2(n10850), .ZN(n14774) );
  OR2_X1 U9183 ( .A1(n14756), .A2(n14752), .ZN(n7032) );
  NAND2_X1 U9184 ( .A1(n10838), .A2(n6523), .ZN(n14758) );
  AND2_X1 U9185 ( .A1(n7030), .A2(n7028), .ZN(n7027) );
  NAND2_X1 U9186 ( .A1(n7026), .A2(n7025), .ZN(n11185) );
  INV_X1 U9187 ( .A(n11184), .ZN(n7024) );
  NOR2_X1 U9188 ( .A1(n10894), .A2(n7421), .ZN(n10944) );
  NOR2_X1 U9189 ( .A1(n10894), .A2(n7422), .ZN(n10930) );
  AOI21_X1 U9190 ( .B1(n10894), .B2(n7420), .A(n6583), .ZN(n10919) );
  NAND2_X1 U9191 ( .A1(n7421), .A2(n7420), .ZN(n7419) );
  INV_X1 U9192 ( .A(n7041), .ZN(n10960) );
  AOI21_X1 U9193 ( .B1(n7045), .B2(n6433), .A(n7044), .ZN(n7041) );
  NAND2_X1 U9194 ( .A1(n7045), .A2(n7047), .ZN(n10952) );
  AND2_X1 U9195 ( .A1(n7418), .A2(n6508), .ZN(n10965) );
  NAND2_X1 U9196 ( .A1(n7418), .A2(n7417), .ZN(n11134) );
  OAI21_X1 U9197 ( .B1(n7045), .B2(n7044), .A(n7042), .ZN(n11141) );
  INV_X1 U9198 ( .A(n7043), .ZN(n7042) );
  OAI21_X1 U9199 ( .B1(n6433), .B2(n7044), .A(n10959), .ZN(n7043) );
  NAND2_X1 U9200 ( .A1(n11466), .A2(n11465), .ZN(n11681) );
  XNOR2_X1 U9201 ( .A(n7409), .B(n15476), .ZN(n15474) );
  NAND2_X1 U9202 ( .A1(n14779), .A2(n6643), .ZN(n14783) );
  NAND2_X1 U9203 ( .A1(n7037), .A2(n14788), .ZN(n14795) );
  OR2_X1 U9204 ( .A1(n14790), .A2(n14789), .ZN(n7037) );
  NOR2_X1 U9205 ( .A1(n14869), .A2(n14868), .ZN(n14871) );
  NAND2_X1 U9206 ( .A1(n10337), .A2(n10336), .ZN(n14916) );
  AND2_X1 U9207 ( .A1(n7853), .A2(n7851), .ZN(n14911) );
  NAND2_X1 U9208 ( .A1(n14986), .A2(n10386), .ZN(n14965) );
  NAND2_X1 U9209 ( .A1(n10385), .A2(n10384), .ZN(n14984) );
  NAND2_X1 U9210 ( .A1(n15008), .A2(n10331), .ZN(n14988) );
  AND2_X1 U9211 ( .A1(n8531), .A2(n8530), .ZN(n15064) );
  NAND2_X1 U9212 ( .A1(n7483), .A2(n10377), .ZN(n15053) );
  NAND2_X1 U9213 ( .A1(n7486), .A2(n7485), .ZN(n7483) );
  NAND2_X1 U9214 ( .A1(n8202), .A2(n8201), .ZN(n12724) );
  NAND2_X1 U9215 ( .A1(n7006), .A2(n7004), .ZN(n12308) );
  INV_X1 U9216 ( .A(n7005), .ZN(n7004) );
  INV_X1 U9217 ( .A(n15519), .ZN(n15015) );
  AND2_X1 U9218 ( .A1(n12835), .A2(n10310), .ZN(n7966) );
  INV_X1 U9219 ( .A(n15096), .ZN(n15515) );
  NAND2_X1 U9220 ( .A1(n7956), .A2(n12677), .ZN(n11823) );
  AND2_X1 U9221 ( .A1(n15513), .A2(n11833), .ZN(n15100) );
  AND2_X1 U9222 ( .A1(n15513), .A2(n11828), .ZN(n15519) );
  AND2_X1 U9223 ( .A1(n10106), .A2(n10756), .ZN(n15531) );
  AND2_X2 U9224 ( .A1(n10115), .A2(n10114), .ZN(n15618) );
  NAND2_X1 U9225 ( .A1(n10093), .A2(n10092), .ZN(n12862) );
  AND2_X1 U9226 ( .A1(n15125), .A2(n15124), .ZN(n15246) );
  INV_X1 U9227 ( .A(n6926), .ZN(n6925) );
  OAI21_X1 U9228 ( .B1(n15134), .B2(n15558), .A(n7495), .ZN(n6926) );
  NAND2_X1 U9229 ( .A1(n6497), .A2(n15572), .ZN(n6668) );
  NOR2_X1 U9230 ( .A1(n14856), .A2(n14857), .ZN(n6669) );
  AOI21_X1 U9231 ( .B1(n15144), .B2(n15572), .A(n6886), .ZN(n6885) );
  NAND2_X1 U9232 ( .A1(n15141), .A2(n15142), .ZN(n6886) );
  NAND2_X1 U9233 ( .A1(n7017), .A2(n7016), .ZN(n7015) );
  INV_X1 U9234 ( .A(n15148), .ZN(n7016) );
  NAND2_X1 U9235 ( .A1(n15309), .A2(n8235), .ZN(n15263) );
  NAND2_X1 U9236 ( .A1(n10865), .A2(n10091), .ZN(n6788) );
  NAND2_X1 U9237 ( .A1(n10756), .A2(n10755), .ZN(n15541) );
  NAND2_X1 U9238 ( .A1(n6664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7248) );
  INV_X1 U9239 ( .A(n8790), .ZN(n15308) );
  INV_X1 U9240 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12283) );
  MUX2_X1 U9241 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8153), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8155) );
  NAND2_X1 U9242 ( .A1(n8793), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8180) );
  INV_X1 U9243 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11706) );
  INV_X1 U9244 ( .A(n8801), .ZN(n12822) );
  INV_X1 U9245 ( .A(n12652), .ZN(n11828) );
  INV_X1 U9246 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11306) );
  INV_X1 U9247 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11121) );
  INV_X1 U9248 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11258) );
  INV_X1 U9249 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11208) );
  INV_X1 U9250 ( .A(n11684), .ZN(n11469) );
  INV_X1 U9251 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10914) );
  INV_X1 U9252 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10866) );
  INV_X1 U9253 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10837) );
  INV_X1 U9254 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10799) );
  INV_X1 U9255 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10765) );
  INV_X1 U9256 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10745) );
  INV_X1 U9257 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10782) );
  AND2_X1 U9258 ( .A1(n6941), .A2(n6940), .ZN(n15884) );
  OAI21_X1 U9259 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15376), .A(n15882), .ZN(
        n15874) );
  NOR2_X1 U9260 ( .A1(n15884), .A2(n15883), .ZN(n15376) );
  XNOR2_X1 U9261 ( .A(n15365), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15875) );
  AND2_X1 U9262 ( .A1(n6877), .A2(n15429), .ZN(n15401) );
  NAND2_X1 U9263 ( .A1(n15448), .A2(n15449), .ZN(n15445) );
  NAND2_X1 U9264 ( .A1(n7868), .A2(n7866), .ZN(n7355) );
  INV_X1 U9265 ( .A(n7869), .ZN(n7356) );
  NAND2_X1 U9266 ( .A1(n15466), .A2(n15467), .ZN(n15465) );
  NAND2_X1 U9267 ( .A1(n15435), .A2(n15433), .ZN(n15441) );
  INV_X1 U9268 ( .A(n15442), .ZN(n6875) );
  AOI21_X1 U9269 ( .B1(n15441), .B2(n15442), .A(n7882), .ZN(n7881) );
  INV_X1 U9270 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U9271 ( .A1(n11523), .A2(n9551), .ZN(n11671) );
  AND2_X1 U9272 ( .A1(n9931), .A2(n8041), .ZN(n7364) );
  NAND2_X1 U9273 ( .A1(n9585), .A2(n9584), .ZN(n12040) );
  XNOR2_X1 U9274 ( .A(n13085), .B(n6956), .ZN(n13091) );
  NAND2_X1 U9275 ( .A1(n6999), .A2(n6998), .ZN(n7677) );
  OAI21_X1 U9276 ( .B1(n13302), .B2(n6451), .A(n13315), .ZN(n6999) );
  NAND2_X1 U9277 ( .A1(n6842), .A2(n6840), .ZN(P3_U3455) );
  NOR2_X1 U9278 ( .A1(n6628), .A2(n6841), .ZN(n6840) );
  OR2_X1 U9279 ( .A1(n13766), .A2(n15858), .ZN(n6842) );
  NOR2_X1 U9280 ( .A1(n15860), .A2(n13765), .ZN(n6841) );
  NAND2_X1 U9281 ( .A1(n10057), .A2(n13986), .ZN(n10063) );
  AOI21_X1 U9282 ( .B1(n14414), .B2(n14399), .A(n10051), .ZN(n10052) );
  MUX2_X1 U9283 ( .A(n14408), .B(n14513), .S(n15778), .Z(n14409) );
  NAND2_X1 U9284 ( .A1(n12934), .A2(n12108), .ZN(n10293) );
  NAND2_X1 U9285 ( .A1(n7183), .A2(n7182), .ZN(P2_U3526) );
  NAND2_X1 U9286 ( .A1(n15775), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U9287 ( .A1(n14522), .A2(n15778), .ZN(n7183) );
  MUX2_X1 U9288 ( .A(n14514), .B(n14513), .S(n15767), .Z(n14515) );
  NAND2_X1 U9289 ( .A1(n7056), .A2(n7055), .ZN(P2_U3496) );
  NAND2_X1 U9290 ( .A1(n15765), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U9291 ( .A1(n14521), .A2(n15767), .ZN(n7056) );
  NAND2_X1 U9292 ( .A1(n12934), .A2(n12114), .ZN(n10299) );
  NAND2_X1 U9293 ( .A1(n7225), .A2(n14685), .ZN(n7222) );
  XNOR2_X1 U9294 ( .A(n7353), .B(n7974), .ZN(n14703) );
  NAND2_X1 U9295 ( .A1(n7413), .A2(n7414), .ZN(n11137) );
  OAI211_X1 U9296 ( .C1(n14819), .C2(n12652), .A(n6709), .B(n6651), .ZN(
        P1_U3262) );
  OAI21_X1 U9297 ( .B1(n7035), .B2(n6710), .A(n12652), .ZN(n6709) );
  OAI21_X1 U9298 ( .B1(n15252), .B2(n15605), .A(n6882), .ZN(P1_U3522) );
  NOR2_X1 U9299 ( .A1(n6884), .A2(n6883), .ZN(n6882) );
  NOR2_X1 U9300 ( .A1(n15606), .A2(n15253), .ZN(n6883) );
  NOR2_X1 U9301 ( .A1(n15254), .A2(n15288), .ZN(n6884) );
  NAND2_X1 U9302 ( .A1(n8168), .A2(n8169), .ZN(n15297) );
  INV_X1 U9303 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9472) );
  AND2_X1 U9304 ( .A1(n7336), .A2(n7330), .ZN(n15427) );
  NAND2_X1 U9305 ( .A1(n15456), .A2(n15455), .ZN(n15454) );
  NAND2_X1 U9306 ( .A1(n7861), .A2(n15450), .ZN(n15456) );
  NAND2_X1 U9307 ( .A1(n15459), .A2(n15460), .ZN(n15458) );
  NAND2_X1 U9308 ( .A1(n7872), .A2(n7870), .ZN(n15462) );
  XNOR2_X1 U9309 ( .A(n7337), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9310 ( .A1(n7339), .A2(n7338), .ZN(n7337) );
  NAND2_X1 U9311 ( .A1(n15441), .A2(n15442), .ZN(n7338) );
  NAND2_X1 U9312 ( .A1(n8771), .A2(n8770), .ZN(n14839) );
  XOR2_X1 U9313 ( .A(n13549), .B(n7457), .Z(n6423) );
  AND2_X1 U9314 ( .A1(n14347), .A2(n7890), .ZN(n6424) );
  AND2_X1 U9315 ( .A1(n10045), .A2(n7888), .ZN(n6425) );
  AND2_X1 U9316 ( .A1(n12797), .A2(n12799), .ZN(n6426) );
  AND2_X1 U9317 ( .A1(n7885), .A2(n7886), .ZN(n6427) );
  INV_X1 U9318 ( .A(n15006), .ZN(n15001) );
  OR2_X1 U9319 ( .A1(n12525), .A2(n12522), .ZN(n6428) );
  AND2_X2 U9320 ( .A1(n7243), .A2(n15517), .ZN(n8292) );
  INV_X1 U9321 ( .A(n13115), .ZN(n13522) );
  NAND2_X1 U9322 ( .A1(n8440), .A2(n8439), .ZN(n6429) );
  INV_X1 U9323 ( .A(n13155), .ZN(n7575) );
  NOR2_X1 U9324 ( .A1(n13190), .A2(n10693), .ZN(n6430) );
  AND2_X1 U9325 ( .A1(n8995), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U9326 ( .A1(n7270), .A2(n6535), .ZN(n6432) );
  AND2_X1 U9327 ( .A1(n7047), .A2(n6659), .ZN(n6433) );
  AND2_X1 U9328 ( .A1(n8988), .A2(n8987), .ZN(n6434) );
  AND2_X1 U9329 ( .A1(n10366), .A2(n7855), .ZN(n6435) );
  AND2_X1 U9330 ( .A1(n14180), .A2(n7790), .ZN(n6436) );
  XNOR2_X1 U9331 ( .A(n13979), .B(n14420), .ZN(n14185) );
  INV_X1 U9332 ( .A(n14185), .ZN(n14180) );
  NAND2_X1 U9333 ( .A1(n10481), .A2(n10470), .ZN(n11437) );
  INV_X1 U9334 ( .A(n12527), .ZN(n7839) );
  INV_X1 U9335 ( .A(n15727), .ZN(n11663) );
  OR2_X1 U9336 ( .A1(n10683), .A2(n15867), .ZN(n6437) );
  INV_X1 U9337 ( .A(n12828), .ZN(n7177) );
  AND2_X1 U9338 ( .A1(n7637), .A2(n15225), .ZN(n6438) );
  OR2_X1 U9339 ( .A1(n7034), .A2(n15512), .ZN(n6439) );
  AND2_X1 U9340 ( .A1(n6579), .A2(n6985), .ZN(n6440) );
  NAND2_X1 U9341 ( .A1(n9103), .A2(n9102), .ZN(n14495) );
  XNOR2_X1 U9342 ( .A(n7125), .B(n14903), .ZN(n14897) );
  INV_X1 U9343 ( .A(n14897), .ZN(n14902) );
  AND2_X1 U9344 ( .A1(n6500), .A2(n7712), .ZN(n6441) );
  AND2_X1 U9345 ( .A1(n14425), .A2(n14006), .ZN(n6442) );
  AND3_X1 U9346 ( .A1(n11974), .A2(n11883), .A3(n11972), .ZN(n6443) );
  AND2_X1 U9347 ( .A1(n15286), .A2(n6438), .ZN(n6444) );
  NAND2_X1 U9348 ( .A1(n9194), .A2(n9193), .ZN(n14321) );
  INV_X1 U9349 ( .A(n14321), .ZN(n7890) );
  AND2_X1 U9350 ( .A1(n7884), .A2(n14233), .ZN(n6445) );
  XNOR2_X1 U9351 ( .A(n15797), .B(n15790), .ZN(n10224) );
  NAND2_X1 U9352 ( .A1(n13215), .A2(n10662), .ZN(n6446) );
  AND2_X1 U9353 ( .A1(n11498), .A2(n6417), .ZN(n6447) );
  INV_X1 U9354 ( .A(n13118), .ZN(n12211) );
  AND2_X1 U9355 ( .A1(n12519), .A2(n12520), .ZN(n6448) );
  AND2_X1 U9356 ( .A1(n7407), .A2(n7180), .ZN(n6449) );
  INV_X1 U9357 ( .A(n14890), .ZN(n15254) );
  NAND2_X1 U9358 ( .A1(n8720), .A2(n8719), .ZN(n14890) );
  AND2_X1 U9359 ( .A1(n10136), .A2(n7747), .ZN(n6450) );
  AND2_X1 U9360 ( .A1(n10671), .A2(n10672), .ZN(n6451) );
  AND2_X1 U9361 ( .A1(n6578), .A2(n7436), .ZN(n6452) );
  NAND2_X1 U9362 ( .A1(n10517), .A2(n10507), .ZN(n6895) );
  AND2_X1 U9363 ( .A1(n9598), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6453) );
  INV_X1 U9364 ( .A(n7621), .ZN(n7618) );
  NAND2_X1 U9365 ( .A1(n6658), .A2(n7624), .ZN(n7621) );
  NAND2_X1 U9366 ( .A1(n9484), .A2(n11033), .ZN(n6454) );
  INV_X1 U9367 ( .A(n14169), .ZN(n14520) );
  NAND2_X1 U9368 ( .A1(n12533), .A2(n12532), .ZN(n14169) );
  OR2_X1 U9369 ( .A1(n14336), .A2(n8007), .ZN(n6455) );
  NAND2_X1 U9370 ( .A1(n10574), .A2(n6417), .ZN(n6456) );
  AND2_X1 U9371 ( .A1(n6646), .A2(n11411), .ZN(n7984) );
  OR2_X1 U9372 ( .A1(n6738), .A2(n6740), .ZN(n6457) );
  INV_X1 U9373 ( .A(n10550), .ZN(n7924) );
  OR2_X1 U9374 ( .A1(n7427), .A2(n14807), .ZN(n6458) );
  NAND2_X1 U9375 ( .A1(n8964), .A2(n8963), .ZN(n12404) );
  AND2_X1 U9376 ( .A1(n7259), .A2(n10379), .ZN(n6459) );
  OR2_X1 U9377 ( .A1(n13057), .A2(n13401), .ZN(n10468) );
  INV_X1 U9378 ( .A(n10468), .ZN(n7509) );
  AND2_X1 U9379 ( .A1(n9867), .A2(n13419), .ZN(n6460) );
  AND2_X1 U9380 ( .A1(n12368), .A2(n6858), .ZN(n6461) );
  OR2_X1 U9381 ( .A1(n12773), .A2(n12774), .ZN(n6462) );
  INV_X1 U9382 ( .A(n7200), .ZN(n13278) );
  OR2_X1 U9383 ( .A1(n7201), .A2(n6595), .ZN(n7200) );
  OR2_X1 U9384 ( .A1(n6864), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6463) );
  INV_X1 U9385 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10780) );
  XNOR2_X1 U9386 ( .A(n15291), .B(n14737), .ZN(n12840) );
  INV_X1 U9387 ( .A(n12840), .ZN(n7010) );
  INV_X1 U9388 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11543) );
  AND2_X1 U9389 ( .A1(n11763), .A2(n6427), .ZN(n6857) );
  AND2_X1 U9390 ( .A1(n6857), .A2(n12368), .ZN(n12153) );
  XOR2_X1 U9391 ( .A(n10082), .B(n10083), .Z(n6464) );
  AND2_X1 U9392 ( .A1(n7073), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6465) );
  AND2_X1 U9393 ( .A1(n15873), .A2(n15789), .ZN(n6466) );
  AND2_X1 U9394 ( .A1(n10403), .A2(n6640), .ZN(n6467) );
  AND2_X1 U9395 ( .A1(n10692), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6468) );
  AND2_X1 U9396 ( .A1(n10542), .A2(n10541), .ZN(n6469) );
  AND2_X1 U9397 ( .A1(n7562), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6470) );
  INV_X1 U9398 ( .A(n14717), .ZN(n14685) );
  AND2_X1 U9399 ( .A1(n7076), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6471) );
  AND2_X1 U9400 ( .A1(n15809), .A2(n10592), .ZN(n6472) );
  OR2_X1 U9401 ( .A1(n15058), .A2(n7633), .ZN(n6473) );
  NAND2_X2 U9402 ( .A1(n8171), .A2(n8170), .ZN(n8267) );
  INV_X1 U9403 ( .A(n12599), .ZN(n8028) );
  NOR2_X1 U9404 ( .A1(n13379), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U9405 ( .A1(n12350), .A2(n10371), .ZN(n7486) );
  INV_X1 U9406 ( .A(n9001), .ZN(n9162) );
  NAND2_X2 U9407 ( .A1(n14273), .A2(n12630), .ZN(n9166) );
  INV_X1 U9408 ( .A(n8484), .ZN(n7262) );
  INV_X2 U9409 ( .A(n12768), .ZN(n12691) );
  XNOR2_X1 U9410 ( .A(n8180), .B(P1_IR_REG_22__SCAN_IN), .ZN(n12651) );
  XNOR2_X1 U9411 ( .A(n9610), .B(n9609), .ZN(n11869) );
  INV_X1 U9412 ( .A(n11869), .ZN(n7623) );
  INV_X1 U9413 ( .A(n11033), .ZN(n7206) );
  INV_X1 U9414 ( .A(n14868), .ZN(n7955) );
  INV_X1 U9415 ( .A(n14696), .ZN(n7974) );
  INV_X1 U9416 ( .A(n9498), .ZN(n7912) );
  NAND2_X1 U9417 ( .A1(n7434), .A2(n8509), .ZN(n14715) );
  INV_X1 U9418 ( .A(n13935), .ZN(n7743) );
  NOR2_X1 U9419 ( .A1(n7484), .A2(n10370), .ZN(n15068) );
  AND2_X1 U9420 ( .A1(n14288), .A2(n7884), .ZN(n6475) );
  OR2_X1 U9421 ( .A1(n9628), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U9422 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  OR2_X1 U9423 ( .A1(n8844), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6477) );
  NOR2_X1 U9424 ( .A1(n9405), .A2(n9404), .ZN(n9451) );
  AND2_X1 U9425 ( .A1(n14936), .A2(n7639), .ZN(n6478) );
  NAND4_X1 U9426 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n13334) );
  INV_X1 U9427 ( .A(n13334), .ZN(n7457) );
  INV_X1 U9428 ( .A(n6671), .ZN(n8553) );
  NAND2_X1 U9429 ( .A1(n6672), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6671) );
  INV_X1 U9430 ( .A(n15188), .ZN(n15032) );
  NAND2_X1 U9431 ( .A1(n8366), .A2(n8365), .ZN(n15597) );
  INV_X1 U9432 ( .A(n7383), .ZN(n7384) );
  AND2_X1 U9433 ( .A1(n7594), .A2(n7600), .ZN(n6479) );
  NOR2_X1 U9434 ( .A1(n12775), .A2(n12777), .ZN(n7900) );
  AND2_X1 U9435 ( .A1(n12501), .A2(n7820), .ZN(n6480) );
  NAND2_X1 U9436 ( .A1(n8125), .A2(n8124), .ZN(n8592) );
  NOR2_X1 U9437 ( .A1(n11155), .A2(n7134), .ZN(n6481) );
  AND2_X1 U9438 ( .A1(n10013), .A2(n10012), .ZN(n6482) );
  INV_X1 U9439 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13694) );
  OR2_X1 U9440 ( .A1(n9965), .A2(n7163), .ZN(n6483) );
  OR2_X1 U9441 ( .A1(n12519), .A2(n12520), .ZN(n6484) );
  OR2_X1 U9442 ( .A1(n8235), .A2(n10848), .ZN(n6485) );
  AND2_X1 U9443 ( .A1(n10899), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6486) );
  AND2_X1 U9444 ( .A1(n7732), .A2(n9174), .ZN(n6487) );
  AND3_X1 U9445 ( .A1(n7744), .A2(n9478), .A3(n9479), .ZN(n6488) );
  AND2_X1 U9446 ( .A1(n7568), .A2(n7569), .ZN(n6489) );
  XNOR2_X1 U9447 ( .A(n14434), .B(n14256), .ZN(n14236) );
  INV_X1 U9448 ( .A(n14236), .ZN(n6689) );
  OR3_X1 U9449 ( .A1(n13497), .A2(n13479), .A3(n10564), .ZN(n6490) );
  AND2_X1 U9450 ( .A1(n6794), .A2(n7229), .ZN(n14657) );
  AND2_X1 U9451 ( .A1(n15460), .A2(n15408), .ZN(n6491) );
  AND2_X1 U9452 ( .A1(n7307), .A2(n7306), .ZN(n6492) );
  NAND2_X1 U9453 ( .A1(n7709), .A2(n10145), .ZN(n13476) );
  NOR2_X1 U9454 ( .A1(n12404), .A2(n14020), .ZN(n6493) );
  INV_X1 U9455 ( .A(n8087), .ZN(n6688) );
  OR2_X1 U9456 ( .A1(n12802), .A2(n12800), .ZN(n6494) );
  NAND2_X1 U9457 ( .A1(n9705), .A2(n9704), .ZN(n9718) );
  OR2_X1 U9458 ( .A1(n12320), .A2(n6777), .ZN(n6495) );
  INV_X1 U9459 ( .A(n7687), .ZN(n7683) );
  AND2_X1 U9460 ( .A1(n10788), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7687) );
  INV_X1 U9461 ( .A(n11238), .ZN(n10684) );
  NAND2_X1 U9462 ( .A1(n15064), .A2(n14707), .ZN(n6496) );
  AND2_X1 U9463 ( .A1(n14850), .A2(n10395), .ZN(n6497) );
  INV_X1 U9464 ( .A(n7528), .ZN(n7527) );
  INV_X1 U9465 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7777) );
  OR2_X1 U9466 ( .A1(n14186), .A2(n14185), .ZN(n6498) );
  AND2_X1 U9467 ( .A1(n6482), .A2(n12604), .ZN(n6499) );
  INV_X2 U9468 ( .A(n11109), .ZN(n12896) );
  OR2_X1 U9469 ( .A1(n13497), .A2(n13113), .ZN(n6500) );
  INV_X1 U9470 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15364) );
  AND2_X1 U9471 ( .A1(n12604), .A2(n8034), .ZN(n6501) );
  NAND2_X1 U9472 ( .A1(n9430), .A2(n9429), .ZN(n9442) );
  INV_X1 U9473 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U9474 ( .A1(n8946), .A2(n8947), .ZN(n12396) );
  INV_X1 U9475 ( .A(n12396), .ZN(n7888) );
  NAND2_X1 U9476 ( .A1(n8707), .A2(n8706), .ZN(n14723) );
  INV_X1 U9477 ( .A(n14723), .ZN(n7125) );
  INV_X1 U9478 ( .A(n10851), .ZN(n7034) );
  OR2_X1 U9479 ( .A1(n7839), .A2(n12526), .ZN(n6502) );
  AND2_X1 U9480 ( .A1(n12849), .A2(n10334), .ZN(n6503) );
  INV_X1 U9481 ( .A(n10946), .ZN(n6706) );
  NOR4_X1 U9482 ( .A1(n14203), .A2(n14236), .A3(n12619), .A4(n12618), .ZN(
        n6504) );
  NAND2_X1 U9483 ( .A1(n8930), .A2(n8941), .ZN(n14031) );
  AND2_X1 U9484 ( .A1(n9551), .A2(n11363), .ZN(n6505) );
  OR2_X1 U9485 ( .A1(n8735), .A2(n8734), .ZN(n6506) );
  AND2_X1 U9486 ( .A1(n6502), .A2(n12528), .ZN(n6507) );
  INV_X1 U9487 ( .A(n12711), .ZN(n7904) );
  NAND2_X1 U9488 ( .A1(n10961), .A2(n13696), .ZN(n6508) );
  OR2_X1 U9489 ( .A1(n12463), .A2(n6515), .ZN(n6509) );
  INV_X1 U9490 ( .A(n12851), .ZN(n14917) );
  XNOR2_X1 U9491 ( .A(n14724), .B(n14921), .ZN(n12851) );
  OAI211_X1 U9492 ( .C1(n10776), .C2(n8301), .A(n6485), .B(n7242), .ZN(n7244)
         );
  NAND2_X1 U9493 ( .A1(n9985), .A2(n9984), .ZN(n14415) );
  INV_X1 U9494 ( .A(n14415), .ZN(n7894) );
  OR2_X1 U9495 ( .A1(n15058), .A2(n7632), .ZN(n6510) );
  NAND2_X1 U9496 ( .A1(n8480), .A2(n8481), .ZN(n7216) );
  AND2_X1 U9497 ( .A1(n7191), .A2(n7188), .ZN(n6511) );
  NAND2_X1 U9498 ( .A1(n8655), .A2(n8654), .ZN(n14940) );
  AND3_X1 U9499 ( .A1(n13598), .A2(n8148), .A3(n8157), .ZN(n6512) );
  AND2_X1 U9500 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(n8169), .ZN(n6513) );
  AND3_X1 U9501 ( .A1(n9604), .A2(n9602), .A3(n9603), .ZN(n6514) );
  AOI21_X1 U9502 ( .B1(n7675), .B2(n7315), .A(n7313), .ZN(n7673) );
  INV_X1 U9503 ( .A(n7673), .ZN(n7672) );
  NAND2_X1 U9504 ( .A1(n9511), .A2(n11440), .ZN(n9514) );
  INV_X1 U9505 ( .A(n12488), .ZN(n7837) );
  AND2_X1 U9506 ( .A1(n12459), .A2(n12458), .ZN(n6515) );
  NOR2_X1 U9507 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n6516) );
  AND2_X1 U9508 ( .A1(n9716), .A2(n13522), .ZN(n6517) );
  INV_X1 U9509 ( .A(n15234), .ZN(n10064) );
  INV_X1 U9510 ( .A(n12835), .ZN(n11718) );
  AND2_X1 U9511 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6518) );
  AND2_X1 U9512 ( .A1(n14500), .A2(n14012), .ZN(n6519) );
  INV_X1 U9513 ( .A(n15271), .ZN(n14994) );
  NOR2_X1 U9514 ( .A1(n13211), .A2(n6991), .ZN(n6520) );
  NOR2_X1 U9515 ( .A1(n11993), .A2(n7279), .ZN(n6521) );
  AND2_X1 U9516 ( .A1(n6425), .A2(n15759), .ZN(n6522) );
  OR2_X1 U9517 ( .A1(n10848), .A2(n10839), .ZN(n6523) );
  NOR2_X1 U9518 ( .A1(n12201), .A2(n13118), .ZN(n6524) );
  NOR3_X1 U9519 ( .A1(n10432), .A2(n10433), .A3(n10434), .ZN(n6525) );
  OR2_X1 U9520 ( .A1(n11183), .A2(n10842), .ZN(n6526) );
  INV_X1 U9521 ( .A(n10390), .ZN(n7489) );
  INV_X1 U9522 ( .A(n13332), .ZN(n13329) );
  NAND2_X1 U9523 ( .A1(n10577), .A2(n10239), .ZN(n13332) );
  INV_X1 U9524 ( .A(n10124), .ZN(n6836) );
  AND2_X1 U9525 ( .A1(n7409), .A2(n12077), .ZN(n6527) );
  INV_X1 U9526 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8157) );
  AND2_X1 U9527 ( .A1(n10668), .A2(n6997), .ZN(n6528) );
  AND2_X1 U9528 ( .A1(n7397), .A2(n7395), .ZN(n6529) );
  AND2_X1 U9529 ( .A1(n13484), .A2(n13112), .ZN(n6530) );
  NAND2_X1 U9530 ( .A1(n10565), .A2(n10150), .ZN(n10563) );
  INV_X1 U9531 ( .A(n10563), .ZN(n13399) );
  AND2_X1 U9532 ( .A1(n7872), .A2(n7871), .ZN(n6531) );
  AND2_X1 U9533 ( .A1(n9508), .A2(n9507), .ZN(n6532) );
  AND2_X1 U9534 ( .A1(n7497), .A2(n10508), .ZN(n6533) );
  OR2_X1 U9535 ( .A1(n7327), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U9536 ( .A1(n9008), .A2(n9007), .ZN(n6535) );
  AND2_X1 U9537 ( .A1(n7130), .A2(n11238), .ZN(n6536) );
  INV_X1 U9538 ( .A(n14434), .ZN(n14233) );
  NAND2_X1 U9539 ( .A1(n9249), .A2(n9248), .ZN(n14434) );
  AND2_X1 U9540 ( .A1(n6496), .A2(n10371), .ZN(n6537) );
  INV_X1 U9541 ( .A(n14773), .ZN(n7031) );
  AND2_X1 U9542 ( .A1(n7127), .A2(n7560), .ZN(n6538) );
  AND2_X1 U9543 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(n8163), .ZN(n6539) );
  INV_X1 U9544 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15367) );
  NAND2_X1 U9545 ( .A1(n7788), .A2(n6690), .ZN(n10279) );
  INV_X1 U9546 ( .A(n10279), .ZN(n6685) );
  AND2_X1 U9547 ( .A1(n8881), .A2(n8888), .ZN(n6540) );
  INV_X1 U9548 ( .A(n7521), .ZN(n7520) );
  AND2_X1 U9549 ( .A1(n6589), .A2(n8125), .ZN(n7521) );
  NOR2_X1 U9550 ( .A1(n15291), .A2(n14737), .ZN(n6541) );
  NOR2_X1 U9551 ( .A1(n12506), .A2(n12508), .ZN(n6542) );
  INV_X1 U9552 ( .A(n7424), .ZN(n7422) );
  NAND2_X1 U9553 ( .A1(n10895), .A2(n10896), .ZN(n7424) );
  NOR2_X1 U9554 ( .A1(n14495), .A2(n14011), .ZN(n6543) );
  AND2_X1 U9555 ( .A1(n8121), .A2(SI_18_), .ZN(n6544) );
  NOR2_X1 U9556 ( .A1(n14743), .A2(n15580), .ZN(n6545) );
  NOR2_X1 U9557 ( .A1(n14974), .A2(n14726), .ZN(n6546) );
  NOR2_X1 U9558 ( .A1(n14233), .A2(n14007), .ZN(n6547) );
  NOR2_X1 U9559 ( .A1(n14190), .A2(n14196), .ZN(n6548) );
  NOR2_X1 U9560 ( .A1(n13037), .A2(n13457), .ZN(n6549) );
  NOR2_X1 U9561 ( .A1(n14190), .A2(n13979), .ZN(n6550) );
  INV_X1 U9562 ( .A(n11602), .ZN(n11600) );
  OR2_X1 U9563 ( .A1(n8421), .A2(n8420), .ZN(n6551) );
  INV_X1 U9564 ( .A(n12504), .ZN(n7816) );
  INV_X1 U9565 ( .A(n7519), .ZN(n7518) );
  OAI21_X1 U9566 ( .B1(n7523), .B2(n7520), .A(n8619), .ZN(n7519) );
  AND2_X1 U9567 ( .A1(n13452), .A2(n10542), .ZN(n13467) );
  AND2_X1 U9568 ( .A1(n11437), .A2(n11503), .ZN(n6552) );
  INV_X1 U9569 ( .A(n12709), .ZN(n6986) );
  NOR2_X1 U9570 ( .A1(n14807), .A2(n7426), .ZN(n6553) );
  INV_X1 U9571 ( .A(n12492), .ZN(n6749) );
  AND2_X1 U9572 ( .A1(n7968), .A2(n6888), .ZN(n6554) );
  INV_X1 U9573 ( .A(n7662), .ZN(n7661) );
  OAI21_X1 U9574 ( .B1(n7663), .B2(n7665), .A(n13482), .ZN(n7662) );
  NOR2_X1 U9575 ( .A1(n10543), .A2(n10541), .ZN(n6555) );
  AND2_X1 U9576 ( .A1(n8492), .A2(n6804), .ZN(n6556) );
  INV_X1 U9577 ( .A(n7065), .ZN(n7064) );
  NAND2_X1 U9578 ( .A1(n10025), .A2(n7066), .ZN(n7065) );
  INV_X1 U9579 ( .A(n7195), .ZN(n7194) );
  NAND2_X1 U9580 ( .A1(n10039), .A2(n7196), .ZN(n7195) );
  INV_X1 U9581 ( .A(n7404), .ZN(n7403) );
  NAND2_X1 U9582 ( .A1(n7405), .A2(n10342), .ZN(n7404) );
  INV_X1 U9583 ( .A(n7640), .ZN(n7639) );
  NAND2_X1 U9584 ( .A1(n7642), .A2(n7641), .ZN(n7640) );
  INV_X1 U9585 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9419) );
  AND2_X1 U9586 ( .A1(n12710), .A2(n7904), .ZN(n6557) );
  AND2_X1 U9587 ( .A1(n7952), .A2(n7953), .ZN(n6558) );
  NOR2_X1 U9588 ( .A1(n13549), .A2(n7457), .ZN(n6559) );
  OR2_X1 U9589 ( .A1(n7623), .A2(n10690), .ZN(n6560) );
  AND2_X1 U9590 ( .A1(n7746), .A2(n9510), .ZN(n6561) );
  AND2_X1 U9591 ( .A1(n6761), .A2(n9941), .ZN(n6562) );
  OR2_X1 U9592 ( .A1(n8054), .A2(n6544), .ZN(n6563) );
  INV_X1 U9593 ( .A(n7893), .ZN(n7892) );
  NAND2_X1 U9594 ( .A1(n7895), .A2(n7894), .ZN(n7893) );
  AND2_X1 U9595 ( .A1(n10741), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6564) );
  XNOR2_X1 U9596 ( .A(n8633), .B(SI_21_), .ZN(n8631) );
  INV_X1 U9597 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10747) );
  AND2_X1 U9598 ( .A1(n10377), .A2(n6537), .ZN(n6565) );
  AND2_X1 U9599 ( .A1(n10160), .A2(n13104), .ZN(n6566) );
  INV_X1 U9600 ( .A(n14746), .ZN(n7840) );
  AND2_X1 U9601 ( .A1(n10320), .A2(n10319), .ZN(n12842) );
  INV_X1 U9602 ( .A(n12842), .ZN(n7008) );
  AND2_X1 U9603 ( .A1(n6469), .A2(n6902), .ZN(n6567) );
  INV_X1 U9604 ( .A(n7936), .ZN(n7935) );
  OAI21_X1 U9605 ( .B1(n9733), .B2(n7937), .A(n9753), .ZN(n7936) );
  AND2_X1 U9606 ( .A1(n10745), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6568) );
  AND2_X1 U9607 ( .A1(n10799), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U9608 ( .A1(n13553), .A2(n13350), .ZN(n6570) );
  INV_X1 U9609 ( .A(n6978), .ZN(n6977) );
  NAND2_X1 U9610 ( .A1(n6979), .A2(n6695), .ZN(n6978) );
  NAND2_X1 U9611 ( .A1(n7972), .A2(n6506), .ZN(n6571) );
  NAND2_X1 U9612 ( .A1(n9533), .A2(n10793), .ZN(n6572) );
  OAI21_X1 U9613 ( .B1(n7989), .B2(n7987), .A(n8630), .ZN(n7986) );
  OAI21_X1 U9614 ( .B1(n12806), .B2(n12807), .A(n7448), .ZN(n7447) );
  OAI21_X1 U9615 ( .B1(n10028), .B2(n8007), .A(n12591), .ZN(n8006) );
  INV_X1 U9616 ( .A(n7574), .ZN(n7573) );
  OAI21_X1 U9617 ( .B1(n13154), .B2(n13155), .A(n7576), .ZN(n7574) );
  INV_X1 U9618 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U9619 ( .A1(n8568), .A2(n8117), .ZN(n6573) );
  AND2_X1 U9620 ( .A1(n10351), .A2(n10350), .ZN(n6574) );
  AND2_X1 U9621 ( .A1(n7623), .A2(n7622), .ZN(n6575) );
  NOR2_X1 U9622 ( .A1(n11135), .A2(n11136), .ZN(n6576) );
  AND2_X1 U9623 ( .A1(n7563), .A2(n6437), .ZN(n6577) );
  OR2_X1 U9624 ( .A1(n12799), .A2(n12797), .ZN(n6578) );
  AOI21_X1 U9625 ( .B1(n12525), .B2(n12522), .A(n12521), .ZN(n12523) );
  OR2_X1 U9626 ( .A1(n7904), .A2(n12710), .ZN(n6579) );
  OR2_X1 U9627 ( .A1(n8039), .A2(n8545), .ZN(n6580) );
  AND2_X1 U9628 ( .A1(n8938), .A2(n8937), .ZN(n6581) );
  INV_X1 U9629 ( .A(n7407), .ZN(n7406) );
  NOR2_X1 U9630 ( .A1(n10343), .A2(n7408), .ZN(n7407) );
  AND2_X1 U9631 ( .A1(n10427), .A2(n10426), .ZN(n10586) );
  INV_X1 U9632 ( .A(n10224), .ZN(n10440) );
  OR2_X1 U9633 ( .A1(n14967), .A2(n7857), .ZN(n6582) );
  NAND2_X1 U9634 ( .A1(n7423), .A2(n7419), .ZN(n6583) );
  INV_X1 U9635 ( .A(n12795), .ZN(n7438) );
  NAND2_X1 U9636 ( .A1(n7507), .A2(n7508), .ZN(n13387) );
  NAND2_X1 U9637 ( .A1(n8940), .A2(n10071), .ZN(n8926) );
  AND2_X1 U9638 ( .A1(n13477), .A2(n6441), .ZN(n6584) );
  AND3_X1 U9639 ( .A1(n7600), .A2(n11343), .A3(n11026), .ZN(n6585) );
  INV_X1 U9640 ( .A(n12796), .ZN(n7437) );
  AND2_X1 U9641 ( .A1(n10566), .A2(n10567), .ZN(n6586) );
  AND2_X1 U9642 ( .A1(n14537), .A2(n14008), .ZN(n6587) );
  AND2_X1 U9643 ( .A1(n12898), .A2(n13074), .ZN(n6588) );
  NOR2_X1 U9644 ( .A1(n15105), .A2(n15525), .ZN(n12826) );
  OR2_X1 U9645 ( .A1(n8618), .A2(SI_20_), .ZN(n6589) );
  AND3_X1 U9646 ( .A1(n12595), .A2(n12594), .A3(n6767), .ZN(n6590) );
  NOR2_X1 U9647 ( .A1(n14921), .A2(n14724), .ZN(n6591) );
  NAND2_X1 U9648 ( .A1(n14288), .A2(n6859), .ZN(n6861) );
  AND2_X1 U9649 ( .A1(n7291), .A2(n10170), .ZN(n6592) );
  INV_X1 U9650 ( .A(n14308), .ZN(n14456) );
  AND2_X1 U9651 ( .A1(n9206), .A2(n9205), .ZN(n14308) );
  NOR2_X1 U9652 ( .A1(n12949), .A2(n7764), .ZN(n6593) );
  INV_X1 U9653 ( .A(n6895), .ZN(n11883) );
  AND2_X1 U9654 ( .A1(n9974), .A2(n9972), .ZN(n14266) );
  INV_X1 U9655 ( .A(n14266), .ZN(n7386) );
  AND2_X1 U9656 ( .A1(n12209), .A2(n7939), .ZN(n6594) );
  NAND2_X1 U9657 ( .A1(n7246), .A2(n6997), .ZN(n10614) );
  INV_X1 U9658 ( .A(n10614), .ZN(n7129) );
  NOR2_X1 U9659 ( .A1(n7204), .A2(n10976), .ZN(n6595) );
  NOR2_X1 U9660 ( .A1(n7803), .A2(n7802), .ZN(n6596) );
  AND2_X1 U9661 ( .A1(n15381), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6597) );
  OR2_X1 U9662 ( .A1(n11183), .A2(n10853), .ZN(n6598) );
  OR2_X1 U9663 ( .A1(n12530), .A2(n7823), .ZN(n6599) );
  AND2_X1 U9664 ( .A1(n13827), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n6600) );
  AND2_X1 U9665 ( .A1(n7953), .A2(n14831), .ZN(n6601) );
  NOR2_X1 U9666 ( .A1(n6455), .A2(n7065), .ZN(n7061) );
  AND2_X1 U9667 ( .A1(n12530), .A2(n7823), .ZN(n6602) );
  INV_X1 U9668 ( .A(n15286), .ZN(n12738) );
  AND2_X1 U9669 ( .A1(n8469), .A2(n8468), .ZN(n15286) );
  INV_X1 U9670 ( .A(n14086), .ZN(n6719) );
  OR2_X1 U9671 ( .A1(n7733), .A2(n7731), .ZN(n6603) );
  AND2_X1 U9672 ( .A1(n8146), .A2(n6512), .ZN(n6604) );
  AND2_X1 U9673 ( .A1(n7684), .A2(n7683), .ZN(n6605) );
  AND2_X1 U9674 ( .A1(n7527), .A2(n10972), .ZN(n6606) );
  AND2_X1 U9675 ( .A1(n6487), .A2(n12361), .ZN(n6607) );
  NAND3_X1 U9676 ( .A1(n12742), .A2(n12741), .A3(n12740), .ZN(n6608) );
  INV_X1 U9677 ( .A(n7747), .ZN(n7285) );
  NOR2_X1 U9678 ( .A1(n7748), .A2(n6524), .ZN(n7747) );
  AND2_X1 U9679 ( .A1(n8884), .A2(n8864), .ZN(n8912) );
  AND2_X1 U9680 ( .A1(n7444), .A2(n7443), .ZN(n6609) );
  NOR2_X1 U9681 ( .A1(n7675), .A2(n7676), .ZN(n7674) );
  AND2_X1 U9682 ( .A1(n12678), .A2(n8052), .ZN(n6610) );
  AND2_X1 U9683 ( .A1(n12759), .A2(n12758), .ZN(n6611) );
  AND2_X1 U9684 ( .A1(n7832), .A2(n12466), .ZN(n6612) );
  INV_X1 U9685 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U9686 ( .A1(n12580), .A2(n6599), .ZN(n6613) );
  OR2_X1 U9687 ( .A1(n13411), .A2(n13419), .ZN(n10565) );
  AND2_X1 U9688 ( .A1(n12891), .A2(n12894), .ZN(n6614) );
  AND2_X1 U9689 ( .A1(n6481), .A2(n10791), .ZN(n6615) );
  INV_X1 U9690 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10741) );
  INV_X1 U9691 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8161) );
  INV_X1 U9692 ( .A(n6429), .ZN(n7213) );
  INV_X1 U9693 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U9694 ( .A1(n12785), .A2(n6973), .ZN(n6616) );
  INV_X1 U9695 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8184) );
  INV_X1 U9696 ( .A(n10219), .ZN(n10220) );
  INV_X1 U9697 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8185) );
  INV_X1 U9698 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10743) );
  AND2_X2 U9699 ( .A1(n10254), .A2(n11312), .ZN(n15873) );
  AND2_X2 U9700 ( .A1(n10046), .A2(n14385), .ZN(n14352) );
  INV_X1 U9701 ( .A(n8292), .ZN(n8643) );
  AND2_X2 U9702 ( .A1(n10264), .A2(n10263), .ZN(n15860) );
  INV_X1 U9703 ( .A(n15045), .ZN(n7636) );
  INV_X1 U9704 ( .A(n14903), .ZN(n7641) );
  AND2_X1 U9705 ( .A1(n10914), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n6618) );
  INV_X1 U9706 ( .A(n10697), .ZN(n6997) );
  INV_X1 U9707 ( .A(n9918), .ZN(n10564) );
  AND2_X1 U9708 ( .A1(n9444), .A2(n9443), .ZN(n13817) );
  INV_X1 U9709 ( .A(n13879), .ZN(n6782) );
  NAND2_X1 U9710 ( .A1(n13197), .A2(n6520), .ZN(n6992) );
  OR2_X1 U9711 ( .A1(n15423), .A2(n15424), .ZN(n7336) );
  NAND2_X1 U9712 ( .A1(n12168), .A2(n6438), .ZN(n12313) );
  AND2_X1 U9713 ( .A1(n11762), .A2(n11896), .ZN(n11763) );
  NAND2_X1 U9714 ( .A1(n15782), .A2(n10440), .ZN(n11435) );
  OR2_X1 U9715 ( .A1(n12163), .A2(n7962), .ZN(n12179) );
  AND2_X1 U9716 ( .A1(n6468), .A2(n7144), .ZN(n6619) );
  AND2_X1 U9717 ( .A1(n9821), .A2(n9817), .ZN(n6620) );
  NAND2_X1 U9718 ( .A1(n8673), .A2(SI_23_), .ZN(n6621) );
  INV_X1 U9719 ( .A(n11925), .ZN(n7400) );
  OAI21_X1 U9720 ( .B1(n12996), .B2(n6916), .A(n6914), .ZN(n13016) );
  AND2_X1 U9721 ( .A1(n7312), .A2(n7311), .ZN(n6622) );
  NAND2_X1 U9722 ( .A1(n7475), .A2(n7474), .ZN(n15506) );
  OAI21_X1 U9723 ( .B1(n11878), .B2(n10233), .A(n10232), .ZN(n11971) );
  NAND2_X1 U9724 ( .A1(n6849), .A2(n10141), .ZN(n13518) );
  NAND2_X1 U9725 ( .A1(n6663), .A2(n7949), .ZN(n11951) );
  NAND2_X1 U9726 ( .A1(n10143), .A2(n10142), .ZN(n13503) );
  INV_X1 U9727 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7749) );
  INV_X1 U9728 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7134) );
  INV_X1 U9729 ( .A(n6917), .ZN(n12958) );
  NAND2_X1 U9730 ( .A1(n12996), .A2(n9656), .ZN(n6917) );
  INV_X1 U9731 ( .A(n8692), .ZN(n8693) );
  NAND2_X1 U9732 ( .A1(n10165), .A2(n10164), .ZN(n13553) );
  INV_X1 U9733 ( .A(n13553), .ZN(n7369) );
  NAND2_X1 U9734 ( .A1(n8183), .A2(n7490), .ZN(n8528) );
  INV_X1 U9735 ( .A(n10665), .ZN(n7247) );
  AND2_X1 U9736 ( .A1(n10191), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n6623) );
  OR2_X1 U9737 ( .A1(n15785), .A2(n6903), .ZN(n6624) );
  NAND2_X1 U9738 ( .A1(n7967), .A2(n10310), .ZN(n11717) );
  AOI21_X1 U9739 ( .B1(n7455), .B2(n9717), .A(n7936), .ZN(n7454) );
  INV_X1 U9740 ( .A(n7896), .ZN(n9082) );
  NOR2_X1 U9741 ( .A1(n12162), .A2(n12837), .ZN(n12163) );
  AND2_X1 U9742 ( .A1(n11789), .A2(n6726), .ZN(n6625) );
  INV_X1 U9743 ( .A(n7537), .ZN(n7536) );
  NOR2_X1 U9744 ( .A1(n9982), .A2(n7538), .ZN(n7537) );
  AND2_X1 U9745 ( .A1(n8445), .A2(n8444), .ZN(n11285) );
  INV_X1 U9746 ( .A(n11285), .ZN(n7019) );
  NAND2_X1 U9747 ( .A1(n7629), .A2(n7630), .ZN(n7631) );
  NAND2_X1 U9748 ( .A1(n11763), .A2(n6427), .ZN(n7887) );
  INV_X1 U9749 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6676) );
  INV_X1 U9750 ( .A(n9959), .ZN(n7786) );
  AND2_X1 U9751 ( .A1(n7769), .A2(n7767), .ZN(n6626) );
  AND2_X1 U9752 ( .A1(n8695), .A2(SI_24_), .ZN(n6627) );
  NOR2_X1 U9753 ( .A1(n13767), .A2(n13815), .ZN(n6628) );
  NAND2_X1 U9754 ( .A1(n8850), .A2(n9132), .ZN(n6629) );
  AND2_X1 U9755 ( .A1(n11306), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6630) );
  AND2_X1 U9756 ( .A1(n9768), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n6631) );
  INV_X1 U9757 ( .A(n7451), .ZN(n7450) );
  OAI21_X1 U9758 ( .B1(n6620), .B2(n7452), .A(n9841), .ZN(n7451) );
  OR2_X1 U9759 ( .A1(n10086), .A2(n10082), .ZN(n6632) );
  OR2_X1 U9760 ( .A1(n13767), .A2(n13750), .ZN(n6633) );
  OR2_X1 U9761 ( .A1(n13030), .A2(n6903), .ZN(n6634) );
  NAND2_X1 U9762 ( .A1(n8844), .A2(n8846), .ZN(n12626) );
  NOR2_X1 U9763 ( .A1(n15873), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6635) );
  AND2_X1 U9764 ( .A1(n12094), .A2(n10525), .ZN(n6636) );
  INV_X1 U9765 ( .A(SI_14_), .ZN(n10972) );
  AND2_X1 U9766 ( .A1(n9836), .A2(n9852), .ZN(n6637) );
  OR2_X1 U9767 ( .A1(n13778), .A2(n7648), .ZN(n6638) );
  INV_X1 U9768 ( .A(n7269), .ZN(n11693) );
  AND2_X1 U9769 ( .A1(n13003), .A2(n9866), .ZN(n9873) );
  NAND2_X1 U9770 ( .A1(n10935), .A2(n7046), .ZN(n7045) );
  INV_X1 U9771 ( .A(n15801), .ZN(n15789) );
  NAND2_X1 U9772 ( .A1(n9646), .A2(n9645), .ZN(n12201) );
  INV_X1 U9773 ( .A(n12201), .ZN(n7110) );
  NAND2_X1 U9774 ( .A1(n9711), .A2(n9710), .ZN(n13510) );
  INV_X1 U9775 ( .A(n13510), .ZN(n7713) );
  INV_X1 U9776 ( .A(n13999), .ZN(n6858) );
  INV_X1 U9777 ( .A(n14379), .ZN(n14302) );
  NOR2_X1 U9778 ( .A1(n10887), .A2(n10723), .ZN(n15479) );
  XNOR2_X1 U9779 ( .A(n10313), .B(n15242), .ZN(n12837) );
  INV_X1 U9780 ( .A(n12837), .ZN(n7011) );
  NAND2_X1 U9781 ( .A1(n10347), .A2(n10346), .ZN(n15604) );
  NAND2_X1 U9782 ( .A1(n6522), .A2(n11643), .ZN(n6639) );
  NAND2_X1 U9783 ( .A1(n11647), .A2(n12598), .ZN(n11587) );
  AND2_X1 U9784 ( .A1(n9851), .A2(n9850), .ZN(n13419) );
  AND2_X2 U9785 ( .A1(n10295), .A2(n15721), .ZN(n15767) );
  AND2_X1 U9786 ( .A1(n9909), .A2(n10263), .ZN(n13074) );
  INV_X1 U9787 ( .A(n13074), .ZN(n13100) );
  OR2_X1 U9788 ( .A1(n15606), .A2(n13655), .ZN(n6640) );
  INV_X1 U9789 ( .A(n15778), .ZN(n15775) );
  AND2_X2 U9790 ( .A1(n10295), .A2(n10289), .ZN(n15778) );
  NAND2_X1 U9791 ( .A1(n9087), .A2(n9086), .ZN(n14500) );
  INV_X1 U9792 ( .A(n14500), .ZN(n7885) );
  INV_X1 U9793 ( .A(n11662), .ZN(n10003) );
  INV_X1 U9794 ( .A(n13307), .ZN(n7561) );
  INV_X1 U9795 ( .A(n9836), .ZN(n7452) );
  NAND2_X1 U9796 ( .A1(n7723), .A2(n7727), .ZN(n13959) );
  NAND2_X1 U9797 ( .A1(n9834), .A2(n9833), .ZN(n13107) );
  INV_X1 U9798 ( .A(n13107), .ZN(n13401) );
  AND2_X1 U9799 ( .A1(n7600), .A2(n11026), .ZN(n6641) );
  NOR2_X1 U9800 ( .A1(n10944), .A2(n6486), .ZN(n6642) );
  OR2_X1 U9801 ( .A1(n14781), .A2(n14780), .ZN(n6643) );
  AND2_X1 U9802 ( .A1(n7320), .A2(n11363), .ZN(n6644) );
  OR2_X1 U9803 ( .A1(n14797), .A2(n15047), .ZN(n6645) );
  NAND2_X1 U9804 ( .A1(n8360), .A2(n8359), .ZN(n6646) );
  INV_X1 U9805 ( .A(n13419), .ZN(n13106) );
  AND2_X1 U9806 ( .A1(n7722), .A2(n7727), .ZN(n6647) );
  NAND2_X1 U9807 ( .A1(n8343), .A2(n8342), .ZN(n6648) );
  NAND2_X1 U9808 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6649) );
  AND2_X1 U9809 ( .A1(n12947), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6650) );
  AND2_X1 U9810 ( .A1(n7431), .A2(n14820), .ZN(n6651) );
  INV_X1 U9811 ( .A(n11066), .ZN(n6718) );
  INV_X1 U9812 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15339) );
  OR2_X1 U9813 ( .A1(n15618), .A2(n8807), .ZN(n6652) );
  AND2_X1 U9814 ( .A1(n7075), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6653) );
  OR2_X1 U9815 ( .A1(n10615), .A2(n10976), .ZN(n6654) );
  NAND2_X1 U9816 ( .A1(n12283), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U9817 ( .A1(n10203), .A2(n7948), .ZN(n7947) );
  AND2_X1 U9818 ( .A1(n6470), .A2(n7561), .ZN(n6656) );
  AND2_X1 U9819 ( .A1(n7572), .A2(n7575), .ZN(n6657) );
  INV_X1 U9820 ( .A(n8043), .ZN(n7763) );
  INV_X1 U9821 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7363) );
  OR2_X1 U9822 ( .A1(n11490), .A2(n10654), .ZN(n6658) );
  OR2_X1 U9823 ( .A1(n6706), .A2(n12010), .ZN(n6659) );
  INV_X1 U9824 ( .A(n8171), .ZN(n8172) );
  NAND2_X1 U9825 ( .A1(n7029), .A2(n7027), .ZN(n6660) );
  AND2_X1 U9826 ( .A1(n7147), .A2(n7682), .ZN(n6661) );
  AND2_X1 U9827 ( .A1(n7753), .A2(n6852), .ZN(n13819) );
  INV_X1 U9828 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n7300) );
  INV_X1 U9829 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7036) );
  INV_X1 U9830 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7399) );
  INV_X1 U9831 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7745) );
  INV_X1 U9832 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7877) );
  INV_X1 U9833 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6955) );
  INV_X1 U9834 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6891) );
  INV_X1 U9835 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7798) );
  INV_X1 U9836 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n7706) );
  AOI22_X1 U9837 ( .A1(n14196), .A2(n14374), .B1(n14376), .B2(n14226), .ZN(
        n7347) );
  INV_X1 U9838 ( .A(n14374), .ZN(n14331) );
  NAND2_X1 U9839 ( .A1(n12307), .A2(n10320), .ZN(n12346) );
  AND2_X2 U9840 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  NAND2_X2 U9841 ( .A1(n6662), .A2(n14967), .ZN(n14970) );
  NAND2_X1 U9842 ( .A1(n14966), .A2(n14968), .ZN(n6662) );
  NAND2_X1 U9843 ( .A1(n11951), .A2(n12833), .ZN(n10308) );
  NAND2_X1 U9844 ( .A1(n7176), .A2(n10304), .ZN(n6663) );
  NAND4_X1 U9845 ( .A1(n8183), .A2(n8141), .A3(n6604), .A4(n8138), .ZN(n6664)
         );
  NAND2_X2 U9846 ( .A1(n12162), .A2(n7961), .ZN(n7958) );
  NAND2_X1 U9847 ( .A1(n11947), .A2(n12834), .ZN(n7967) );
  NAND3_X1 U9848 ( .A1(n6667), .A2(n6666), .A3(n7126), .ZN(n6665) );
  INV_X1 U9849 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U9850 ( .A1(n9975), .A2(n7807), .ZN(n6681) );
  OAI21_X2 U9851 ( .B1(n7122), .B2(n6691), .A(n7120), .ZN(n8593) );
  OAI211_X2 U9852 ( .C1(n8384), .C2(n6688), .A(n6687), .B(n8088), .ZN(n8091)
         );
  OR2_X2 U9853 ( .A1(n10279), .A2(n10270), .ZN(n10280) );
  OAI21_X1 U9854 ( .B1(n6691), .B2(n8003), .A(n6416), .ZN(n8569) );
  OAI21_X1 U9855 ( .B1(n6691), .B2(n8522), .A(n8521), .ZN(n8524) );
  XNOR2_X2 U9856 ( .A(n8650), .B(SI_22_), .ZN(n9218) );
  OAI21_X1 U9857 ( .B1(n6694), .B2(n12805), .A(n7445), .ZN(n6693) );
  INV_X1 U9858 ( .A(n12808), .ZN(n6695) );
  NAND2_X1 U9859 ( .A1(n12781), .A2(n12780), .ZN(n6697) );
  INV_X1 U9860 ( .A(n12781), .ZN(n6698) );
  NAND3_X1 U9861 ( .A1(n12767), .A2(n12766), .A3(n6702), .ZN(n6701) );
  NAND2_X1 U9862 ( .A1(n6611), .A2(n12755), .ZN(n6702) );
  AND2_X1 U9863 ( .A1(n15041), .A2(n12750), .ZN(n12755) );
  NAND3_X1 U9864 ( .A1(n12793), .A2(n7435), .A3(n12794), .ZN(n6704) );
  NAND2_X2 U9865 ( .A1(n14947), .A2(n10335), .ZN(n14929) );
  OAI21_X1 U9866 ( .B1(n10840), .B2(n8254), .A(n14757), .ZN(n14770) );
  NAND3_X1 U9867 ( .A1(n6716), .A2(n6715), .A3(n6712), .ZN(n15663) );
  NAND3_X1 U9868 ( .A1(n6713), .A2(n11067), .A3(n14086), .ZN(n6712) );
  NOR2_X1 U9869 ( .A1(n14162), .A2(n14161), .ZN(n14163) );
  NAND2_X1 U9870 ( .A1(n14159), .A2(n14158), .ZN(n6727) );
  NAND3_X1 U9871 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U9872 ( .B1(n6733), .B2(n12457), .A(n6509), .ZN(n6732) );
  OAI21_X1 U9873 ( .B1(n12452), .B2(n12451), .A(n12450), .ZN(n6733) );
  NAND2_X1 U9874 ( .A1(n6734), .A2(n7821), .ZN(n7541) );
  NAND3_X1 U9875 ( .A1(n6737), .A2(n6736), .A3(n6735), .ZN(n6734) );
  NAND2_X1 U9876 ( .A1(n6743), .A2(n6738), .ZN(n6735) );
  NAND2_X1 U9877 ( .A1(n6741), .A2(n6740), .ZN(n6737) );
  NAND2_X1 U9878 ( .A1(n6428), .A2(n6502), .ZN(n6741) );
  INV_X1 U9879 ( .A(n12528), .ZN(n6742) );
  NAND2_X1 U9880 ( .A1(n6745), .A2(n6744), .ZN(n12498) );
  NAND2_X1 U9881 ( .A1(n6748), .A2(n12499), .ZN(n12500) );
  OAI21_X1 U9882 ( .B1(n6750), .B2(n12436), .A(n12435), .ZN(n12437) );
  NAND4_X1 U9883 ( .A1(n12415), .A2(n6753), .A3(n6752), .A4(n12414), .ZN(n6751) );
  OR2_X1 U9884 ( .A1(n12413), .A2(n12412), .ZN(n6753) );
  INV_X1 U9885 ( .A(n12509), .ZN(n12512) );
  NAND2_X2 U9886 ( .A1(n8940), .A2(n10769), .ZN(n9191) );
  NAND2_X2 U9887 ( .A1(n8883), .A2(n8887), .ZN(n11054) );
  NAND2_X1 U9888 ( .A1(n11590), .A2(n6759), .ZN(n11591) );
  NAND2_X1 U9889 ( .A1(n7801), .A2(n7799), .ZN(n6759) );
  NAND3_X1 U9890 ( .A1(n9932), .A2(n11577), .A3(n9933), .ZN(n11576) );
  INV_X1 U9891 ( .A(n11577), .ZN(n6766) );
  NAND2_X1 U9892 ( .A1(n9932), .A2(n9933), .ZN(n6768) );
  NAND2_X1 U9893 ( .A1(n6764), .A2(n10002), .ZN(n11640) );
  NAND2_X1 U9894 ( .A1(n6768), .A2(n11662), .ZN(n6764) );
  NAND2_X1 U9895 ( .A1(n11576), .A2(n6765), .ZN(n11582) );
  NAND2_X1 U9896 ( .A1(n6766), .A2(n6768), .ZN(n6765) );
  NOR2_X1 U9897 ( .A1(n6768), .A2(n12626), .ZN(n6767) );
  XNOR2_X1 U9898 ( .A(n6768), .B(n10003), .ZN(n15736) );
  NAND2_X1 U9899 ( .A1(n8219), .A2(n9009), .ZN(n6769) );
  OR2_X2 U9900 ( .A1(n14261), .A2(n7386), .ZN(n14263) );
  NAND2_X1 U9902 ( .A1(n7724), .A2(n7721), .ZN(n7723) );
  NAND2_X1 U9903 ( .A1(n11325), .A2(n8958), .ZN(n11384) );
  NAND2_X1 U9904 ( .A1(n6774), .A2(n6775), .ZN(n12362) );
  NAND2_X1 U9905 ( .A1(n12362), .A2(n6607), .ZN(n7280) );
  INV_X1 U9906 ( .A(n13852), .ZN(n6779) );
  INV_X1 U9908 ( .A(n13944), .ZN(n13850) );
  INV_X1 U9909 ( .A(n13851), .ZN(n6783) );
  NAND2_X1 U9910 ( .A1(n12550), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8886) );
  NAND3_X1 U9911 ( .A1(n7481), .A2(n10378), .A3(n6787), .ZN(n15037) );
  NAND2_X2 U9912 ( .A1(n6788), .A2(n8446), .ZN(n15291) );
  NAND2_X1 U9913 ( .A1(n6789), .A2(n6652), .ZN(P1_U3557) );
  NAND2_X1 U9914 ( .A1(n15250), .A2(n15618), .ZN(n6789) );
  NAND2_X1 U9915 ( .A1(n6790), .A2(n6925), .ZN(n15250) );
  NAND2_X1 U9916 ( .A1(n15133), .A2(n15572), .ZN(n6790) );
  NAND3_X1 U9917 ( .A1(n8091), .A2(n7996), .A3(n7527), .ZN(n6797) );
  NAND3_X1 U9918 ( .A1(n8091), .A2(n7996), .A3(n6606), .ZN(n6795) );
  NAND2_X1 U9919 ( .A1(n8091), .A2(n7996), .ZN(n7992) );
  NAND3_X1 U9920 ( .A1(n6799), .A2(n6797), .A3(SI_14_), .ZN(n6798) );
  OAI21_X1 U9921 ( .B1(n7198), .B2(n6802), .A(n6800), .ZN(n6803) );
  INV_X1 U9922 ( .A(n8691), .ZN(n6801) );
  NAND2_X1 U9923 ( .A1(n14618), .A2(n7970), .ZN(n7969) );
  NAND2_X1 U9924 ( .A1(n6803), .A2(n14574), .ZN(n8834) );
  XNOR2_X1 U9925 ( .A(n6805), .B(n10397), .ZN(n8495) );
  NAND3_X1 U9926 ( .A1(n7977), .A2(n7216), .A3(n7215), .ZN(n6806) );
  NAND2_X1 U9927 ( .A1(n6817), .A2(n6815), .ZN(n6814) );
  NAND2_X1 U9928 ( .A1(n6819), .A2(n6814), .ZN(n6818) );
  NAND2_X1 U9929 ( .A1(n6818), .A2(n7460), .ZN(n7927) );
  NAND3_X1 U9930 ( .A1(n10565), .A2(n10150), .A3(n7509), .ZN(n6828) );
  NAND2_X1 U9931 ( .A1(n10123), .A2(n6830), .ZN(n6832) );
  INV_X1 U9932 ( .A(n10122), .ZN(n6831) );
  NAND2_X1 U9933 ( .A1(n6832), .A2(n6833), .ZN(n11442) );
  NAND2_X1 U9934 ( .A1(n6552), .A2(n11442), .ZN(n6835) );
  NAND2_X1 U9935 ( .A1(n6835), .A2(n6834), .ZN(n11401) );
  NAND2_X2 U9936 ( .A1(n6838), .A2(n6839), .ZN(n13127) );
  NAND3_X1 U9937 ( .A1(n6461), .A2(n6857), .A3(n12248), .ZN(n14381) );
  INV_X1 U9938 ( .A(n6861), .ZN(n14197) );
  NAND2_X2 U9939 ( .A1(n12936), .A2(n10281), .ZN(n7158) );
  NAND3_X1 U9940 ( .A1(n7861), .A2(n15450), .A3(n6463), .ZN(n6863) );
  AND2_X2 U9941 ( .A1(n6863), .A2(n6862), .ZN(n15459) );
  INV_X1 U9942 ( .A(n15459), .ZN(n7357) );
  NOR2_X2 U9943 ( .A1(n15420), .A2(n15421), .ZN(n15419) );
  NAND3_X1 U9944 ( .A1(n6865), .A2(n6868), .A3(n6866), .ZN(n15420) );
  NAND2_X1 U9945 ( .A1(n15876), .A2(n6597), .ZN(n6865) );
  NAND2_X1 U9946 ( .A1(n15878), .A2(n15877), .ZN(n15876) );
  NAND2_X1 U9947 ( .A1(n15878), .A2(n6867), .ZN(n6866) );
  NAND2_X1 U9948 ( .A1(n15876), .A2(n15381), .ZN(n15383) );
  NAND2_X1 U9949 ( .A1(n6869), .A2(n15382), .ZN(n6868) );
  INV_X1 U9950 ( .A(n15381), .ZN(n6869) );
  NAND2_X1 U9951 ( .A1(n15366), .A2(n7328), .ZN(n7326) );
  NAND2_X1 U9952 ( .A1(n7324), .A2(n7326), .ZN(n6871) );
  NAND2_X1 U9953 ( .A1(n6873), .A2(n15366), .ZN(n6872) );
  NAND3_X1 U9954 ( .A1(n15435), .A2(n15433), .A3(n6875), .ZN(n7339) );
  INV_X1 U9955 ( .A(n7339), .ZN(n6874) );
  INV_X1 U9956 ( .A(n15438), .ZN(n6876) );
  NAND2_X1 U9957 ( .A1(n7335), .A2(n15425), .ZN(n15430) );
  NAND3_X1 U9958 ( .A1(n6877), .A2(n15429), .A3(n15400), .ZN(n15448) );
  NAND3_X1 U9959 ( .A1(n7335), .A2(n15425), .A3(n6879), .ZN(n6878) );
  XNOR2_X2 U9960 ( .A(n6880), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8170) );
  OR2_X2 U9961 ( .A1(n8168), .A2(n15296), .ZN(n6880) );
  AND4_X2 U9962 ( .A1(n7491), .A2(n6881), .A3(n6604), .A4(n7490), .ZN(n8168)
         );
  NAND2_X1 U9963 ( .A1(n10337), .A2(n7180), .ZN(n14914) );
  NAND2_X2 U9964 ( .A1(n12929), .A2(n8172), .ZN(n6892) );
  XNOR2_X2 U9965 ( .A(n7316), .B(P3_IR_REG_29__SCAN_IN), .ZN(n6893) );
  NAND3_X1 U9966 ( .A1(n6893), .A2(n9413), .A3(P3_REG3_REG_0__SCAN_IN), .ZN(
        n9463) );
  NAND2_X1 U9967 ( .A1(n13516), .A2(n6899), .ZN(n6896) );
  NAND2_X1 U9968 ( .A1(n6896), .A2(n6897), .ZN(n13496) );
  NAND3_X1 U9969 ( .A1(n11988), .A2(n11987), .A3(n6634), .ZN(n11989) );
  XNOR2_X1 U9970 ( .A(n10405), .B(n10240), .ZN(n12926) );
  AOI21_X1 U9971 ( .B1(n12926), .B2(n15851), .A(n10220), .ZN(n7729) );
  NAND3_X1 U9972 ( .A1(n7729), .A2(n7510), .A3(n15873), .ZN(n7728) );
  NAND3_X1 U9973 ( .A1(n6907), .A2(n6905), .A3(n7364), .ZN(P3_U3169) );
  NAND2_X1 U9974 ( .A1(n6908), .A2(n6906), .ZN(n6905) );
  NAND2_X1 U9975 ( .A1(n6908), .A2(n6911), .ZN(n6907) );
  INV_X1 U9976 ( .A(n13007), .ZN(n6912) );
  NAND2_X1 U9977 ( .A1(n6460), .A2(n7756), .ZN(n7757) );
  NAND2_X2 U9978 ( .A1(n12975), .A2(n9780), .ZN(n13034) );
  NAND2_X2 U9979 ( .A1(n7760), .A2(n7758), .ZN(n12973) );
  OR2_X2 U9980 ( .A1(n9870), .A2(n9871), .ZN(n7365) );
  NAND2_X2 U9981 ( .A1(n12982), .A2(n9814), .ZN(n9870) );
  NAND2_X2 U9982 ( .A1(n7776), .A2(n7775), .ZN(n12982) );
  NAND2_X2 U9983 ( .A1(n12915), .A2(n13831), .ZN(n9422) );
  NAND2_X4 U9984 ( .A1(n7343), .A2(n7609), .ZN(n13831) );
  XNOR2_X2 U9985 ( .A(n6913), .B(n9418), .ZN(n12915) );
  NAND2_X4 U9986 ( .A1(n9455), .A2(n9454), .ZN(n11109) );
  NAND2_X1 U9987 ( .A1(n9585), .A2(n7770), .ZN(n12038) );
  OAI21_X1 U9988 ( .B1(n9585), .B2(n6921), .A(n6919), .ZN(n6922) );
  INV_X1 U9989 ( .A(n6920), .ZN(n6919) );
  OAI21_X1 U9990 ( .B1(n6921), .B2(n7770), .A(n9638), .ZN(n6920) );
  NAND2_X1 U9991 ( .A1(n12038), .A2(n9621), .ZN(n11983) );
  NAND2_X2 U9992 ( .A1(n9654), .A2(n12994), .ZN(n12996) );
  NAND2_X1 U9993 ( .A1(n11745), .A2(n11746), .ZN(n9585) );
  NAND2_X1 U9994 ( .A1(n11396), .A2(n10488), .ZN(n11612) );
  NAND3_X1 U9995 ( .A1(n7105), .A2(n7498), .A3(n6594), .ZN(n7107) );
  NAND2_X1 U9996 ( .A1(n11063), .A2(n11062), .ZN(n14068) );
  NAND2_X1 U9997 ( .A1(n14158), .A2(n14137), .ZN(n14139) );
  INV_X1 U9998 ( .A(n11974), .ZN(n7503) );
  NAND2_X1 U9999 ( .A1(n7499), .A2(n10508), .ZN(n7498) );
  NAND3_X1 U10000 ( .A1(n7729), .A2(n15860), .A3(n7730), .ZN(n10266) );
  NAND2_X1 U10001 ( .A1(n11001), .A2(n10603), .ZN(n10990) );
  INV_X1 U10002 ( .A(n6938), .ZN(n6937) );
  NAND2_X1 U10003 ( .A1(n7234), .A2(n13192), .ZN(n13191) );
  NAND2_X1 U10004 ( .A1(n7942), .A2(n7940), .ZN(n10405) );
  NAND2_X1 U10005 ( .A1(n7200), .A2(n6656), .ZN(n7553) );
  NOR2_X1 U10006 ( .A1(n11866), .A2(n7133), .ZN(n10608) );
  INV_X1 U10007 ( .A(n11218), .ZN(n6928) );
  NAND2_X2 U10008 ( .A1(n13034), .A2(n13035), .ZN(n7776) );
  NAND4_X1 U10009 ( .A1(n9494), .A2(n6928), .A3(n11295), .A4(n13127), .ZN(
        n9495) );
  NAND2_X1 U10010 ( .A1(n7368), .A2(n7367), .ZN(n11218) );
  NAND2_X1 U10011 ( .A1(n7318), .A2(n9514), .ZN(n7319) );
  NAND3_X1 U10012 ( .A1(n9496), .A2(n9497), .A3(n9495), .ZN(n7318) );
  NAND2_X1 U10013 ( .A1(n12237), .A2(n9435), .ZN(n9440) );
  NAND4_X1 U10014 ( .A1(n7440), .A2(n7439), .A3(n7441), .A4(n6929), .ZN(n7898)
         );
  NAND3_X1 U10015 ( .A1(n12754), .A2(n6462), .A3(n6608), .ZN(n6929) );
  INV_X1 U10016 ( .A(n8353), .ZN(n7250) );
  NAND2_X1 U10017 ( .A1(n7249), .A2(n8082), .ZN(n8362) );
  NAND2_X1 U10018 ( .A1(n6981), .A2(n6494), .ZN(n6980) );
  INV_X1 U10019 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U10020 ( .A1(n15037), .A2(n12762), .ZN(n7259) );
  INV_X1 U10021 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10022 ( .A1(n8080), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U10023 ( .A1(n8194), .A2(n8100), .ZN(n8462) );
  NAND2_X1 U10024 ( .A1(n7266), .A2(n7265), .ZN(n14955) );
  NOR2_X1 U10025 ( .A1(n7015), .A2(n15147), .ZN(n15255) );
  NAND2_X1 U10026 ( .A1(n15149), .A2(n15572), .ZN(n7017) );
  AOI22_X1 U10027 ( .A1(n12514), .A2(n12513), .B1(n12512), .B2(n12511), .ZN(
        n12518) );
  NOR2_X2 U10028 ( .A1(n9905), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U10029 ( .A1(n12967), .A2(n13106), .ZN(n6932) );
  NAND2_X1 U10030 ( .A1(n7319), .A2(n6933), .ZN(n7322) );
  NAND2_X1 U10031 ( .A1(n9430), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U10032 ( .A1(n13061), .A2(n13060), .ZN(n12993) );
  AOI21_X1 U10033 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(n12955) );
  AOI21_X1 U10034 ( .B1(n12888), .B2(n12887), .A(n12886), .ZN(n12890) );
  NAND2_X1 U10035 ( .A1(n11294), .A2(n15784), .ZN(n9494) );
  INV_X1 U10036 ( .A(n12883), .ZN(n12888) );
  INV_X1 U10037 ( .A(n7772), .ZN(n7771) );
  NAND2_X1 U10038 ( .A1(n6946), .A2(n6614), .ZN(n7765) );
  INV_X4 U10039 ( .A(n12896), .ZN(n12895) );
  OAI211_X1 U10040 ( .C1(n7539), .C2(n12650), .A(n6934), .B(n12649), .ZN(
        P2_U3328) );
  NAND2_X1 U10041 ( .A1(n7539), .A2(n12629), .ZN(n6934) );
  NAND2_X1 U10042 ( .A1(n7897), .A2(n7896), .ZN(n8880) );
  NAND2_X1 U10043 ( .A1(n7833), .A2(n7835), .ZN(n12494) );
  NAND2_X1 U10044 ( .A1(n7107), .A2(n6937), .ZN(n13516) );
  OAI21_X1 U10045 ( .B1(n12205), .B2(n7108), .A(n10516), .ZN(n6938) );
  AOI21_X2 U10046 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(n15466) );
  NAND2_X1 U10047 ( .A1(n15373), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n6940) );
  INV_X1 U10048 ( .A(n15415), .ZN(n6941) );
  INV_X1 U10049 ( .A(n7330), .ZN(n15394) );
  NAND2_X1 U10050 ( .A1(n6943), .A2(n6942), .ZN(n7330) );
  INV_X1 U10051 ( .A(n15393), .ZN(n6943) );
  NAND2_X1 U10052 ( .A1(n7333), .A2(n7331), .ZN(n7335) );
  NOR2_X1 U10053 ( .A1(n15887), .A2(n15888), .ZN(n15886) );
  XNOR2_X1 U10054 ( .A(n15371), .B(n15632), .ZN(n15887) );
  NAND2_X1 U10055 ( .A1(n7738), .A2(n7737), .ZN(n13878) );
  NAND3_X1 U10056 ( .A1(n7280), .A2(n6603), .A3(n7281), .ZN(n13968) );
  AND2_X1 U10057 ( .A1(n7730), .A2(n10219), .ZN(n12919) );
  NAND2_X1 U10058 ( .A1(n7587), .A2(n7586), .ZN(n9426) );
  NAND2_X1 U10059 ( .A1(n7714), .A2(n6584), .ZN(n7296) );
  NAND2_X1 U10060 ( .A1(n13348), .A2(n10199), .ZN(n13331) );
  INV_X1 U10061 ( .A(n13008), .ZN(n6946) );
  OR2_X2 U10062 ( .A1(n9426), .A2(n9427), .ZN(n9905) );
  OAI21_X1 U10063 ( .B1(n10402), .B2(n15605), .A(n6467), .ZN(P1_U3524) );
  NAND2_X1 U10064 ( .A1(n7649), .A2(n6638), .ZN(n10570) );
  INV_X1 U10065 ( .A(n10478), .ZN(n7647) );
  NOR2_X1 U10066 ( .A1(n10487), .A2(n11399), .ZN(n10506) );
  OAI21_X1 U10067 ( .B1(n10485), .B2(n11503), .A(n10484), .ZN(n10486) );
  NOR4_X1 U10068 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n13519), .ZN(
        n7660) );
  NAND2_X1 U10069 ( .A1(n7251), .A2(n8079), .ZN(n8354) );
  INV_X1 U10070 ( .A(n7485), .ZN(n7482) );
  OAI211_X1 U10071 ( .C1(n12948), .C2(n12907), .A(n6949), .B(n12906), .ZN(
        P3_U3160) );
  NAND2_X1 U10072 ( .A1(n12948), .A2(n6588), .ZN(n6949) );
  BUF_X4 U10073 ( .A(n9744), .Z(n10207) );
  NAND2_X1 U10074 ( .A1(n6950), .A2(n6612), .ZN(n12472) );
  BUF_X4 U10075 ( .A(n6617), .Z(n12547) );
  NAND2_X1 U10076 ( .A1(n7541), .A2(n7540), .ZN(n7539) );
  AND2_X2 U10077 ( .A1(n7754), .A2(n6477), .ZN(n12534) );
  NAND2_X1 U10078 ( .A1(n15361), .A2(n15360), .ZN(n15331) );
  NAND2_X1 U10079 ( .A1(n15384), .A2(n15385), .ZN(n15326) );
  XNOR2_X1 U10080 ( .A(n7880), .B(n7879), .ZN(SUB_1596_U4) );
  NAND3_X1 U10081 ( .A1(n6959), .A2(n6958), .A3(n6957), .ZN(n7909) );
  NAND4_X1 U10082 ( .A1(n6967), .A2(n15507), .A3(n6966), .A4(n6965), .ZN(
        n12688) );
  NAND3_X1 U10083 ( .A1(n12683), .A2(n12682), .A3(n12829), .ZN(n6966) );
  NAND2_X1 U10084 ( .A1(n6610), .A2(n12829), .ZN(n6967) );
  NAND2_X1 U10085 ( .A1(n6970), .A2(n6972), .ZN(n7432) );
  NAND3_X1 U10086 ( .A1(n12783), .A2(n12782), .A3(n6616), .ZN(n6970) );
  NAND4_X1 U10087 ( .A1(n7490), .A2(n8131), .A3(n8463), .A4(n8184), .ZN(n8549)
         );
  AND2_X2 U10088 ( .A1(n8131), .A2(n8463), .ZN(n8183) );
  NAND2_X1 U10089 ( .A1(n12708), .A2(n6440), .ZN(n6984) );
  NAND2_X2 U10090 ( .A1(n6989), .A2(n6988), .ZN(n12768) );
  INV_X1 U10091 ( .A(n6992), .ZN(n13209) );
  NAND4_X1 U10092 ( .A1(n13609), .A2(n7511), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .A4(P1_ADDR_REG_19__SCAN_IN), .ZN(n7001) );
  NAND4_X1 U10093 ( .A1(n8065), .A2(n8063), .A3(n8064), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U10094 ( .A1(n7003), .A2(n7007), .ZN(n12307) );
  NAND3_X1 U10095 ( .A1(n7958), .A2(n7959), .A3(n10317), .ZN(n7003) );
  NAND2_X1 U10096 ( .A1(n7009), .A2(n12840), .ZN(n12269) );
  NAND2_X1 U10097 ( .A1(n7958), .A2(n7959), .ZN(n7009) );
  NAND2_X2 U10098 ( .A1(n8407), .A2(n8406), .ZN(n15242) );
  INV_X1 U10099 ( .A(n14772), .ZN(n7030) );
  NAND3_X1 U10100 ( .A1(n7026), .A2(n7025), .A3(n7024), .ZN(n7033) );
  NAND2_X1 U10101 ( .A1(n7033), .A2(n6598), .ZN(n10854) );
  NOR2_X1 U10102 ( .A1(n12071), .A2(n7038), .ZN(n14790) );
  NAND2_X1 U10103 ( .A1(n15470), .A2(n12069), .ZN(n12071) );
  INV_X1 U10104 ( .A(n10915), .ZN(n7050) );
  OAI21_X1 U10105 ( .B1(n8016), .B2(n7054), .A(n12240), .ZN(n7053) );
  NAND2_X1 U10106 ( .A1(n14476), .A2(n7061), .ZN(n7058) );
  NAND2_X1 U10107 ( .A1(n7058), .A2(n7059), .ZN(n14298) );
  NAND2_X1 U10108 ( .A1(n14242), .A2(n10036), .ZN(n7070) );
  NAND2_X2 U10109 ( .A1(n8850), .A2(n8872), .ZN(n8863) );
  AND4_X2 U10110 ( .A1(n7787), .A2(n8839), .A3(n8866), .A4(n7749), .ZN(n8850)
         );
  AND2_X2 U10111 ( .A1(n8838), .A2(n8837), .ZN(n8866) );
  AND3_X2 U10112 ( .A1(n8865), .A2(n8835), .A3(n8929), .ZN(n7787) );
  NAND3_X1 U10113 ( .A1(n7159), .A2(n10283), .A3(n15778), .ZN(n10292) );
  INV_X1 U10114 ( .A(n12940), .ZN(n7072) );
  NAND2_X1 U10115 ( .A1(n10272), .A2(n10273), .ZN(n12940) );
  INV_X1 U10116 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U10117 ( .A1(n9221), .A2(n6653), .ZN(n9250) );
  NAND2_X1 U10118 ( .A1(n9221), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U10119 ( .A1(n9275), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U10120 ( .A1(n7082), .A2(n6637), .ZN(n7080) );
  INV_X1 U10121 ( .A(n7453), .ZN(n7084) );
  OAI21_X1 U10122 ( .B1(n7084), .B2(n7086), .A(n7085), .ZN(n9782) );
  INV_X1 U10123 ( .A(n7454), .ZN(n7090) );
  NAND2_X1 U10124 ( .A1(n7092), .A2(n6472), .ZN(n7095) );
  INV_X1 U10125 ( .A(n10588), .ZN(n7092) );
  NAND4_X1 U10126 ( .A1(n7095), .A2(n10595), .A3(n7094), .A4(n7093), .ZN(
        P3_U3296) );
  NAND3_X1 U10127 ( .A1(n10588), .A2(n10592), .A3(n10589), .ZN(n7093) );
  NAND3_X1 U10128 ( .A1(n7100), .A2(n7096), .A3(n10580), .ZN(n7283) );
  OAI211_X1 U10129 ( .C1(n7671), .C2(n13332), .A(n10579), .B(n7097), .ZN(n7096) );
  NAND2_X1 U10130 ( .A1(n7099), .A2(n7673), .ZN(n7097) );
  OAI21_X1 U10131 ( .B1(n7472), .B2(n7674), .A(n7098), .ZN(n7100) );
  NOR2_X1 U10132 ( .A1(n7672), .A2(n10581), .ZN(n7098) );
  NOR2_X1 U10133 ( .A1(n10575), .A2(n13332), .ZN(n7099) );
  NAND2_X1 U10134 ( .A1(n6600), .A2(n12371), .ZN(n9415) );
  NAND2_X1 U10135 ( .A1(n10416), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U10136 ( .A1(n7728), .A2(n7104), .ZN(n7354) );
  AOI21_X1 U10137 ( .B1(n7729), .B2(n6466), .A(n6635), .ZN(n7104) );
  INV_X1 U10138 ( .A(n11878), .ZN(n7106) );
  NAND3_X1 U10139 ( .A1(n7105), .A2(n7939), .A3(n7498), .ZN(n7109) );
  NAND2_X1 U10140 ( .A1(n7109), .A2(n7108), .ZN(n12206) );
  NAND3_X1 U10141 ( .A1(n7511), .A2(n13609), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7112) );
  NAND3_X1 U10142 ( .A1(n8064), .A2(n8063), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7113) );
  NAND2_X1 U10143 ( .A1(n10608), .A2(n10658), .ZN(n7578) );
  NAND2_X1 U10144 ( .A1(n13258), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U10145 ( .A1(n13185), .A2(n13184), .ZN(n7143) );
  OAI21_X1 U10146 ( .B1(n10692), .B2(n6430), .A(n7139), .ZN(n7142) );
  AOI21_X1 U10147 ( .B1(n13184), .B2(P3_REG2_REG_11__SCAN_IN), .A(n6430), .ZN(
        n7140) );
  NAND2_X1 U10148 ( .A1(n7144), .A2(n10692), .ZN(n13169) );
  INV_X1 U10149 ( .A(n10691), .ZN(n7145) );
  NAND2_X1 U10150 ( .A1(n10682), .A2(n11349), .ZN(n7146) );
  NAND4_X1 U10151 ( .A1(n7146), .A2(n7147), .A3(n7682), .A4(
        P3_REG2_REG_5__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U10152 ( .A1(n6615), .A2(n11018), .ZN(n7147) );
  NAND3_X1 U10153 ( .A1(n7150), .A2(n7778), .A3(P3_IR_REG_4__SCAN_IN), .ZN(
        n7149) );
  NAND2_X1 U10154 ( .A1(n7153), .A2(n7152), .ZN(n9519) );
  NAND2_X2 U10155 ( .A1(n12149), .A2(n9958), .ZN(n12241) );
  NAND3_X1 U10156 ( .A1(n10283), .A2(n7159), .A3(n15767), .ZN(n10298) );
  NAND2_X1 U10157 ( .A1(n11035), .A2(n12595), .ZN(n11034) );
  NAND2_X2 U10158 ( .A1(n7780), .A2(n7165), .ZN(n14373) );
  NAND3_X1 U10159 ( .A1(n8887), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_29__SCAN_IN), .ZN(n7169) );
  NAND3_X1 U10160 ( .A1(n7897), .A2(n7896), .A3(n8881), .ZN(n8887) );
  AOI21_X1 U10161 ( .B1(n14869), .B2(n7173), .A(n7172), .ZN(n7171) );
  NOR2_X1 U10162 ( .A1(n7177), .A2(n7951), .ZN(n7176) );
  NAND2_X1 U10163 ( .A1(n7178), .A2(n10305), .ZN(n15485) );
  NAND2_X1 U10164 ( .A1(n11962), .A2(n7178), .ZN(n11964) );
  INV_X1 U10165 ( .A(n10302), .ZN(n10301) );
  NAND3_X1 U10166 ( .A1(n7179), .A2(n8214), .A3(n8215), .ZN(n10302) );
  AND3_X2 U10167 ( .A1(n7787), .A2(n8912), .A3(n8866), .ZN(n7896) );
  NAND2_X1 U10168 ( .A1(n10010), .A2(n10009), .ZN(n11626) );
  NAND2_X1 U10169 ( .A1(n7193), .A2(n7192), .ZN(n8026) );
  NAND2_X1 U10170 ( .A1(n14646), .A2(n14647), .ZN(n7198) );
  NAND2_X1 U10171 ( .A1(n14591), .A2(n14592), .ZN(n7199) );
  NAND2_X1 U10172 ( .A1(n7200), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13276) );
  NAND3_X1 U10173 ( .A1(n7205), .A2(n10976), .A3(n7547), .ZN(n7203) );
  NAND2_X1 U10174 ( .A1(n7205), .A2(n7547), .ZN(n13270) );
  OAI211_X1 U10175 ( .C1(n7205), .C2(n6654), .A(n7203), .B(n7202), .ZN(n7201)
         );
  NAND2_X1 U10176 ( .A1(n11019), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U10177 ( .A1(n11907), .A2(n7212), .ZN(n7210) );
  NAND2_X1 U10178 ( .A1(n11907), .A2(n7208), .ZN(n7207) );
  NAND2_X1 U10179 ( .A1(n6429), .A2(n12218), .ZN(n7209) );
  NAND2_X1 U10180 ( .A1(n12217), .A2(n12218), .ZN(n12252) );
  NAND2_X1 U10181 ( .A1(n7210), .A2(n7211), .ZN(n12217) );
  NAND2_X1 U10182 ( .A1(n12300), .A2(n12299), .ZN(n7215) );
  NAND2_X1 U10183 ( .A1(n7217), .A2(n8248), .ZN(n11122) );
  NAND2_X1 U10184 ( .A1(n7219), .A2(n8225), .ZN(n8248) );
  NAND2_X1 U10185 ( .A1(n7360), .A2(n7218), .ZN(n7217) );
  INV_X1 U10186 ( .A(n7219), .ZN(n7218) );
  NAND2_X1 U10187 ( .A1(n7969), .A2(n7221), .ZN(n7220) );
  OAI211_X1 U10188 ( .C1(n7969), .C2(n7222), .A(n7220), .B(n14579), .ZN(
        P1_U3214) );
  NOR2_X1 U10189 ( .A1(n14574), .A2(n6571), .ZN(n7226) );
  NAND2_X1 U10190 ( .A1(n6571), .A2(n14574), .ZN(n7227) );
  INV_X1 U10191 ( .A(n14574), .ZN(n7228) );
  NAND2_X1 U10192 ( .A1(n7577), .A2(n7235), .ZN(n7234) );
  INV_X1 U10193 ( .A(n13194), .ZN(n7235) );
  NAND3_X1 U10194 ( .A1(n7241), .A2(n9483), .A3(n10674), .ZN(n7237) );
  NAND3_X1 U10195 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7240), .A3(
        P3_IR_REG_2__SCAN_IN), .ZN(n7239) );
  INV_X1 U10196 ( .A(n8645), .ZN(n7243) );
  NAND3_X1 U10197 ( .A1(n7580), .A2(n7579), .A3(n10665), .ZN(n7246) );
  NAND2_X1 U10198 ( .A1(n7580), .A2(n7579), .ZN(n13235) );
  XNOR2_X2 U10199 ( .A(n7248), .B(n8166), .ZN(n8811) );
  NAND2_X1 U10200 ( .A1(n8354), .A2(n7250), .ZN(n7249) );
  NAND2_X1 U10201 ( .A1(n7361), .A2(n8077), .ZN(n7251) );
  OAI211_X1 U10202 ( .C1(n8080), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n7253), .B(
        SI_1_), .ZN(n7252) );
  NAND2_X1 U10203 ( .A1(n8080), .A2(n10748), .ZN(n7253) );
  NAND2_X1 U10204 ( .A1(n8216), .A2(n7255), .ZN(n7254) );
  OAI211_X1 U10205 ( .C1(n8080), .C2(n10776), .A(n7256), .B(n10775), .ZN(n7255) );
  NAND2_X1 U10206 ( .A1(n7259), .A2(n7257), .ZN(n10383) );
  NAND2_X1 U10207 ( .A1(n14935), .A2(n10389), .ZN(n7853) );
  NAND2_X1 U10208 ( .A1(n7992), .A2(n7993), .ZN(n8192) );
  NAND2_X1 U10209 ( .A1(n15000), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U10210 ( .A1(n11893), .A2(n9049), .ZN(n11994) );
  INV_X1 U10211 ( .A(n9115), .ZN(n7282) );
  NAND2_X1 U10212 ( .A1(n12362), .A2(n12361), .ZN(n12360) );
  NAND2_X1 U10213 ( .A1(n7283), .A2(n10584), .ZN(n10587) );
  NAND2_X1 U10214 ( .A1(n11882), .A2(n6450), .ZN(n7284) );
  NAND2_X1 U10215 ( .A1(n11884), .A2(n10136), .ZN(n7286) );
  OR2_X2 U10216 ( .A1(n13388), .A2(n10152), .ZN(n7293) );
  NAND3_X1 U10217 ( .A1(n7301), .A2(n9525), .A3(n9524), .ZN(n9562) );
  AND2_X1 U10218 ( .A1(n9725), .A2(n9724), .ZN(n9742) );
  NAND3_X1 U10219 ( .A1(n6423), .A2(n10573), .A3(n13368), .ZN(n7315) );
  NAND2_X1 U10220 ( .A1(n7321), .A2(n9514), .ZN(n7320) );
  NAND2_X1 U10221 ( .A1(n11246), .A2(n9514), .ZN(n11362) );
  NAND2_X1 U10222 ( .A1(n7755), .A2(n11247), .ZN(n11246) );
  NAND2_X1 U10223 ( .A1(n7322), .A2(n7771), .ZN(n9571) );
  OAI21_X1 U10224 ( .B1(n15880), .B2(n15881), .A(n7323), .ZN(SUB_1596_U56) );
  NAND2_X1 U10225 ( .A1(n7323), .A2(n15391), .ZN(n15393) );
  NAND2_X1 U10226 ( .A1(n15881), .A2(n15880), .ZN(n7323) );
  NAND2_X1 U10227 ( .A1(n7326), .A2(n7327), .ZN(n15318) );
  NOR2_X1 U10228 ( .A1(n7325), .A2(n15317), .ZN(n7324) );
  OR2_X1 U10229 ( .A1(n15423), .A2(n7332), .ZN(n7331) );
  OR2_X1 U10230 ( .A1(n15426), .A2(n15424), .ZN(n7332) );
  AOI21_X1 U10231 ( .B1(n15394), .B2(n7334), .A(P2_ADDR_REG_9__SCAN_IN), .ZN(
        n7333) );
  INV_X1 U10232 ( .A(n15426), .ZN(n7334) );
  INV_X1 U10233 ( .A(n7336), .ZN(n15422) );
  XNOR2_X1 U10234 ( .A(n15366), .B(n7341), .ZN(n15417) );
  XNOR2_X1 U10235 ( .A(n15368), .B(n15369), .ZN(n15371) );
  NAND2_X1 U10236 ( .A1(n15874), .A2(n15875), .ZN(n7859) );
  NAND2_X1 U10237 ( .A1(n7496), .A2(n10482), .ZN(n11396) );
  OAI22_X2 U10238 ( .A1(n13416), .A2(n10149), .B1(n13782), .B2(n13401), .ZN(
        n13400) );
  OAI211_X1 U10239 ( .C1(n13333), .C2(n13332), .A(n13331), .B(n15801), .ZN(
        n13339) );
  NOR2_X2 U10240 ( .A1(n9405), .A2(n9399), .ZN(n7587) );
  NAND2_X1 U10241 ( .A1(n11983), .A2(n9640), .ZN(n13063) );
  NAND3_X1 U10242 ( .A1(n9424), .A2(n9423), .A3(n9425), .ZN(n10121) );
  NAND3_X1 U10243 ( .A1(n7979), .A2(n7377), .A3(n7981), .ZN(n7376) );
  NAND2_X1 U10244 ( .A1(n8223), .A2(n8224), .ZN(n7350) );
  INV_X1 U10245 ( .A(n7352), .ZN(n8156) );
  INV_X1 U10246 ( .A(n7351), .ZN(n8152) );
  NAND2_X1 U10247 ( .A1(n7352), .A2(n8157), .ZN(n7351) );
  INV_X1 U10248 ( .A(n14202), .ZN(n8023) );
  NAND2_X1 U10249 ( .A1(n8038), .A2(n7584), .ZN(n9410) );
  INV_X4 U10250 ( .A(n8080), .ZN(n10769) );
  OAI21_X1 U10251 ( .B1(n7849), .B2(n7489), .A(n14883), .ZN(n7488) );
  NAND2_X1 U10252 ( .A1(n7354), .A2(n10256), .ZN(P3_U3488) );
  AOI22_X1 U10253 ( .A1(n9494), .A2(n9493), .B1(n9492), .B2(n13126), .ZN(n9496) );
  INV_X1 U10254 ( .A(n7502), .ZN(n7499) );
  XNOR2_X1 U10255 ( .A(n15388), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15881) );
  INV_X1 U10256 ( .A(n10121), .ZN(n15807) );
  NAND2_X1 U10257 ( .A1(n10143), .A2(n7715), .ZN(n7714) );
  NAND2_X1 U10258 ( .A1(n11195), .A2(n11197), .ZN(n11196) );
  OAI21_X1 U10259 ( .B1(n8461), .B2(n8460), .A(n12253), .ZN(n12300) );
  NAND2_X1 U10260 ( .A1(n11123), .A2(n8248), .ZN(n11195) );
  NAND3_X1 U10261 ( .A1(n8303), .A2(n8074), .A3(n8304), .ZN(n7361) );
  OAI21_X1 U10262 ( .B1(n7774), .B2(n7773), .A(n11670), .ZN(n7772) );
  NAND2_X1 U10263 ( .A1(n11401), .A2(n10128), .ZN(n11615) );
  NAND2_X1 U10264 ( .A1(n13548), .A2(n6633), .ZN(P3_U3487) );
  INV_X1 U10265 ( .A(n9908), .ZN(n13834) );
  INV_X1 U10266 ( .A(n10166), .ZN(n10167) );
  INV_X1 U10267 ( .A(n15446), .ZN(n15447) );
  NAND2_X1 U10268 ( .A1(n15714), .A2(n15436), .ZN(n15433) );
  XNOR2_X2 U10269 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n15368) );
  NAND2_X1 U10270 ( .A1(n15447), .A2(n15445), .ZN(n15452) );
  XNOR2_X1 U10271 ( .A(n15393), .B(n15392), .ZN(n15423) );
  NAND2_X1 U10272 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n7374), .ZN(n7373) );
  INV_X1 U10273 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7374) );
  NAND2_X1 U10274 ( .A1(n15315), .A2(n15368), .ZN(n7878) );
  NAND2_X1 U10275 ( .A1(n15362), .A2(n10845), .ZN(n15324) );
  INV_X1 U10276 ( .A(n11422), .ZN(n7721) );
  NAND2_X1 U10277 ( .A1(n9204), .A2(n7739), .ZN(n7738) );
  NAND2_X1 U10278 ( .A1(n11327), .A2(n11326), .ZN(n11325) );
  NOR2_X1 U10279 ( .A1(n13922), .A2(n13921), .ZN(n13926) );
  AND2_X2 U10280 ( .A1(n7376), .A2(n8382), .ZN(n11907) );
  NAND2_X1 U10281 ( .A1(n8362), .A2(n8083), .ZN(n7380) );
  MUX2_X1 U10282 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n10769), .Z(n8217) );
  NAND2_X1 U10283 ( .A1(n7804), .A2(n7385), .ZN(n7383) );
  NAND2_X1 U10284 ( .A1(n7389), .A2(n7393), .ZN(n14282) );
  NAND2_X1 U10285 ( .A1(n14313), .A2(n7395), .ZN(n7389) );
  OAI21_X1 U10286 ( .B1(n7392), .B2(n14313), .A(n7390), .ZN(n9971) );
  AOI21_X1 U10287 ( .B1(n7393), .B2(n7391), .A(n6587), .ZN(n7390) );
  INV_X1 U10288 ( .A(n7395), .ZN(n7391) );
  INV_X1 U10289 ( .A(n7393), .ZN(n7392) );
  OAI21_X1 U10290 ( .B1(n8080), .B2(n7399), .A(n7398), .ZN(n8078) );
  NAND2_X1 U10291 ( .A1(n8080), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U10292 ( .A1(n7402), .A2(n7401), .ZN(n7952) );
  NAND2_X2 U10293 ( .A1(n8235), .A2(n10071), .ZN(n8301) );
  NAND2_X4 U10294 ( .A1(n10101), .A2(n8811), .ZN(n8235) );
  NAND2_X2 U10295 ( .A1(n8143), .A2(n8167), .ZN(n10101) );
  NAND3_X1 U10296 ( .A1(n6604), .A2(n8183), .A3(n8138), .ZN(n8150) );
  NOR2_X2 U10297 ( .A1(n8329), .A2(n8137), .ZN(n8138) );
  INV_X1 U10298 ( .A(n10897), .ZN(n7423) );
  MUX2_X1 U10299 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10840), .S(n14751), .Z(
        n14759) );
  INV_X1 U10300 ( .A(n7428), .ZN(n7426) );
  INV_X1 U10301 ( .A(n14809), .ZN(n7429) );
  INV_X1 U10302 ( .A(n14798), .ZN(n7430) );
  NAND2_X1 U10303 ( .A1(n7432), .A2(n12789), .ZN(n12787) );
  INV_X1 U10304 ( .A(n12785), .ZN(n7433) );
  NAND2_X1 U10305 ( .A1(n11257), .A2(n10091), .ZN(n7434) );
  NAND2_X1 U10306 ( .A1(n12795), .A2(n7437), .ZN(n7436) );
  NAND4_X1 U10307 ( .A1(n12754), .A2(n12732), .A3(n12731), .A4(n6462), .ZN(
        n7440) );
  NAND2_X1 U10308 ( .A1(n9642), .A2(n9641), .ZN(n7449) );
  NAND2_X1 U10309 ( .A1(n9705), .A2(n7455), .ZN(n7453) );
  NAND2_X1 U10310 ( .A1(n10154), .A2(n12230), .ZN(n7944) );
  NAND2_X1 U10311 ( .A1(n7471), .A2(n7469), .ZN(n10173) );
  NAND2_X1 U10312 ( .A1(n7473), .A2(n10352), .ZN(n11968) );
  NAND3_X1 U10313 ( .A1(n7482), .A2(n10377), .A3(n6496), .ZN(n7481) );
  INV_X1 U10314 ( .A(n8329), .ZN(n7490) );
  AND2_X2 U10315 ( .A1(n8172), .A2(n8170), .ZN(n8226) );
  NAND3_X1 U10316 ( .A1(n8172), .A2(n8170), .A3(P1_REG1_REG_2__SCAN_IN), .ZN(
        n7494) );
  NAND2_X1 U10317 ( .A1(n10225), .A2(n10226), .ZN(n7496) );
  NAND3_X1 U10318 ( .A1(n7501), .A2(n7500), .A3(n10508), .ZN(n12092) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8080), .Z(n8075) );
  OAI21_X2 U10320 ( .B1(n8191), .B2(n7529), .A(n8051), .ZN(n7528) );
  NAND2_X1 U10321 ( .A1(n7821), .A2(n6613), .ZN(n7540) );
  NAND3_X1 U10322 ( .A1(n10090), .A2(n10089), .A3(n7543), .ZN(n14557) );
  NAND3_X1 U10323 ( .A1(n7557), .A2(n7554), .A3(n7553), .ZN(n13301) );
  NAND3_X1 U10324 ( .A1(n7558), .A2(n13307), .A3(n13278), .ZN(n7557) );
  XNOR2_X1 U10325 ( .A(n10605), .B(n10791), .ZN(n11340) );
  OR2_X1 U10326 ( .A1(n10605), .A2(n11349), .ZN(n7563) );
  AND4_X2 U10327 ( .A1(n7569), .A2(n7568), .A3(n7566), .A4(n7565), .ZN(n11487)
         );
  NAND3_X1 U10328 ( .A1(n7573), .A2(n13156), .A3(n10688), .ZN(n7565) );
  NAND2_X1 U10329 ( .A1(n13231), .A2(n13232), .ZN(n7580) );
  NAND3_X1 U10330 ( .A1(n7582), .A2(n7581), .A3(n10611), .ZN(n7579) );
  INV_X1 U10331 ( .A(n10610), .ZN(n7583) );
  INV_X1 U10332 ( .A(n9410), .ZN(n7585) );
  INV_X1 U10333 ( .A(n9427), .ZN(n7584) );
  NAND3_X1 U10334 ( .A1(n7585), .A2(n7587), .A3(n7586), .ZN(n9438) );
  INV_X1 U10335 ( .A(n7590), .ZN(n13261) );
  NAND2_X1 U10336 ( .A1(n11028), .A2(n6585), .ZN(n7591) );
  NAND2_X1 U10337 ( .A1(n7596), .A2(n11163), .ZN(n7595) );
  NAND2_X1 U10338 ( .A1(n7598), .A2(n7597), .ZN(n11345) );
  OR2_X1 U10339 ( .A1(n9420), .A2(n7604), .ZN(n7603) );
  NAND2_X1 U10340 ( .A1(n7609), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U10341 ( .A1(n13163), .A2(n7611), .ZN(n7610) );
  NAND2_X1 U10342 ( .A1(n7610), .A2(n7613), .ZN(n13172) );
  INV_X1 U10343 ( .A(n15498), .ZN(n7629) );
  NAND3_X1 U10344 ( .A1(n7630), .A2(n7629), .A3(n7628), .ZN(n11722) );
  INV_X1 U10345 ( .A(n7631), .ZN(n11956) );
  NAND3_X1 U10346 ( .A1(n7646), .A2(n7645), .A3(n10481), .ZN(n7644) );
  NAND3_X1 U10347 ( .A1(n10477), .A2(n10476), .A3(n10564), .ZN(n7645) );
  OR2_X1 U10348 ( .A1(n7677), .A2(n10717), .ZN(P3_U3200) );
  AND2_X1 U10349 ( .A1(n10696), .A2(n10697), .ZN(n7692) );
  NAND2_X1 U10350 ( .A1(n11859), .A2(n11858), .ZN(n7696) );
  AND2_X1 U10351 ( .A1(n10689), .A2(n10688), .ZN(n7707) );
  NAND2_X1 U10352 ( .A1(n7702), .A2(n11858), .ZN(n11862) );
  NAND2_X1 U10353 ( .A1(n7705), .A2(n7704), .ZN(n7702) );
  INV_X1 U10354 ( .A(n11858), .ZN(n7703) );
  NOR2_X4 U10355 ( .A1(n11722), .A2(n15242), .ZN(n12168) );
  NOR2_X2 U10356 ( .A1(n10095), .A2(n15517), .ZN(n14821) );
  NAND2_X1 U10357 ( .A1(n7746), .A2(n7745), .ZN(n7744) );
  AOI211_X1 U10358 ( .C1(n10570), .C2(n6586), .A(n10569), .B(n13375), .ZN(
        n10575) );
  CLKBUF_X1 U10359 ( .A(n7714), .Z(n7708) );
  NAND2_X1 U10360 ( .A1(n10131), .A2(n10132), .ZN(n7717) );
  OAI21_X1 U10361 ( .B1(n10132), .B2(n7366), .A(n10131), .ZN(n7719) );
  NAND3_X1 U10362 ( .A1(n7718), .A2(n7717), .A3(n10133), .ZN(n10135) );
  NAND2_X1 U10363 ( .A1(n11615), .A2(n10131), .ZN(n7718) );
  XNOR2_X1 U10364 ( .A(n7719), .B(n11877), .ZN(n11772) );
  NAND2_X1 U10365 ( .A1(n7726), .A2(n7725), .ZN(n7724) );
  INV_X1 U10366 ( .A(n8898), .ZN(n7726) );
  NAND2_X1 U10367 ( .A1(n10221), .A2(n15801), .ZN(n7730) );
  INV_X1 U10368 ( .A(n11299), .ZN(n11448) );
  NAND3_X1 U10369 ( .A1(n7787), .A2(n8839), .A3(n8866), .ZN(n9099) );
  INV_X1 U10370 ( .A(n9366), .ZN(n10062) );
  INV_X1 U10371 ( .A(n9426), .ZN(n7753) );
  OAI21_X1 U10372 ( .B1(n11247), .B2(n7755), .A(n11246), .ZN(n11248) );
  OR2_X2 U10373 ( .A1(n9844), .A2(n9874), .ZN(n7756) );
  NOR2_X1 U10374 ( .A1(n13008), .A2(n12892), .ZN(n13085) );
  NAND2_X1 U10375 ( .A1(n7765), .A2(n7766), .ZN(n12950) );
  NAND3_X1 U10376 ( .A1(n9501), .A2(n9451), .A3(n9520), .ZN(n9720) );
  NAND4_X1 U10377 ( .A1(n9501), .A2(n9451), .A3(n9520), .A4(n7779), .ZN(n9736)
         );
  NAND2_X1 U10378 ( .A1(n11733), .A2(n9943), .ZN(n9946) );
  NAND2_X1 U10379 ( .A1(n12241), .A2(n7783), .ZN(n7780) );
  NAND2_X1 U10380 ( .A1(n8893), .A2(n7797), .ZN(n7796) );
  NAND2_X1 U10381 ( .A1(n11034), .A2(n6596), .ZN(n7801) );
  NAND2_X1 U10382 ( .A1(n12500), .A2(n7810), .ZN(n7809) );
  NAND2_X1 U10383 ( .A1(n7809), .A2(n7813), .ZN(n12507) );
  INV_X1 U10384 ( .A(n12531), .ZN(n7823) );
  INV_X1 U10385 ( .A(n7824), .ZN(n12482) );
  AOI21_X1 U10386 ( .B1(n12477), .B2(n7827), .A(n7825), .ZN(n7824) );
  AND2_X1 U10387 ( .A1(n12395), .A2(n7831), .ZN(n12409) );
  NAND3_X1 U10388 ( .A1(n12485), .A2(n7834), .A3(n12484), .ZN(n7833) );
  NAND2_X2 U10389 ( .A1(n7840), .A2(n10303), .ZN(n12667) );
  OAI21_X1 U10390 ( .B1(n15874), .B2(n15875), .A(n7859), .ZN(SUB_1596_U59) );
  NAND3_X1 U10391 ( .A1(n15447), .A2(n15445), .A3(n7863), .ZN(n7862) );
  INV_X1 U10392 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7864) );
  XNOR2_X2 U10393 ( .A(n15320), .B(n7865), .ZN(n15363) );
  NAND3_X1 U10394 ( .A1(n6522), .A2(n11552), .A3(n11643), .ZN(n11533) );
  AND2_X1 U10395 ( .A1(n14197), .A2(n7892), .ZN(n14176) );
  NAND2_X1 U10396 ( .A1(n14197), .A2(n7891), .ZN(n14175) );
  NAND2_X1 U10397 ( .A1(n14197), .A2(n7895), .ZN(n8060) );
  AND4_X2 U10398 ( .A1(n8872), .A2(n8873), .A3(n8871), .A4(n8870), .ZN(n7897)
         );
  NAND2_X1 U10399 ( .A1(n7898), .A2(n7899), .ZN(n12781) );
  NAND2_X1 U10400 ( .A1(n12727), .A2(n12728), .ZN(n12726) );
  INV_X1 U10401 ( .A(n12772), .ZN(n7905) );
  NAND2_X1 U10402 ( .A1(n7909), .A2(n7908), .ZN(n12708) );
  NAND2_X1 U10403 ( .A1(n12703), .A2(n12705), .ZN(n7908) );
  NAND2_X1 U10404 ( .A1(n9469), .A2(n9468), .ZN(n9471) );
  NAND2_X1 U10405 ( .A1(n9482), .A2(n9473), .ZN(n7913) );
  NAND2_X1 U10406 ( .A1(n10229), .A2(n7915), .ZN(n7914) );
  XNOR2_X1 U10407 ( .A(n7917), .B(n11600), .ZN(n15846) );
  OAI21_X1 U10408 ( .B1(n13451), .B2(n7922), .A(n7920), .ZN(n13427) );
  NAND2_X1 U10409 ( .A1(n7919), .A2(n7918), .ZN(n10236) );
  NAND2_X1 U10410 ( .A1(n7927), .A2(n7928), .ZN(n9625) );
  INV_X1 U10411 ( .A(n10576), .ZN(n7943) );
  OAI21_X1 U10412 ( .B1(n7943), .B2(n6423), .A(n10577), .ZN(n7941) );
  NAND2_X1 U10413 ( .A1(n13357), .A2(n10576), .ZN(n7942) );
  NAND2_X1 U10414 ( .A1(n7944), .A2(n10156), .ZN(n10161) );
  NAND2_X1 U10415 ( .A1(n10186), .A2(n7947), .ZN(n7945) );
  OAI21_X1 U10416 ( .B1(n10186), .B2(n10185), .A(n10187), .ZN(n10204) );
  NAND4_X1 U10417 ( .A1(n7956), .A2(n12677), .A3(n12668), .A4(n12667), .ZN(
        n11821) );
  INV_X1 U10418 ( .A(n12826), .ZN(n7957) );
  INV_X2 U10419 ( .A(n8226), .ZN(n12660) );
  NAND2_X1 U10420 ( .A1(n14618), .A2(n14619), .ZN(n7975) );
  NAND2_X1 U10421 ( .A1(n8317), .A2(n8320), .ZN(n8313) );
  NAND2_X1 U10422 ( .A1(n7985), .A2(n7984), .ZN(n7983) );
  NAND2_X1 U10423 ( .A1(n7980), .A2(n8322), .ZN(n7985) );
  NAND2_X1 U10424 ( .A1(n8322), .A2(n11372), .ZN(n11413) );
  AND2_X1 U10425 ( .A1(n8614), .A2(n8615), .ZN(n7991) );
  INV_X1 U10426 ( .A(n8672), .ZN(n8002) );
  NAND3_X1 U10427 ( .A1(n8005), .A2(n8004), .A3(n8069), .ZN(n8234) );
  NOR2_X2 U10428 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8884) );
  NAND2_X1 U10429 ( .A1(n12118), .A2(n8017), .ZN(n8014) );
  AOI21_X1 U10430 ( .B1(n11397), .B2(n11503), .A(n10126), .ZN(n10127) );
  NOR2_X2 U10431 ( .A1(n15091), .A2(n15212), .ZN(n15076) );
  INV_X1 U10432 ( .A(n8899), .ZN(n9014) );
  AND2_X1 U10433 ( .A1(n11051), .A2(n11054), .ZN(n14374) );
  OAI21_X1 U10434 ( .B1(n10063), .B2(n10062), .A(n8047), .ZN(P2_U3186) );
  OR2_X1 U10435 ( .A1(n10054), .A2(n10053), .ZN(P2_U3236) );
  NAND2_X1 U10436 ( .A1(n10414), .A2(n10413), .ZN(n10458) );
  OAI21_X1 U10437 ( .B1(n12672), .B2(n12816), .A(n12671), .ZN(n12673) );
  OAI211_X1 U10438 ( .C1(SI_2_), .C2(n8073), .A(n8071), .B(n8274), .ZN(n8304)
         );
  NAND2_X1 U10439 ( .A1(n12673), .A2(n12691), .ZN(n12675) );
  NAND2_X1 U10440 ( .A1(n12826), .A2(n12768), .ZN(n12674) );
  NAND2_X1 U10441 ( .A1(n15795), .A2(n10475), .ZN(n10223) );
  NAND2_X1 U10442 ( .A1(n8317), .A2(n8321), .ZN(n11372) );
  AOI21_X1 U10443 ( .B1(n14835), .B2(n14834), .A(n15517), .ZN(n14836) );
  INV_X1 U10444 ( .A(n15517), .ZN(n15500) );
  XNOR2_X1 U10445 ( .A(n8737), .B(n8718), .ZN(n14568) );
  INV_X1 U10446 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9344) );
  AND2_X1 U10447 ( .A1(n10597), .A2(n10761), .ZN(n10756) );
  NAND4_X4 U10448 ( .A1(n8231), .A2(n8230), .A3(n8229), .A4(n8228), .ZN(n15105) );
  OR2_X1 U10449 ( .A1(n12381), .A2(n12380), .ZN(n12383) );
  OR2_X1 U10450 ( .A1(n12380), .A2(n10044), .ZN(n9932) );
  INV_X1 U10451 ( .A(n15798), .ZN(n9465) );
  INV_X4 U10452 ( .A(n10769), .ZN(n10768) );
  NAND2_X1 U10453 ( .A1(n7746), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9416) );
  INV_X1 U10454 ( .A(n12601), .ZN(n10013) );
  AND2_X1 U10455 ( .A1(n9419), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8037) );
  INV_X1 U10456 ( .A(n12608), .ZN(n10020) );
  AND3_X1 U10457 ( .A1(n14626), .A2(n14628), .A3(n14704), .ZN(n8039) );
  XOR2_X1 U10458 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n8040) );
  INV_X1 U10459 ( .A(n15228), .ZN(n10399) );
  INV_X4 U10460 ( .A(n10769), .ZN(n10071) );
  OR2_X1 U10461 ( .A1(n13774), .A2(n13083), .ZN(n8041) );
  NOR2_X1 U10462 ( .A1(n10354), .A2(n12830), .ZN(n8042) );
  AND2_X1 U10463 ( .A1(n9751), .A2(n13112), .ZN(n8043) );
  OR2_X1 U10464 ( .A1(n13347), .A2(n13358), .ZN(n8044) );
  NAND2_X1 U10465 ( .A1(n10280), .A2(n9990), .ZN(n8045) );
  AND2_X1 U10466 ( .A1(n9132), .A2(n9133), .ZN(n8046) );
  AND2_X1 U10467 ( .A1(n10061), .A2(n10060), .ZN(n8047) );
  NAND2_X2 U10468 ( .A1(n14842), .A2(n15511), .ZN(n15513) );
  INV_X1 U10469 ( .A(n15288), .ZN(n10118) );
  AND2_X1 U10470 ( .A1(n8856), .A2(n8855), .ZN(n8048) );
  INV_X1 U10471 ( .A(n14987), .ZN(n10333) );
  NAND2_X1 U10472 ( .A1(n10301), .A2(n7244), .ZN(n12676) );
  INV_X1 U10473 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15397) );
  OR2_X1 U10474 ( .A1(n14281), .A2(n14240), .ZN(n8049) );
  NAND2_X1 U10475 ( .A1(n14308), .A2(n14315), .ZN(n8050) );
  AND2_X1 U10476 ( .A1(n8104), .A2(n8103), .ZN(n8051) );
  NOR2_X1 U10477 ( .A1(n10243), .A2(n11660), .ZN(n9918) );
  AND2_X1 U10478 ( .A1(n12676), .A2(n12677), .ZN(n8052) );
  AND3_X1 U10479 ( .A1(n12687), .A2(n12686), .A3(n12828), .ZN(n8053) );
  OR3_X1 U10480 ( .A1(n9383), .A2(n11051), .A3(n15750), .ZN(n13984) );
  NOR2_X1 U10481 ( .A1(n8120), .A2(n8570), .ZN(n8054) );
  AND2_X1 U10482 ( .A1(n10423), .A2(SI_30_), .ZN(n8055) );
  AND2_X1 U10483 ( .A1(n10085), .A2(n10083), .ZN(n8056) );
  INV_X1 U10484 ( .A(n12862), .ZN(n14825) );
  OR4_X1 U10485 ( .A1(n12621), .A2(n9997), .A3(n14302), .A4(n12934), .ZN(n8057) );
  XNOR2_X1 U10486 ( .A(n14415), .B(n14004), .ZN(n12621) );
  INV_X1 U10487 ( .A(n12606), .ZN(n10015) );
  AND2_X1 U10488 ( .A1(n12455), .A2(n14015), .ZN(n8058) );
  AND2_X1 U10489 ( .A1(n15242), .A2(n10313), .ZN(n8059) );
  INV_X1 U10490 ( .A(n12168), .ZN(n12184) );
  INV_X1 U10491 ( .A(n12620), .ZN(n10270) );
  INV_X1 U10492 ( .A(n12804), .ZN(n14861) );
  NOR3_X1 U10493 ( .A1(n14230), .A2(n14229), .A3(n14380), .ZN(n8061) );
  NAND2_X1 U10494 ( .A1(n14025), .A2(n12381), .ZN(n12374) );
  AND2_X1 U10495 ( .A1(n12547), .A2(n12404), .ZN(n12403) );
  INV_X1 U10496 ( .A(n12448), .ZN(n12444) );
  NAND2_X1 U10497 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  NAND2_X1 U10498 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  NOR2_X1 U10499 ( .A1(n10501), .A2(n6895), .ZN(n10502) );
  AND2_X1 U10500 ( .A1(n10503), .A2(n10502), .ZN(n10504) );
  OAI21_X1 U10501 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(n10518) );
  OAI21_X1 U10502 ( .B1(n7943), .B2(n10564), .A(n10577), .ZN(n10578) );
  AND2_X1 U10503 ( .A1(n11974), .A2(n11972), .ZN(n10136) );
  OR2_X1 U10504 ( .A1(n12934), .A2(n9997), .ZN(n9987) );
  INV_X1 U10505 ( .A(n10578), .ZN(n10579) );
  NAND2_X1 U10506 ( .A1(n9987), .A2(n14379), .ZN(n9988) );
  INV_X1 U10507 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n13598) );
  AOI211_X1 U10508 ( .C1(n10583), .C2(n13322), .A(n10429), .B(n13758), .ZN(
        n10430) );
  NAND2_X1 U10509 ( .A1(n11602), .A2(n10129), .ZN(n10132) );
  NOR2_X1 U10510 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  INV_X1 U10511 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8881) );
  OAI21_X1 U10512 ( .B1(n14628), .B2(n14704), .A(n14626), .ZN(n8541) );
  INV_X1 U10513 ( .A(n12190), .ZN(n8420) );
  INV_X1 U10514 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8532) );
  AND2_X1 U10515 ( .A1(n8791), .A2(n10757), .ZN(n8813) );
  AND2_X1 U10516 ( .A1(n10583), .A2(n10582), .ZN(n10584) );
  INV_X1 U10517 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9724) );
  INV_X1 U10518 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9406) );
  INV_X1 U10519 ( .A(n10033), .ZN(n10030) );
  INV_X1 U10520 ( .A(n14625), .ZN(n8545) );
  INV_X1 U10521 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8472) );
  AND2_X1 U10522 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8163) );
  INV_X1 U10523 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8554) );
  INV_X1 U10524 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10525 ( .A1(n12724), .A2(n10318), .ZN(n10320) );
  INV_X1 U10526 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n13695) );
  NAND2_X1 U10527 ( .A1(n8101), .A2(n10891), .ZN(n8104) );
  OR2_X1 U10528 ( .A1(n9871), .A2(n13401), .ZN(n9869) );
  INV_X1 U10529 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9679) );
  INV_X1 U10530 ( .A(n10791), .ZN(n11349) );
  INV_X1 U10531 ( .A(n11490), .ZN(n10688) );
  OR2_X1 U10532 ( .A1(n13190), .A2(n12202), .ZN(n10609) );
  INV_X1 U10533 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9524) );
  INV_X1 U10534 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15316) );
  INV_X1 U10535 ( .A(n9822), .ZN(n9821) );
  INV_X1 U10536 ( .A(n14336), .ZN(n10026) );
  INV_X1 U10537 ( .A(n10034), .ZN(n10035) );
  OR2_X1 U10538 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  AND2_X1 U10539 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  INV_X1 U10540 ( .A(n14839), .ZN(n14851) );
  INV_X1 U10541 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U10542 ( .A1(n8080), .A2(n13590), .ZN(n8066) );
  INV_X1 U10543 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15332) );
  INV_X1 U10544 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15408) );
  INV_X1 U10545 ( .A(n13027), .ZN(n13079) );
  INV_X1 U10546 ( .A(n13350), .ZN(n13010) );
  NAND2_X1 U10547 ( .A1(n11487), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11864) );
  AND2_X1 U10548 ( .A1(n10713), .A2(n10624), .ZN(n10708) );
  NAND2_X1 U10549 ( .A1(n13350), .A2(n15799), .ZN(n13351) );
  OR2_X1 U10550 ( .A1(n10451), .A2(n10450), .ZN(n13454) );
  INV_X1 U10551 ( .A(n11438), .ZN(n15809) );
  INV_X1 U10552 ( .A(n6423), .ZN(n13358) );
  AND2_X1 U10553 ( .A1(n10245), .A2(n10244), .ZN(n15805) );
  INV_X1 U10554 ( .A(n10059), .ZN(n10060) );
  INV_X1 U10555 ( .A(n14015), .ZN(n11847) );
  INV_X1 U10556 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14097) );
  INV_X1 U10557 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13914) );
  INV_X1 U10558 ( .A(n12619), .ZN(n14209) );
  INV_X1 U10559 ( .A(n12614), .ZN(n12333) );
  INV_X1 U10560 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10290) );
  INV_X1 U10561 ( .A(n12600), .ZN(n11534) );
  XNOR2_X1 U10562 ( .A(n9345), .B(n9344), .ZN(n11050) );
  OR2_X1 U10563 ( .A1(n9338), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9340) );
  AND2_X1 U10564 ( .A1(n8827), .A2(n14685), .ZN(n8828) );
  NAND2_X1 U10565 ( .A1(n8247), .A2(n8246), .ZN(n11123) );
  INV_X1 U10566 ( .A(n14698), .ZN(n14712) );
  AND2_X1 U10567 ( .A1(n12825), .A2(n12820), .ZN(n12818) );
  INV_X1 U10568 ( .A(n8267), .ZN(n8803) );
  INV_X1 U10569 ( .A(n12849), .ZN(n14954) );
  INV_X1 U10570 ( .A(n15070), .ZN(n15073) );
  NAND2_X1 U10571 ( .A1(n15589), .A2(n15588), .ZN(n15572) );
  INV_X1 U10572 ( .A(n15598), .ZN(n15579) );
  NAND2_X1 U10573 ( .A1(n10084), .A2(n8056), .ZN(n10090) );
  INV_X1 U10574 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15313) );
  AND2_X1 U10575 ( .A1(n13086), .A2(n15796), .ZN(n13027) );
  NOR2_X1 U10576 ( .A1(n10260), .A2(n10591), .ZN(n13086) );
  INV_X1 U10577 ( .A(n13319), .ZN(n13290) );
  AND2_X1 U10578 ( .A1(n10708), .A2(n13831), .ZN(n13300) );
  NAND2_X1 U10579 ( .A1(n10241), .A2(n10433), .ZN(n15801) );
  INV_X1 U10580 ( .A(n15812), .ZN(n13532) );
  INV_X1 U10581 ( .A(n15805), .ZN(n15843) );
  INV_X1 U10582 ( .A(n15841), .ZN(n15856) );
  AND2_X1 U10583 ( .A1(n15860), .A2(n15836), .ZN(n13759) );
  NAND2_X1 U10584 ( .A1(n9906), .A2(n9905), .ZN(n10621) );
  INV_X1 U10585 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9412) );
  INV_X1 U10586 ( .A(n13984), .ZN(n13986) );
  INV_X1 U10587 ( .A(n15690), .ZN(n15701) );
  AND2_X1 U10588 ( .A1(n11101), .A2(n12942), .ZN(n15690) );
  AND2_X1 U10589 ( .A1(n11076), .A2(n11075), .ZN(n15707) );
  NAND2_X1 U10590 ( .A1(n15722), .A2(n9372), .ZN(n14385) );
  INV_X1 U10591 ( .A(n14368), .ZN(n14401) );
  AND2_X1 U10592 ( .A1(n15778), .A2(n15750), .ZN(n12108) );
  AND2_X1 U10593 ( .A1(n14337), .A2(n12373), .ZN(n15748) );
  INV_X1 U10594 ( .A(n15748), .ZN(n15764) );
  AND2_X1 U10595 ( .A1(n15723), .A2(n10288), .ZN(n10295) );
  INV_X1 U10596 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8990) );
  AND2_X1 U10597 ( .A1(n14689), .A2(n15598), .ZN(n14714) );
  NAND2_X1 U10598 ( .A1(n8226), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8231) );
  INV_X1 U10599 ( .A(n15475), .ZN(n14765) );
  NOR2_X1 U10600 ( .A1(n10887), .A2(n10881), .ZN(n15475) );
  INV_X1 U10601 ( .A(n14817), .ZN(n15478) );
  AOI21_X1 U10602 ( .B1(n15487), .B2(n10355), .A(n8042), .ZN(n11950) );
  INV_X1 U10603 ( .A(n15549), .ZN(n15117) );
  AND2_X1 U10604 ( .A1(n8792), .A2(n10760), .ZN(n10114) );
  INV_X1 U10605 ( .A(n15604), .ZN(n15558) );
  INV_X1 U10606 ( .A(n10114), .ZN(n11825) );
  XNOR2_X1 U10607 ( .A(n8795), .B(n8794), .ZN(n10719) );
  INV_X1 U10608 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8169) );
  INV_X1 U10609 ( .A(n15378), .ZN(n15379) );
  AND2_X1 U10610 ( .A1(n10713), .A2(n10712), .ZN(n15779) );
  NAND2_X1 U10611 ( .A1(n9930), .A2(n11316), .ZN(n13083) );
  AND2_X1 U10612 ( .A1(n9921), .A2(n9920), .ZN(n13088) );
  INV_X1 U10613 ( .A(n10200), .ZN(n13349) );
  INV_X1 U10614 ( .A(n13315), .ZN(n13282) );
  INV_X1 U10615 ( .A(n13300), .ZN(n13293) );
  OR2_X1 U10616 ( .A1(n10711), .A2(n10709), .ZN(n13319) );
  INV_X1 U10617 ( .A(n13537), .ZN(n13528) );
  NAND2_X2 U10618 ( .A1(n11318), .A2(n13532), .ZN(n15813) );
  INV_X1 U10619 ( .A(n13340), .ZN(n13767) );
  INV_X1 U10620 ( .A(n15860), .ZN(n15858) );
  INV_X1 U10621 ( .A(n13759), .ZN(n13815) );
  INV_X1 U10622 ( .A(n12160), .ZN(n11781) );
  INV_X1 U10623 ( .A(SI_13_), .ZN(n10891) );
  INV_X1 U10624 ( .A(n13822), .ZN(n13838) );
  NOR2_X1 U10625 ( .A1(n10596), .A2(n12099), .ZN(n11053) );
  INV_X1 U10626 ( .A(n13873), .ZN(n13993) );
  OR2_X1 U10627 ( .A1(n13952), .A2(n14331), .ZN(n13991) );
  INV_X1 U10628 ( .A(n13998), .ZN(n13973) );
  AND4_X1 U10629 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12649) );
  NAND2_X1 U10630 ( .A1(n9298), .A2(n9297), .ZN(n14006) );
  INV_X1 U10631 ( .A(n15634), .ZN(n15715) );
  NAND2_X1 U10632 ( .A1(n14396), .A2(n10043), .ZN(n14371) );
  OR2_X1 U10633 ( .A1(n14352), .A2(n11569), .ZN(n14348) );
  INV_X1 U10634 ( .A(n12108), .ZN(n14487) );
  INV_X1 U10635 ( .A(n14277), .ZN(n14533) );
  INV_X1 U10636 ( .A(n12114), .ZN(n14551) );
  INV_X1 U10637 ( .A(n15767), .ZN(n15765) );
  NOR2_X1 U10638 ( .A1(n15724), .A2(n15716), .ZN(n15718) );
  INV_X1 U10639 ( .A(n15718), .ZN(n15719) );
  INV_X1 U10640 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11206) );
  CLKBUF_X1 U10641 ( .A(n14569), .Z(n12913) );
  NAND2_X1 U10642 ( .A1(n8799), .A2(n8798), .ZN(n14717) );
  INV_X1 U10643 ( .A(n14677), .ZN(n14728) );
  INV_X1 U10644 ( .A(n15479), .ZN(n14805) );
  NAND2_X1 U10645 ( .A1(n15513), .A2(n11829), .ZN(n15096) );
  INV_X1 U10646 ( .A(n15100), .ZN(n15529) );
  INV_X1 U10647 ( .A(n15618), .ZN(n15615) );
  INV_X1 U10648 ( .A(n14826), .ZN(n15249) );
  INV_X1 U10649 ( .A(n14715), .ZN(n15281) );
  INV_X1 U10650 ( .A(n15606), .ZN(n15605) );
  AND2_X2 U10651 ( .A1(n10115), .A2(n11825), .ZN(n15606) );
  AND2_X1 U10652 ( .A1(n10719), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10761) );
  XNOR2_X1 U10653 ( .A(n8158), .B(n8157), .ZN(n12229) );
  INV_X1 U10654 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11410) );
  INV_X1 U10655 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10980) );
  AND2_X2 U10656 ( .A1(n10600), .A2(n13816), .ZN(P3_U3897) );
  AND2_X1 U10657 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11053), .ZN(P2_U3947) );
  NAND2_X1 U10658 ( .A1(n8073), .A2(SI_2_), .ZN(n8275) );
  INV_X1 U10659 ( .A(SI_3_), .ZN(n10792) );
  NAND2_X1 U10660 ( .A1(n8275), .A2(n10792), .ZN(n8067) );
  INV_X1 U10661 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10784) );
  MUX2_X1 U10662 ( .A(n10784), .B(n10741), .S(n8080), .Z(n8068) );
  INV_X1 U10663 ( .A(n8068), .ZN(n8278) );
  NAND2_X1 U10664 ( .A1(n8067), .A2(n8278), .ZN(n8303) );
  NAND2_X1 U10665 ( .A1(n8068), .A2(n10792), .ZN(n8071) );
  AND2_X1 U10666 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8069) );
  AND2_X1 U10667 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8070) );
  INV_X1 U10668 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10776) );
  INV_X1 U10669 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10748) );
  AND2_X1 U10670 ( .A1(SI_2_), .A2(SI_3_), .ZN(n8072) );
  NAND2_X1 U10671 ( .A1(n8073), .A2(n8072), .ZN(n8302) );
  XNOR2_X1 U10672 ( .A(n8078), .B(SI_5_), .ZN(n8335) );
  NOR2_X1 U10673 ( .A1(n8075), .A2(SI_4_), .ZN(n8076) );
  NOR2_X1 U10674 ( .A1(n8335), .A2(n8076), .ZN(n8077) );
  NAND2_X1 U10675 ( .A1(n8078), .A2(SI_5_), .ZN(n8079) );
  NAND2_X1 U10676 ( .A1(n8081), .A2(SI_6_), .ZN(n8082) );
  MUX2_X1 U10677 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10768), .Z(n8084) );
  XNOR2_X1 U10678 ( .A(n8084), .B(SI_7_), .ZN(n8361) );
  INV_X1 U10679 ( .A(n8361), .ZN(n8083) );
  NAND2_X1 U10680 ( .A1(n8084), .A2(SI_7_), .ZN(n8085) );
  MUX2_X1 U10681 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10071), .Z(n8086) );
  NAND2_X1 U10682 ( .A1(n8086), .A2(SI_8_), .ZN(n8087) );
  MUX2_X1 U10683 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10071), .Z(n8089) );
  INV_X1 U10684 ( .A(n8401), .ZN(n8088) );
  NAND2_X1 U10685 ( .A1(n8089), .A2(SI_9_), .ZN(n8090) );
  MUX2_X1 U10686 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10071), .Z(n8423) );
  INV_X1 U10687 ( .A(SI_10_), .ZN(n10871) );
  NAND2_X1 U10688 ( .A1(n8423), .A2(SI_10_), .ZN(n8092) );
  MUX2_X1 U10689 ( .A(n10866), .B(n10867), .S(n10768), .Z(n8093) );
  NAND2_X1 U10690 ( .A1(n8093), .A2(n10863), .ZN(n8096) );
  INV_X1 U10691 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U10692 ( .A1(n8094), .A2(SI_11_), .ZN(n8095) );
  NAND2_X1 U10693 ( .A1(n8096), .A2(n8095), .ZN(n8442) );
  MUX2_X1 U10694 ( .A(n10914), .B(n10912), .S(n10768), .Z(n8097) );
  NAND2_X1 U10695 ( .A1(n8097), .A2(n10860), .ZN(n8100) );
  INV_X1 U10696 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U10697 ( .A1(n8098), .A2(SI_12_), .ZN(n8099) );
  MUX2_X1 U10698 ( .A(n10980), .B(n13593), .S(n10768), .Z(n8101) );
  INV_X1 U10699 ( .A(n8101), .ZN(n8102) );
  NAND2_X1 U10700 ( .A1(n8102), .A2(SI_13_), .ZN(n8103) );
  MUX2_X1 U10701 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10071), .Z(n8501) );
  INV_X1 U10702 ( .A(n8522), .ZN(n8105) );
  MUX2_X1 U10703 ( .A(n11258), .B(n11308), .S(n10768), .Z(n8106) );
  INV_X1 U10704 ( .A(n8106), .ZN(n8107) );
  NAND2_X1 U10705 ( .A1(n8107), .A2(SI_15_), .ZN(n8108) );
  NAND2_X1 U10706 ( .A1(n8523), .A2(n8108), .ZN(n8503) );
  INV_X1 U10707 ( .A(n8501), .ZN(n8109) );
  NOR2_X1 U10708 ( .A1(n8109), .A2(n10972), .ZN(n8110) );
  INV_X1 U10709 ( .A(n8521), .ZN(n8114) );
  MUX2_X1 U10710 ( .A(n11121), .B(n11132), .S(n10071), .Z(n8111) );
  NAND2_X1 U10711 ( .A1(n8111), .A2(n10957), .ZN(n8546) );
  INV_X1 U10712 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U10713 ( .A1(n8112), .A2(SI_16_), .ZN(n8113) );
  NAND2_X1 U10714 ( .A1(n8546), .A2(n8113), .ZN(n8525) );
  MUX2_X1 U10715 ( .A(n11306), .B(n11323), .S(n10768), .Z(n8118) );
  INV_X1 U10716 ( .A(SI_17_), .ZN(n8116) );
  NAND2_X1 U10717 ( .A1(n8118), .A2(n8116), .ZN(n8547) );
  MUX2_X1 U10718 ( .A(n9768), .B(n11360), .S(n10768), .Z(n8572) );
  INV_X1 U10719 ( .A(n8120), .ZN(n8117) );
  INV_X1 U10720 ( .A(n8118), .ZN(n8119) );
  MUX2_X1 U10721 ( .A(n11410), .B(n11408), .S(n10071), .Z(n8122) );
  INV_X1 U10722 ( .A(n8122), .ZN(n8123) );
  NAND2_X1 U10723 ( .A1(n8123), .A2(SI_19_), .ZN(n8124) );
  MUX2_X1 U10724 ( .A(n11543), .B(n11541), .S(n10768), .Z(n8616) );
  XNOR2_X1 U10725 ( .A(n8616), .B(SI_20_), .ZN(n8126) );
  XNOR2_X1 U10726 ( .A(n8617), .B(n8126), .ZN(n11540) );
  NOR2_X1 U10727 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8129) );
  NOR2_X2 U10728 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8128) );
  NOR2_X2 U10729 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8127) );
  AND4_X2 U10730 ( .A1(n8129), .A2(n8128), .A3(n8127), .A4(n8331), .ZN(n8131)
         );
  NOR2_X2 U10731 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8197) );
  AND2_X2 U10732 ( .A1(n8197), .A2(n8130), .ZN(n8463) );
  NOR2_X2 U10733 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8134) );
  NAND4_X2 U10734 ( .A1(n8134), .A2(n11181), .A3(n8133), .A4(n8132), .ZN(n8329) );
  NAND4_X1 U10735 ( .A1(n8136), .A2(n8185), .A3(n8184), .A4(n8135), .ZN(n8137)
         );
  INV_X1 U10736 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10737 ( .A1(n8150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10738 ( .A1(n11540), .A2(n10091), .ZN(n8145) );
  NAND2_X1 U10739 ( .A1(n6422), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8144) );
  AND2_X2 U10740 ( .A1(n8145), .A2(n8144), .ZN(n15271) );
  INV_X1 U10741 ( .A(n8146), .ZN(n8147) );
  NAND2_X1 U10742 ( .A1(n8152), .A2(n8148), .ZN(n8154) );
  NAND2_X1 U10743 ( .A1(n8154), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U10744 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8149), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8151) );
  NAND2_X1 U10745 ( .A1(n7351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10746 ( .A1(n8155), .A2(n8154), .ZN(n12284) );
  NAND2_X1 U10747 ( .A1(n8156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10748 ( .A1(n8178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8159) );
  XNOR2_X2 U10749 ( .A(n8159), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U10750 ( .A1(n8160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8162) );
  INV_X1 U10751 ( .A(n12670), .ZN(n12816) );
  OR2_X1 U10752 ( .A1(n15271), .A2(n8644), .ZN(n8182) );
  INV_X1 U10753 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8597) );
  INV_X1 U10754 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10755 ( .A1(n8600), .A2(n8164), .ZN(n8165) );
  NAND2_X1 U10756 ( .A1(n8636), .A2(n8165), .ZN(n14992) );
  INV_X1 U10757 ( .A(n14992), .ZN(n14653) );
  NAND2_X1 U10758 ( .A1(n14653), .A2(n8803), .ZN(n8177) );
  INV_X1 U10759 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U10760 ( .A1(n12656), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10761 ( .A1(n12657), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8173) );
  OAI211_X1 U10762 ( .C1(n12660), .C2(n15177), .A(n8174), .B(n8173), .ZN(n8175) );
  INV_X1 U10763 ( .A(n8175), .ZN(n8176) );
  INV_X1 U10764 ( .A(n14611), .ZN(n14727) );
  INV_X1 U10765 ( .A(n12651), .ZN(n8188) );
  OR2_X4 U10766 ( .A1(n12814), .A2(n8801), .ZN(n15517) );
  NAND2_X1 U10767 ( .A1(n14727), .A2(n8292), .ZN(n8181) );
  NAND2_X1 U10768 ( .A1(n8182), .A2(n8181), .ZN(n8615) );
  OAI22_X1 U10769 ( .A1(n15271), .A2(n8645), .B1(n14611), .B2(n8644), .ZN(
        n8190) );
  OR2_X1 U10770 ( .A1(n8188), .A2(n12652), .ZN(n8189) );
  XNOR2_X1 U10771 ( .A(n8190), .B(n8755), .ZN(n8614) );
  NAND2_X1 U10772 ( .A1(n8194), .A2(n8193), .ZN(n10911) );
  NAND2_X1 U10773 ( .A1(n10911), .A2(n10091), .ZN(n8202) );
  NAND2_X1 U10774 ( .A1(n7490), .A2(n8331), .ZN(n8351) );
  INV_X1 U10775 ( .A(n8363), .ZN(n8196) );
  NAND2_X1 U10776 ( .A1(n8196), .A2(n8195), .ZN(n8385) );
  INV_X1 U10777 ( .A(n8197), .ZN(n8198) );
  NAND2_X1 U10778 ( .A1(n8198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U10779 ( .A1(n8465), .A2(n8199), .ZN(n8443) );
  NAND2_X1 U10780 ( .A1(n8445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U10781 ( .A(n8200), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U10782 ( .A1(n6422), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11460), 
        .B2(n8594), .ZN(n8201) );
  NAND2_X1 U10783 ( .A1(n12657), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8208) );
  INV_X1 U10784 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8203) );
  OR2_X1 U10785 ( .A1(n12660), .A2(n8203), .ZN(n8207) );
  NAND2_X1 U10786 ( .A1(n8450), .A2(n13649), .ZN(n8204) );
  NAND2_X1 U10787 ( .A1(n8473), .A2(n8204), .ZN(n12311) );
  OR2_X1 U10788 ( .A1(n8267), .A2(n12311), .ZN(n8206) );
  INV_X1 U10789 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12312) );
  OR2_X1 U10790 ( .A1(n8296), .A2(n12312), .ZN(n8205) );
  NAND4_X1 U10791 ( .A1(n8208), .A2(n8207), .A3(n8206), .A4(n8205), .ZN(n14736) );
  AND2_X1 U10792 ( .A1(n14736), .A2(n8292), .ZN(n8209) );
  AOI21_X1 U10793 ( .B1(n12724), .B2(n8732), .A(n8209), .ZN(n8461) );
  NAND2_X1 U10794 ( .A1(n12724), .A2(n8775), .ZN(n8211) );
  NAND2_X1 U10795 ( .A1(n14736), .A2(n6415), .ZN(n8210) );
  NAND2_X1 U10796 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  XNOR2_X1 U10797 ( .A(n8212), .B(n8755), .ZN(n8457) );
  INV_X1 U10798 ( .A(n8457), .ZN(n8460) );
  INV_X1 U10799 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15115) );
  OR2_X1 U10800 ( .A1(n8267), .A2(n15115), .ZN(n8214) );
  INV_X1 U10801 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8213) );
  INV_X1 U10802 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10839) );
  NAND2_X1 U10803 ( .A1(n14747), .A2(n8292), .ZN(n8222) );
  INV_X1 U10804 ( .A(SI_1_), .ZN(n10775) );
  XNOR2_X1 U10805 ( .A(n8216), .B(n10775), .ZN(n8218) );
  XNOR2_X1 U10806 ( .A(n8218), .B(n8217), .ZN(n10777) );
  INV_X1 U10807 ( .A(n10777), .ZN(n8219) );
  NAND2_X1 U10808 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8220) );
  XNOR2_X1 U10809 ( .A(n8220), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10730) );
  OR2_X1 U10810 ( .A1(n15549), .A2(n8644), .ZN(n8221) );
  NAND2_X1 U10811 ( .A1(n10302), .A2(n6415), .ZN(n8224) );
  INV_X1 U10812 ( .A(n11122), .ZN(n8247) );
  INV_X1 U10813 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10885) );
  OR2_X1 U10814 ( .A1(n8267), .A2(n10885), .ZN(n8230) );
  INV_X1 U10815 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10879) );
  OR2_X1 U10816 ( .A1(n8227), .A2(n10879), .ZN(n8229) );
  NAND2_X1 U10817 ( .A1(n15105), .A2(n8292), .ZN(n8238) );
  INV_X1 U10818 ( .A(SI_0_), .ZN(n8232) );
  INV_X1 U10819 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9456) );
  OAI21_X1 U10820 ( .B1(n10071), .B2(n8232), .A(n9456), .ZN(n8233) );
  NAND2_X1 U10821 ( .A1(n8234), .A2(n8233), .ZN(n15310) );
  OAI22_X1 U10822 ( .A1(n15525), .A2(n8644), .B1(n11181), .B2(n10597), .ZN(
        n8236) );
  INV_X1 U10823 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U10824 ( .A1(n8238), .A2(n8237), .ZN(n11172) );
  NAND2_X1 U10825 ( .A1(n15105), .A2(n6415), .ZN(n8243) );
  INV_X1 U10826 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8240) );
  OAI22_X1 U10827 ( .A1(n15525), .A2(n8645), .B1(n8240), .B2(n10597), .ZN(
        n8241) );
  INV_X1 U10828 ( .A(n8241), .ZN(n8242) );
  NAND2_X1 U10829 ( .A1(n8243), .A2(n8242), .ZN(n11171) );
  NAND2_X1 U10830 ( .A1(n8245), .A2(n8244), .ZN(n11125) );
  INV_X1 U10831 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10849) );
  OR2_X1 U10832 ( .A1(n8296), .A2(n10849), .ZN(n8250) );
  INV_X1 U10833 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U10834 ( .A1(n8470), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10835 ( .A1(n14746), .A2(n6415), .ZN(n8259) );
  XNOR2_X1 U10836 ( .A(n8251), .B(SI_2_), .ZN(n8273) );
  XNOR2_X1 U10837 ( .A(n8274), .B(n8273), .ZN(n10778) );
  INV_X1 U10838 ( .A(n10778), .ZN(n8252) );
  NAND2_X1 U10839 ( .A1(n8355), .A2(n8252), .ZN(n8257) );
  NAND2_X1 U10840 ( .A1(n6420), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8256) );
  INV_X1 U10841 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8253) );
  INV_X1 U10842 ( .A(n14751), .ZN(n8254) );
  AND3_X2 U10843 ( .A1(n8257), .A2(n8256), .A3(n8255), .ZN(n11204) );
  OR2_X1 U10844 ( .A1(n11204), .A2(n8645), .ZN(n8258) );
  NAND2_X1 U10845 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  XNOR2_X1 U10846 ( .A(n8260), .B(n10397), .ZN(n8265) );
  NAND2_X1 U10847 ( .A1(n14746), .A2(n8292), .ZN(n8262) );
  OR2_X1 U10848 ( .A1(n11204), .A2(n8644), .ZN(n8261) );
  NAND2_X1 U10849 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XNOR2_X1 U10850 ( .A(n8265), .B(n8263), .ZN(n11197) );
  INV_X1 U10851 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U10852 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  NAND2_X1 U10853 ( .A1(n8226), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8272) );
  OR2_X1 U10854 ( .A1(n8267), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8271) );
  INV_X1 U10855 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n15512) );
  OR2_X1 U10856 ( .A1(n8296), .A2(n15512), .ZN(n8270) );
  INV_X1 U10857 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8268) );
  OR2_X1 U10858 ( .A1(n10097), .A2(n8268), .ZN(n8269) );
  NAND2_X1 U10859 ( .A1(n14745), .A2(n6415), .ZN(n8290) );
  INV_X1 U10860 ( .A(n8273), .ZN(n8277) );
  INV_X1 U10861 ( .A(n8274), .ZN(n8276) );
  OAI21_X1 U10862 ( .B1(n8277), .B2(n8276), .A(n8275), .ZN(n8280) );
  XNOR2_X1 U10863 ( .A(n8278), .B(SI_3_), .ZN(n8279) );
  XNOR2_X1 U10864 ( .A(n8280), .B(n8279), .ZN(n10740) );
  NAND2_X1 U10865 ( .A1(n8355), .A2(n10740), .ZN(n8288) );
  INV_X1 U10866 ( .A(n8281), .ZN(n8283) );
  INV_X1 U10867 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U10868 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  NAND2_X1 U10869 ( .A1(n8285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8284) );
  MUX2_X1 U10870 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8284), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8286) );
  OR2_X1 U10871 ( .A1(n8285), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8307) );
  AND2_X1 U10872 ( .A1(n8286), .A2(n8307), .ZN(n10851) );
  NAND2_X1 U10873 ( .A1(n8594), .A2(n10851), .ZN(n8287) );
  OAI211_X2 U10874 ( .C1(n8301), .C2(n10784), .A(n8288), .B(n8287), .ZN(n15564) );
  NAND2_X1 U10875 ( .A1(n15564), .A2(n8775), .ZN(n8289) );
  NAND2_X1 U10876 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  XNOR2_X1 U10877 ( .A(n8291), .B(n8755), .ZN(n8293) );
  AOI22_X1 U10878 ( .A1(n14745), .A2(n8292), .B1(n6415), .B2(n15564), .ZN(
        n8294) );
  XNOR2_X1 U10879 ( .A(n8293), .B(n8294), .ZN(n11210) );
  INV_X1 U10880 ( .A(n8293), .ZN(n8295) );
  OR2_X1 U10881 ( .A1(n8295), .A2(n8294), .ZN(n8320) );
  NAND2_X1 U10882 ( .A1(n12657), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8300) );
  INV_X1 U10883 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10842) );
  OAI21_X1 U10884 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8323), .ZN(n11965) );
  OR2_X1 U10885 ( .A1(n8267), .A2(n11965), .ZN(n8298) );
  INV_X1 U10886 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10853) );
  OR2_X1 U10887 ( .A1(n8296), .A2(n10853), .ZN(n8297) );
  NAND4_X2 U10888 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n14744) );
  NAND2_X1 U10889 ( .A1(n14744), .A2(n8292), .ZN(n8312) );
  NAND3_X1 U10890 ( .A1(n8304), .A2(n8303), .A3(n8302), .ZN(n8333) );
  XNOR2_X1 U10891 ( .A(n8305), .B(SI_4_), .ZN(n8332) );
  INV_X1 U10892 ( .A(n8332), .ZN(n8306) );
  XNOR2_X1 U10893 ( .A(n8333), .B(n8306), .ZN(n10742) );
  NAND2_X1 U10894 ( .A1(n8355), .A2(n10742), .ZN(n8310) );
  NAND2_X1 U10895 ( .A1(n8307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U10896 ( .A(n8308), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U10897 ( .A1(n8594), .A2(n10852), .ZN(n8309) );
  NAND2_X1 U10898 ( .A1(n15569), .A2(n8239), .ZN(n8311) );
  NAND2_X1 U10899 ( .A1(n8312), .A2(n8311), .ZN(n8318) );
  NAND2_X1 U10900 ( .A1(n14744), .A2(n6415), .ZN(n8315) );
  NAND2_X1 U10901 ( .A1(n15569), .A2(n8775), .ZN(n8314) );
  NAND2_X1 U10902 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  XNOR2_X1 U10903 ( .A(n8316), .B(n10397), .ZN(n11373) );
  INV_X1 U10904 ( .A(n8318), .ZN(n8319) );
  AND2_X1 U10905 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  NAND2_X1 U10906 ( .A1(n12657), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10907 ( .A1(n8323), .A2(n6676), .ZN(n8324) );
  NAND2_X1 U10908 ( .A1(n8345), .A2(n8324), .ZN(n15493) );
  OR2_X1 U10909 ( .A1(n8267), .A2(n15493), .ZN(n8327) );
  INV_X1 U10910 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10847) );
  OR2_X1 U10911 ( .A1(n8296), .A2(n10847), .ZN(n8326) );
  INV_X1 U10912 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10896) );
  OR2_X1 U10913 ( .A1(n12660), .A2(n10896), .ZN(n8325) );
  NAND2_X1 U10914 ( .A1(n14743), .A2(n6415), .ZN(n8340) );
  NAND2_X1 U10915 ( .A1(n8329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8330) );
  XNOR2_X1 U10916 ( .A(n8331), .B(n8330), .ZN(n10895) );
  NAND2_X1 U10917 ( .A1(n8333), .A2(n8332), .ZN(n8334) );
  XNOR2_X1 U10918 ( .A(n8336), .B(n8335), .ZN(n10752) );
  NAND2_X1 U10919 ( .A1(n10752), .A2(n8355), .ZN(n8338) );
  NAND2_X1 U10920 ( .A1(n6420), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8337) );
  OAI211_X2 U10921 ( .C1(n8235), .C2(n10895), .A(n8338), .B(n8337), .ZN(n15495) );
  NAND2_X1 U10922 ( .A1(n15495), .A2(n8775), .ZN(n8339) );
  NAND2_X1 U10923 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  XNOR2_X1 U10924 ( .A(n8341), .B(n10397), .ZN(n8343) );
  AOI22_X1 U10925 ( .A1(n14743), .A2(n8292), .B1(n8732), .B2(n15495), .ZN(
        n8342) );
  OR2_X1 U10926 ( .A1(n8343), .A2(n8342), .ZN(n11411) );
  NAND2_X1 U10927 ( .A1(n8226), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8350) );
  INV_X1 U10928 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8344) );
  OR2_X1 U10929 ( .A1(n10097), .A2(n8344), .ZN(n8349) );
  NAND2_X1 U10930 ( .A1(n8345), .A2(n6677), .ZN(n8346) );
  NAND2_X1 U10931 ( .A1(n8369), .A2(n8346), .ZN(n14690) );
  OR2_X1 U10932 ( .A1(n8267), .A2(n14690), .ZN(n8348) );
  INV_X1 U10933 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11955) );
  OR2_X1 U10934 ( .A1(n8296), .A2(n11955), .ZN(n8347) );
  NAND2_X1 U10935 ( .A1(n8351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8352) );
  XNOR2_X1 U10936 ( .A(n8352), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U10937 ( .A1(n6422), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8594), .B2(
        n10899), .ZN(n8357) );
  XNOR2_X1 U10938 ( .A(n8354), .B(n8353), .ZN(n10746) );
  NAND2_X1 U10939 ( .A1(n10746), .A2(n8355), .ZN(n8356) );
  OAI22_X1 U10940 ( .A1(n12699), .A2(n8644), .B1(n14688), .B2(n8645), .ZN(
        n8358) );
  XNOR2_X1 U10941 ( .A(n8358), .B(n8755), .ZN(n8360) );
  OAI22_X1 U10942 ( .A1(n12699), .A2(n8643), .B1(n14688), .B2(n8644), .ZN(
        n8359) );
  OR2_X1 U10943 ( .A1(n8360), .A2(n8359), .ZN(n14682) );
  XNOR2_X1 U10944 ( .A(n8362), .B(n8361), .ZN(n10744) );
  NAND2_X1 U10945 ( .A1(n10744), .A2(n10091), .ZN(n8366) );
  NAND2_X1 U10946 ( .A1(n8363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8364) );
  XNOR2_X1 U10947 ( .A(n8364), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U10948 ( .A1(n6422), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8594), .B2(
        n10920), .ZN(n8365) );
  NAND2_X1 U10949 ( .A1(n15597), .A2(n8775), .ZN(n8376) );
  NAND2_X1 U10950 ( .A1(n8226), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8374) );
  INV_X1 U10951 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8367) );
  OR2_X1 U10952 ( .A1(n10097), .A2(n8367), .ZN(n8373) );
  NAND2_X1 U10953 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U10954 ( .A1(n8391), .A2(n8370), .ZN(n11944) );
  OR2_X1 U10955 ( .A1(n8267), .A2(n11944), .ZN(n8372) );
  INV_X1 U10956 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11942) );
  OR2_X1 U10957 ( .A1(n8296), .A2(n11942), .ZN(n8371) );
  NAND4_X1 U10958 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n14741) );
  NAND2_X1 U10959 ( .A1(n14741), .A2(n8239), .ZN(n8375) );
  NAND2_X1 U10960 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  XNOR2_X1 U10961 ( .A(n8377), .B(n8755), .ZN(n8381) );
  NAND2_X1 U10962 ( .A1(n15597), .A2(n8239), .ZN(n8379) );
  NAND2_X1 U10963 ( .A1(n14741), .A2(n8292), .ZN(n8378) );
  NAND2_X1 U10964 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  XNOR2_X1 U10965 ( .A(n8381), .B(n8380), .ZN(n11707) );
  NAND2_X1 U10966 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  XNOR2_X1 U10967 ( .A(n8384), .B(n8383), .ZN(n10764) );
  NAND2_X1 U10968 ( .A1(n10764), .A2(n10091), .ZN(n8389) );
  NAND2_X1 U10969 ( .A1(n8385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8386) );
  MUX2_X1 U10970 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8386), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n8387) );
  AND2_X1 U10971 ( .A1(n8387), .A2(n8507), .ZN(n10946) );
  AOI22_X1 U10972 ( .A1(n6422), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8594), .B2(
        n10946), .ZN(n8388) );
  NAND2_X1 U10973 ( .A1(n8389), .A2(n8388), .ZN(n12706) );
  NAND2_X1 U10974 ( .A1(n12706), .A2(n8775), .ZN(n8398) );
  NAND2_X1 U10975 ( .A1(n12657), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8396) );
  INV_X1 U10976 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12010) );
  OR2_X1 U10977 ( .A1(n8296), .A2(n12010), .ZN(n8395) );
  NAND2_X1 U10978 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  NAND2_X1 U10979 ( .A1(n8408), .A2(n8392), .ZN(n12012) );
  OR2_X1 U10980 ( .A1(n8267), .A2(n12012), .ZN(n8394) );
  INV_X1 U10981 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10921) );
  OR2_X1 U10982 ( .A1(n12660), .A2(n10921), .ZN(n8393) );
  NAND4_X1 U10983 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n14740) );
  NAND2_X1 U10984 ( .A1(n14740), .A2(n8732), .ZN(n8397) );
  NAND2_X1 U10985 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  XNOR2_X1 U10986 ( .A(n8399), .B(n10397), .ZN(n11904) );
  AND2_X1 U10987 ( .A1(n14740), .A2(n8292), .ZN(n8400) );
  AOI21_X1 U10988 ( .B1(n12706), .B2(n8732), .A(n8400), .ZN(n11905) );
  NOR2_X1 U10989 ( .A1(n11904), .A2(n11905), .ZN(n8421) );
  XNOR2_X1 U10990 ( .A(n8402), .B(n8401), .ZN(n10796) );
  NAND2_X1 U10991 ( .A1(n10796), .A2(n10091), .ZN(n8407) );
  NAND2_X1 U10992 ( .A1(n8403), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8405) );
  INV_X1 U10993 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U10994 ( .A1(n8465), .A2(n8404), .ZN(n8425) );
  AOI22_X1 U10995 ( .A1(n6422), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8594), .B2(
        n10949), .ZN(n8406) );
  NAND2_X1 U10996 ( .A1(n15242), .A2(n8775), .ZN(n8416) );
  NAND2_X1 U10997 ( .A1(n12657), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8414) );
  INV_X1 U10998 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n13696) );
  OR2_X1 U10999 ( .A1(n12660), .A2(n13696), .ZN(n8413) );
  NAND2_X1 U11000 ( .A1(n8408), .A2(n13694), .ZN(n8409) );
  NAND2_X1 U11001 ( .A1(n8449), .A2(n8409), .ZN(n12169) );
  OR2_X1 U11002 ( .A1(n8267), .A2(n12169), .ZN(n8412) );
  INV_X1 U11003 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8410) );
  OR2_X1 U11004 ( .A1(n8296), .A2(n8410), .ZN(n8411) );
  NAND4_X1 U11005 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(n14739) );
  NAND2_X1 U11006 ( .A1(n14739), .A2(n8732), .ZN(n8415) );
  NAND2_X1 U11007 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  XNOR2_X1 U11008 ( .A(n8417), .B(n8755), .ZN(n12054) );
  NAND2_X1 U11009 ( .A1(n15242), .A2(n8732), .ZN(n8419) );
  NAND2_X1 U11010 ( .A1(n14739), .A2(n8292), .ZN(n8418) );
  NAND2_X1 U11011 ( .A1(n8419), .A2(n8418), .ZN(n8422) );
  NAND2_X1 U11012 ( .A1(n12054), .A2(n8422), .ZN(n12190) );
  INV_X1 U11013 ( .A(n8422), .ZN(n12053) );
  NAND2_X1 U11014 ( .A1(n11904), .A2(n11905), .ZN(n12055) );
  INV_X1 U11015 ( .A(n12055), .ZN(n12051) );
  AOI21_X1 U11016 ( .B1(n8422), .B2(n12055), .A(n12054), .ZN(n8437) );
  XNOR2_X1 U11017 ( .A(n8423), .B(SI_10_), .ZN(n8424) );
  NAND2_X1 U11018 ( .A1(n10833), .A2(n10091), .ZN(n8428) );
  NAND2_X1 U11019 ( .A1(n8425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8426) );
  XNOR2_X1 U11020 ( .A(n8426), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U11021 ( .A1(n6422), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8594), 
        .B2(n11139), .ZN(n8427) );
  NAND2_X2 U11022 ( .A1(n8428), .A2(n8427), .ZN(n15234) );
  NAND2_X1 U11023 ( .A1(n8226), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8433) );
  INV_X1 U11024 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8429) );
  OR2_X1 U11025 ( .A1(n10097), .A2(n8429), .ZN(n8432) );
  INV_X1 U11026 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U11027 ( .A(n8449), .B(n8448), .ZN(n12196) );
  OR2_X1 U11028 ( .A1(n8267), .A2(n12196), .ZN(n8431) );
  INV_X1 U11029 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12183) );
  OR2_X1 U11030 ( .A1(n8296), .A2(n12183), .ZN(n8430) );
  NAND4_X1 U11031 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n14738) );
  AOI22_X1 U11032 ( .A1(n15234), .A2(n6415), .B1(n8292), .B2(n14738), .ZN(
        n8438) );
  NAND2_X1 U11033 ( .A1(n15234), .A2(n8775), .ZN(n8435) );
  NAND2_X1 U11034 ( .A1(n14738), .A2(n8732), .ZN(n8434) );
  NAND2_X1 U11035 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  XNOR2_X1 U11036 ( .A(n8436), .B(n8755), .ZN(n8440) );
  XOR2_X1 U11037 ( .A(n8438), .B(n8440), .Z(n12193) );
  AOI211_X1 U11038 ( .C1(n12053), .C2(n12051), .A(n8437), .B(n12193), .ZN(
        n8441) );
  INV_X1 U11039 ( .A(n8438), .ZN(n8439) );
  NAND2_X1 U11040 ( .A1(n8443), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8444) );
  AOI22_X1 U11041 ( .A1(n6422), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8594), 
        .B2(n11285), .ZN(n8446) );
  NAND2_X1 U11042 ( .A1(n12657), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8455) );
  INV_X1 U11043 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11283) );
  OR2_X1 U11044 ( .A1(n12660), .A2(n11283), .ZN(n8454) );
  INV_X1 U11045 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8447) );
  OAI21_X1 U11046 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8451) );
  NAND2_X1 U11047 ( .A1(n8451), .A2(n8450), .ZN(n12275) );
  OR2_X1 U11048 ( .A1(n8267), .A2(n12275), .ZN(n8453) );
  INV_X1 U11049 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12276) );
  OR2_X1 U11050 ( .A1(n8296), .A2(n12276), .ZN(n8452) );
  NAND4_X1 U11051 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n14737) );
  AOI22_X1 U11052 ( .A1(n15291), .A2(n8732), .B1(n8292), .B2(n14737), .ZN(
        n8458) );
  AOI22_X1 U11053 ( .A1(n15291), .A2(n8775), .B1(n8732), .B2(n14737), .ZN(
        n8456) );
  XNOR2_X1 U11054 ( .A(n8456), .B(n8755), .ZN(n8459) );
  XOR2_X1 U11055 ( .A(n8458), .B(n8459), .Z(n12218) );
  XNOR2_X1 U11056 ( .A(n8457), .B(n8461), .ZN(n12254) );
  NAND2_X1 U11057 ( .A1(n8459), .A2(n8458), .ZN(n12251) );
  XNOR2_X1 U11058 ( .A(n8462), .B(n8051), .ZN(n10979) );
  NAND2_X1 U11059 ( .A1(n10979), .A2(n10091), .ZN(n8469) );
  INV_X1 U11060 ( .A(n8463), .ZN(n8505) );
  NAND2_X1 U11061 ( .A1(n8505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U11062 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U11063 ( .A1(n8466), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n8467) );
  AOI22_X1 U11064 ( .A1(n6422), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8594), 
        .B2(n11684), .ZN(n8468) );
  NAND2_X1 U11065 ( .A1(n12657), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8478) );
  INV_X1 U11066 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11463) );
  OR2_X1 U11067 ( .A1(n8296), .A2(n11463), .ZN(n8477) );
  INV_X1 U11068 ( .A(n8471), .ZN(n8486) );
  NAND2_X1 U11069 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  NAND2_X1 U11070 ( .A1(n8486), .A2(n8474), .ZN(n12353) );
  OR2_X1 U11071 ( .A1(n8267), .A2(n12353), .ZN(n8476) );
  INV_X1 U11072 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15220) );
  OR2_X1 U11073 ( .A1(n12660), .A2(n15220), .ZN(n8475) );
  OAI22_X1 U11074 ( .A1(n15286), .A2(n8644), .B1(n14584), .B2(n8643), .ZN(
        n8481) );
  OAI22_X1 U11075 ( .A1(n15286), .A2(n8645), .B1(n14584), .B2(n8644), .ZN(
        n8479) );
  XNOR2_X1 U11076 ( .A(n8479), .B(n8755), .ZN(n8480) );
  XOR2_X1 U11077 ( .A(n8481), .B(n8480), .Z(n12299) );
  XNOR2_X1 U11078 ( .A(n8502), .B(n8501), .ZN(n11205) );
  NAND2_X1 U11079 ( .A1(n8482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8483) );
  AOI22_X1 U11080 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n6422), .B1(n12076), 
        .B2(n8594), .ZN(n8484) );
  NAND2_X1 U11081 ( .A1(n12656), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8491) );
  INV_X1 U11082 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n13636) );
  OR2_X1 U11083 ( .A1(n10097), .A2(n13636), .ZN(n8490) );
  INV_X1 U11084 ( .A(n8485), .ZN(n8511) );
  INV_X1 U11085 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n13679) );
  NAND2_X1 U11086 ( .A1(n8486), .A2(n13679), .ZN(n8487) );
  NAND2_X1 U11087 ( .A1(n8511), .A2(n8487), .ZN(n15093) );
  OR2_X1 U11088 ( .A1(n15093), .A2(n8267), .ZN(n8489) );
  INV_X1 U11089 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11682) );
  OR2_X1 U11090 ( .A1(n12660), .A2(n11682), .ZN(n8488) );
  INV_X1 U11091 ( .A(n10323), .ZN(n14734) );
  NAND2_X1 U11092 ( .A1(n14734), .A2(n8732), .ZN(n8492) );
  INV_X1 U11093 ( .A(n8495), .ZN(n8497) );
  NOR2_X1 U11094 ( .A1(n10323), .A2(n8643), .ZN(n8493) );
  AOI21_X1 U11095 ( .B1(n15212), .B2(n8732), .A(n8493), .ZN(n8494) );
  INV_X1 U11096 ( .A(n8494), .ZN(n8496) );
  AND2_X1 U11097 ( .A1(n8495), .A2(n8494), .ZN(n8498) );
  AOI21_X1 U11098 ( .B1(n8497), .B2(n8496), .A(n8498), .ZN(n14582) );
  INV_X1 U11099 ( .A(n8498), .ZN(n8499) );
  INV_X1 U11100 ( .A(n8503), .ZN(n8504) );
  OR3_X1 U11101 ( .A1(n8505), .A2(P1_IR_REG_13__SCAN_IN), .A3(
        P1_IR_REG_14__SCAN_IN), .ZN(n8506) );
  OAI21_X1 U11102 ( .B1(n8507), .B2(n8506), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8508) );
  XNOR2_X1 U11103 ( .A(n8508), .B(P1_IR_REG_15__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U11104 ( .A1(n6422), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8594), 
        .B2(n15476), .ZN(n8509) );
  NAND2_X1 U11105 ( .A1(n14715), .A2(n8775), .ZN(n8518) );
  INV_X1 U11106 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U11107 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NAND2_X1 U11108 ( .A1(n8533), .A2(n8512), .ZN(n15078) );
  OR2_X1 U11109 ( .A1(n15078), .A2(n8267), .ZN(n8516) );
  INV_X1 U11110 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15473) );
  OR2_X1 U11111 ( .A1(n12660), .A2(n15473), .ZN(n8515) );
  INV_X1 U11112 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15279) );
  OR2_X1 U11113 ( .A1(n10097), .A2(n15279), .ZN(n8514) );
  INV_X1 U11114 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15471) );
  OR2_X1 U11115 ( .A1(n8296), .A2(n15471), .ZN(n8513) );
  INV_X1 U11116 ( .A(n14586), .ZN(n14732) );
  NAND2_X1 U11117 ( .A1(n14732), .A2(n8239), .ZN(n8517) );
  NAND2_X1 U11118 ( .A1(n8518), .A2(n8517), .ZN(n8519) );
  XNOR2_X1 U11119 ( .A(n8519), .B(n10397), .ZN(n14628) );
  NOR2_X1 U11120 ( .A1(n14586), .A2(n8643), .ZN(n8520) );
  AOI21_X1 U11121 ( .B1(n14715), .B2(n8732), .A(n8520), .ZN(n14704) );
  NAND2_X1 U11122 ( .A1(n8524), .A2(n8523), .ZN(n8527) );
  INV_X1 U11123 ( .A(n8525), .ZN(n8526) );
  XNOR2_X1 U11124 ( .A(n8527), .B(n8526), .ZN(n11120) );
  NAND2_X1 U11125 ( .A1(n11120), .A2(n10091), .ZN(n8531) );
  NAND2_X1 U11126 ( .A1(n8528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U11127 ( .A(n8529), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U11128 ( .A1(n6422), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8594), 
        .B2(n12078), .ZN(n8530) );
  NAND2_X1 U11129 ( .A1(n8533), .A2(n8532), .ZN(n8534) );
  AND2_X1 U11130 ( .A1(n8555), .A2(n8534), .ZN(n15061) );
  NAND2_X1 U11131 ( .A1(n15061), .A2(n8803), .ZN(n8539) );
  NAND2_X1 U11132 ( .A1(n8226), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U11133 ( .A1(n12657), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8535) );
  AND2_X1 U11134 ( .A1(n8536), .A2(n8535), .ZN(n8538) );
  NAND2_X1 U11135 ( .A1(n12656), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8537) );
  OAI22_X1 U11136 ( .A1(n15064), .A2(n8645), .B1(n14707), .B2(n8644), .ZN(
        n8540) );
  XNOR2_X1 U11137 ( .A(n8540), .B(n8755), .ZN(n8544) );
  OAI22_X1 U11138 ( .A1(n15064), .A2(n8644), .B1(n14707), .B2(n8643), .ZN(
        n8543) );
  NAND2_X1 U11139 ( .A1(n8544), .A2(n8543), .ZN(n14626) );
  INV_X1 U11140 ( .A(n8541), .ZN(n8542) );
  OR2_X1 U11141 ( .A1(n8544), .A2(n8543), .ZN(n14625) );
  AND2_X1 U11142 ( .A1(n8547), .A2(n8570), .ZN(n8548) );
  NAND2_X1 U11143 ( .A1(n11305), .A2(n10091), .ZN(n8552) );
  NAND2_X1 U11144 ( .A1(n8549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8550) );
  XNOR2_X1 U11145 ( .A(n8550), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U11146 ( .A1(n6422), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8594), 
        .B2(n14787), .ZN(n8551) );
  NAND2_X2 U11147 ( .A1(n8552), .A2(n8551), .ZN(n15045) );
  NAND2_X1 U11148 ( .A1(n15045), .A2(n8775), .ZN(n8560) );
  INV_X1 U11149 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U11150 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  NAND2_X1 U11151 ( .A1(n6671), .A2(n8556), .ZN(n15046) );
  OR2_X1 U11152 ( .A1(n15046), .A2(n8267), .ZN(n8558) );
  AOI22_X1 U11153 ( .A1(n8226), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n12657), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n8557) );
  OAI211_X1 U11154 ( .C1(n8296), .C2(n15047), .A(n8558), .B(n8557), .ZN(n14730) );
  NAND2_X1 U11155 ( .A1(n14730), .A2(n8732), .ZN(n8559) );
  NAND2_X1 U11156 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  XNOR2_X1 U11157 ( .A(n8561), .B(n8755), .ZN(n8564) );
  NAND2_X1 U11158 ( .A1(n15045), .A2(n8732), .ZN(n8563) );
  NAND2_X1 U11159 ( .A1(n14730), .A2(n8292), .ZN(n8562) );
  NAND2_X1 U11160 ( .A1(n8563), .A2(n8562), .ZN(n8565) );
  NAND2_X1 U11161 ( .A1(n8564), .A2(n8565), .ZN(n14638) );
  INV_X1 U11162 ( .A(n8564), .ZN(n8567) );
  INV_X1 U11163 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U11164 ( .A1(n8567), .A2(n8566), .ZN(n14640) );
  NAND2_X1 U11165 ( .A1(n14636), .A2(n14640), .ZN(n14672) );
  NAND2_X1 U11166 ( .A1(n8569), .A2(n8568), .ZN(n8571) );
  XNOR2_X1 U11167 ( .A(n8572), .B(SI_18_), .ZN(n8573) );
  NAND2_X1 U11168 ( .A1(n11309), .A2(n10091), .ZN(n8578) );
  NAND2_X1 U11169 ( .A1(n8575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8576) );
  XNOR2_X1 U11170 ( .A(n8576), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U11171 ( .A1(n6422), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8594), 
        .B2(n14809), .ZN(n8577) );
  INV_X1 U11172 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U11173 ( .A1(n6671), .A2(n8579), .ZN(n8580) );
  NAND2_X1 U11174 ( .A1(n8598), .A2(n8580), .ZN(n15029) );
  OR2_X1 U11175 ( .A1(n15029), .A2(n8267), .ZN(n8585) );
  INV_X1 U11176 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U11177 ( .A1(n12656), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U11178 ( .A1(n12657), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8581) );
  OAI211_X1 U11179 ( .C1(n12660), .C2(n14799), .A(n8582), .B(n8581), .ZN(n8583) );
  INV_X1 U11180 ( .A(n8583), .ZN(n8584) );
  NAND2_X1 U11181 ( .A1(n8585), .A2(n8584), .ZN(n14729) );
  INV_X1 U11182 ( .A(n14729), .ZN(n14599) );
  OAI22_X1 U11183 ( .A1(n15032), .A2(n8644), .B1(n14599), .B2(n8643), .ZN(
        n8589) );
  NAND2_X1 U11184 ( .A1(n15188), .A2(n8775), .ZN(n8587) );
  NAND2_X1 U11185 ( .A1(n14729), .A2(n6415), .ZN(n8586) );
  NAND2_X1 U11186 ( .A1(n8587), .A2(n8586), .ZN(n8588) );
  XNOR2_X1 U11187 ( .A(n8588), .B(n8755), .ZN(n8590) );
  XOR2_X1 U11188 ( .A(n8589), .B(n8590), .Z(n14673) );
  XNOR2_X1 U11189 ( .A(n8593), .B(n8592), .ZN(n11407) );
  NAND2_X1 U11190 ( .A1(n11407), .A2(n10091), .ZN(n8596) );
  AOI22_X1 U11191 ( .A1(n6422), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12652), 
        .B2(n8594), .ZN(n8595) );
  NAND2_X1 U11192 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U11193 ( .A1(n8600), .A2(n8599), .ZN(n15010) );
  OR2_X1 U11194 ( .A1(n15010), .A2(n8267), .ZN(n8605) );
  INV_X1 U11195 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U11196 ( .A1(n12656), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11197 ( .A1(n12657), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U11198 ( .C1(n12660), .C2(n14808), .A(n8602), .B(n8601), .ZN(n8603) );
  INV_X1 U11199 ( .A(n8603), .ZN(n8604) );
  NOR2_X1 U11200 ( .A1(n14677), .A2(n8643), .ZN(n8606) );
  AOI21_X1 U11201 ( .B1(n15012), .B2(n8732), .A(n8606), .ZN(n8610) );
  NAND2_X1 U11202 ( .A1(n15012), .A2(n8775), .ZN(n8608) );
  NAND2_X1 U11203 ( .A1(n14728), .A2(n8239), .ZN(n8607) );
  NAND2_X1 U11204 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  XNOR2_X1 U11205 ( .A(n8609), .B(n8755), .ZN(n8612) );
  XOR2_X1 U11206 ( .A(n8610), .B(n8612), .Z(n14603) );
  INV_X1 U11207 ( .A(n8610), .ZN(n8611) );
  XNOR2_X1 U11208 ( .A(n8614), .B(n8615), .ZN(n14656) );
  NAND2_X1 U11209 ( .A1(n8618), .A2(SI_20_), .ZN(n8619) );
  MUX2_X1 U11210 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10071), .Z(n8633) );
  XNOR2_X1 U11211 ( .A(n8632), .B(n8631), .ZN(n11705) );
  NAND2_X1 U11212 ( .A1(n11705), .A2(n10091), .ZN(n8621) );
  NAND2_X1 U11213 ( .A1(n6422), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8620) );
  XNOR2_X1 U11214 ( .A(n8636), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n14978) );
  NAND2_X1 U11215 ( .A1(n14978), .A2(n8803), .ZN(n8626) );
  INV_X1 U11216 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U11217 ( .A1(n12656), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11218 ( .A1(n12657), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8622) );
  OAI211_X1 U11219 ( .C1(n12660), .C2(n15171), .A(n8623), .B(n8622), .ZN(n8624) );
  INV_X1 U11220 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U11221 ( .A1(n8626), .A2(n8625), .ZN(n14726) );
  AOI22_X1 U11222 ( .A1(n14974), .A2(n8732), .B1(n8292), .B2(n14726), .ZN(
        n8628) );
  AOI22_X1 U11223 ( .A1(n14974), .A2(n8775), .B1(n8732), .B2(n14726), .ZN(
        n8627) );
  XNOR2_X1 U11224 ( .A(n8627), .B(n8755), .ZN(n8629) );
  XOR2_X1 U11225 ( .A(n8628), .B(n8629), .Z(n14609) );
  NAND2_X1 U11226 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  NAND2_X1 U11227 ( .A1(n8633), .A2(SI_21_), .ZN(n8634) );
  OR2_X1 U11228 ( .A1(n9218), .A2(n10071), .ZN(n8635) );
  XNOR2_X1 U11229 ( .A(n8635), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15309) );
  INV_X1 U11230 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14613) );
  INV_X1 U11231 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14667) );
  OAI21_X1 U11232 ( .B1(n8636), .B2(n14613), .A(n14667), .ZN(n8637) );
  NAND2_X1 U11233 ( .A1(n8656), .A2(n8637), .ZN(n14958) );
  OR2_X1 U11234 ( .A1(n14958), .A2(n8267), .ZN(n8642) );
  INV_X1 U11235 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U11236 ( .A1(n8226), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11237 ( .A1(n12656), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8638) );
  OAI211_X1 U11238 ( .C1(n10097), .C2(n15261), .A(n8639), .B(n8638), .ZN(n8640) );
  INV_X1 U11239 ( .A(n8640), .ZN(n8641) );
  OAI22_X1 U11240 ( .A1(n15263), .A2(n8644), .B1(n14612), .B2(n8643), .ZN(
        n8647) );
  OAI22_X1 U11241 ( .A1(n15263), .A2(n8645), .B1(n14612), .B2(n8644), .ZN(
        n8646) );
  XNOR2_X1 U11242 ( .A(n8646), .B(n8755), .ZN(n8648) );
  XOR2_X1 U11243 ( .A(n8647), .B(n8648), .Z(n14663) );
  NAND2_X1 U11244 ( .A1(n14662), .A2(n14663), .ZN(n14661) );
  OR2_X1 U11245 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U11246 ( .A1(n14661), .A2(n8649), .ZN(n14591) );
  MUX2_X1 U11247 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10071), .Z(n9217) );
  INV_X1 U11248 ( .A(n9217), .ZN(n8652) );
  NAND2_X1 U11249 ( .A1(n8650), .A2(SI_22_), .ZN(n8651) );
  MUX2_X1 U11250 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10768), .Z(n8673) );
  XNOR2_X1 U11251 ( .A(n8673), .B(SI_23_), .ZN(n8653) );
  NAND2_X1 U11252 ( .A1(n12098), .A2(n10091), .ZN(n8655) );
  NAND2_X1 U11253 ( .A1(n6422), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U11254 ( .A1(n14940), .A2(n8775), .ZN(n8665) );
  INV_X1 U11255 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U11256 ( .A1(n8656), .A2(n13611), .ZN(n8657) );
  NAND2_X1 U11257 ( .A1(n8677), .A2(n8657), .ZN(n14594) );
  INV_X1 U11258 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11259 ( .A1(n12657), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11260 ( .A1(n12656), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8658) );
  OAI211_X1 U11261 ( .C1(n8660), .C2(n12660), .A(n8659), .B(n8658), .ZN(n8661)
         );
  INV_X1 U11262 ( .A(n8661), .ZN(n8662) );
  NAND2_X1 U11263 ( .A1(n14725), .A2(n8732), .ZN(n8664) );
  NAND2_X1 U11264 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  XNOR2_X1 U11265 ( .A(n8666), .B(n8755), .ZN(n8667) );
  AOI22_X1 U11266 ( .A1(n14940), .A2(n8732), .B1(n8292), .B2(n14725), .ZN(
        n8668) );
  XNOR2_X1 U11267 ( .A(n8667), .B(n8668), .ZN(n14592) );
  INV_X1 U11268 ( .A(n8667), .ZN(n8669) );
  NAND2_X1 U11269 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  INV_X1 U11270 ( .A(n8673), .ZN(n8671) );
  INV_X1 U11271 ( .A(SI_23_), .ZN(n11785) );
  NAND2_X1 U11272 ( .A1(n8671), .A2(n11785), .ZN(n8672) );
  MUX2_X1 U11273 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10071), .Z(n8695) );
  XNOR2_X1 U11274 ( .A(n8695), .B(SI_24_), .ZN(n8692) );
  NAND2_X1 U11275 ( .A1(n12228), .A2(n10091), .ZN(n8675) );
  NAND2_X1 U11276 ( .A1(n6422), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11277 ( .A1(n14921), .A2(n8775), .ZN(n8686) );
  INV_X1 U11278 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11279 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  AND2_X1 U11280 ( .A1(n8701), .A2(n8678), .ZN(n14922) );
  NAND2_X1 U11281 ( .A1(n14922), .A2(n8803), .ZN(n8684) );
  INV_X1 U11282 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11283 ( .A1(n12657), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11284 ( .A1(n12656), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U11285 ( .C1(n12660), .C2(n8681), .A(n8680), .B(n8679), .ZN(n8682)
         );
  INV_X1 U11286 ( .A(n8682), .ZN(n8683) );
  NAND2_X1 U11287 ( .A1(n14724), .A2(n8732), .ZN(n8685) );
  NAND2_X1 U11288 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  XNOR2_X1 U11289 ( .A(n8687), .B(n8755), .ZN(n8688) );
  AOI22_X1 U11290 ( .A1(n14921), .A2(n8732), .B1(n8292), .B2(n14724), .ZN(
        n8689) );
  XNOR2_X1 U11291 ( .A(n8688), .B(n8689), .ZN(n14647) );
  INV_X1 U11292 ( .A(n8688), .ZN(n8690) );
  NAND2_X1 U11293 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  MUX2_X1 U11294 ( .A(n12283), .B(n12285), .S(n10071), .Z(n8696) );
  INV_X1 U11295 ( .A(SI_25_), .ZN(n12235) );
  NAND2_X1 U11296 ( .A1(n8696), .A2(n12235), .ZN(n8715) );
  INV_X1 U11297 ( .A(n8696), .ZN(n8697) );
  NAND2_X1 U11298 ( .A1(n8697), .A2(SI_25_), .ZN(n8698) );
  NAND2_X1 U11299 ( .A1(n8715), .A2(n8698), .ZN(n8716) );
  XNOR2_X1 U11300 ( .A(n8717), .B(n8716), .ZN(n12282) );
  NAND2_X1 U11301 ( .A1(n6422), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U11302 ( .A1(n14903), .A2(n8775), .ZN(n8709) );
  INV_X1 U11303 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U11304 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  NAND2_X1 U11305 ( .A1(n8722), .A2(n8702), .ZN(n14620) );
  OR2_X1 U11306 ( .A1(n14620), .A2(n8267), .ZN(n8707) );
  INV_X1 U11307 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U11308 ( .A1(n12656), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11309 ( .A1(n12657), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8703) );
  OAI211_X1 U11310 ( .C1(n12660), .C2(n15150), .A(n8704), .B(n8703), .ZN(n8705) );
  INV_X1 U11311 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U11312 ( .A1(n14723), .A2(n8732), .ZN(n8708) );
  NAND2_X1 U11313 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  XNOR2_X1 U11314 ( .A(n8710), .B(n8755), .ZN(n8711) );
  AOI22_X1 U11315 ( .A1(n14903), .A2(n8732), .B1(n8292), .B2(n14723), .ZN(
        n8712) );
  XNOR2_X1 U11316 ( .A(n8711), .B(n8712), .ZN(n14619) );
  INV_X1 U11317 ( .A(n8711), .ZN(n8713) );
  NAND2_X1 U11318 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  INV_X1 U11319 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15306) );
  INV_X1 U11320 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14570) );
  MUX2_X1 U11321 ( .A(n15306), .B(n14570), .S(n10768), .Z(n8736) );
  XNOR2_X1 U11322 ( .A(n8736), .B(SI_26_), .ZN(n8718) );
  NAND2_X1 U11323 ( .A1(n14568), .A2(n10091), .ZN(n8720) );
  NAND2_X1 U11324 ( .A1(n6422), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11325 ( .A1(n14890), .A2(n8775), .ZN(n8730) );
  INV_X1 U11326 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11327 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  NAND2_X1 U11328 ( .A1(n14885), .A2(n8803), .ZN(n8728) );
  INV_X1 U11329 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15145) );
  NAND2_X1 U11330 ( .A1(n12656), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11331 ( .A1(n12657), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8724) );
  OAI211_X1 U11332 ( .C1(n12660), .C2(n15145), .A(n8725), .B(n8724), .ZN(n8726) );
  INV_X1 U11333 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U11334 ( .A1(n14722), .A2(n8732), .ZN(n8729) );
  NAND2_X1 U11335 ( .A1(n8730), .A2(n8729), .ZN(n8731) );
  XNOR2_X1 U11336 ( .A(n8731), .B(n8755), .ZN(n8735) );
  AOI22_X1 U11337 ( .A1(n14890), .A2(n8732), .B1(n8292), .B2(n14722), .ZN(
        n8733) );
  XNOR2_X1 U11338 ( .A(n8735), .B(n8733), .ZN(n14696) );
  INV_X1 U11339 ( .A(n8733), .ZN(n8734) );
  INV_X1 U11340 ( .A(SI_26_), .ZN(n13837) );
  NAND2_X1 U11341 ( .A1(n8737), .A2(n13837), .ZN(n8738) );
  MUX2_X1 U11342 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10071), .Z(n8760) );
  INV_X1 U11343 ( .A(n8760), .ZN(n8740) );
  XNOR2_X1 U11344 ( .A(n8740), .B(SI_27_), .ZN(n8741) );
  NAND2_X1 U11345 ( .A1(n12941), .A2(n10091), .ZN(n8743) );
  NAND2_X1 U11346 ( .A1(n6422), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11347 ( .A1(n14880), .A2(n8775), .ZN(n8754) );
  INV_X1 U11348 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11349 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U11350 ( .A1(n14844), .A2(n8747), .ZN(n14875) );
  OR2_X1 U11351 ( .A1(n14875), .A2(n8267), .ZN(n8752) );
  INV_X1 U11352 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U11353 ( .A1(n8226), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11354 ( .A1(n12657), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8748) );
  OAI211_X1 U11355 ( .C1(n14874), .C2(n8296), .A(n8749), .B(n8748), .ZN(n8750)
         );
  INV_X1 U11356 ( .A(n8750), .ZN(n8751) );
  NAND2_X1 U11357 ( .A1(n14721), .A2(n8732), .ZN(n8753) );
  NAND2_X1 U11358 ( .A1(n8754), .A2(n8753), .ZN(n8756) );
  XNOR2_X1 U11359 ( .A(n8756), .B(n8755), .ZN(n8824) );
  AND2_X1 U11360 ( .A1(n14721), .A2(n8292), .ZN(n8757) );
  AOI21_X1 U11361 ( .B1(n14880), .B2(n8732), .A(n8757), .ZN(n8822) );
  XNOR2_X1 U11362 ( .A(n8824), .B(n8822), .ZN(n14574) );
  NOR2_X1 U11363 ( .A1(n8760), .A2(SI_27_), .ZN(n8758) );
  NAND2_X1 U11364 ( .A1(n8760), .A2(SI_27_), .ZN(n8761) );
  INV_X1 U11365 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12947) );
  INV_X1 U11366 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U11367 ( .A(n12947), .B(n10202), .S(n10071), .Z(n8762) );
  INV_X1 U11368 ( .A(SI_28_), .ZN(n12917) );
  NAND2_X1 U11369 ( .A1(n8762), .A2(n12917), .ZN(n9981) );
  INV_X1 U11370 ( .A(n8762), .ZN(n8763) );
  NAND2_X1 U11371 ( .A1(n8763), .A2(SI_28_), .ZN(n8764) );
  NAND2_X1 U11372 ( .A1(n9981), .A2(n8764), .ZN(n9982) );
  NAND2_X1 U11373 ( .A1(n12945), .A2(n10091), .ZN(n8766) );
  NAND2_X1 U11374 ( .A1(n6422), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8765) );
  NAND2_X2 U11375 ( .A1(n8766), .A2(n8765), .ZN(n12804) );
  NAND2_X1 U11376 ( .A1(n12804), .A2(n8732), .ZN(n8773) );
  NAND2_X1 U11377 ( .A1(n14858), .A2(n8803), .ZN(n8771) );
  INV_X1 U11378 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n13655) );
  NAND2_X1 U11379 ( .A1(n8226), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11380 ( .A1(n12656), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8767) );
  OAI211_X1 U11381 ( .C1(n10097), .C2(n13655), .A(n8768), .B(n8767), .ZN(n8769) );
  INV_X1 U11382 ( .A(n8769), .ZN(n8770) );
  NAND2_X1 U11383 ( .A1(n14839), .A2(n8292), .ZN(n8772) );
  NAND2_X1 U11384 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  XNOR2_X1 U11385 ( .A(n8774), .B(n10397), .ZN(n8777) );
  AOI22_X1 U11386 ( .A1(n12804), .A2(n8775), .B1(n8732), .B2(n14839), .ZN(
        n8776) );
  XNOR2_X1 U11387 ( .A(n8777), .B(n8776), .ZN(n8829) );
  INV_X1 U11388 ( .A(n8829), .ZN(n8800) );
  INV_X1 U11389 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10759) );
  NOR4_X1 U11390 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8786) );
  NOR4_X1 U11391 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8785) );
  INV_X1 U11392 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15535) );
  INV_X1 U11393 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15539) );
  INV_X1 U11394 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15537) );
  INV_X1 U11395 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15536) );
  NAND4_X1 U11396 ( .A1(n15535), .A2(n15539), .A3(n15537), .A4(n15536), .ZN(
        n8783) );
  NOR4_X1 U11397 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n8781) );
  NOR4_X1 U11398 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n8780) );
  NOR4_X1 U11399 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n8779) );
  NOR4_X1 U11400 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n8778) );
  NAND4_X1 U11401 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(n8782)
         );
  NOR4_X1 U11402 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        n8783), .A4(n8782), .ZN(n8784) );
  NAND3_X1 U11403 ( .A1(n8786), .A2(n8785), .A3(n8784), .ZN(n10104) );
  AND2_X1 U11404 ( .A1(n12229), .A2(P1_B_REG_SCAN_IN), .ZN(n8788) );
  NOR2_X1 U11405 ( .A1(n12229), .A2(P1_B_REG_SCAN_IN), .ZN(n8787) );
  AOI21_X1 U11406 ( .B1(n12284), .B2(n8788), .A(n8787), .ZN(n8789) );
  AND2_X1 U11407 ( .A1(n8790), .A2(n8789), .ZN(n10754) );
  OAI21_X1 U11408 ( .B1(n10759), .B2(n10104), .A(n10754), .ZN(n8791) );
  NAND2_X1 U11409 ( .A1(n15308), .A2(n12284), .ZN(n10757) );
  INV_X1 U11410 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U11411 ( .A1(n10754), .A2(n10763), .ZN(n8792) );
  NAND2_X1 U11412 ( .A1(n15308), .A2(n12229), .ZN(n10760) );
  NAND2_X1 U11413 ( .A1(n8813), .A2(n10114), .ZN(n8816) );
  INV_X1 U11414 ( .A(n8816), .ZN(n8796) );
  NAND2_X1 U11415 ( .A1(n8796), .A2(n10756), .ZN(n8802) );
  INV_X1 U11416 ( .A(n8802), .ZN(n8799) );
  INV_X1 U11417 ( .A(n15524), .ZN(n8797) );
  NAND2_X1 U11418 ( .A1(n11828), .A2(n15526), .ZN(n8812) );
  NAND2_X1 U11419 ( .A1(n12651), .A2(n8801), .ZN(n12815) );
  AND2_X1 U11420 ( .A1(n15579), .A2(n12815), .ZN(n8798) );
  NAND2_X1 U11421 ( .A1(n8800), .A2(n14685), .ZN(n8833) );
  NOR2_X1 U11422 ( .A1(n15588), .A2(n8801), .ZN(n10106) );
  NAND2_X1 U11423 ( .A1(n8802), .A2(n15511), .ZN(n14689) );
  NAND2_X1 U11424 ( .A1(n8803), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8804) );
  OR2_X1 U11425 ( .A1(n14844), .A2(n8804), .ZN(n8810) );
  INV_X1 U11426 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11427 ( .A1(n12657), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U11428 ( .A1(n12656), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8805) );
  OAI211_X1 U11429 ( .C1(n12660), .C2(n8807), .A(n8806), .B(n8805), .ZN(n8808)
         );
  INV_X1 U11430 ( .A(n8808), .ZN(n8809) );
  INV_X1 U11431 ( .A(n8811), .ZN(n10881) );
  OR2_X1 U11432 ( .A1(n12815), .A2(n8811), .ZN(n14675) );
  AOI22_X1 U11433 ( .A1(n14720), .A2(n14697), .B1(n14721), .B2(n15111), .ZN(
        n10348) );
  INV_X1 U11434 ( .A(n12815), .ZN(n10720) );
  NAND2_X1 U11435 ( .A1(n10720), .A2(n8812), .ZN(n11126) );
  NAND3_X1 U11436 ( .A1(n10597), .A2(n11126), .A3(n10719), .ZN(n8817) );
  INV_X1 U11437 ( .A(n8813), .ZN(n8814) );
  NAND2_X1 U11438 ( .A1(n11826), .A2(n10114), .ZN(n14700) );
  INV_X1 U11439 ( .A(n10106), .ZN(n8815) );
  NAND2_X1 U11440 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  INV_X1 U11441 ( .A(n8817), .ZN(n8818) );
  NAND2_X1 U11442 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  AOI22_X1 U11443 ( .A1(n14858), .A2(n14698), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n8821) );
  OAI21_X1 U11444 ( .B1(n10348), .B2(n14700), .A(n8821), .ZN(n8826) );
  INV_X1 U11445 ( .A(n8822), .ZN(n8823) );
  OR2_X1 U11446 ( .A1(n8824), .A2(n8823), .ZN(n8827) );
  NOR3_X1 U11447 ( .A1(n8829), .A2(n14717), .A3(n8827), .ZN(n8825) );
  AOI211_X1 U11448 ( .C1(n14714), .C2(n12804), .A(n8826), .B(n8825), .ZN(n8832) );
  AND2_X1 U11449 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  NAND2_X1 U11450 ( .A1(n8834), .A2(n8830), .ZN(n8831) );
  OAI211_X1 U11451 ( .C1(n8834), .C2(n8833), .A(n8832), .B(n8831), .ZN(
        P1_U3220) );
  NOR2_X2 U11452 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8835) );
  NAND2_X1 U11453 ( .A1(n8844), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11454 ( .A1(n8863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8845) );
  MUX2_X1 U11455 ( .A(n8845), .B(P2_IR_REG_31__SCAN_IN), .S(n13610), .Z(n8846)
         );
  NAND2_X1 U11456 ( .A1(n6477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8847) );
  INV_X1 U11457 ( .A(n9334), .ZN(n9343) );
  INV_X1 U11458 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11459 ( .A1(n9143), .A2(n8851), .ZN(n9154) );
  AND2_X1 U11460 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8852) );
  INV_X1 U11461 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8854) );
  INV_X1 U11462 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8853) );
  NAND3_X1 U11463 ( .A1(n8854), .A2(n8853), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n8856) );
  XNOR2_X1 U11464 ( .A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n8855) );
  NAND2_X2 U11465 ( .A1(n8860), .A2(n12630), .ZN(n14337) );
  INV_X1 U11466 ( .A(n12582), .ZN(n8861) );
  INV_X1 U11467 ( .A(n8871), .ZN(n8862) );
  NOR3_X1 U11468 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .A3(P2_IR_REG_27__SCAN_IN), .ZN(n8870) );
  INV_X1 U11469 ( .A(n8873), .ZN(n8876) );
  NOR2_X1 U11470 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n8874) );
  AOI21_X1 U11471 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n8877) );
  AND2_X1 U11472 ( .A1(n8880), .A2(n8877), .ZN(n8878) );
  NAND2_X1 U11473 ( .A1(n8880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8882) );
  MUX2_X1 U11474 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8882), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8883) );
  INV_X1 U11475 ( .A(n8884), .ZN(n8910) );
  INV_X1 U11476 ( .A(n15619), .ZN(n11082) );
  NAND2_X1 U11477 ( .A1(n11049), .A2(n11082), .ZN(n8885) );
  XNOR2_X1 U11478 ( .A(n8899), .B(n11574), .ZN(n8898) );
  NAND2_X1 U11479 ( .A1(n9001), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8893) );
  INV_X1 U11480 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8892) );
  AND2_X1 U11481 ( .A1(n8895), .A2(n12626), .ZN(n8896) );
  AND2_X2 U11482 ( .A1(n12625), .A2(n8896), .ZN(n14273) );
  NAND2_X1 U11483 ( .A1(n14024), .A2(n9166), .ZN(n8897) );
  NAND2_X1 U11484 ( .A1(n10071), .A2(SI_0_), .ZN(n8900) );
  NAND2_X1 U11485 ( .A1(n8900), .A2(n9421), .ZN(n8902) );
  NAND2_X1 U11486 ( .A1(n8902), .A2(n8901), .ZN(n14572) );
  MUX2_X1 U11487 ( .A(n8903), .B(n14572), .S(n8940), .Z(n15727) );
  NAND2_X1 U11488 ( .A1(n9014), .A2(n15727), .ZN(n8909) );
  NAND2_X1 U11489 ( .A1(n9374), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U11490 ( .A1(n6474), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8907) );
  INV_X1 U11491 ( .A(n12539), .ZN(n8904) );
  NAND2_X1 U11492 ( .A1(n8904), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U11493 ( .A1(n9001), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11494 ( .A1(n14025), .A2(n11663), .ZN(n11662) );
  NAND2_X1 U11495 ( .A1(n10003), .A2(n9166), .ZN(n11390) );
  NAND2_X1 U11496 ( .A1(n8909), .A2(n11390), .ZN(n11422) );
  NAND2_X1 U11497 ( .A1(n12550), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11498 ( .A1(n8910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8911) );
  INV_X1 U11499 ( .A(n8912), .ZN(n8927) );
  NAND2_X1 U11500 ( .A1(n8913), .A2(n8927), .ZN(n15639) );
  INV_X1 U11501 ( .A(n15639), .ZN(n11084) );
  NAND2_X1 U11502 ( .A1(n11049), .A2(n11084), .ZN(n8914) );
  INV_X1 U11503 ( .A(n14400), .ZN(n11039) );
  XNOR2_X1 U11504 ( .A(n8899), .B(n11039), .ZN(n8920) );
  NAND2_X1 U11505 ( .A1(n9374), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11506 ( .A1(n6474), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11507 ( .A1(n9001), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11508 ( .A1(n8904), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11509 ( .A1(n14023), .A2(n9166), .ZN(n8921) );
  NAND2_X1 U11510 ( .A1(n8920), .A2(n8921), .ZN(n8925) );
  INV_X1 U11511 ( .A(n8920), .ZN(n8923) );
  INV_X1 U11512 ( .A(n8921), .ZN(n8922) );
  NAND2_X1 U11513 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  AND2_X1 U11514 ( .A1(n8925), .A2(n8924), .ZN(n13961) );
  NAND2_X1 U11515 ( .A1(n8927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U11516 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8928), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8930) );
  INV_X1 U11517 ( .A(n8943), .ZN(n8941) );
  XNOR2_X1 U11518 ( .A(n8899), .B(n10045), .ZN(n8935) );
  INV_X1 U11519 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U11520 ( .A1(n9374), .A2(n11652), .ZN(n8934) );
  NAND2_X1 U11521 ( .A1(n6474), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U11522 ( .A1(n8904), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11523 ( .A1(n9001), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U11524 ( .A1(n14022), .A2(n9166), .ZN(n8936) );
  XNOR2_X1 U11525 ( .A(n8935), .B(n8936), .ZN(n13863) );
  INV_X1 U11526 ( .A(n13863), .ZN(n8939) );
  INV_X1 U11527 ( .A(n8935), .ZN(n8938) );
  INV_X1 U11528 ( .A(n8936), .ZN(n8937) );
  NAND2_X1 U11529 ( .A1(n10742), .A2(n9009), .ZN(n8947) );
  NAND2_X1 U11530 ( .A1(n8941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U11531 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8942), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8944) );
  NAND2_X1 U11532 ( .A1(n8943), .A2(n13592), .ZN(n8960) );
  NAND2_X1 U11533 ( .A1(n8944), .A2(n8960), .ZN(n11088) );
  OAI22_X1 U11534 ( .A1(n9191), .A2(n10743), .B1(n8940), .B2(n11088), .ZN(
        n8945) );
  INV_X1 U11535 ( .A(n8945), .ZN(n8946) );
  XNOR2_X1 U11536 ( .A(n8899), .B(n7888), .ZN(n8953) );
  INV_X1 U11537 ( .A(n8965), .ZN(n8967) );
  OAI21_X1 U11538 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8967), .ZN(n11595) );
  INV_X1 U11539 ( .A(n11595), .ZN(n8948) );
  NAND2_X1 U11540 ( .A1(n9374), .A2(n8948), .ZN(n8952) );
  NAND2_X1 U11541 ( .A1(n6474), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11542 ( .A1(n9001), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11543 ( .A1(n14021), .A2(n9166), .ZN(n8954) );
  NAND2_X1 U11544 ( .A1(n8953), .A2(n8954), .ZN(n8958) );
  INV_X1 U11545 ( .A(n8953), .ZN(n8956) );
  INV_X1 U11546 ( .A(n8954), .ZN(n8955) );
  NAND2_X1 U11547 ( .A1(n8956), .A2(n8955), .ZN(n8957) );
  AND2_X1 U11548 ( .A1(n8958), .A2(n8957), .ZN(n11326) );
  NAND2_X1 U11549 ( .A1(n10752), .A2(n9009), .ZN(n8964) );
  NAND2_X1 U11550 ( .A1(n8960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8959) );
  MUX2_X1 U11551 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8959), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8961) );
  NAND2_X1 U11552 ( .A1(n8961), .A2(n8989), .ZN(n14045) );
  OAI22_X1 U11553 ( .A1(n9191), .A2(n10753), .B1(n8940), .B2(n14045), .ZN(
        n8962) );
  INV_X1 U11554 ( .A(n8962), .ZN(n8963) );
  INV_X1 U11555 ( .A(n12404), .ZN(n15759) );
  XNOR2_X1 U11556 ( .A(n8899), .B(n15759), .ZN(n8973) );
  INV_X1 U11557 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11558 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  AND2_X1 U11559 ( .A1(n8999), .A2(n8968), .ZN(n11382) );
  NAND2_X1 U11560 ( .A1(n9374), .A2(n11382), .ZN(n8972) );
  NAND2_X1 U11561 ( .A1(n6474), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11562 ( .A1(n9001), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11563 ( .A1(n14020), .A2(n9166), .ZN(n8974) );
  NAND2_X1 U11564 ( .A1(n8973), .A2(n8974), .ZN(n8978) );
  INV_X1 U11565 ( .A(n8973), .ZN(n8976) );
  INV_X1 U11566 ( .A(n8974), .ZN(n8975) );
  NAND2_X1 U11567 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  AND2_X1 U11568 ( .A1(n8978), .A2(n8977), .ZN(n11385) );
  NAND2_X1 U11569 ( .A1(n10746), .A2(n9009), .ZN(n8982) );
  NAND2_X1 U11570 ( .A1(n8989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U11571 ( .A(n8979), .B(n8990), .ZN(n14058) );
  OAI22_X1 U11572 ( .A1(n9191), .A2(n10747), .B1(n8940), .B2(n14058), .ZN(
        n8980) );
  INV_X1 U11573 ( .A(n8980), .ZN(n8981) );
  XNOR2_X1 U11574 ( .A(n8899), .B(n12420), .ZN(n8988) );
  XNOR2_X1 U11575 ( .A(n8999), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U11576 ( .A1(n9374), .A2(n11550), .ZN(n8986) );
  NAND2_X1 U11577 ( .A1(n6474), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11578 ( .A1(n9991), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U11579 ( .A1(n9001), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8983) );
  AND2_X1 U11580 ( .A1(n14019), .A2(n9166), .ZN(n8987) );
  XNOR2_X1 U11581 ( .A(n8988), .B(n8987), .ZN(n11427) );
  NAND2_X1 U11582 ( .A1(n10744), .A2(n9302), .ZN(n8994) );
  INV_X4 U11583 ( .A(n9191), .ZN(n12550) );
  INV_X1 U11584 ( .A(n8989), .ZN(n8991) );
  NAND2_X1 U11585 ( .A1(n8991), .A2(n8990), .ZN(n9010) );
  NAND2_X1 U11586 ( .A1(n9010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8992) );
  XNOR2_X1 U11587 ( .A(n8992), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U11588 ( .A1(n12550), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11049), 
        .B2(n14074), .ZN(n8993) );
  XNOR2_X1 U11589 ( .A(n12428), .B(n8899), .ZN(n9008) );
  INV_X1 U11590 ( .A(n8999), .ZN(n8996) );
  INV_X1 U11591 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8998) );
  INV_X1 U11592 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8997) );
  OAI21_X1 U11593 ( .B1(n8999), .B2(n8998), .A(n8997), .ZN(n9000) );
  AND2_X1 U11594 ( .A1(n9016), .A2(n9000), .ZN(n11697) );
  NAND2_X1 U11595 ( .A1(n9374), .A2(n11697), .ZN(n9005) );
  NAND2_X1 U11596 ( .A1(n6474), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11597 ( .A1(n9991), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11598 ( .A1(n9375), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9002) );
  NAND4_X1 U11599 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n14018) );
  NAND2_X1 U11600 ( .A1(n14018), .A2(n9166), .ZN(n9006) );
  XNOR2_X1 U11601 ( .A(n9008), .B(n9006), .ZN(n11694) );
  INV_X1 U11602 ( .A(n9006), .ZN(n9007) );
  NAND2_X1 U11603 ( .A1(n10764), .A2(n9302), .ZN(n9013) );
  NAND2_X1 U11604 ( .A1(n9028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U11605 ( .A(n9011), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U11606 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n12550), .B1(n14084), 
        .B2(n11049), .ZN(n9012) );
  XNOR2_X1 U11607 ( .A(n14509), .B(n9305), .ZN(n9022) );
  NAND2_X1 U11608 ( .A1(n6474), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9021) );
  INV_X1 U11609 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11610 ( .A1(n9016), .A2(n9015), .ZN(n9017) );
  AND2_X1 U11611 ( .A1(n9038), .A2(n9017), .ZN(n11849) );
  NAND2_X1 U11612 ( .A1(n9374), .A2(n11849), .ZN(n9020) );
  NAND2_X1 U11613 ( .A1(n9375), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11614 ( .A1(n9991), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9018) );
  NAND4_X1 U11615 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(n9018), .ZN(n14017) );
  NAND2_X1 U11616 ( .A1(n14017), .A2(n9166), .ZN(n9023) );
  NAND2_X1 U11617 ( .A1(n9022), .A2(n9023), .ZN(n9027) );
  INV_X1 U11618 ( .A(n9022), .ZN(n9025) );
  INV_X1 U11619 ( .A(n9023), .ZN(n9024) );
  NAND2_X1 U11620 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  AND2_X1 U11621 ( .A1(n9027), .A2(n9026), .ZN(n11845) );
  NAND2_X1 U11622 ( .A1(n11844), .A2(n9027), .ZN(n11894) );
  NAND2_X1 U11623 ( .A1(n10796), .A2(n9302), .ZN(n9036) );
  NAND2_X1 U11624 ( .A1(n9030), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9029) );
  MUX2_X1 U11625 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9029), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9033) );
  INV_X1 U11626 ( .A(n9030), .ZN(n9032) );
  INV_X1 U11627 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U11628 ( .A1(n9032), .A2(n9031), .ZN(n9065) );
  NAND2_X1 U11629 ( .A1(n9033), .A2(n9065), .ZN(n15675) );
  INV_X1 U11630 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10797) );
  OAI22_X1 U11631 ( .A1(n15675), .A2(n8940), .B1(n10797), .B2(n9191), .ZN(
        n9034) );
  INV_X1 U11632 ( .A(n9034), .ZN(n9035) );
  XNOR2_X1 U11633 ( .A(n12455), .B(n9305), .ZN(n9044) );
  NAND2_X1 U11634 ( .A1(n6474), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11635 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  AND2_X1 U11636 ( .A1(n9054), .A2(n9039), .ZN(n11897) );
  NAND2_X1 U11637 ( .A1(n9374), .A2(n11897), .ZN(n9042) );
  INV_X2 U11638 ( .A(n9162), .ZN(n9375) );
  NAND2_X1 U11639 ( .A1(n9375), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11640 ( .A1(n9991), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9040) );
  NAND4_X1 U11641 ( .A1(n9043), .A2(n9042), .A3(n9041), .A4(n9040), .ZN(n14015) );
  NAND2_X1 U11642 ( .A1(n14015), .A2(n9166), .ZN(n9045) );
  NAND2_X1 U11643 ( .A1(n9044), .A2(n9045), .ZN(n9049) );
  INV_X1 U11644 ( .A(n9044), .ZN(n9047) );
  INV_X1 U11645 ( .A(n9045), .ZN(n9046) );
  NAND2_X1 U11646 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  AND2_X1 U11647 ( .A1(n9049), .A2(n9048), .ZN(n11895) );
  NAND2_X1 U11648 ( .A1(n11894), .A2(n11895), .ZN(n11893) );
  NAND2_X1 U11649 ( .A1(n10833), .A2(n9302), .ZN(n9052) );
  NAND2_X1 U11650 ( .A1(n9065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U11651 ( .A(n9050), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U11652 ( .A1(n11267), .A2(n11049), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n12550), .ZN(n9051) );
  XNOR2_X1 U11653 ( .A(n12460), .B(n9305), .ZN(n9060) );
  INV_X1 U11654 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n13604) );
  NAND2_X1 U11655 ( .A1(n9054), .A2(n13604), .ZN(n9055) );
  AND2_X1 U11656 ( .A1(n9070), .A2(n9055), .ZN(n12032) );
  NAND2_X1 U11657 ( .A1(n9374), .A2(n12032), .ZN(n9059) );
  NAND2_X1 U11658 ( .A1(n6474), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11659 ( .A1(n9991), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11660 ( .A1(n9375), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9056) );
  NAND4_X1 U11661 ( .A1(n9059), .A2(n9058), .A3(n9057), .A4(n9056), .ZN(n14014) );
  NAND2_X1 U11662 ( .A1(n14014), .A2(n9166), .ZN(n9061) );
  XNOR2_X1 U11663 ( .A(n9060), .B(n9061), .ZN(n11993) );
  INV_X1 U11664 ( .A(n9060), .ZN(n9063) );
  INV_X1 U11665 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U11666 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  NAND2_X1 U11667 ( .A1(n10865), .A2(n9302), .ZN(n9068) );
  OAI21_X1 U11668 ( .B1(n9065), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9066) );
  XNOR2_X1 U11669 ( .A(n9066), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U11670 ( .A1(n11798), .A2(n11049), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n12550), .ZN(n9067) );
  XNOR2_X1 U11671 ( .A(n14504), .B(n9305), .ZN(n9076) );
  NAND2_X1 U11672 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  AND2_X1 U11673 ( .A1(n9090), .A2(n9071), .ZN(n12292) );
  NAND2_X1 U11674 ( .A1(n9374), .A2(n12292), .ZN(n9075) );
  NAND2_X1 U11675 ( .A1(n6474), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U11676 ( .A1(n9375), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11677 ( .A1(n9991), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9072) );
  NAND4_X1 U11678 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n14013) );
  NAND2_X1 U11679 ( .A1(n14013), .A2(n9166), .ZN(n9077) );
  NAND2_X1 U11680 ( .A1(n9076), .A2(n9077), .ZN(n9081) );
  INV_X1 U11681 ( .A(n9076), .ZN(n9079) );
  INV_X1 U11682 ( .A(n9077), .ZN(n9078) );
  NAND2_X1 U11683 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NAND2_X1 U11684 ( .A1(n9081), .A2(n9080), .ZN(n12290) );
  NAND2_X1 U11685 ( .A1(n10911), .A2(n9302), .ZN(n9087) );
  NAND2_X1 U11686 ( .A1(n9082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  XNOR2_X1 U11687 ( .A(n9084), .B(n9083), .ZN(n15695) );
  OAI22_X1 U11688 ( .A1(n9191), .A2(n10912), .B1(n8940), .B2(n15695), .ZN(
        n9085) );
  INV_X1 U11689 ( .A(n9085), .ZN(n9086) );
  XNOR2_X1 U11690 ( .A(n14500), .B(n9305), .ZN(n9095) );
  INV_X1 U11691 ( .A(n9090), .ZN(n9088) );
  INV_X1 U11692 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11693 ( .A1(n9090), .A2(n9089), .ZN(n9091) );
  NAND2_X1 U11694 ( .A1(n9104), .A2(n9091), .ZN(n12325) );
  INV_X1 U11695 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11800) );
  OAI22_X1 U11696 ( .A1(n9326), .A2(n12325), .B1(n9379), .B2(n11800), .ZN(
        n9094) );
  INV_X1 U11697 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9092) );
  INV_X1 U11698 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11788) );
  OAI22_X1 U11699 ( .A1(n12539), .A2(n9092), .B1(n9162), .B2(n11788), .ZN(
        n9093) );
  NAND2_X1 U11700 ( .A1(n14012), .A2(n9166), .ZN(n9096) );
  AND2_X1 U11701 ( .A1(n9095), .A2(n9096), .ZN(n12320) );
  INV_X1 U11702 ( .A(n9095), .ZN(n9098) );
  INV_X1 U11703 ( .A(n9096), .ZN(n9097) );
  NAND2_X1 U11704 ( .A1(n9098), .A2(n9097), .ZN(n12321) );
  NAND2_X1 U11705 ( .A1(n10979), .A2(n9302), .ZN(n9103) );
  NAND2_X1 U11706 ( .A1(n9099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9100) );
  XNOR2_X1 U11707 ( .A(n9100), .B(n7749), .ZN(n11803) );
  OAI22_X1 U11708 ( .A1(n9191), .A2(n13593), .B1(n8940), .B2(n11803), .ZN(
        n9101) );
  INV_X1 U11709 ( .A(n9101), .ZN(n9102) );
  XNOR2_X1 U11710 ( .A(n14495), .B(n8899), .ZN(n9110) );
  NAND2_X1 U11711 ( .A1(n9104), .A2(n14097), .ZN(n9105) );
  AND2_X1 U11712 ( .A1(n9121), .A2(n9105), .ZN(n12365) );
  NAND2_X1 U11713 ( .A1(n9374), .A2(n12365), .ZN(n9109) );
  NAND2_X1 U11714 ( .A1(n6474), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11715 ( .A1(n9991), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11716 ( .A1(n9375), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9106) );
  NAND4_X1 U11717 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n14011) );
  AND2_X1 U11718 ( .A1(n14011), .A2(n9166), .ZN(n9111) );
  NAND2_X1 U11719 ( .A1(n9110), .A2(n9111), .ZN(n9115) );
  INV_X1 U11720 ( .A(n9110), .ZN(n9113) );
  INV_X1 U11721 ( .A(n9111), .ZN(n9112) );
  NAND2_X1 U11722 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  AND2_X1 U11723 ( .A1(n9115), .A2(n9114), .ZN(n12361) );
  NAND2_X1 U11724 ( .A1(n11205), .A2(n9302), .ZN(n9120) );
  INV_X1 U11725 ( .A(n8850), .ZN(n9116) );
  NAND2_X1 U11726 ( .A1(n9116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9117) );
  XNOR2_X1 U11727 ( .A(n9117), .B(n9132), .ZN(n11806) );
  OAI22_X1 U11728 ( .A1(n9191), .A2(n11206), .B1(n8940), .B2(n11806), .ZN(
        n9118) );
  INV_X1 U11729 ( .A(n9118), .ZN(n9119) );
  XNOR2_X1 U11730 ( .A(n14490), .B(n9305), .ZN(n9130) );
  NAND2_X1 U11731 ( .A1(n9121), .A2(n13603), .ZN(n9122) );
  NAND2_X1 U11732 ( .A1(n9139), .A2(n9122), .ZN(n13844) );
  INV_X1 U11733 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9123) );
  OAI22_X1 U11734 ( .A1(n13844), .A2(n9326), .B1(n12539), .B2(n9123), .ZN(
        n9126) );
  INV_X1 U11735 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11805) );
  INV_X1 U11736 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9124) );
  OAI22_X1 U11737 ( .A1(n9379), .A2(n11805), .B1(n9162), .B2(n9124), .ZN(n9125) );
  NAND2_X1 U11738 ( .A1(n14010), .A2(n9166), .ZN(n9129) );
  XNOR2_X1 U11739 ( .A(n9130), .B(n9129), .ZN(n13843) );
  INV_X1 U11740 ( .A(n13843), .ZN(n9127) );
  NAND2_X1 U11741 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  NAND2_X1 U11742 ( .A1(n11257), .A2(n9302), .ZN(n9137) );
  NAND2_X1 U11743 ( .A1(n6629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9134) );
  XNOR2_X1 U11744 ( .A(n9134), .B(n9133), .ZN(n11808) );
  OAI22_X1 U11745 ( .A1(n9191), .A2(n11308), .B1(n8940), .B2(n11808), .ZN(
        n9135) );
  INV_X1 U11746 ( .A(n9135), .ZN(n9136) );
  XNOR2_X1 U11747 ( .A(n13999), .B(n8899), .ZN(n13896) );
  INV_X1 U11748 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14485) );
  INV_X1 U11749 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n14122) );
  NAND2_X1 U11750 ( .A1(n9139), .A2(n14122), .ZN(n9140) );
  NAND2_X1 U11751 ( .A1(n9148), .A2(n9140), .ZN(n13992) );
  OR2_X1 U11752 ( .A1(n13992), .A2(n9326), .ZN(n9142) );
  AOI22_X1 U11753 ( .A1(n9991), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n9375), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n9141) );
  OAI211_X1 U11754 ( .C1(n9379), .C2(n14485), .A(n9142), .B(n9141), .ZN(n14377) );
  AND2_X1 U11755 ( .A1(n14377), .A2(n9166), .ZN(n13988) );
  NAND2_X1 U11756 ( .A1(n11120), .A2(n9302), .ZN(n9147) );
  INV_X1 U11757 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U11758 ( .A1(n9144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9145) );
  XNOR2_X1 U11759 ( .A(n9145), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U11760 ( .A1(n12550), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n11049), 
        .B2(n14143), .ZN(n9146) );
  XNOR2_X1 U11761 ( .A(n14477), .B(n9305), .ZN(n13895) );
  INV_X1 U11762 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U11763 ( .A1(n9148), .A2(n7074), .ZN(n9149) );
  NAND2_X1 U11764 ( .A1(n9158), .A2(n9149), .ZN(n14384) );
  OR2_X1 U11765 ( .A1(n14384), .A2(n9326), .ZN(n9151) );
  AOI22_X1 U11766 ( .A1(n9991), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n9375), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n9150) );
  OAI211_X1 U11767 ( .C1(n9379), .C2(n11811), .A(n9151), .B(n9150), .ZN(n14359) );
  NAND2_X1 U11768 ( .A1(n14359), .A2(n9166), .ZN(n13894) );
  NAND2_X1 U11769 ( .A1(n13895), .A2(n13894), .ZN(n13907) );
  OAI21_X1 U11770 ( .B1(n13896), .B2(n13988), .A(n13907), .ZN(n9170) );
  NAND2_X1 U11771 ( .A1(n13896), .A2(n13988), .ZN(n9168) );
  NAND2_X1 U11772 ( .A1(n9168), .A2(n13894), .ZN(n9153) );
  INV_X1 U11773 ( .A(n13895), .ZN(n9152) );
  NAND2_X1 U11774 ( .A1(n9153), .A2(n9152), .ZN(n9167) );
  NAND2_X1 U11775 ( .A1(n11305), .A2(n9302), .ZN(n9157) );
  NAND2_X1 U11776 ( .A1(n9154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9155) );
  XNOR2_X1 U11777 ( .A(n9155), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15706) );
  AOI22_X1 U11778 ( .A1(n15706), .A2(n11049), .B1(n12550), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n9156) );
  XNOR2_X1 U11779 ( .A(n14546), .B(n8899), .ZN(n9173) );
  NAND2_X1 U11780 ( .A1(n9158), .A2(n13914), .ZN(n9159) );
  AND2_X1 U11781 ( .A1(n9180), .A2(n9159), .ZN(n14365) );
  NAND2_X1 U11782 ( .A1(n14365), .A2(n9374), .ZN(n9165) );
  INV_X1 U11783 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U11784 ( .A1(n6474), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11785 ( .A1(n9991), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9160) );
  OAI211_X1 U11786 ( .C1(n9162), .C2(n14134), .A(n9161), .B(n9160), .ZN(n9163)
         );
  INV_X1 U11787 ( .A(n9163), .ZN(n9164) );
  INV_X1 U11788 ( .A(n9166), .ZN(n9315) );
  NOR2_X1 U11789 ( .A1(n14330), .A2(n9315), .ZN(n9171) );
  XNOR2_X1 U11790 ( .A(n9173), .B(n9171), .ZN(n13908) );
  OAI211_X1 U11791 ( .C1(n13894), .C2(n9168), .A(n9167), .B(n13908), .ZN(n9169) );
  INV_X1 U11792 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U11793 ( .A1(n9173), .A2(n9172), .ZN(n9174) );
  NAND2_X1 U11794 ( .A1(n11309), .A2(n9302), .ZN(n9177) );
  OAI21_X1 U11795 ( .B1(n9154), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9175) );
  XNOR2_X1 U11796 ( .A(n9175), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U11797 ( .A1(n14147), .A2(n11049), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n12550), .ZN(n9176) );
  XNOR2_X1 U11798 ( .A(n14466), .B(n8899), .ZN(n9189) );
  INV_X1 U11799 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11800 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U11801 ( .A1(n9209), .A2(n9181), .ZN(n14344) );
  OR2_X1 U11802 ( .A1(n14344), .A2(n9326), .ZN(n9186) );
  INV_X1 U11803 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U11804 ( .A1(n9991), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11805 ( .A1(n9375), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9182) );
  OAI211_X1 U11806 ( .C1(n14150), .C2(n9379), .A(n9183), .B(n9182), .ZN(n9184)
         );
  INV_X1 U11807 ( .A(n9184), .ZN(n9185) );
  NAND2_X1 U11808 ( .A1(n14360), .A2(n9166), .ZN(n9187) );
  XNOR2_X1 U11809 ( .A(n9189), .B(n9187), .ZN(n13967) );
  INV_X1 U11810 ( .A(n9187), .ZN(n9188) );
  NAND2_X1 U11811 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  NAND2_X1 U11812 ( .A1(n11407), .A2(n9302), .ZN(n9194) );
  OAI22_X1 U11813 ( .A1(n12630), .A2(n8940), .B1(n9191), .B2(n11408), .ZN(
        n9192) );
  INV_X1 U11814 ( .A(n9192), .ZN(n9193) );
  XNOR2_X1 U11815 ( .A(n14321), .B(n9305), .ZN(n9200) );
  XNOR2_X1 U11816 ( .A(n9209), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U11817 ( .A1(n14322), .A2(n9374), .ZN(n9199) );
  INV_X1 U11818 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U11819 ( .A1(n9991), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U11820 ( .A1(n9375), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9195) );
  OAI211_X1 U11821 ( .C1(n14463), .C2(n9379), .A(n9196), .B(n9195), .ZN(n9197)
         );
  INV_X1 U11822 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U11823 ( .A1(n9199), .A2(n9198), .ZN(n14009) );
  NAND2_X1 U11824 ( .A1(n14009), .A2(n9166), .ZN(n9201) );
  NAND2_X1 U11825 ( .A1(n9200), .A2(n9201), .ZN(n13870) );
  NAND2_X1 U11826 ( .A1(n13871), .A2(n13870), .ZN(n9204) );
  INV_X1 U11827 ( .A(n9200), .ZN(n9203) );
  INV_X1 U11828 ( .A(n9201), .ZN(n9202) );
  NAND2_X1 U11829 ( .A1(n9203), .A2(n9202), .ZN(n13869) );
  NAND2_X1 U11830 ( .A1(n11540), .A2(n9302), .ZN(n9206) );
  NAND2_X1 U11831 ( .A1(n12550), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9205) );
  XNOR2_X1 U11832 ( .A(n14308), .B(n9305), .ZN(n13935) );
  INV_X1 U11833 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9207) );
  INV_X1 U11834 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13938) );
  OAI21_X1 U11835 ( .B1(n9209), .B2(n9207), .A(n13938), .ZN(n9210) );
  NAND2_X1 U11836 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9208) );
  AND2_X1 U11837 ( .A1(n9210), .A2(n9231), .ZN(n14305) );
  NAND2_X1 U11838 ( .A1(n14305), .A2(n9374), .ZN(n9216) );
  INV_X1 U11839 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U11840 ( .A1(n9991), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11841 ( .A1(n9375), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9211) );
  OAI211_X1 U11842 ( .C1(n9213), .C2(n9379), .A(n9212), .B(n9211), .ZN(n9214)
         );
  INV_X1 U11843 ( .A(n9214), .ZN(n9215) );
  INV_X1 U11844 ( .A(n14315), .ZN(n14284) );
  NAND2_X1 U11845 ( .A1(n14284), .A2(n9166), .ZN(n13934) );
  XNOR2_X1 U11846 ( .A(n9218), .B(n9217), .ZN(n11874) );
  NAND2_X1 U11847 ( .A1(n11874), .A2(n9302), .ZN(n9220) );
  NAND2_X1 U11848 ( .A1(n12550), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9219) );
  XNOR2_X1 U11849 ( .A(n14277), .B(n8899), .ZN(n13947) );
  INV_X1 U11850 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13951) );
  NAND2_X1 U11851 ( .A1(n9233), .A2(n13951), .ZN(n9222) );
  NAND2_X1 U11852 ( .A1(n9239), .A2(n9222), .ZN(n14270) );
  OR2_X1 U11853 ( .A1(n14270), .A2(n9326), .ZN(n9227) );
  INV_X1 U11854 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U11855 ( .A1(n9375), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11856 ( .A1(n9991), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9223) );
  OAI211_X1 U11857 ( .C1(n14447), .C2(n9379), .A(n9224), .B(n9223), .ZN(n9225)
         );
  INV_X1 U11858 ( .A(n9225), .ZN(n9226) );
  NAND2_X1 U11859 ( .A1(n9227), .A2(n9226), .ZN(n14285) );
  AND2_X1 U11860 ( .A1(n14285), .A2(n9166), .ZN(n13946) );
  NAND2_X1 U11861 ( .A1(n11705), .A2(n9302), .ZN(n9229) );
  NAND2_X1 U11862 ( .A1(n12550), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9228) );
  XNOR2_X1 U11863 ( .A(n14537), .B(n9305), .ZN(n9258) );
  INV_X1 U11864 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U11865 ( .A1(n9231), .A2(n9230), .ZN(n9232) );
  NAND2_X1 U11866 ( .A1(n9233), .A2(n9232), .ZN(n14291) );
  OR2_X1 U11867 ( .A1(n14291), .A2(n9326), .ZN(n9238) );
  INV_X1 U11868 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14452) );
  NAND2_X1 U11869 ( .A1(n9991), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U11870 ( .A1(n9375), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9234) );
  OAI211_X1 U11871 ( .C1(n14452), .C2(n9379), .A(n9235), .B(n9234), .ZN(n9236)
         );
  INV_X1 U11872 ( .A(n9236), .ZN(n9237) );
  NOR2_X1 U11873 ( .A1(n14303), .A2(n9315), .ZN(n9259) );
  AND2_X1 U11874 ( .A1(n9258), .A2(n9259), .ZN(n13945) );
  AOI21_X1 U11875 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n13852) );
  INV_X1 U11876 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13857) );
  NAND2_X1 U11877 ( .A1(n9239), .A2(n13857), .ZN(n9240) );
  NAND2_X1 U11878 ( .A1(n9250), .A2(n9240), .ZN(n14257) );
  INV_X1 U11879 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11880 ( .A1(n9375), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U11881 ( .A1(n9991), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9241) );
  OAI211_X1 U11882 ( .C1(n9379), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9244)
         );
  INV_X1 U11883 ( .A(n9244), .ZN(n9245) );
  AND2_X1 U11884 ( .A1(n14227), .A2(n9166), .ZN(n13854) );
  NAND2_X1 U11885 ( .A1(n12550), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9247) );
  XNOR2_X1 U11886 ( .A(n14440), .B(n8899), .ZN(n13919) );
  NAND2_X1 U11887 ( .A1(n12228), .A2(n9302), .ZN(n9249) );
  NAND2_X1 U11888 ( .A1(n12550), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9248) );
  XNOR2_X1 U11889 ( .A(n14233), .B(n8899), .ZN(n9266) );
  INV_X1 U11890 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U11891 ( .A1(n9250), .A2(n13927), .ZN(n9251) );
  AND2_X1 U11892 ( .A1(n9276), .A2(n9251), .ZN(n14231) );
  NAND2_X1 U11893 ( .A1(n14231), .A2(n9374), .ZN(n9257) );
  INV_X1 U11894 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11895 ( .A1(n9375), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11896 ( .A1(n9991), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9252) );
  OAI211_X1 U11897 ( .C1(n9379), .C2(n9254), .A(n9253), .B(n9252), .ZN(n9255)
         );
  INV_X1 U11898 ( .A(n9255), .ZN(n9256) );
  OR2_X1 U11899 ( .A1(n14256), .A2(n9315), .ZN(n9267) );
  NAND2_X1 U11900 ( .A1(n9266), .A2(n9267), .ZN(n13924) );
  INV_X1 U11901 ( .A(n9258), .ZN(n9261) );
  INV_X1 U11902 ( .A(n9259), .ZN(n9260) );
  XNOR2_X1 U11903 ( .A(n9261), .B(n9260), .ZN(n13879) );
  INV_X1 U11904 ( .A(n13947), .ZN(n9263) );
  INV_X1 U11905 ( .A(n13946), .ZN(n9262) );
  AND2_X1 U11906 ( .A1(n9263), .A2(n9262), .ZN(n13851) );
  AOI21_X1 U11907 ( .B1(n13852), .B2(n13879), .A(n13851), .ZN(n9264) );
  OAI211_X1 U11908 ( .C1(n13854), .C2(n13919), .A(n13924), .B(n9264), .ZN(
        n9265) );
  AOI21_X1 U11909 ( .B1(n13878), .B2(n13852), .A(n9265), .ZN(n9272) );
  NAND3_X1 U11910 ( .A1(n13924), .A2(n13854), .A3(n13919), .ZN(n9270) );
  INV_X1 U11911 ( .A(n9266), .ZN(n9269) );
  INV_X1 U11912 ( .A(n9267), .ZN(n9268) );
  NAND2_X1 U11913 ( .A1(n9269), .A2(n9268), .ZN(n13923) );
  NAND2_X1 U11914 ( .A1(n9270), .A2(n13923), .ZN(n9271) );
  NAND2_X1 U11915 ( .A1(n12282), .A2(n9302), .ZN(n9274) );
  NAND2_X1 U11916 ( .A1(n12550), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9273) );
  XNOR2_X1 U11917 ( .A(n14527), .B(n9305), .ZN(n9283) );
  INV_X1 U11918 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U11919 ( .A1(n9276), .A2(n13888), .ZN(n9277) );
  NAND2_X1 U11920 ( .A1(n9291), .A2(n9277), .ZN(n14218) );
  INV_X1 U11921 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U11922 ( .A1(n9991), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11923 ( .A1(n9375), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9278) );
  OAI211_X1 U11924 ( .C1(n14432), .C2(n9379), .A(n9279), .B(n9278), .ZN(n9280)
         );
  INV_X1 U11925 ( .A(n9280), .ZN(n9281) );
  NOR2_X1 U11926 ( .A1(n13980), .A2(n9315), .ZN(n9284) );
  NAND2_X1 U11927 ( .A1(n9283), .A2(n9284), .ZN(n9288) );
  INV_X1 U11928 ( .A(n9283), .ZN(n9286) );
  INV_X1 U11929 ( .A(n9284), .ZN(n9285) );
  NAND2_X1 U11930 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  AND2_X1 U11931 ( .A1(n9288), .A2(n9287), .ZN(n13886) );
  NAND2_X1 U11932 ( .A1(n14568), .A2(n9302), .ZN(n9290) );
  NAND2_X1 U11933 ( .A1(n12550), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U11934 ( .A(n14425), .B(n9305), .ZN(n9300) );
  INV_X1 U11935 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U11936 ( .A1(n9291), .A2(n13978), .ZN(n9292) );
  NAND2_X1 U11937 ( .A1(n9307), .A2(n9292), .ZN(n14201) );
  INV_X1 U11938 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U11939 ( .A1(n9991), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11940 ( .A1(n9375), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9293) );
  OAI211_X1 U11941 ( .C1(n9295), .C2(n9379), .A(n9294), .B(n9293), .ZN(n9296)
         );
  INV_X1 U11942 ( .A(n9296), .ZN(n9297) );
  NAND2_X1 U11943 ( .A1(n14006), .A2(n9166), .ZN(n9299) );
  XNOR2_X1 U11944 ( .A(n9300), .B(n9299), .ZN(n13977) );
  NAND2_X1 U11945 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  NAND2_X1 U11946 ( .A1(n12941), .A2(n9302), .ZN(n9304) );
  NAND2_X1 U11947 ( .A1(n12550), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9303) );
  AND2_X2 U11948 ( .A1(n9304), .A2(n9303), .ZN(n14190) );
  XNOR2_X1 U11949 ( .A(n14190), .B(n9305), .ZN(n9316) );
  INV_X1 U11950 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U11951 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  NAND2_X1 U11952 ( .A1(n14188), .A2(n9374), .ZN(n9314) );
  INV_X1 U11953 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11954 ( .A1(n9991), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11955 ( .A1(n9375), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9309) );
  OAI211_X1 U11956 ( .C1(n9311), .C2(n9379), .A(n9310), .B(n9309), .ZN(n9312)
         );
  INV_X1 U11957 ( .A(n9312), .ZN(n9313) );
  NOR2_X1 U11958 ( .A1(n13979), .A2(n9315), .ZN(n9317) );
  NAND2_X1 U11959 ( .A1(n9316), .A2(n9317), .ZN(n9368) );
  INV_X1 U11960 ( .A(n9316), .ZN(n9319) );
  INV_X1 U11961 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U11962 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  NAND2_X1 U11963 ( .A1(n9368), .A2(n9320), .ZN(n10055) );
  NAND2_X1 U11964 ( .A1(n12945), .A2(n9302), .ZN(n9322) );
  NAND2_X1 U11965 ( .A1(n12550), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9321) );
  INV_X1 U11966 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9389) );
  INV_X1 U11967 ( .A(n10049), .ZN(n9325) );
  NAND2_X1 U11968 ( .A1(n9323), .A2(n9389), .ZN(n9324) );
  NAND2_X1 U11969 ( .A1(n9325), .A2(n9324), .ZN(n12932) );
  NAND2_X1 U11970 ( .A1(n9991), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11971 ( .A1(n9375), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9327) );
  OAI211_X1 U11972 ( .C1(n10290), .C2(n9379), .A(n9328), .B(n9327), .ZN(n9329)
         );
  INV_X1 U11973 ( .A(n9329), .ZN(n9330) );
  NAND2_X1 U11974 ( .A1(n14005), .A2(n9166), .ZN(n9332) );
  XNOR2_X1 U11975 ( .A(n9332), .B(n8899), .ZN(n9333) );
  XNOR2_X1 U11976 ( .A(n12934), .B(n9333), .ZN(n9367) );
  NAND2_X1 U11977 ( .A1(n9334), .A2(n9344), .ZN(n9338) );
  NAND2_X1 U11978 ( .A1(n9340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9337) );
  XNOR2_X1 U11979 ( .A(n9337), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11980 ( .A1(n9338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9339) );
  MUX2_X1 U11981 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9339), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9341) );
  NAND2_X1 U11982 ( .A1(n9355), .A2(n9363), .ZN(n9342) );
  NAND2_X1 U11983 ( .A1(n9343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9345) );
  NOR4_X1 U11984 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9354) );
  OR4_X1 U11985 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n9351) );
  NOR4_X1 U11986 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9349) );
  NOR4_X1 U11987 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9348) );
  NOR4_X1 U11988 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9347) );
  NOR4_X1 U11989 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9346) );
  NAND4_X1 U11990 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n9350)
         );
  NOR4_X1 U11991 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9351), .A4(n9350), .ZN(n9353) );
  NOR4_X1 U11992 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9352) );
  NAND3_X1 U11993 ( .A1(n9354), .A2(n9353), .A3(n9352), .ZN(n9359) );
  INV_X1 U11994 ( .A(n14571), .ZN(n9358) );
  INV_X1 U11995 ( .A(P2_B_REG_SCAN_IN), .ZN(n9995) );
  XNOR2_X1 U11996 ( .A(n9363), .B(n9995), .ZN(n9356) );
  INV_X1 U11997 ( .A(n9355), .ZN(n12287) );
  NAND2_X1 U11998 ( .A1(n9356), .A2(n12287), .ZN(n9357) );
  NAND2_X1 U11999 ( .A1(n9359), .A2(n15716), .ZN(n10287) );
  NAND2_X1 U12000 ( .A1(n15722), .A2(n10287), .ZN(n9362) );
  INV_X1 U12001 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15725) );
  NAND2_X1 U12002 ( .A1(n15716), .A2(n15725), .ZN(n9361) );
  NAND2_X1 U12003 ( .A1(n14571), .A2(n12287), .ZN(n9360) );
  NAND2_X1 U12004 ( .A1(n9361), .A2(n9360), .ZN(n10284) );
  NOR2_X1 U12005 ( .A1(n9362), .A2(n10284), .ZN(n10001) );
  INV_X1 U12006 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15720) );
  NAND2_X1 U12007 ( .A1(n15716), .A2(n15720), .ZN(n9365) );
  INV_X1 U12008 ( .A(n9363), .ZN(n12233) );
  NAND2_X1 U12009 ( .A1(n14571), .A2(n12233), .ZN(n9364) );
  NAND2_X1 U12010 ( .A1(n10001), .A2(n10289), .ZN(n9383) );
  NAND2_X1 U12011 ( .A1(n12630), .A2(n12626), .ZN(n12640) );
  NAND4_X1 U12012 ( .A1(n9366), .A2(n9367), .A3(n9368), .A4(n13986), .ZN(n9395) );
  INV_X1 U12013 ( .A(n9367), .ZN(n9369) );
  NAND3_X1 U12014 ( .A1(n10062), .A2(n13986), .A3(n9369), .ZN(n9394) );
  INV_X1 U12015 ( .A(n9368), .ZN(n9370) );
  NAND3_X1 U12016 ( .A1(n9370), .A2(n13986), .A3(n9369), .ZN(n9393) );
  INV_X1 U12017 ( .A(n12626), .ZN(n12636) );
  AND3_X1 U12018 ( .A1(n12625), .A2(n12636), .A3(n8895), .ZN(n10048) );
  INV_X1 U12019 ( .A(n10048), .ZN(n9371) );
  OR2_X1 U12020 ( .A1(n9383), .A2(n9371), .ZN(n9373) );
  NAND2_X1 U12021 ( .A1(n14273), .A2(n14386), .ZN(n10286) );
  INV_X1 U12022 ( .A(n10286), .ZN(n9372) );
  INV_X1 U12023 ( .A(n11054), .ZN(n11074) );
  NAND2_X1 U12024 ( .A1(n10049), .A2(n9374), .ZN(n9382) );
  INV_X1 U12025 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U12026 ( .A1(n9991), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U12027 ( .A1(n9375), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9376) );
  OAI211_X1 U12028 ( .C1(n9379), .C2(n9378), .A(n9377), .B(n9376), .ZN(n9380)
         );
  INV_X1 U12029 ( .A(n9380), .ZN(n9381) );
  NAND2_X1 U12030 ( .A1(n9382), .A2(n9381), .ZN(n14004) );
  AOI22_X1 U12031 ( .A1(n14196), .A2(n14376), .B1(n14374), .B2(n14004), .ZN(
        n10281) );
  NOR2_X1 U12032 ( .A1(n10281), .A2(n13952), .ZN(n9391) );
  INV_X1 U12033 ( .A(n10284), .ZN(n9384) );
  NAND3_X1 U12034 ( .A1(n10289), .A2(n9384), .A3(n10287), .ZN(n9385) );
  NAND2_X1 U12035 ( .A1(n9385), .A2(n10286), .ZN(n9388) );
  NAND2_X1 U12036 ( .A1(n11051), .A2(n12640), .ZN(n10285) );
  AND2_X1 U12037 ( .A1(n9386), .A2(n10285), .ZN(n9387) );
  NAND2_X1 U12038 ( .A1(n9388), .A2(n9387), .ZN(n11392) );
  OAI22_X1 U12039 ( .A1(n12932), .A2(n13993), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9389), .ZN(n9390) );
  AOI211_X1 U12040 ( .C1(n12934), .C2(n13998), .A(n9391), .B(n9390), .ZN(n9392) );
  NAND4_X1 U12041 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(
        P2_U3192) );
  NOR2_X1 U12042 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n9398) );
  NAND4_X1 U12043 ( .A1(n9398), .A2(n9397), .A3(n9396), .A4(n9476), .ZN(n9399)
         );
  NOR2_X1 U12044 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n9402) );
  NAND4_X1 U12045 ( .A1(n9402), .A2(n9401), .A3(n9400), .A4(n9554), .ZN(n9405)
         );
  NAND4_X1 U12046 ( .A1(n9609), .A2(n9403), .A3(n9593), .A4(n9552), .ZN(n9404)
         );
  NAND2_X1 U12047 ( .A1(n9598), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9414) );
  XNOR2_X1 U12048 ( .A(n9469), .B(n9468), .ZN(n10773) );
  NAND2_X1 U12049 ( .A1(n9533), .A2(n10773), .ZN(n9425) );
  NAND2_X1 U12050 ( .A1(n9484), .A2(n10676), .ZN(n9423) );
  NAND2_X1 U12051 ( .A1(n13127), .A2(n15807), .ZN(n10475) );
  INV_X1 U12052 ( .A(n9433), .ZN(n9430) );
  NAND2_X1 U12053 ( .A1(n9905), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9428) );
  MUX2_X1 U12054 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9428), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9429) );
  XNOR2_X1 U12055 ( .A(n9442), .B(P3_B_REG_SCAN_IN), .ZN(n9435) );
  NAND2_X1 U12056 ( .A1(n9433), .A2(n9432), .ZN(n9436) );
  NAND2_X1 U12057 ( .A1(n9436), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9437) );
  INV_X1 U12059 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U12060 ( .A1(n9878), .A2(n9441), .ZN(n9444) );
  NAND2_X1 U12061 ( .A1(n13834), .A2(n9442), .ZN(n9443) );
  NAND2_X1 U12062 ( .A1(n9446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U12063 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9445), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9447) );
  NAND2_X1 U12064 ( .A1(n9426), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9449) );
  INV_X1 U12065 ( .A(n11454), .ZN(n10212) );
  NAND2_X1 U12066 ( .A1(n11660), .A2(n10212), .ZN(n10464) );
  INV_X1 U12067 ( .A(n10464), .ZN(n9450) );
  XNOR2_X2 U12068 ( .A(n9453), .B(n9452), .ZN(n13312) );
  INV_X1 U12069 ( .A(n11660), .ZN(n10213) );
  OAI21_X1 U12070 ( .B1(n13312), .B2(n10213), .A(n11454), .ZN(n9454) );
  INV_X1 U12071 ( .A(n9468), .ZN(n9458) );
  NAND2_X1 U12072 ( .A1(n9456), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U12073 ( .A1(n9458), .A2(n9457), .ZN(n9459) );
  MUX2_X1 U12074 ( .A(n9459), .B(SI_0_), .S(n10071), .Z(n13839) );
  MUX2_X1 U12075 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13839), .S(n10622), .Z(n9466)
         );
  INV_X1 U12076 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9460) );
  OR2_X1 U12077 ( .A1(n9506), .A2(n9460), .ZN(n9464) );
  NAND2_X1 U12078 ( .A1(n9598), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U12079 ( .A1(n15798), .A2(n9466), .ZN(n15800) );
  NAND2_X1 U12080 ( .A1(n12896), .A2(n15800), .ZN(n9467) );
  AND2_X1 U12081 ( .A1(n10223), .A2(n9467), .ZN(n11107) );
  NAND2_X1 U12082 ( .A1(n10423), .A2(n10792), .ZN(n9477) );
  NAND2_X1 U12083 ( .A1(n10748), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12084 ( .A1(n9471), .A2(n9470), .ZN(n9482) );
  INV_X1 U12085 ( .A(n9481), .ZN(n9473) );
  NAND2_X1 U12086 ( .A1(n13590), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9474) );
  XNOR2_X1 U12087 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .ZN(n9498) );
  XNOR2_X1 U12088 ( .A(n9499), .B(n7912), .ZN(n10793) );
  XNOR2_X1 U12089 ( .A(n11448), .B(n11109), .ZN(n11294) );
  NAND2_X1 U12090 ( .A1(n9744), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9480) );
  INV_X1 U12091 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15864) );
  OR2_X1 U12092 ( .A1(n9506), .A2(n15864), .ZN(n9478) );
  XNOR2_X1 U12093 ( .A(n9482), .B(n9481), .ZN(n10795) );
  NAND2_X1 U12094 ( .A1(n9533), .A2(n10795), .ZN(n9486) );
  NAND2_X1 U12095 ( .A1(n9484), .A2(n10999), .ZN(n9485) );
  INV_X1 U12096 ( .A(n15790), .ZN(n10479) );
  XNOR2_X1 U12097 ( .A(n11109), .B(n10479), .ZN(n11216) );
  INV_X1 U12098 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9487) );
  INV_X1 U12099 ( .A(n15797), .ZN(n11441) );
  NAND4_X1 U12100 ( .A1(n11218), .A2(n11107), .A3(n9494), .A4(n11295), .ZN(
        n9497) );
  INV_X1 U12101 ( .A(n11294), .ZN(n9492) );
  XNOR2_X1 U12102 ( .A(n10780), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n9515) );
  XNOR2_X1 U12103 ( .A(n9517), .B(n9515), .ZN(n10787) );
  NAND2_X1 U12104 ( .A1(n9533), .A2(n10787), .ZN(n9503) );
  NAND2_X1 U12105 ( .A1(n9484), .A2(n10788), .ZN(n9502) );
  INV_X1 U12106 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9505) );
  AND2_X1 U12107 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9509) );
  NOR2_X1 U12108 ( .A1(n9525), .A2(n9509), .ZN(n11510) );
  INV_X1 U12109 ( .A(n11510), .ZN(n9510) );
  INV_X1 U12110 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U12111 ( .A1(n9512), .A2(n11365), .ZN(n9513) );
  INV_X1 U12112 ( .A(n9515), .ZN(n9516) );
  NAND2_X1 U12113 ( .A1(n10743), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9518) );
  XNOR2_X1 U12114 ( .A(n10753), .B(P2_DATAO_REG_5__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U12115 ( .A(n9536), .B(n9534), .ZN(n10790) );
  NAND2_X1 U12116 ( .A1(n9533), .A2(n10790), .ZN(n9523) );
  NAND2_X1 U12117 ( .A1(n9519), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U12118 ( .A(n9521), .B(n9520), .ZN(n10791) );
  NAND2_X1 U12119 ( .A1(n9484), .A2(n10791), .ZN(n9522) );
  OAI211_X1 U12120 ( .C1(n9708), .C2(SI_5_), .A(n9523), .B(n9522), .ZN(n11547)
         );
  INV_X2 U12121 ( .A(n9506), .ZN(n10415) );
  NAND2_X1 U12122 ( .A1(n10415), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U12123 ( .A1(n9744), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9529) );
  OR2_X1 U12124 ( .A1(n9525), .A2(n9524), .ZN(n9526) );
  NAND2_X1 U12125 ( .A1(n9544), .A2(n9526), .ZN(n11518) );
  NAND2_X1 U12126 ( .A1(n10180), .A2(n11518), .ZN(n9528) );
  INV_X1 U12127 ( .A(n13125), .ZN(n11243) );
  NAND2_X1 U12128 ( .A1(n9531), .A2(n11243), .ZN(n9532) );
  INV_X1 U12129 ( .A(n9534), .ZN(n9535) );
  NAND2_X1 U12130 ( .A1(n10753), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9537) );
  XNOR2_X1 U12131 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9538) );
  XNOR2_X1 U12132 ( .A(n9557), .B(n9538), .ZN(n10770) );
  NAND2_X1 U12133 ( .A1(n10424), .A2(n10770), .ZN(n9543) );
  NAND2_X1 U12134 ( .A1(n10423), .A2(SI_6_), .ZN(n9542) );
  INV_X1 U12135 ( .A(n9553), .ZN(n9539) );
  NAND2_X1 U12136 ( .A1(n9539), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9540) );
  XNOR2_X1 U12137 ( .A(n9540), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10683) );
  NAND2_X1 U12138 ( .A1(n9484), .A2(n10683), .ZN(n9541) );
  XNOR2_X1 U12139 ( .A(n11109), .B(n10130), .ZN(n9550) );
  NAND2_X1 U12140 ( .A1(n10415), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12141 ( .A1(n9744), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U12142 ( .A1(n9544), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U12143 ( .A1(n9562), .A2(n9545), .ZN(n11621) );
  NAND2_X1 U12144 ( .A1(n10180), .A2(n11621), .ZN(n9547) );
  NAND2_X1 U12145 ( .A1(n10416), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9546) );
  NAND4_X1 U12146 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n13124) );
  INV_X1 U12147 ( .A(n13124), .ZN(n11673) );
  XNOR2_X1 U12148 ( .A(n9550), .B(n11673), .ZN(n11524) );
  NAND2_X1 U12149 ( .A1(n9550), .A2(n13124), .ZN(n9551) );
  INV_X1 U12150 ( .A(SI_7_), .ZN(n13591) );
  NAND2_X1 U12151 ( .A1(n9553), .A2(n9552), .ZN(n9574) );
  NAND2_X1 U12152 ( .A1(n9574), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9555) );
  XNOR2_X1 U12153 ( .A(n9554), .B(n9555), .ZN(n11238) );
  AOI22_X1 U12154 ( .A1(n10423), .A2(n13591), .B1(n9484), .B2(n11238), .ZN(
        n9560) );
  NAND2_X1 U12155 ( .A1(n10782), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9558) );
  XNOR2_X1 U12156 ( .A(n9573), .B(n9572), .ZN(n10876) );
  NAND2_X1 U12157 ( .A1(n10876), .A2(n10424), .ZN(n9559) );
  XNOR2_X1 U12158 ( .A(n11109), .B(n11607), .ZN(n9568) );
  NAND2_X1 U12159 ( .A1(n10207), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U12160 ( .A1(n10191), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9566) );
  INV_X1 U12161 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15869) );
  OR2_X1 U12162 ( .A1(n9506), .A2(n15869), .ZN(n9565) );
  AND2_X1 U12163 ( .A1(n9562), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9563) );
  NOR2_X1 U12164 ( .A1(n9599), .A2(n9563), .ZN(n11608) );
  OR2_X1 U12165 ( .A1(n9561), .A2(n11608), .ZN(n9564) );
  XNOR2_X1 U12166 ( .A(n9568), .B(n13123), .ZN(n11670) );
  INV_X1 U12167 ( .A(n9568), .ZN(n9569) );
  NAND2_X1 U12168 ( .A1(n9569), .A2(n13123), .ZN(n9570) );
  NAND2_X1 U12169 ( .A1(n9571), .A2(n9570), .ZN(n11745) );
  XNOR2_X1 U12170 ( .A(n10765), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n9586) );
  XNOR2_X1 U12171 ( .A(n9588), .B(n9586), .ZN(n10873) );
  NAND2_X1 U12172 ( .A1(n10873), .A2(n10424), .ZN(n9577) );
  NAND2_X1 U12173 ( .A1(n9590), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9575) );
  XNOR2_X1 U12174 ( .A(n9575), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U12175 ( .A1(n6931), .A2(SI_8_), .B1(n9484), .B2(n10687), .ZN(n9576) );
  NAND2_X1 U12176 ( .A1(n9577), .A2(n9576), .ZN(n11775) );
  XNOR2_X1 U12177 ( .A(n12895), .B(n11775), .ZN(n9582) );
  NAND2_X1 U12178 ( .A1(n10207), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U12179 ( .A1(n10191), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9580) );
  XNOR2_X1 U12180 ( .A(n9599), .B(n11747), .ZN(n11776) );
  NAND2_X1 U12181 ( .A1(n10180), .A2(n11776), .ZN(n9579) );
  NAND2_X1 U12182 ( .A1(n10415), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U12183 ( .A(n9582), .B(n13122), .ZN(n11746) );
  INV_X1 U12184 ( .A(n9582), .ZN(n9583) );
  NAND2_X1 U12185 ( .A1(n9583), .A2(n13122), .ZN(n9584) );
  INV_X1 U12186 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12187 ( .A1(n10765), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9589) );
  XNOR2_X1 U12188 ( .A(n9608), .B(n9607), .ZN(n10878) );
  NAND2_X1 U12189 ( .A1(n10878), .A2(n10424), .ZN(n9597) );
  INV_X1 U12190 ( .A(n9594), .ZN(n9591) );
  NAND2_X1 U12191 ( .A1(n9591), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U12192 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9592), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9595) );
  NAND2_X1 U12193 ( .A1(n9594), .A2(n9593), .ZN(n9628) );
  NAND2_X1 U12194 ( .A1(n9595), .A2(n9628), .ZN(n11490) );
  INV_X1 U12195 ( .A(SI_9_), .ZN(n10877) );
  AOI22_X1 U12196 ( .A1(n9484), .A2(n11490), .B1(n10423), .B2(n10877), .ZN(
        n9596) );
  NAND2_X1 U12197 ( .A1(n9597), .A2(n9596), .ZN(n12107) );
  XNOR2_X1 U12198 ( .A(n12107), .B(n12895), .ZN(n9620) );
  NAND2_X1 U12199 ( .A1(n10207), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U12200 ( .A1(n10415), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12201 ( .A1(n10416), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9603) );
  OR2_X1 U12202 ( .A1(n9600), .A2(n11488), .ZN(n9601) );
  AND2_X1 U12203 ( .A1(n9614), .A2(n9601), .ZN(n12046) );
  OR2_X1 U12204 ( .A1(n9561), .A2(n12046), .ZN(n9602) );
  XNOR2_X1 U12205 ( .A(n9620), .B(n13121), .ZN(n12041) );
  INV_X1 U12206 ( .A(n12041), .ZN(n9606) );
  XNOR2_X1 U12207 ( .A(n9625), .B(n9624), .ZN(n10872) );
  NAND2_X1 U12208 ( .A1(n10872), .A2(n10424), .ZN(n9613) );
  NAND2_X1 U12209 ( .A1(n9628), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9610) );
  NOR2_X1 U12210 ( .A1(n9708), .A2(SI_10_), .ZN(n9611) );
  AOI21_X1 U12211 ( .B1(n11869), .B2(n9484), .A(n9611), .ZN(n9612) );
  NAND2_X1 U12212 ( .A1(n9613), .A2(n9612), .ZN(n12143) );
  XNOR2_X1 U12213 ( .A(n12143), .B(n12896), .ZN(n9622) );
  NAND2_X1 U12214 ( .A1(n9744), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U12215 ( .A1(n10415), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12216 ( .A1(n9614), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U12217 ( .A1(n9631), .A2(n9615), .ZN(n12136) );
  NAND2_X1 U12218 ( .A1(n10180), .A2(n12136), .ZN(n9617) );
  NAND2_X1 U12219 ( .A1(n10416), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9616) );
  NAND4_X1 U12220 ( .A1(n9619), .A2(n9618), .A3(n9617), .A4(n9616), .ZN(n13120) );
  XNOR2_X1 U12221 ( .A(n9622), .B(n13120), .ZN(n11984) );
  OR2_X1 U12222 ( .A1(n9620), .A2(n13121), .ZN(n11985) );
  AND2_X1 U12223 ( .A1(n11984), .A2(n11985), .ZN(n9621) );
  INV_X1 U12224 ( .A(n9622), .ZN(n9623) );
  NAND2_X1 U12225 ( .A1(n9623), .A2(n13120), .ZN(n9638) );
  NAND2_X1 U12226 ( .A1(n9625), .A2(n9624), .ZN(n9627) );
  NAND2_X1 U12227 ( .A1(n10837), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9626) );
  XNOR2_X1 U12228 ( .A(n9642), .B(n9641), .ZN(n10864) );
  NAND2_X1 U12229 ( .A1(n6476), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9629) );
  XNOR2_X1 U12230 ( .A(n9629), .B(P3_IR_REG_11__SCAN_IN), .ZN(n10658) );
  OAI22_X1 U12231 ( .A1(n10658), .A2(n10622), .B1(SI_11_), .B2(n9708), .ZN(
        n9630) );
  AOI21_X2 U12232 ( .B1(n10864), .B2(n10424), .A(n9630), .ZN(n13753) );
  XNOR2_X1 U12233 ( .A(n13753), .B(n12896), .ZN(n9637) );
  NAND2_X1 U12234 ( .A1(n10415), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12235 ( .A1(n9744), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12236 ( .A1(n9631), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12237 ( .A1(n9647), .A2(n9632), .ZN(n13065) );
  NAND2_X1 U12238 ( .A1(n10180), .A2(n13065), .ZN(n9634) );
  NAND2_X1 U12239 ( .A1(n10191), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9633) );
  NAND4_X1 U12240 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), .ZN(n13119) );
  INV_X1 U12241 ( .A(n13119), .ZN(n13060) );
  INV_X1 U12242 ( .A(n9637), .ZN(n9639) );
  AND2_X1 U12243 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  NAND2_X1 U12244 ( .A1(n12993), .A2(n13063), .ZN(n9654) );
  NAND2_X1 U12245 ( .A1(n10866), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9643) );
  XNOR2_X1 U12246 ( .A(n10914), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U12247 ( .A(n9659), .B(n9657), .ZN(n10859) );
  NAND2_X1 U12248 ( .A1(n10859), .A2(n10424), .ZN(n9646) );
  XNOR2_X2 U12249 ( .A(n9644), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U12250 ( .A1(n13190), .A2(n9484), .B1(n10423), .B2(SI_12_), .ZN(
        n9645) );
  XNOR2_X1 U12251 ( .A(n12201), .B(n12895), .ZN(n9655) );
  NAND2_X1 U12252 ( .A1(n10415), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U12253 ( .A1(n10207), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9652) );
  INV_X1 U12254 ( .A(n9680), .ZN(n9649) );
  NAND2_X1 U12255 ( .A1(n9647), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U12256 ( .A1(n9649), .A2(n9648), .ZN(n13531) );
  NAND2_X1 U12257 ( .A1(n10180), .A2(n13531), .ZN(n9651) );
  NAND2_X1 U12258 ( .A1(n10191), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9650) );
  NAND4_X1 U12259 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n13118) );
  XNOR2_X1 U12260 ( .A(n9655), .B(n13118), .ZN(n12994) );
  NAND2_X1 U12261 ( .A1(n9655), .A2(n12211), .ZN(n9656) );
  INV_X1 U12262 ( .A(n9657), .ZN(n9658) );
  XNOR2_X1 U12263 ( .A(n9701), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U12264 ( .A1(n9687), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12265 ( .A1(n9701), .A2(n10980), .ZN(n9660) );
  NAND2_X1 U12266 ( .A1(n9661), .A2(n9660), .ZN(n9663) );
  XNOR2_X1 U12267 ( .A(n11206), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n9662) );
  XNOR2_X1 U12268 ( .A(n9663), .B(n9662), .ZN(n10971) );
  NAND2_X1 U12269 ( .A1(n10971), .A2(n10424), .ZN(n9672) );
  INV_X1 U12270 ( .A(n9664), .ZN(n9666) );
  INV_X1 U12271 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U12272 ( .A1(n9666), .A2(n9665), .ZN(n9688) );
  INV_X1 U12273 ( .A(n9688), .ZN(n9668) );
  INV_X1 U12274 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U12275 ( .A1(n9668), .A2(n9667), .ZN(n9706) );
  NAND2_X1 U12276 ( .A1(n9706), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9669) );
  NOR2_X1 U12277 ( .A1(n9708), .A2(n10972), .ZN(n9670) );
  AOI21_X1 U12278 ( .B1(n13230), .B2(n9484), .A(n9670), .ZN(n9671) );
  XNOR2_X1 U12279 ( .A(n13523), .B(n12896), .ZN(n12959) );
  NAND2_X1 U12280 ( .A1(n10207), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U12281 ( .A1(n10191), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9673) );
  AND2_X1 U12282 ( .A1(n9674), .A2(n9673), .ZN(n9678) );
  NAND2_X1 U12283 ( .A1(n9682), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12284 ( .A1(n9712), .A2(n9675), .ZN(n13524) );
  NAND2_X1 U12285 ( .A1(n13524), .A2(n10180), .ZN(n9677) );
  NAND2_X1 U12286 ( .A1(n10415), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U12287 ( .A1(n10415), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12288 ( .A1(n10207), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9685) );
  OR2_X1 U12289 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U12290 ( .A1(n9682), .A2(n9681), .ZN(n13048) );
  NAND2_X1 U12291 ( .A1(n10180), .A2(n13048), .ZN(n9684) );
  NAND2_X1 U12292 ( .A1(n10191), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9683) );
  NAND4_X1 U12293 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n13117) );
  XNOR2_X1 U12294 ( .A(n9687), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U12295 ( .A1(n10892), .A2(n10424), .ZN(n9693) );
  NAND2_X1 U12296 ( .A1(n9688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9689) );
  MUX2_X1 U12297 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9689), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9690) );
  NAND2_X1 U12298 ( .A1(n9690), .A2(n9706), .ZN(n10893) );
  NOR2_X1 U12299 ( .A1(n9708), .A2(SI_13_), .ZN(n9691) );
  AOI21_X1 U12300 ( .B1(n10893), .B2(n9484), .A(n9691), .ZN(n9692) );
  XNOR2_X1 U12301 ( .A(n13814), .B(n12895), .ZN(n13042) );
  OAI22_X1 U12302 ( .A1(n12959), .A2(n13116), .B1(n13117), .B2(n13042), .ZN(
        n9694) );
  INV_X1 U12303 ( .A(n9694), .ZN(n9695) );
  INV_X1 U12304 ( .A(n13042), .ZN(n12956) );
  INV_X1 U12305 ( .A(n13117), .ZN(n13521) );
  OAI21_X1 U12306 ( .B1(n12956), .B2(n13521), .A(n13045), .ZN(n9697) );
  NOR2_X1 U12307 ( .A1(n13045), .A2(n13521), .ZN(n9696) );
  AOI22_X1 U12308 ( .A1(n9697), .A2(n12959), .B1(n9696), .B2(n13042), .ZN(
        n9698) );
  NAND2_X1 U12309 ( .A1(n11206), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U12310 ( .A1(n13593), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9699) );
  AND2_X1 U12311 ( .A1(n9702), .A2(n9699), .ZN(n9700) );
  AND2_X1 U12312 ( .A1(n10980), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U12313 ( .A1(n9703), .A2(n9702), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n11208), .ZN(n9704) );
  XNOR2_X1 U12314 ( .A(n11258), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n9717) );
  XNOR2_X1 U12315 ( .A(n9718), .B(n9717), .ZN(n10909) );
  NAND2_X1 U12316 ( .A1(n10909), .A2(n10424), .ZN(n9711) );
  OAI21_X1 U12317 ( .B1(n9706), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9707) );
  XNOR2_X1 U12318 ( .A(n9707), .B(P3_IR_REG_15__SCAN_IN), .ZN(n10697) );
  NOR2_X1 U12319 ( .A1(n9708), .A2(n13693), .ZN(n9709) );
  AOI21_X1 U12320 ( .B1(n10697), .B2(n9484), .A(n9709), .ZN(n9710) );
  XNOR2_X1 U12321 ( .A(n13510), .B(n12895), .ZN(n9716) );
  INV_X1 U12322 ( .A(n10191), .ZN(n9806) );
  INV_X1 U12323 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13805) );
  AND2_X1 U12324 ( .A1(n9712), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9713) );
  OR2_X1 U12325 ( .A1(n9713), .A2(n9725), .ZN(n13511) );
  NAND2_X1 U12326 ( .A1(n13511), .A2(n10180), .ZN(n9715) );
  AOI22_X1 U12327 ( .A1(n10207), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n10415), 
        .B2(P3_REG1_REG_15__SCAN_IN), .ZN(n9714) );
  OAI211_X1 U12328 ( .C1(n9806), .C2(n13805), .A(n9715), .B(n9714), .ZN(n13115) );
  XNOR2_X1 U12329 ( .A(n9716), .B(n13522), .ZN(n13093) );
  NAND2_X1 U12330 ( .A1(n11258), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9719) );
  XNOR2_X1 U12331 ( .A(n11121), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n9732) );
  XNOR2_X1 U12332 ( .A(n9734), .B(n9732), .ZN(n10956) );
  NAND2_X1 U12333 ( .A1(n10956), .A2(n10424), .ZN(n9723) );
  NAND2_X1 U12334 ( .A1(n9720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9721) );
  XNOR2_X1 U12335 ( .A(n9721), .B(P3_IR_REG_16__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U12336 ( .A1(n6931), .A2(SI_16_), .B1(n9484), .B2(n10699), .ZN(
        n9722) );
  XNOR2_X1 U12337 ( .A(n13497), .B(n12896), .ZN(n9729) );
  INV_X1 U12338 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13801) );
  NOR2_X1 U12339 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  OR2_X1 U12340 ( .A1(n9742), .A2(n9726), .ZN(n13498) );
  NAND2_X1 U12341 ( .A1(n13498), .A2(n10180), .ZN(n9728) );
  AOI22_X1 U12342 ( .A1(n10207), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n10415), 
        .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n9727) );
  OAI211_X1 U12343 ( .C1(n9806), .C2(n13801), .A(n9728), .B(n9727), .ZN(n13113) );
  NAND2_X1 U12344 ( .A1(n9729), .A2(n13113), .ZN(n13017) );
  INV_X1 U12345 ( .A(n9729), .ZN(n9730) );
  INV_X1 U12346 ( .A(n13113), .ZN(n13479) );
  NAND2_X1 U12347 ( .A1(n9730), .A2(n13479), .ZN(n13018) );
  INV_X1 U12348 ( .A(n9732), .ZN(n9733) );
  NAND2_X1 U12349 ( .A1(n11121), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9735) );
  XNOR2_X1 U12350 ( .A(n11306), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n9752) );
  XNOR2_X1 U12351 ( .A(n9754), .B(n9752), .ZN(n10975) );
  NAND2_X1 U12352 ( .A1(n10975), .A2(n10424), .ZN(n9740) );
  NAND2_X1 U12353 ( .A1(n9736), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9737) );
  MUX2_X1 U12354 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9737), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9738) );
  AND2_X1 U12355 ( .A1(n9738), .A2(n9755), .ZN(n10976) );
  AOI22_X1 U12356 ( .A1(n6931), .A2(SI_17_), .B1(n10976), .B2(n9484), .ZN(
        n9739) );
  XNOR2_X1 U12357 ( .A(n13484), .B(n12895), .ZN(n9750) );
  OR2_X1 U12358 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  NAND2_X1 U12359 ( .A1(n9759), .A2(n9743), .ZN(n13485) );
  NAND2_X1 U12360 ( .A1(n13485), .A2(n10180), .ZN(n9749) );
  INV_X1 U12361 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U12362 ( .A1(n10415), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12363 ( .A1(n10207), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9745) );
  OAI211_X1 U12364 ( .C1(n13797), .C2(n9806), .A(n9746), .B(n9745), .ZN(n9747)
         );
  INV_X1 U12365 ( .A(n9747), .ZN(n9748) );
  XNOR2_X1 U12366 ( .A(n9750), .B(n13469), .ZN(n13025) );
  INV_X1 U12367 ( .A(n9750), .ZN(n9751) );
  INV_X1 U12368 ( .A(n9752), .ZN(n9753) );
  XNOR2_X1 U12369 ( .A(n9768), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n9766) );
  XNOR2_X1 U12370 ( .A(n9767), .B(n9766), .ZN(n11116) );
  NAND2_X1 U12371 ( .A1(n11116), .A2(n10424), .ZN(n9758) );
  NAND2_X1 U12372 ( .A1(n9755), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9756) );
  XNOR2_X1 U12373 ( .A(n9756), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U12374 ( .A1(n6931), .A2(SI_18_), .B1(n13303), .B2(n9484), .ZN(
        n9757) );
  XNOR2_X1 U12375 ( .A(n13587), .B(n12895), .ZN(n9777) );
  NAND2_X1 U12376 ( .A1(n9759), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12377 ( .A1(n9771), .A2(n9760), .ZN(n13471) );
  NAND2_X1 U12378 ( .A1(n13471), .A2(n10180), .ZN(n9765) );
  INV_X1 U12379 ( .A(n10207), .ZN(n9860) );
  INV_X1 U12380 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U12381 ( .A1(n10415), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U12382 ( .A1(n10191), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9761) );
  OAI211_X1 U12383 ( .C1(n9860), .C2(n10702), .A(n9762), .B(n9761), .ZN(n9763)
         );
  INV_X1 U12384 ( .A(n9763), .ZN(n9764) );
  XNOR2_X1 U12385 ( .A(n9777), .B(n13111), .ZN(n13072) );
  XNOR2_X1 U12386 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .ZN(n9781) );
  XNOR2_X1 U12387 ( .A(n9782), .B(n9781), .ZN(n11194) );
  NAND2_X1 U12388 ( .A1(n11194), .A2(n10424), .ZN(n9770) );
  AOI22_X1 U12389 ( .A1(n13312), .A2(n9484), .B1(n10423), .B2(n11193), .ZN(
        n9769) );
  XNOR2_X1 U12390 ( .A(n13794), .B(n12895), .ZN(n9779) );
  AND2_X1 U12391 ( .A1(n9771), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9772) );
  OR2_X1 U12392 ( .A1(n9772), .A2(n9787), .ZN(n13458) );
  INV_X1 U12393 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12394 ( .A1(n10415), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U12395 ( .A1(n10191), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9773) );
  OAI211_X1 U12396 ( .C1(n9860), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9776)
         );
  XNOR2_X1 U12397 ( .A(n9779), .B(n13470), .ZN(n12976) );
  NAND2_X1 U12398 ( .A1(n9777), .A2(n13480), .ZN(n12974) );
  AND2_X1 U12399 ( .A1(n12976), .A2(n12974), .ZN(n9778) );
  INV_X1 U12400 ( .A(n13470), .ZN(n13110) );
  NAND2_X1 U12401 ( .A1(n9779), .A2(n13110), .ZN(n9780) );
  NAND2_X1 U12402 ( .A1(n9782), .A2(n9781), .ZN(n9784) );
  NAND2_X1 U12403 ( .A1(n11410), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9783) );
  XNOR2_X1 U12404 ( .A(n9797), .B(n11543), .ZN(n11452) );
  NAND2_X1 U12405 ( .A1(n11452), .A2(n10424), .ZN(n9786) );
  NAND2_X1 U12406 ( .A1(n10423), .A2(SI_20_), .ZN(n9785) );
  XNOR2_X1 U12407 ( .A(n13037), .B(n12895), .ZN(n9794) );
  NOR2_X1 U12408 ( .A1(n9787), .A2(n13036), .ZN(n9788) );
  OR2_X1 U12409 ( .A1(n9802), .A2(n9788), .ZN(n13446) );
  NAND2_X1 U12410 ( .A1(n13446), .A2(n10180), .ZN(n9793) );
  INV_X1 U12411 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U12412 ( .A1(n10415), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U12413 ( .A1(n10207), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9789) );
  OAI211_X1 U12414 ( .C1(n13788), .C2(n9806), .A(n9790), .B(n9789), .ZN(n9791)
         );
  INV_X1 U12415 ( .A(n9791), .ZN(n9792) );
  XNOR2_X1 U12416 ( .A(n9794), .B(n13109), .ZN(n13035) );
  INV_X1 U12417 ( .A(n9794), .ZN(n9795) );
  NAND2_X1 U12418 ( .A1(n9795), .A2(n13109), .ZN(n9796) );
  NAND2_X1 U12419 ( .A1(n9798), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9799) );
  XNOR2_X1 U12420 ( .A(n11706), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n9815) );
  XNOR2_X1 U12421 ( .A(n9816), .B(n9815), .ZN(n11658) );
  NAND2_X1 U12422 ( .A1(n11658), .A2(n10424), .ZN(n9801) );
  NAND2_X1 U12423 ( .A1(n10423), .A2(SI_21_), .ZN(n9800) );
  XNOR2_X1 U12424 ( .A(n12988), .B(n12895), .ZN(n9810) );
  OR2_X1 U12425 ( .A1(n9802), .A2(n12986), .ZN(n9803) );
  NAND2_X1 U12426 ( .A1(n9827), .A2(n9803), .ZN(n13435) );
  NAND2_X1 U12427 ( .A1(n13435), .A2(n10180), .ZN(n9809) );
  INV_X1 U12428 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U12429 ( .A1(n10415), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U12430 ( .A1(n10207), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9804) );
  OAI211_X1 U12431 ( .C1(n13784), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9807)
         );
  INV_X1 U12432 ( .A(n9807), .ZN(n9808) );
  NAND2_X1 U12433 ( .A1(n9810), .A2(n13418), .ZN(n9814) );
  INV_X1 U12434 ( .A(n9810), .ZN(n9811) );
  NAND2_X1 U12435 ( .A1(n9811), .A2(n13108), .ZN(n9812) );
  NAND2_X1 U12436 ( .A1(n9814), .A2(n9812), .ZN(n12985) );
  INV_X1 U12437 ( .A(n12985), .ZN(n9813) );
  NAND2_X1 U12438 ( .A1(n11706), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9817) );
  INV_X1 U12439 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U12440 ( .A1(n11875), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9836) );
  INV_X1 U12441 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U12442 ( .A1(n9819), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U12443 ( .A1(n9836), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U12444 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  NAND2_X1 U12445 ( .A1(n9837), .A2(n9824), .ZN(n11701) );
  NAND2_X1 U12446 ( .A1(n11701), .A2(n10424), .ZN(n9826) );
  NAND2_X1 U12447 ( .A1(n6931), .A2(SI_22_), .ZN(n9825) );
  XNOR2_X1 U12448 ( .A(n13057), .B(n12895), .ZN(n9871) );
  NAND2_X1 U12449 ( .A1(n9827), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12450 ( .A1(n9845), .A2(n9828), .ZN(n13422) );
  NAND2_X1 U12451 ( .A1(n13422), .A2(n10180), .ZN(n9834) );
  INV_X1 U12452 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12453 ( .A1(n10416), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12454 ( .A1(n10415), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9829) );
  OAI211_X1 U12455 ( .C1(n9860), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9832)
         );
  INV_X1 U12456 ( .A(n9832), .ZN(n9833) );
  INV_X1 U12457 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12458 ( .A1(n9838), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9852) );
  INV_X1 U12459 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U12460 ( .A1(n9839), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9840) );
  AND2_X1 U12461 ( .A1(n9852), .A2(n9840), .ZN(n9841) );
  NAND2_X1 U12462 ( .A1(n6931), .A2(SI_23_), .ZN(n9842) );
  NAND2_X1 U12463 ( .A1(n9845), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12464 ( .A1(n9856), .A2(n9846), .ZN(n13406) );
  NAND2_X1 U12465 ( .A1(n13406), .A2(n10180), .ZN(n9851) );
  INV_X1 U12466 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U12467 ( .A1(n10191), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U12468 ( .A1(n10415), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9847) );
  OAI211_X1 U12469 ( .C1(n9860), .C2(n13407), .A(n9848), .B(n9847), .ZN(n9849)
         );
  INV_X1 U12470 ( .A(n9849), .ZN(n9850) );
  XNOR2_X1 U12471 ( .A(n10154), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U12472 ( .A1(n12158), .A2(n10424), .ZN(n9855) );
  NAND2_X1 U12473 ( .A1(n10423), .A2(SI_24_), .ZN(n9854) );
  XNOR2_X1 U12474 ( .A(n10238), .B(n12895), .ZN(n9864) );
  NAND2_X1 U12475 ( .A1(n9856), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U12476 ( .A1(n9857), .A2(n9923), .ZN(n9911) );
  NAND2_X1 U12477 ( .A1(n9911), .A2(n10180), .ZN(n9863) );
  INV_X1 U12478 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13393) );
  NAND2_X1 U12479 ( .A1(n10415), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12480 ( .A1(n10416), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9858) );
  OAI211_X1 U12481 ( .C1(n9860), .C2(n13393), .A(n9859), .B(n9858), .ZN(n9861)
         );
  INV_X1 U12482 ( .A(n9861), .ZN(n9862) );
  NAND2_X1 U12483 ( .A1(n9864), .A2(n13402), .ZN(n13003) );
  INV_X1 U12484 ( .A(n9864), .ZN(n9865) );
  NAND2_X1 U12485 ( .A1(n9865), .A2(n13105), .ZN(n9866) );
  INV_X1 U12486 ( .A(n9867), .ZN(n9868) );
  AND2_X1 U12487 ( .A1(n9871), .A2(n13401), .ZN(n9872) );
  AOI21_X1 U12488 ( .B1(n9874), .B2(n13419), .A(n9872), .ZN(n12884) );
  INV_X1 U12489 ( .A(n9873), .ZN(n9877) );
  INV_X1 U12490 ( .A(n9874), .ZN(n9875) );
  AND2_X1 U12491 ( .A1(n9875), .A2(n13106), .ZN(n9876) );
  AOI21_X1 U12492 ( .B1(n12883), .B2(n12884), .A(n12885), .ZN(n13007) );
  INV_X1 U12493 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U12494 ( .A1(n10800), .A2(n10739), .ZN(n9880) );
  NAND2_X1 U12495 ( .A1(n13834), .A2(n12237), .ZN(n9879) );
  INV_X1 U12496 ( .A(n11315), .ZN(n10737) );
  NOR2_X1 U12497 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n9884) );
  NOR4_X1 U12498 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9883) );
  NOR4_X1 U12499 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9882) );
  NOR4_X1 U12500 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9881) );
  NAND4_X1 U12501 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n9890)
         );
  NOR4_X1 U12502 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9888) );
  NOR4_X1 U12503 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9887) );
  NOR4_X1 U12504 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9886) );
  NOR4_X1 U12505 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9885) );
  NAND4_X1 U12506 ( .A1(n9888), .A2(n9887), .A3(n9886), .A4(n9885), .ZN(n9889)
         );
  OAI21_X1 U12507 ( .B1(n9890), .B2(n9889), .A(n10800), .ZN(n10251) );
  NAND3_X1 U12508 ( .A1(n10737), .A2(n13817), .A3(n10251), .ZN(n10261) );
  NAND2_X1 U12509 ( .A1(n9893), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9891) );
  MUX2_X1 U12510 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9891), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9892) );
  NAND2_X1 U12511 ( .A1(n11702), .A2(n11454), .ZN(n9895) );
  NAND2_X1 U12512 ( .A1(n10429), .A2(n9895), .ZN(n9896) );
  NAND2_X1 U12513 ( .A1(n9896), .A2(n11660), .ZN(n9898) );
  NAND2_X1 U12514 ( .A1(n11660), .A2(n11454), .ZN(n10248) );
  NAND2_X1 U12515 ( .A1(n10243), .A2(n10248), .ZN(n9897) );
  NAND2_X1 U12516 ( .A1(n9898), .A2(n9897), .ZN(n10258) );
  NAND2_X1 U12517 ( .A1(n10258), .A2(n15806), .ZN(n9901) );
  INV_X1 U12518 ( .A(n13817), .ZN(n9899) );
  NAND2_X1 U12519 ( .A1(n11315), .A2(n9899), .ZN(n10253) );
  INV_X1 U12520 ( .A(n10251), .ZN(n9900) );
  NAND2_X1 U12521 ( .A1(n10429), .A2(n11702), .ZN(n10241) );
  OR2_X1 U12522 ( .A1(n10241), .A2(n10464), .ZN(n10257) );
  OAI22_X1 U12523 ( .A1(n10261), .A2(n9901), .B1(n10260), .B2(n10257), .ZN(
        n9909) );
  INV_X1 U12524 ( .A(n9902), .ZN(n9903) );
  NAND2_X1 U12525 ( .A1(n9903), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9904) );
  MUX2_X1 U12526 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9904), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9906) );
  NOR2_X1 U12527 ( .A1(n12237), .A2(n9442), .ZN(n9907) );
  NAND2_X1 U12528 ( .A1(n9908), .A2(n9907), .ZN(n10599) );
  NAND2_X1 U12529 ( .A1(n13312), .A2(n11454), .ZN(n10242) );
  INV_X1 U12530 ( .A(n10242), .ZN(n10589) );
  NAND2_X1 U12531 ( .A1(n10589), .A2(n10263), .ZN(n10591) );
  INV_X1 U12532 ( .A(n13831), .ZN(n13305) );
  INV_X1 U12533 ( .A(n12915), .ZN(n10214) );
  NAND2_X1 U12534 ( .A1(n13305), .A2(n10214), .ZN(n10709) );
  NAND2_X1 U12535 ( .A1(n10709), .A2(n10622), .ZN(n9922) );
  INV_X1 U12536 ( .A(n9922), .ZN(n9910) );
  INV_X1 U12537 ( .A(n9911), .ZN(n13394) );
  NAND2_X1 U12538 ( .A1(n10261), .A2(n10258), .ZN(n9916) );
  INV_X1 U12539 ( .A(n10257), .ZN(n9912) );
  NAND2_X1 U12540 ( .A1(n10260), .A2(n9912), .ZN(n9915) );
  AND2_X1 U12541 ( .A1(n10242), .A2(n6417), .ZN(n10247) );
  NAND2_X1 U12542 ( .A1(n10599), .A2(n10621), .ZN(n9913) );
  NOR2_X1 U12543 ( .A1(n10247), .A2(n9913), .ZN(n9914) );
  NAND3_X1 U12544 ( .A1(n9916), .A2(n9915), .A3(n9914), .ZN(n9917) );
  NAND2_X1 U12545 ( .A1(n9917), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9921) );
  OR2_X1 U12546 ( .A1(n10242), .A2(n10564), .ZN(n11251) );
  INV_X1 U12547 ( .A(n10263), .ZN(n10620) );
  NOR2_X1 U12548 ( .A1(n11251), .A2(n10620), .ZN(n9919) );
  NAND2_X1 U12549 ( .A1(n10260), .A2(n9919), .ZN(n9920) );
  NAND2_X1 U12550 ( .A1(n10415), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U12551 ( .A1(n10207), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12552 ( .A1(n10191), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9925) );
  AOI21_X1 U12553 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n9923), .A(n10166), .ZN(
        n13377) );
  OR2_X1 U12554 ( .A1(n9561), .A2(n13377), .ZN(n9924) );
  INV_X1 U12555 ( .A(n13389), .ZN(n13104) );
  AOI22_X1 U12556 ( .A1(n13027), .A2(n13104), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9928) );
  OAI21_X1 U12557 ( .B1(n13394), .B2(n13088), .A(n9928), .ZN(n9929) );
  AOI21_X1 U12558 ( .B1(n13076), .B2(n13106), .A(n9929), .ZN(n9931) );
  INV_X1 U12559 ( .A(n10238), .ZN(n13774) );
  NAND2_X1 U12560 ( .A1(n10429), .A2(n11454), .ZN(n11438) );
  NAND2_X1 U12561 ( .A1(n10261), .A2(n11438), .ZN(n9930) );
  NAND2_X1 U12562 ( .A1(n12380), .A2(n10044), .ZN(n9933) );
  NOR2_X1 U12563 ( .A1(n14025), .A2(n15727), .ZN(n11577) );
  NAND2_X1 U12564 ( .A1(n11578), .A2(n6421), .ZN(n9935) );
  NAND2_X1 U12565 ( .A1(n14023), .A2(n11039), .ZN(n9934) );
  NAND2_X1 U12566 ( .A1(n11330), .A2(n15742), .ZN(n11588) );
  AND2_X1 U12567 ( .A1(n11588), .A2(n9936), .ZN(n12598) );
  XNOR2_X1 U12568 ( .A(n14021), .B(n12396), .ZN(n12596) );
  INV_X1 U12569 ( .A(n14021), .ZN(n10008) );
  NAND2_X1 U12570 ( .A1(n10008), .A2(n12396), .ZN(n9937) );
  NAND2_X1 U12571 ( .A1(n15759), .A2(n14020), .ZN(n11625) );
  NAND2_X1 U12572 ( .A1(n11631), .A2(n11625), .ZN(n9938) );
  INV_X1 U12573 ( .A(n14020), .ZN(n11329) );
  NAND2_X1 U12574 ( .A1(n11329), .A2(n12404), .ZN(n11624) );
  NAND2_X1 U12575 ( .A1(n9938), .A2(n11624), .ZN(n11475) );
  XNOR2_X1 U12576 ( .A(n12420), .B(n14019), .ZN(n12599) );
  INV_X1 U12577 ( .A(n14019), .ZN(n9939) );
  NAND2_X1 U12578 ( .A1(n9939), .A2(n12420), .ZN(n9940) );
  INV_X1 U12579 ( .A(n14018), .ZN(n11848) );
  OR2_X1 U12580 ( .A1(n11848), .A2(n12428), .ZN(n9941) );
  NAND2_X1 U12581 ( .A1(n12428), .A2(n11848), .ZN(n9942) );
  INV_X1 U12582 ( .A(n14017), .ZN(n9944) );
  OR2_X1 U12583 ( .A1(n14509), .A2(n9944), .ZN(n9943) );
  NAND2_X1 U12584 ( .A1(n14509), .A2(n9944), .ZN(n9945) );
  NAND2_X1 U12585 ( .A1(n9946), .A2(n9945), .ZN(n11755) );
  XNOR2_X1 U12586 ( .A(n14504), .B(n14013), .ZN(n12605) );
  OR2_X1 U12587 ( .A1(n12455), .A2(n11847), .ZN(n12022) );
  INV_X1 U12588 ( .A(n14014), .ZN(n12462) );
  NAND2_X1 U12589 ( .A1(n12022), .A2(n12462), .ZN(n9949) );
  NAND2_X1 U12590 ( .A1(n14014), .A2(n14015), .ZN(n9947) );
  NOR2_X1 U12591 ( .A1(n12455), .A2(n9947), .ZN(n9948) );
  AOI21_X1 U12592 ( .B1(n12120), .B2(n9949), .A(n9948), .ZN(n9950) );
  NAND2_X1 U12593 ( .A1(n11755), .A2(n11926), .ZN(n9955) );
  XNOR2_X1 U12594 ( .A(n14500), .B(n14012), .ZN(n12608) );
  INV_X1 U12595 ( .A(n14013), .ZN(n9951) );
  NAND2_X1 U12596 ( .A1(n14504), .A2(n9951), .ZN(n11928) );
  AND2_X1 U12597 ( .A1(n12608), .A2(n11928), .ZN(n9953) );
  AOI22_X1 U12598 ( .A1(n12460), .A2(n12462), .B1(n11847), .B2(n12455), .ZN(
        n11925) );
  INV_X1 U12599 ( .A(n14012), .ZN(n9956) );
  OR2_X1 U12600 ( .A1(n14500), .A2(n9956), .ZN(n9957) );
  INV_X1 U12601 ( .A(n14011), .ZN(n13845) );
  XNOR2_X1 U12602 ( .A(n14495), .B(n13845), .ZN(n12610) );
  INV_X1 U12603 ( .A(n12610), .ZN(n12150) );
  OR2_X1 U12604 ( .A1(n14495), .A2(n13845), .ZN(n9958) );
  INV_X1 U12605 ( .A(n14010), .ZN(n13994) );
  NAND2_X1 U12606 ( .A1(n14490), .A2(n13994), .ZN(n9959) );
  OR2_X1 U12607 ( .A1(n14490), .A2(n13994), .ZN(n9960) );
  INV_X1 U12608 ( .A(n14377), .ZN(n13902) );
  XNOR2_X1 U12609 ( .A(n13999), .B(n13902), .ZN(n12614) );
  OR2_X1 U12610 ( .A1(n13999), .A2(n13902), .ZN(n9961) );
  XNOR2_X1 U12611 ( .A(n14477), .B(n14359), .ZN(n14389) );
  INV_X1 U12612 ( .A(n14359), .ZN(n13990) );
  OR2_X1 U12613 ( .A1(n14477), .A2(n13990), .ZN(n9962) );
  INV_X1 U12614 ( .A(n14360), .ZN(n14314) );
  OR2_X1 U12615 ( .A1(n14364), .A2(n14330), .ZN(n12593) );
  OAI21_X1 U12616 ( .B1(n14466), .B2(n14314), .A(n12593), .ZN(n9965) );
  NAND2_X1 U12617 ( .A1(n14364), .A2(n14330), .ZN(n12592) );
  INV_X1 U12618 ( .A(n12592), .ZN(n14327) );
  NAND2_X1 U12619 ( .A1(n12592), .A2(n14360), .ZN(n9963) );
  AOI22_X1 U12620 ( .A1(n14314), .A2(n14327), .B1(n9963), .B2(n14466), .ZN(
        n9964) );
  INV_X1 U12621 ( .A(n14009), .ZN(n14332) );
  AND2_X1 U12622 ( .A1(n14321), .A2(n14332), .ZN(n9966) );
  OR2_X1 U12623 ( .A1(n14321), .A2(n14332), .ZN(n9967) );
  NAND2_X1 U12624 ( .A1(n14456), .A2(n14315), .ZN(n9969) );
  OR2_X1 U12625 ( .A1(n14456), .A2(n14315), .ZN(n9968) );
  NAND2_X1 U12626 ( .A1(n9969), .A2(n9968), .ZN(n14300) );
  OR2_X1 U12627 ( .A1(n14537), .A2(n14008), .ZN(n9970) );
  NAND2_X1 U12628 ( .A1(n9971), .A2(n9970), .ZN(n14261) );
  NAND2_X1 U12629 ( .A1(n14277), .A2(n14255), .ZN(n9972) );
  INV_X1 U12630 ( .A(n14227), .ZN(n13929) );
  NAND2_X1 U12631 ( .A1(n14440), .A2(n13929), .ZN(n9975) );
  OR2_X1 U12632 ( .A1(n14440), .A2(n13929), .ZN(n9976) );
  INV_X1 U12633 ( .A(n14256), .ZN(n14007) );
  INV_X1 U12634 ( .A(n14527), .ZN(n14217) );
  XNOR2_X1 U12635 ( .A(n14217), .B(n13980), .ZN(n12619) );
  OR2_X1 U12636 ( .A1(n14527), .A2(n14226), .ZN(n9977) );
  INV_X1 U12637 ( .A(n14006), .ZN(n12587) );
  OR2_X1 U12638 ( .A1(n14425), .A2(n12587), .ZN(n9978) );
  NAND2_X1 U12639 ( .A1(n14425), .A2(n12587), .ZN(n9979) );
  INV_X2 U12640 ( .A(n14190), .ZN(n14420) );
  NAND2_X1 U12641 ( .A1(n12934), .A2(n14005), .ZN(n10042) );
  OR2_X1 U12642 ( .A1(n12934), .A2(n14005), .ZN(n9980) );
  NAND2_X1 U12643 ( .A1(n10042), .A2(n9980), .ZN(n12620) );
  INV_X1 U12644 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12930) );
  INV_X1 U12645 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14561) );
  MUX2_X1 U12646 ( .A(n12930), .B(n14561), .S(n10071), .Z(n10070) );
  XNOR2_X1 U12647 ( .A(n10070), .B(SI_29_), .ZN(n10068) );
  NAND2_X1 U12648 ( .A1(n12928), .A2(n9302), .ZN(n9985) );
  NAND2_X1 U12649 ( .A1(n12550), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9984) );
  INV_X1 U12650 ( .A(n12621), .ZN(n9989) );
  INV_X1 U12651 ( .A(n14005), .ZN(n9997) );
  NOR2_X1 U12652 ( .A1(n12625), .A2(n12630), .ZN(n12536) );
  NOR2_X1 U12653 ( .A1(n8895), .A2(n12626), .ZN(n9986) );
  OR2_X2 U12654 ( .A1(n12536), .A2(n9986), .ZN(n14379) );
  NAND2_X1 U12655 ( .A1(n6474), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12656 ( .A1(n9375), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U12657 ( .A1(n9991), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9992) );
  AND3_X1 U12658 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(n12543) );
  OR2_X1 U12659 ( .A1(n12942), .A2(n9995), .ZN(n9996) );
  NAND2_X1 U12660 ( .A1(n14374), .A2(n9996), .ZN(n14172) );
  OAI22_X1 U12661 ( .A1(n9997), .A2(n14329), .B1(n12543), .B2(n14172), .ZN(
        n9998) );
  INV_X1 U12662 ( .A(n9998), .ZN(n9999) );
  AND2_X1 U12663 ( .A1(n15721), .A2(n10285), .ZN(n10000) );
  NAND2_X1 U12664 ( .A1(n10001), .A2(n10000), .ZN(n10046) );
  NOR2_X1 U12665 ( .A1(n14417), .A2(n14352), .ZN(n10054) );
  NAND2_X1 U12666 ( .A1(n12380), .A2(n11574), .ZN(n10002) );
  NAND2_X1 U12667 ( .A1(n11578), .A2(n11039), .ZN(n10004) );
  INV_X1 U12668 ( .A(n10004), .ZN(n11638) );
  INV_X1 U12669 ( .A(n12598), .ZN(n11641) );
  NAND2_X1 U12670 ( .A1(n12595), .A2(n10004), .ZN(n10005) );
  OAI211_X1 U12671 ( .C1(n11640), .C2(n11638), .A(n11641), .B(n10005), .ZN(
        n10007) );
  NAND2_X1 U12672 ( .A1(n11330), .A2(n10045), .ZN(n10006) );
  NAND2_X1 U12673 ( .A1(n10007), .A2(n10006), .ZN(n11586) );
  INV_X1 U12674 ( .A(n12596), .ZN(n11589) );
  NAND2_X1 U12675 ( .A1(n11586), .A2(n11589), .ZN(n10010) );
  NAND2_X1 U12676 ( .A1(n10008), .A2(n7888), .ZN(n10009) );
  NAND2_X1 U12677 ( .A1(n12404), .A2(n14020), .ZN(n10011) );
  XNOR2_X1 U12678 ( .A(n12428), .B(n14018), .ZN(n12600) );
  OR2_X1 U12679 ( .A1(n12428), .A2(n14018), .ZN(n10012) );
  XNOR2_X1 U12680 ( .A(n14509), .B(n14017), .ZN(n12601) );
  NAND2_X1 U12681 ( .A1(n14509), .A2(n14017), .ZN(n10014) );
  XNOR2_X1 U12682 ( .A(n12455), .B(n11847), .ZN(n12604) );
  XNOR2_X1 U12683 ( .A(n12460), .B(n14014), .ZN(n12606) );
  NAND2_X1 U12684 ( .A1(n12021), .A2(n10015), .ZN(n12020) );
  OR2_X1 U12685 ( .A1(n12460), .A2(n14014), .ZN(n10016) );
  NAND2_X1 U12686 ( .A1(n12020), .A2(n10016), .ZN(n12118) );
  NAND2_X1 U12687 ( .A1(n14504), .A2(n14013), .ZN(n10019) );
  OR2_X1 U12688 ( .A1(n14504), .A2(n14013), .ZN(n10017) );
  INV_X1 U12689 ( .A(n10017), .ZN(n10018) );
  NAND2_X1 U12690 ( .A1(n14495), .A2(n14011), .ZN(n10021) );
  OR2_X1 U12691 ( .A1(n14490), .A2(n14010), .ZN(n12240) );
  NAND2_X1 U12692 ( .A1(n14490), .A2(n14010), .ZN(n12239) );
  NAND2_X1 U12693 ( .A1(n14477), .A2(n14359), .ZN(n10023) );
  NAND2_X1 U12694 ( .A1(n14546), .A2(n14330), .ZN(n10024) );
  OR2_X1 U12695 ( .A1(n14546), .A2(n14330), .ZN(n10025) );
  XNOR2_X1 U12696 ( .A(n14466), .B(n14360), .ZN(n14336) );
  OR2_X1 U12697 ( .A1(n14466), .A2(n14360), .ZN(n10028) );
  NAND2_X1 U12698 ( .A1(n14321), .A2(n14009), .ZN(n12590) );
  OR2_X1 U12699 ( .A1(n14321), .A2(n14009), .ZN(n12591) );
  NAND2_X1 U12700 ( .A1(n10029), .A2(n8050), .ZN(n14242) );
  NAND2_X1 U12701 ( .A1(n14440), .A2(n14227), .ZN(n12588) );
  NAND2_X1 U12702 ( .A1(n14277), .A2(n14285), .ZN(n14245) );
  AND2_X1 U12703 ( .A1(n12588), .A2(n14245), .ZN(n10033) );
  INV_X1 U12704 ( .A(n14537), .ZN(n14290) );
  XNOR2_X1 U12705 ( .A(n14290), .B(n14008), .ZN(n14281) );
  NOR2_X1 U12706 ( .A1(n14308), .A2(n14315), .ZN(n14240) );
  AND2_X1 U12707 ( .A1(n14537), .A2(n14303), .ZN(n14243) );
  OR2_X1 U12708 ( .A1(n14266), .A2(n14243), .ZN(n10032) );
  OR2_X1 U12709 ( .A1(n14440), .A2(n14227), .ZN(n12589) );
  INV_X1 U12710 ( .A(n12589), .ZN(n10031) );
  AOI21_X1 U12711 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10034) );
  OR2_X1 U12712 ( .A1(n14233), .A2(n14256), .ZN(n10037) );
  NAND2_X1 U12713 ( .A1(n14527), .A2(n13980), .ZN(n10038) );
  OR2_X1 U12714 ( .A1(n14527), .A2(n13980), .ZN(n10039) );
  OR2_X1 U12715 ( .A1(n14425), .A2(n14006), .ZN(n10040) );
  INV_X1 U12716 ( .A(n10040), .ZN(n10041) );
  NAND2_X1 U12717 ( .A1(n10269), .A2(n10270), .ZN(n10273) );
  NAND2_X1 U12718 ( .A1(n12582), .A2(n14386), .ZN(n11569) );
  NAND2_X1 U12719 ( .A1(n14337), .A2(n11569), .ZN(n10043) );
  INV_X1 U12720 ( .A(n12420), .ZN(n11552) );
  INV_X1 U12721 ( .A(n12455), .ZN(n11896) );
  INV_X1 U12722 ( .A(n14495), .ZN(n12368) );
  INV_X1 U12723 ( .A(n14490), .ZN(n12248) );
  NOR2_X4 U12724 ( .A1(n14382), .A2(n14364), .ZN(n14363) );
  INV_X1 U12725 ( .A(n14466), .ZN(n14347) );
  AND2_X2 U12726 ( .A1(n14304), .A2(n14537), .ZN(n14288) );
  AOI211_X1 U12727 ( .C1(n14415), .C2(n8060), .A(n14380), .B(n14176), .ZN(
        n14414) );
  INV_X1 U12728 ( .A(n10046), .ZN(n10047) );
  AND2_X2 U12729 ( .A1(n10047), .A2(n12630), .ZN(n14399) );
  NAND2_X2 U12730 ( .A1(n14396), .A2(n10048), .ZN(n14368) );
  INV_X1 U12731 ( .A(n14385), .ZN(n14397) );
  AOI22_X1 U12732 ( .A1(n10049), .A2(n14397), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14352), .ZN(n10050) );
  OAI21_X1 U12733 ( .B1(n7894), .B2(n14368), .A(n10050), .ZN(n10051) );
  OAI21_X1 U12734 ( .B1(n14418), .B2(n14371), .A(n10052), .ZN(n10053) );
  NAND2_X1 U12735 ( .A1(n14420), .A2(n13998), .ZN(n10061) );
  AOI22_X1 U12736 ( .A1(n14005), .A2(n14374), .B1(n14376), .B2(n14006), .ZN(
        n14182) );
  AOI22_X1 U12737 ( .A1(n14188), .A2(n13873), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10058) );
  OAI21_X1 U12738 ( .B1(n14182), .B2(n13952), .A(n10058), .ZN(n10059) );
  INV_X1 U12739 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10111) );
  INV_X1 U12740 ( .A(n15569), .ZN(n12689) );
  NAND2_X1 U12741 ( .A1(n15516), .A2(n12689), .ZN(n15498) );
  INV_X1 U12742 ( .A(n15597), .ZN(n11940) );
  INV_X1 U12743 ( .A(n12706), .ZN(n11914) );
  INV_X1 U12744 ( .A(n12724), .ZN(n15225) );
  NAND2_X1 U12745 ( .A1(n15076), .A2(n15281), .ZN(n15057) );
  OR2_X2 U12746 ( .A1(n15057), .A2(n15200), .ZN(n15058) );
  INV_X1 U12747 ( .A(n15012), .ZN(n15182) );
  INV_X1 U12748 ( .A(n14940), .ZN(n14944) );
  INV_X1 U12749 ( .A(n10065), .ZN(n14876) );
  NAND2_X1 U12750 ( .A1(n12928), .A2(n10091), .ZN(n10067) );
  NAND2_X1 U12751 ( .A1(n6420), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10066) );
  AND2_X2 U12752 ( .A1(n14833), .A2(n15131), .ZN(n14838) );
  INV_X1 U12753 ( .A(SI_29_), .ZN(n13828) );
  NAND2_X1 U12754 ( .A1(n10070), .A2(n13828), .ZN(n10078) );
  NAND2_X1 U12755 ( .A1(n10088), .A2(n10078), .ZN(n10075) );
  MUX2_X1 U12756 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10071), .Z(n10072) );
  NAND2_X1 U12757 ( .A1(n10072), .A2(SI_30_), .ZN(n10083) );
  INV_X1 U12758 ( .A(n10072), .ZN(n10073) );
  INV_X1 U12759 ( .A(SI_30_), .ZN(n12370) );
  NAND2_X1 U12760 ( .A1(n10073), .A2(n12370), .ZN(n10079) );
  AND2_X1 U12761 ( .A1(n10083), .A2(n10079), .ZN(n10074) );
  NAND2_X1 U12762 ( .A1(n12910), .A2(n10091), .ZN(n10077) );
  NAND2_X1 U12763 ( .A1(n6420), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U12764 ( .A1(n14838), .A2(n15249), .ZN(n10094) );
  NAND2_X1 U12765 ( .A1(n10079), .A2(n10078), .ZN(n10086) );
  MUX2_X1 U12766 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10768), .Z(n10081) );
  INV_X1 U12767 ( .A(SI_31_), .ZN(n10080) );
  XNOR2_X1 U12768 ( .A(n10081), .B(n10080), .ZN(n10085) );
  INV_X1 U12769 ( .A(n10085), .ZN(n10082) );
  INV_X1 U12770 ( .A(n10088), .ZN(n10084) );
  NOR2_X1 U12771 ( .A1(n10086), .A2(n10085), .ZN(n10087) );
  NAND2_X1 U12772 ( .A1(n10088), .A2(n10087), .ZN(n10089) );
  NAND2_X1 U12773 ( .A1(n14557), .A2(n10091), .ZN(n10093) );
  NAND2_X1 U12774 ( .A1(n6422), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10092) );
  XNOR2_X1 U12775 ( .A(n10094), .B(n12862), .ZN(n10095) );
  NOR2_X1 U12776 ( .A1(n12660), .A2(n10111), .ZN(n10100) );
  INV_X1 U12777 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U12778 ( .A1(n8296), .A2(n10096), .ZN(n10099) );
  INV_X1 U12779 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U12780 ( .A1(n10097), .A2(n10117), .ZN(n10098) );
  INV_X1 U12781 ( .A(P1_B_REG_SCAN_IN), .ZN(n10102) );
  NOR2_X1 U12782 ( .A1(n10101), .A2(n10102), .ZN(n10103) );
  NOR2_X1 U12783 ( .A1(n14706), .A2(n10103), .ZN(n14840) );
  AND2_X1 U12784 ( .A1(n14719), .A2(n14840), .ZN(n14822) );
  NOR2_X1 U12785 ( .A1(n14821), .A2(n14822), .ZN(n10116) );
  INV_X1 U12786 ( .A(n12878), .ZN(n10110) );
  AND2_X1 U12787 ( .A1(n10754), .A2(n10104), .ZN(n10105) );
  NOR2_X1 U12788 ( .A1(n10106), .A2(n10105), .ZN(n10109) );
  NAND2_X1 U12789 ( .A1(n10754), .A2(n10759), .ZN(n10107) );
  NAND2_X1 U12790 ( .A1(n10107), .A2(n10757), .ZN(n10108) );
  MUX2_X1 U12791 ( .A(n10111), .B(n10116), .S(n15618), .Z(n10113) );
  NAND2_X1 U12792 ( .A1(n15618), .A2(n15598), .ZN(n15228) );
  NAND2_X1 U12793 ( .A1(n12862), .A2(n10399), .ZN(n10112) );
  NAND2_X1 U12794 ( .A1(n10113), .A2(n10112), .ZN(P1_U3559) );
  MUX2_X1 U12795 ( .A(n10117), .B(n10116), .S(n15606), .Z(n10120) );
  NAND2_X1 U12796 ( .A1(n15606), .A2(n15598), .ZN(n15288) );
  NAND2_X1 U12797 ( .A1(n12862), .A2(n10118), .ZN(n10119) );
  NAND2_X1 U12798 ( .A1(n10120), .A2(n10119), .ZN(P1_U3527) );
  NAND2_X1 U12799 ( .A1(n10442), .A2(n15800), .ZN(n10123) );
  OR2_X1 U12800 ( .A1(n13127), .A2(n10121), .ZN(n10122) );
  NOR2_X1 U12801 ( .A1(n15797), .A2(n10479), .ZN(n10124) );
  INV_X1 U12802 ( .A(n11509), .ZN(n10125) );
  NAND2_X1 U12803 ( .A1(n11365), .A2(n10125), .ZN(n10483) );
  AND2_X1 U12804 ( .A1(n11448), .A2(n13126), .ZN(n11397) );
  NAND2_X1 U12805 ( .A1(n11365), .A2(n11509), .ZN(n11400) );
  NAND2_X1 U12806 ( .A1(n13125), .A2(n11547), .ZN(n10488) );
  OR2_X1 U12807 ( .A1(n13125), .A2(n11519), .ZN(n10128) );
  NAND2_X1 U12808 ( .A1(n11749), .A2(n11607), .ZN(n10496) );
  INV_X1 U12809 ( .A(n11607), .ZN(n11672) );
  NAND2_X1 U12810 ( .A1(n13123), .A2(n11672), .ZN(n10494) );
  OR2_X1 U12811 ( .A1(n13124), .A2(n10130), .ZN(n10227) );
  NAND2_X1 U12812 ( .A1(n13124), .A2(n10130), .ZN(n10493) );
  INV_X1 U12813 ( .A(n10130), .ZN(n15837) );
  AND2_X1 U12814 ( .A1(n13124), .A2(n15837), .ZN(n11601) );
  AOI22_X1 U12815 ( .A1(n11602), .A2(n11601), .B1(n11607), .B2(n13123), .ZN(
        n10131) );
  OR2_X1 U12816 ( .A1(n13122), .A2(n11775), .ZN(n10133) );
  NAND2_X1 U12817 ( .A1(n11775), .A2(n13122), .ZN(n10134) );
  NAND2_X1 U12818 ( .A1(n10135), .A2(n10134), .ZN(n11882) );
  OR2_X1 U12819 ( .A1(n12143), .A2(n13120), .ZN(n10508) );
  NAND2_X1 U12820 ( .A1(n12143), .A2(n13120), .ZN(n10520) );
  NAND2_X1 U12821 ( .A1(n10508), .A2(n10520), .ZN(n11974) );
  INV_X1 U12822 ( .A(n12143), .ZN(n12137) );
  AND2_X1 U12823 ( .A1(n12137), .A2(n13120), .ZN(n12083) );
  AOI21_X1 U12824 ( .B1(n13753), .B2(n13119), .A(n12083), .ZN(n10137) );
  NAND2_X1 U12825 ( .A1(n12107), .A2(n13121), .ZN(n10507) );
  INV_X1 U12826 ( .A(n13753), .ZN(n10234) );
  NAND2_X1 U12827 ( .A1(n10234), .A2(n13060), .ZN(n10138) );
  NAND2_X1 U12828 ( .A1(n12201), .A2(n13118), .ZN(n10140) );
  NAND2_X1 U12829 ( .A1(n13814), .A2(n13117), .ZN(n10512) );
  NAND2_X1 U12830 ( .A1(n10516), .A2(n10512), .ZN(n12205) );
  OR2_X1 U12831 ( .A1(n13814), .A2(n13521), .ZN(n10141) );
  OR2_X1 U12832 ( .A1(n13523), .A2(n13045), .ZN(n10529) );
  NAND2_X1 U12833 ( .A1(n13523), .A2(n13045), .ZN(n10530) );
  NAND2_X1 U12834 ( .A1(n10529), .A2(n10530), .ZN(n13519) );
  NAND2_X1 U12835 ( .A1(n13523), .A2(n13116), .ZN(n10142) );
  AND2_X1 U12836 ( .A1(n13510), .A2(n13115), .ZN(n10144) );
  NAND2_X1 U12837 ( .A1(n13497), .A2(n13113), .ZN(n10145) );
  OR2_X1 U12838 ( .A1(n13484), .A2(n13469), .ZN(n10544) );
  NAND2_X1 U12839 ( .A1(n13484), .A2(n13469), .ZN(n10541) );
  NAND2_X1 U12840 ( .A1(n10544), .A2(n10541), .ZN(n13477) );
  NAND2_X1 U12841 ( .A1(n13587), .A2(n13480), .ZN(n10542) );
  OR2_X1 U12842 ( .A1(n13587), .A2(n13111), .ZN(n10146) );
  AND2_X1 U12843 ( .A1(n13794), .A2(n13470), .ZN(n10450) );
  OR2_X1 U12844 ( .A1(n13794), .A2(n13470), .ZN(n10449) );
  XNOR2_X1 U12845 ( .A(n13037), .B(n13457), .ZN(n13442) );
  NAND2_X1 U12846 ( .A1(n12988), .A2(n13418), .ZN(n10557) );
  NAND2_X1 U12847 ( .A1(n10558), .A2(n10557), .ZN(n13430) );
  NAND2_X1 U12848 ( .A1(n13037), .A2(n13109), .ZN(n13428) );
  AND2_X1 U12849 ( .A1(n13430), .A2(n13428), .ZN(n10147) );
  NAND2_X1 U12850 ( .A1(n13441), .A2(n10147), .ZN(n13429) );
  OR2_X1 U12851 ( .A1(n12988), .A2(n13108), .ZN(n10148) );
  NAND2_X1 U12852 ( .A1(n13429), .A2(n10148), .ZN(n13416) );
  NOR2_X1 U12853 ( .A1(n13057), .A2(n13107), .ZN(n10149) );
  INV_X1 U12854 ( .A(n13057), .ZN(n13782) );
  NAND2_X1 U12855 ( .A1(n13411), .A2(n13419), .ZN(n10150) );
  NAND2_X1 U12856 ( .A1(n13411), .A2(n13106), .ZN(n10151) );
  AND2_X1 U12857 ( .A1(n10238), .A2(n13105), .ZN(n10152) );
  OR2_X1 U12858 ( .A1(n10238), .A2(n13105), .ZN(n10153) );
  INV_X1 U12859 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12230) );
  INV_X1 U12860 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12231) );
  XNOR2_X1 U12861 ( .A(n12283), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n10157) );
  XNOR2_X1 U12862 ( .A(n10161), .B(n10157), .ZN(n12234) );
  NAND2_X1 U12863 ( .A1(n12234), .A2(n10424), .ZN(n10159) );
  NAND2_X1 U12864 ( .A1(n6931), .A2(SI_25_), .ZN(n10158) );
  NAND2_X1 U12865 ( .A1(n10160), .A2(n13389), .ZN(n10571) );
  NAND2_X1 U12866 ( .A1(n12285), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10162) );
  XNOR2_X1 U12867 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n10163) );
  NAND2_X1 U12868 ( .A1(n10423), .A2(SI_26_), .ZN(n10164) );
  NAND2_X1 U12869 ( .A1(n10207), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U12870 ( .A1(n10415), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10168) );
  OR2_X1 U12871 ( .A1(n13553), .A2(n13350), .ZN(n10170) );
  AND2_X1 U12872 ( .A1(n14570), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12873 ( .A1(n15306), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10172) );
  INV_X1 U12874 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15302) );
  XNOR2_X1 U12875 ( .A(n15302), .B(P1_DATAO_REG_27__SCAN_IN), .ZN(n10174) );
  XNOR2_X1 U12876 ( .A(n10186), .B(n10174), .ZN(n13829) );
  NAND2_X1 U12877 ( .A1(n10423), .A2(SI_27_), .ZN(n10175) );
  NAND2_X1 U12878 ( .A1(n10415), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U12879 ( .A1(n10207), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10183) );
  INV_X1 U12880 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U12881 ( .A1(n10176), .A2(n10177), .ZN(n10193) );
  INV_X1 U12882 ( .A(n10177), .ZN(n10178) );
  NAND2_X1 U12883 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n10178), .ZN(n10179) );
  NAND2_X1 U12884 ( .A1(n10193), .A2(n10179), .ZN(n13359) );
  NAND2_X1 U12885 ( .A1(n10180), .A2(n13359), .ZN(n10182) );
  NAND2_X1 U12886 ( .A1(n10416), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10181) );
  AND2_X1 U12887 ( .A1(n15302), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10185) );
  INV_X1 U12888 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13654) );
  NAND2_X1 U12889 ( .A1(n13654), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n10187) );
  XNOR2_X1 U12890 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n10188) );
  XNOR2_X1 U12891 ( .A(n10204), .B(n10188), .ZN(n12914) );
  NAND2_X1 U12892 ( .A1(n12914), .A2(n10424), .ZN(n10190) );
  NAND2_X1 U12893 ( .A1(n6931), .A2(SI_28_), .ZN(n10189) );
  NAND2_X1 U12894 ( .A1(n10207), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U12895 ( .A1(n10191), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U12896 ( .A1(n10415), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10196) );
  INV_X1 U12897 ( .A(n10193), .ZN(n10192) );
  INV_X1 U12898 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13665) );
  NAND2_X1 U12899 ( .A1(n10193), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12900 ( .A1(n13340), .A2(n10200), .ZN(n10239) );
  OR2_X1 U12901 ( .A1(n13549), .A2(n13334), .ZN(n13330) );
  AND2_X1 U12902 ( .A1(n13332), .A2(n13330), .ZN(n10199) );
  NAND2_X1 U12903 ( .A1(n13340), .A2(n13349), .ZN(n10201) );
  NAND2_X1 U12904 ( .A1(n13331), .A2(n10201), .ZN(n10211) );
  AND2_X1 U12905 ( .A1(n10202), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10203) );
  XNOR2_X1 U12906 ( .A(n12930), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n10406) );
  XNOR2_X1 U12907 ( .A(n10408), .B(n10406), .ZN(n13825) );
  NAND2_X1 U12908 ( .A1(n13825), .A2(n10424), .ZN(n10206) );
  NAND2_X1 U12909 ( .A1(n10423), .A2(SI_29_), .ZN(n10205) );
  NAND2_X1 U12910 ( .A1(n10207), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U12911 ( .A1(n10191), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U12912 ( .A1(n10415), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U12913 ( .A1(n10420), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n13103) );
  XNOR2_X1 U12914 ( .A(n12920), .B(n13103), .ZN(n10460) );
  XNOR2_X1 U12915 ( .A(n10211), .B(n10460), .ZN(n10221) );
  NAND2_X1 U12916 ( .A1(n10213), .A2(n10212), .ZN(n10433) );
  AND2_X1 U12917 ( .A1(n10214), .A2(P3_B_REG_SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12918 ( .A1(n15783), .A2(n10215), .ZN(n13321) );
  NAND2_X1 U12919 ( .A1(n10415), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12920 ( .A1(n10207), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U12921 ( .A1(n10191), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U12922 ( .A1(n10420), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n13102) );
  AOI22_X1 U12923 ( .A1(n13321), .A2(n13102), .B1(n13349), .B2(n15799), .ZN(
        n10219) );
  INV_X1 U12924 ( .A(n10481), .ZN(n10222) );
  NOR2_X1 U12925 ( .A1(n11503), .A2(n10222), .ZN(n10226) );
  NAND2_X1 U12926 ( .A1(n10223), .A2(n10472), .ZN(n15782) );
  OR2_X1 U12927 ( .A1(n15797), .A2(n15790), .ZN(n11436) );
  NAND2_X1 U12928 ( .A1(n11435), .A2(n10476), .ZN(n10225) );
  NAND2_X1 U12929 ( .A1(n11611), .A2(n10227), .ZN(n10490) );
  INV_X1 U12930 ( .A(n10490), .ZN(n10228) );
  NAND2_X1 U12931 ( .A1(n12042), .A2(n11775), .ZN(n10499) );
  INV_X1 U12932 ( .A(n11775), .ZN(n11748) );
  NAND2_X1 U12933 ( .A1(n11748), .A2(n13122), .ZN(n11879) );
  NAND2_X1 U12934 ( .A1(n10499), .A2(n11879), .ZN(n11877) );
  AND2_X1 U12935 ( .A1(n11879), .A2(n10507), .ZN(n10230) );
  OR2_X1 U12936 ( .A1(n10234), .A2(n13119), .ZN(n10510) );
  NAND2_X1 U12937 ( .A1(n10234), .A2(n13119), .ZN(n10525) );
  NAND2_X1 U12938 ( .A1(n10510), .A2(n10525), .ZN(n12091) );
  INV_X1 U12939 ( .A(n12205), .ZN(n12209) );
  INV_X1 U12940 ( .A(n13519), .ZN(n13517) );
  OR2_X1 U12941 ( .A1(n13510), .A2(n13522), .ZN(n10532) );
  NAND2_X1 U12942 ( .A1(n13510), .A2(n13522), .ZN(n10536) );
  OR2_X1 U12943 ( .A1(n13497), .A2(n13479), .ZN(n10533) );
  NAND2_X1 U12944 ( .A1(n13497), .A2(n13479), .ZN(n10535) );
  NAND2_X1 U12945 ( .A1(n13496), .A2(n13495), .ZN(n13494) );
  INV_X1 U12946 ( .A(n13477), .ZN(n13482) );
  INV_X1 U12947 ( .A(n10542), .ZN(n10545) );
  NAND2_X1 U12948 ( .A1(n13794), .A2(n13110), .ZN(n10549) );
  AND2_X1 U12949 ( .A1(n10549), .A2(n13452), .ZN(n10540) );
  OR2_X1 U12950 ( .A1(n13794), .A2(n13110), .ZN(n10550) );
  NAND2_X1 U12951 ( .A1(n10236), .A2(n10558), .ZN(n13420) );
  NAND2_X1 U12952 ( .A1(n13057), .A2(n13401), .ZN(n10467) );
  OR2_X1 U12953 ( .A1(n10238), .A2(n13402), .ZN(n10566) );
  NAND2_X1 U12954 ( .A1(n10238), .A2(n13402), .ZN(n10567) );
  NAND2_X1 U12955 ( .A1(n13553), .A2(n13010), .ZN(n10574) );
  NAND2_X1 U12956 ( .A1(n13549), .A2(n7457), .ZN(n13328) );
  AND2_X1 U12957 ( .A1(n10239), .A2(n13328), .ZN(n10576) );
  INV_X1 U12958 ( .A(n10460), .ZN(n10240) );
  NAND3_X1 U12959 ( .A1(n10258), .A2(n10589), .A3(n15806), .ZN(n10245) );
  NAND2_X1 U12960 ( .A1(n10242), .A2(n10241), .ZN(n10249) );
  OR2_X1 U12961 ( .A1(n10249), .A2(n10243), .ZN(n10244) );
  OR2_X1 U12962 ( .A1(n11438), .A2(n11702), .ZN(n15841) );
  NAND2_X1 U12963 ( .A1(n10249), .A2(n11660), .ZN(n10246) );
  NAND2_X1 U12964 ( .A1(n10246), .A2(n11702), .ZN(n11314) );
  OAI211_X1 U12965 ( .C1(n10249), .C2(n10248), .A(n11314), .B(n11315), .ZN(
        n10250) );
  OAI21_X1 U12966 ( .B1(n11311), .B2(n13817), .A(n10250), .ZN(n10254) );
  AND2_X1 U12967 ( .A1(n10251), .A2(n10263), .ZN(n10252) );
  INV_X1 U12968 ( .A(n15873), .ZN(n10255) );
  NAND2_X1 U12969 ( .A1(n12920), .A2(n13754), .ZN(n10256) );
  AND2_X1 U12970 ( .A1(n11251), .A2(n10257), .ZN(n10262) );
  INV_X1 U12971 ( .A(n10258), .ZN(n10259) );
  OAI22_X1 U12972 ( .A1(n10262), .A2(n10261), .B1(n10260), .B2(n10259), .ZN(
        n10264) );
  OR2_X1 U12973 ( .A1(n15860), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12974 ( .A1(n10266), .A2(n10265), .ZN(n10268) );
  NAND2_X1 U12975 ( .A1(n12920), .A2(n13759), .ZN(n10267) );
  NAND2_X1 U12976 ( .A1(n10268), .A2(n10267), .ZN(P3_U3456) );
  INV_X1 U12977 ( .A(n10269), .ZN(n10271) );
  NAND2_X1 U12978 ( .A1(n10271), .A2(n12620), .ZN(n10272) );
  INV_X1 U12979 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12980 ( .A1(n10274), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n10277) );
  INV_X1 U12981 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U12982 ( .A1(n10275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10276) );
  AND2_X1 U12983 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U12984 ( .A1(n10282), .A2(n8060), .ZN(n12936) );
  AND2_X1 U12985 ( .A1(n10284), .A2(n15722), .ZN(n15723) );
  AND3_X1 U12986 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n10288) );
  NAND2_X1 U12987 ( .A1(n15775), .A2(n10290), .ZN(n10291) );
  NAND2_X1 U12988 ( .A1(n10292), .A2(n10291), .ZN(n10294) );
  NAND2_X1 U12989 ( .A1(n10294), .A2(n10293), .ZN(P2_U3527) );
  INV_X1 U12990 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12991 ( .A1(n15765), .A2(n10296), .ZN(n10297) );
  NAND2_X1 U12992 ( .A1(n10298), .A2(n10297), .ZN(n10300) );
  AND2_X1 U12993 ( .A1(n15767), .A2(n15750), .ZN(n12114) );
  NAND2_X1 U12994 ( .A1(n10300), .A2(n10299), .ZN(P2_U3495) );
  INV_X1 U12995 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U12996 ( .A1(n10302), .A2(n15549), .ZN(n12677) );
  NAND2_X1 U12997 ( .A1(n11821), .A2(n12667), .ZN(n15504) );
  XNOR2_X2 U12998 ( .A(n14745), .B(n15564), .ZN(n15507) );
  NAND2_X1 U12999 ( .A1(n15504), .A2(n15507), .ZN(n11960) );
  INV_X1 U13000 ( .A(n15564), .ZN(n12685) );
  NOR2_X1 U13001 ( .A1(n14745), .A2(n12685), .ZN(n12684) );
  INV_X1 U13002 ( .A(n12684), .ZN(n11961) );
  XNOR2_X2 U13003 ( .A(n14744), .B(n15569), .ZN(n12828) );
  OR2_X1 U13004 ( .A1(n14744), .A2(n12689), .ZN(n10305) );
  INV_X1 U13005 ( .A(n15495), .ZN(n15580) );
  INV_X1 U13006 ( .A(n12699), .ZN(n14742) );
  XNOR2_X2 U13007 ( .A(n14742), .B(n12700), .ZN(n12833) );
  NAND2_X1 U13008 ( .A1(n12699), .A2(n12700), .ZN(n10307) );
  NAND2_X1 U13009 ( .A1(n10308), .A2(n10307), .ZN(n11947) );
  XNOR2_X1 U13010 ( .A(n15597), .B(n14741), .ZN(n12834) );
  INV_X1 U13011 ( .A(n14741), .ZN(n10309) );
  NAND2_X1 U13012 ( .A1(n10309), .A2(n15597), .ZN(n10310) );
  XNOR2_X1 U13013 ( .A(n12706), .B(n14740), .ZN(n12835) );
  INV_X1 U13014 ( .A(n14740), .ZN(n10311) );
  OR2_X1 U13015 ( .A1(n12706), .A2(n10311), .ZN(n10312) );
  INV_X1 U13016 ( .A(n14739), .ZN(n10313) );
  INV_X1 U13017 ( .A(n14738), .ZN(n10314) );
  NAND2_X1 U13018 ( .A1(n15234), .A2(n10314), .ZN(n10315) );
  INV_X1 U13019 ( .A(n14737), .ZN(n10316) );
  OR2_X1 U13020 ( .A1(n15291), .A2(n10316), .ZN(n10317) );
  INV_X1 U13021 ( .A(n14736), .ZN(n10318) );
  NAND2_X1 U13022 ( .A1(n12724), .A2(n10318), .ZN(n10319) );
  NAND2_X1 U13023 ( .A1(n12738), .A2(n14584), .ZN(n10321) );
  NAND2_X1 U13024 ( .A1(n10322), .A2(n10321), .ZN(n12844) );
  INV_X1 U13025 ( .A(n12844), .ZN(n12345) );
  NAND2_X1 U13026 ( .A1(n15212), .A2(n10323), .ZN(n12735) );
  NAND2_X1 U13027 ( .A1(n15089), .A2(n12733), .ZN(n15002) );
  NAND2_X1 U13028 ( .A1(n14715), .A2(n14586), .ZN(n12747) );
  AND2_X1 U13029 ( .A1(n15064), .A2(n14731), .ZN(n10326) );
  OR2_X1 U13030 ( .A1(n15045), .A2(n14730), .ZN(n12762) );
  NAND2_X1 U13031 ( .A1(n15045), .A2(n14730), .ZN(n10379) );
  NAND2_X1 U13032 ( .A1(n12762), .A2(n10379), .ZN(n15041) );
  OR2_X1 U13033 ( .A1(n15064), .A2(n14731), .ZN(n15039) );
  OAI211_X1 U13034 ( .C1(n12747), .C2(n10326), .A(n15041), .B(n15039), .ZN(
        n15022) );
  INV_X1 U13035 ( .A(n14730), .ZN(n14676) );
  OR2_X1 U13036 ( .A1(n15045), .A2(n14676), .ZN(n15020) );
  NAND2_X1 U13037 ( .A1(n15022), .A2(n15020), .ZN(n10324) );
  OR2_X1 U13038 ( .A1(n15188), .A2(n14729), .ZN(n10382) );
  NAND2_X1 U13039 ( .A1(n15188), .A2(n14729), .ZN(n10381) );
  NAND2_X1 U13040 ( .A1(n10382), .A2(n10381), .ZN(n15033) );
  NAND2_X1 U13041 ( .A1(n15002), .A2(n10325), .ZN(n10330) );
  INV_X1 U13042 ( .A(n10326), .ZN(n10327) );
  NAND2_X1 U13043 ( .A1(n10372), .A2(n10327), .ZN(n15019) );
  INV_X1 U13044 ( .A(n15020), .ZN(n10328) );
  NOR2_X1 U13045 ( .A1(n15019), .A2(n10328), .ZN(n15004) );
  XNOR2_X1 U13046 ( .A(n15012), .B(n14677), .ZN(n15006) );
  OR2_X1 U13047 ( .A1(n15188), .A2(n14599), .ZN(n15005) );
  NAND2_X1 U13048 ( .A1(n15012), .A2(n14677), .ZN(n10331) );
  NAND2_X1 U13049 ( .A1(n14994), .A2(n14611), .ZN(n10332) );
  NAND2_X1 U13050 ( .A1(n14968), .A2(n10332), .ZN(n14987) );
  XNOR2_X1 U13051 ( .A(n14974), .B(n14726), .ZN(n14967) );
  INV_X1 U13052 ( .A(n14726), .ZN(n14665) );
  OR2_X1 U13053 ( .A1(n14974), .A2(n14665), .ZN(n10334) );
  XNOR2_X1 U13054 ( .A(n15263), .B(n14612), .ZN(n12849) );
  INV_X1 U13055 ( .A(n15263), .ZN(n14957) );
  NAND2_X1 U13056 ( .A1(n14957), .A2(n14612), .ZN(n10335) );
  XNOR2_X1 U13057 ( .A(n14940), .B(n14666), .ZN(n14934) );
  INV_X1 U13058 ( .A(n14934), .ZN(n14928) );
  NAND2_X1 U13059 ( .A1(n14940), .A2(n14666), .ZN(n10336) );
  INV_X1 U13060 ( .A(n14724), .ZN(n10338) );
  OR2_X1 U13061 ( .A1(n14921), .A2(n10338), .ZN(n10339) );
  NAND2_X1 U13062 ( .A1(n14903), .A2(n7125), .ZN(n10340) );
  INV_X1 U13063 ( .A(n14722), .ZN(n10341) );
  AND2_X1 U13064 ( .A1(n14890), .A2(n10341), .ZN(n10343) );
  OR2_X1 U13065 ( .A1(n14890), .A2(n10341), .ZN(n10342) );
  NOR2_X1 U13066 ( .A1(n6419), .A2(n14721), .ZN(n10345) );
  NAND2_X1 U13067 ( .A1(n12804), .A2(n14851), .ZN(n14831) );
  OR2_X1 U13068 ( .A1(n12804), .A2(n14851), .ZN(n10344) );
  NAND2_X1 U13069 ( .A1(n12652), .A2(n12651), .ZN(n10347) );
  INV_X1 U13070 ( .A(n15526), .ZN(n12821) );
  NAND2_X1 U13071 ( .A1(n8801), .A2(n12821), .ZN(n10346) );
  INV_X1 U13072 ( .A(n15525), .ZN(n12672) );
  NAND2_X1 U13073 ( .A1(n15105), .A2(n12672), .ZN(n15104) );
  NAND2_X1 U13074 ( .A1(n10301), .A2(n15104), .ZN(n10349) );
  NAND2_X1 U13075 ( .A1(n10349), .A2(n15117), .ZN(n10351) );
  OR2_X1 U13076 ( .A1(n15104), .A2(n10301), .ZN(n10350) );
  INV_X1 U13077 ( .A(n15507), .ZN(n12831) );
  OR2_X1 U13078 ( .A1(n14745), .A2(n15564), .ZN(n10352) );
  NAND2_X1 U13079 ( .A1(n11968), .A2(n7177), .ZN(n15487) );
  OR2_X1 U13080 ( .A1(n14744), .A2(n15569), .ZN(n15486) );
  OR2_X1 U13081 ( .A1(n14743), .A2(n15495), .ZN(n10353) );
  AND2_X1 U13082 ( .A1(n15486), .A2(n10353), .ZN(n10355) );
  INV_X1 U13083 ( .A(n10353), .ZN(n10354) );
  INV_X1 U13084 ( .A(n15488), .ZN(n12830) );
  INV_X1 U13085 ( .A(n12833), .ZN(n10356) );
  NAND2_X1 U13086 ( .A1(n11950), .A2(n10356), .ZN(n10358) );
  NAND2_X1 U13087 ( .A1(n12699), .A2(n14688), .ZN(n10357) );
  NAND2_X1 U13088 ( .A1(n10358), .A2(n10357), .ZN(n11938) );
  INV_X1 U13089 ( .A(n12834), .ZN(n10359) );
  NAND2_X1 U13090 ( .A1(n11938), .A2(n10359), .ZN(n10361) );
  OR2_X1 U13091 ( .A1(n14741), .A2(n15597), .ZN(n10360) );
  OR2_X1 U13092 ( .A1(n12706), .A2(n14740), .ZN(n10362) );
  OR2_X1 U13093 ( .A1(n15234), .A2(n14738), .ZN(n12264) );
  OR2_X1 U13094 ( .A1(n15242), .A2(n14739), .ZN(n12177) );
  AND2_X1 U13095 ( .A1(n12264), .A2(n12177), .ZN(n10363) );
  INV_X1 U13096 ( .A(n12264), .ZN(n10364) );
  NOR2_X1 U13097 ( .A1(n12839), .A2(n10364), .ZN(n10365) );
  NOR2_X1 U13098 ( .A1(n12840), .A2(n10365), .ZN(n10366) );
  OR2_X1 U13099 ( .A1(n12724), .A2(n14736), .ZN(n12349) );
  NAND2_X1 U13100 ( .A1(n15286), .A2(n14584), .ZN(n10367) );
  AND2_X1 U13101 ( .A1(n12349), .A2(n10367), .ZN(n10371) );
  INV_X1 U13102 ( .A(n10367), .ZN(n10368) );
  OR2_X1 U13103 ( .A1(n10368), .A2(n12844), .ZN(n10369) );
  AND2_X1 U13104 ( .A1(n15212), .A2(n14734), .ZN(n15069) );
  INV_X1 U13105 ( .A(n15069), .ZN(n10374) );
  NAND2_X1 U13106 ( .A1(n15099), .A2(n10374), .ZN(n10375) );
  OAI22_X1 U13107 ( .A1(n15070), .A2(n10375), .B1(n14732), .B2(n14715), .ZN(
        n10376) );
  INV_X1 U13108 ( .A(n10376), .ZN(n10377) );
  OR2_X1 U13109 ( .A1(n15064), .A2(n14707), .ZN(n10378) );
  INV_X1 U13110 ( .A(n10379), .ZN(n10380) );
  NAND2_X1 U13111 ( .A1(n10383), .A2(n10382), .ZN(n15000) );
  OR2_X1 U13112 ( .A1(n15012), .A2(n14728), .ZN(n10384) );
  OR2_X1 U13113 ( .A1(n15271), .A2(n14611), .ZN(n10386) );
  INV_X1 U13114 ( .A(n14967), .ZN(n10387) );
  NAND2_X1 U13115 ( .A1(n14955), .A2(n14954), .ZN(n14953) );
  NAND2_X1 U13116 ( .A1(n15263), .A2(n14612), .ZN(n10388) );
  AND2_X1 U13117 ( .A1(n14934), .A2(n14917), .ZN(n10389) );
  OR2_X1 U13118 ( .A1(n14940), .A2(n14725), .ZN(n14910) );
  NAND2_X1 U13119 ( .A1(n14903), .A2(n14723), .ZN(n10390) );
  XNOR2_X1 U13120 ( .A(n14890), .B(n14722), .ZN(n14891) );
  INV_X1 U13121 ( .A(n14891), .ZN(n14883) );
  NAND2_X1 U13122 ( .A1(n14890), .A2(n14722), .ZN(n10391) );
  OR2_X1 U13123 ( .A1(n14880), .A2(n14721), .ZN(n10392) );
  NAND2_X1 U13124 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  AND2_X1 U13125 ( .A1(n12816), .A2(n12651), .ZN(n10396) );
  NOR2_X1 U13126 ( .A1(n10397), .A2(n10396), .ZN(n11833) );
  NAND2_X1 U13127 ( .A1(n11833), .A2(n11828), .ZN(n15589) );
  AOI211_X1 U13128 ( .C1(n12804), .C2(n14876), .A(n15517), .B(n14833), .ZN(
        n14857) );
  NAND2_X1 U13129 ( .A1(n12804), .A2(n10399), .ZN(n10400) );
  NAND2_X1 U13130 ( .A1(n10401), .A2(n10400), .ZN(P1_U3556) );
  NAND2_X1 U13131 ( .A1(n12804), .A2(n10118), .ZN(n10403) );
  INV_X1 U13132 ( .A(n13103), .ZN(n13336) );
  OR2_X1 U13133 ( .A1(n12920), .A2(n13336), .ZN(n10582) );
  INV_X1 U13134 ( .A(n10582), .ZN(n10404) );
  INV_X1 U13135 ( .A(n10406), .ZN(n10407) );
  NAND2_X1 U13136 ( .A1(n10408), .A2(n10407), .ZN(n10410) );
  NAND2_X1 U13137 ( .A1(n12930), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10409) );
  INV_X1 U13138 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12911) );
  XNOR2_X1 U13139 ( .A(n12911), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n10421) );
  INV_X1 U13140 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12944) );
  OAI22_X1 U13141 ( .A1(n10422), .A2(n10421), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12944), .ZN(n10412) );
  XNOR2_X1 U13142 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n10411) );
  XNOR2_X1 U13143 ( .A(n10412), .B(n10411), .ZN(n13818) );
  NAND2_X1 U13144 ( .A1(n13818), .A2(n10424), .ZN(n10414) );
  NAND2_X1 U13145 ( .A1(n6931), .A2(SI_31_), .ZN(n10413) );
  NAND2_X1 U13146 ( .A1(n10415), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13147 ( .A1(n10207), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U13148 ( .A1(n10416), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10417) );
  OR2_X1 U13149 ( .A1(n10458), .A2(n10457), .ZN(n10427) );
  XNOR2_X1 U13150 ( .A(n10422), .B(n10421), .ZN(n12369) );
  INV_X1 U13151 ( .A(n13102), .ZN(n10425) );
  NAND2_X1 U13152 ( .A1(n13760), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U13153 ( .A1(n12920), .A2(n13336), .ZN(n10580) );
  OAI211_X1 U13154 ( .C1(n13327), .C2(n13322), .A(n13312), .B(n10580), .ZN(
        n10428) );
  AOI211_X1 U13155 ( .C1(n13327), .C2(n10580), .A(n13312), .B(n10458), .ZN(
        n10434) );
  NAND2_X1 U13156 ( .A1(n13327), .A2(n13102), .ZN(n10583) );
  NAND3_X1 U13157 ( .A1(n10583), .A2(n10429), .A3(n13322), .ZN(n10436) );
  INV_X1 U13158 ( .A(n13312), .ZN(n10429) );
  INV_X1 U13159 ( .A(n10430), .ZN(n10431) );
  OAI21_X1 U13160 ( .B1(n10580), .B2(n10436), .A(n10431), .ZN(n10432) );
  INV_X1 U13161 ( .A(n10435), .ZN(n10439) );
  INV_X1 U13162 ( .A(n10436), .ZN(n10437) );
  AOI21_X1 U13163 ( .B1(n13758), .B2(n10429), .A(n10437), .ZN(n10438) );
  AOI21_X1 U13164 ( .B1(n10586), .B2(n10439), .A(n10438), .ZN(n10465) );
  INV_X1 U13165 ( .A(n10583), .ZN(n10456) );
  NAND2_X1 U13166 ( .A1(n10468), .A2(n10467), .ZN(n13421) );
  INV_X1 U13167 ( .A(n13421), .ZN(n13415) );
  INV_X1 U13168 ( .A(n10473), .ZN(n10441) );
  NAND2_X1 U13169 ( .A1(n11110), .A2(n10441), .ZN(n11254) );
  NOR2_X1 U13170 ( .A1(n11254), .A2(n11437), .ZN(n10444) );
  NOR3_X1 U13171 ( .A1(n10442), .A2(n11503), .A3(n11399), .ZN(n10443) );
  NAND4_X1 U13172 ( .A1(n11616), .A2(n15781), .A3(n10444), .A4(n10443), .ZN(
        n10445) );
  OR4_X1 U13173 ( .A1(n10445), .A2(n6895), .A3(n11877), .A4(n11602), .ZN(
        n10446) );
  NOR4_X1 U13174 ( .A1(n10446), .A2(n12091), .A3(n11974), .A4(n12001), .ZN(
        n10447) );
  NAND4_X1 U13175 ( .A1(n10447), .A2(n13508), .A3(n12209), .A4(n13495), .ZN(
        n10448) );
  NOR3_X1 U13176 ( .A1(n10448), .A2(n13477), .A3(n13519), .ZN(n10452) );
  INV_X1 U13177 ( .A(n10449), .ZN(n10451) );
  NAND4_X1 U13178 ( .A1(n13415), .A2(n13467), .A3(n10452), .A4(n13454), .ZN(
        n10453) );
  NOR4_X1 U13179 ( .A1(n10563), .A2(n10453), .A3(n13442), .A4(n13430), .ZN(
        n10454) );
  NAND4_X1 U13180 ( .A1(n13379), .A2(n6586), .A3(n13368), .A4(n10454), .ZN(
        n10455) );
  NOR4_X1 U13181 ( .A1(n10456), .A2(n13358), .A3(n13332), .A4(n10455), .ZN(
        n10461) );
  AND2_X1 U13182 ( .A1(n10458), .A2(n10457), .ZN(n10585) );
  INV_X1 U13183 ( .A(n10585), .ZN(n10459) );
  NAND4_X1 U13184 ( .A1(n10461), .A2(n10586), .A3(n10460), .A4(n10459), .ZN(
        n10462) );
  XNOR2_X1 U13185 ( .A(n10462), .B(n13312), .ZN(n10463) );
  OAI22_X1 U13186 ( .A1(n10466), .A2(n10465), .B1(n10464), .B2(n10463), .ZN(
        n10590) );
  INV_X1 U13187 ( .A(n13411), .ZN(n13778) );
  INV_X1 U13188 ( .A(n10467), .ZN(n10469) );
  MUX2_X1 U13189 ( .A(n10469), .B(n7509), .S(n6417), .Z(n10562) );
  INV_X1 U13190 ( .A(n10470), .ZN(n11498) );
  NAND2_X1 U13191 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  AOI21_X1 U13192 ( .B1(n10475), .B2(n10471), .A(n10224), .ZN(n10478) );
  OAI211_X1 U13193 ( .C1(n10473), .C2(n11660), .A(n11110), .B(n10472), .ZN(
        n10474) );
  NAND3_X1 U13194 ( .A1(n15781), .A2(n10475), .A3(n10474), .ZN(n10477) );
  OAI21_X1 U13195 ( .B1(n11441), .B2(n10479), .A(n10481), .ZN(n10480) );
  MUX2_X1 U13196 ( .A(n10483), .B(n10482), .S(n6417), .Z(n10484) );
  INV_X1 U13197 ( .A(n10486), .ZN(n10487) );
  OAI21_X1 U13198 ( .B1(n10488), .B2(n6417), .A(n10493), .ZN(n10489) );
  AOI211_X1 U13199 ( .C1(n6417), .C2(n10490), .A(n10489), .B(n11602), .ZN(
        n10491) );
  INV_X1 U13200 ( .A(n11877), .ZN(n11770) );
  INV_X1 U13201 ( .A(n10496), .ZN(n10492) );
  AOI211_X1 U13202 ( .C1(n10494), .C2(n10493), .A(n10564), .B(n10492), .ZN(
        n10498) );
  NAND4_X1 U13203 ( .A1(n10494), .A2(n11673), .A3(n15837), .A4(n10564), .ZN(
        n10495) );
  OAI21_X1 U13204 ( .B1(n10496), .B2(n6417), .A(n10495), .ZN(n10497) );
  OAI21_X1 U13205 ( .B1(n10498), .B2(n10497), .A(n11770), .ZN(n10503) );
  MUX2_X1 U13206 ( .A(n11879), .B(n10499), .S(n10564), .Z(n10500) );
  NAND3_X1 U13207 ( .A1(n10518), .A2(n7503), .A3(n10507), .ZN(n10509) );
  AND2_X1 U13208 ( .A1(n10509), .A2(n10508), .ZN(n10511) );
  OAI211_X1 U13209 ( .C1(n10511), .C2(n12091), .A(n10522), .B(n10510), .ZN(
        n10513) );
  NAND4_X1 U13210 ( .A1(n10513), .A2(n10512), .A3(n10524), .A4(n10564), .ZN(
        n10515) );
  NAND3_X1 U13211 ( .A1(n13814), .A2(n6417), .A3(n13117), .ZN(n10514) );
  OAI211_X1 U13212 ( .C1(n6417), .C2(n10516), .A(n10515), .B(n10514), .ZN(
        n10528) );
  NAND3_X1 U13213 ( .A1(n10518), .A2(n7503), .A3(n10517), .ZN(n10521) );
  INV_X1 U13214 ( .A(n12091), .ZN(n12086) );
  NAND3_X1 U13215 ( .A1(n12086), .A2(n6417), .A3(n10522), .ZN(n10519) );
  AOI211_X1 U13216 ( .C1(n10521), .C2(n10520), .A(n12205), .B(n10519), .ZN(
        n10527) );
  NAND2_X1 U13217 ( .A1(n10522), .A2(n6417), .ZN(n10523) );
  AOI211_X1 U13218 ( .C1(n10525), .C2(n10524), .A(n10523), .B(n12205), .ZN(
        n10526) );
  MUX2_X1 U13219 ( .A(n10530), .B(n10529), .S(n10564), .Z(n10531) );
  INV_X1 U13220 ( .A(n13508), .ZN(n13504) );
  AOI21_X1 U13221 ( .B1(n10533), .B2(n10532), .A(n6417), .ZN(n10534) );
  INV_X1 U13222 ( .A(n10535), .ZN(n10538) );
  INV_X1 U13223 ( .A(n10536), .ZN(n10537) );
  OAI21_X1 U13224 ( .B1(n10538), .B2(n10537), .A(n6417), .ZN(n10539) );
  AND2_X1 U13225 ( .A1(n10540), .A2(n6417), .ZN(n10543) );
  NAND3_X1 U13226 ( .A1(n10550), .A2(n10542), .A3(n10564), .ZN(n10547) );
  OAI21_X1 U13227 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(n10546) );
  AOI22_X1 U13228 ( .A1(n10548), .A2(n13467), .B1(n10547), .B2(n10546), .ZN(
        n10553) );
  INV_X1 U13229 ( .A(n10549), .ZN(n10551) );
  MUX2_X1 U13230 ( .A(n10551), .B(n7924), .S(n6417), .Z(n10552) );
  NOR2_X1 U13231 ( .A1(n13457), .A2(n10564), .ZN(n10555) );
  NOR2_X1 U13232 ( .A1(n13109), .A2(n6417), .ZN(n10554) );
  MUX2_X1 U13233 ( .A(n10555), .B(n10554), .S(n13037), .Z(n10556) );
  INV_X1 U13234 ( .A(n10557), .ZN(n10560) );
  INV_X1 U13235 ( .A(n10558), .ZN(n10559) );
  MUX2_X1 U13236 ( .A(n10560), .B(n10559), .S(n10564), .Z(n10561) );
  AOI21_X1 U13237 ( .B1(n10566), .B2(n10565), .A(n6417), .ZN(n10568) );
  MUX2_X1 U13238 ( .A(n6417), .B(n10568), .S(n10567), .Z(n10569) );
  INV_X1 U13239 ( .A(n13379), .ZN(n13375) );
  NAND2_X1 U13240 ( .A1(n13329), .A2(n6417), .ZN(n10581) );
  NOR2_X1 U13241 ( .A1(n10621), .A2(P3_U3151), .ZN(n10592) );
  NOR3_X1 U13242 ( .A1(n10591), .A2(n13305), .A3(n15785), .ZN(n10594) );
  INV_X1 U13243 ( .A(n10592), .ZN(n11783) );
  OAI21_X1 U13244 ( .B1(n11783), .B2(n11702), .A(P3_B_REG_SCAN_IN), .ZN(n10593) );
  OR2_X1 U13245 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  INV_X1 U13246 ( .A(n11050), .ZN(n12099) );
  INV_X1 U13247 ( .A(n10597), .ZN(n10598) );
  AND2_X2 U13248 ( .A1(n10598), .A2(n10761), .ZN(P1_U4016) );
  INV_X1 U13249 ( .A(n10599), .ZN(n10600) );
  INV_X1 U13250 ( .A(n10687), .ZN(n13158) );
  INV_X1 U13251 ( .A(n10683), .ZN(n13134) );
  XNOR2_X1 U13252 ( .A(n10999), .B(n9487), .ZN(n10991) );
  INV_X1 U13253 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13254 ( .A1(n10674), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13255 ( .A1(n10676), .A2(n10601), .ZN(n10602) );
  NAND2_X1 U13256 ( .A1(n6516), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13257 ( .A1(n10602), .A2(n10603), .ZN(n11000) );
  INV_X1 U13258 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15861) );
  OR2_X1 U13259 ( .A1(n11000), .A2(n15861), .ZN(n11001) );
  NAND2_X1 U13260 ( .A1(n10999), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10604) );
  XNOR2_X1 U13261 ( .A(n10788), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n11150) );
  AOI21_X1 U13262 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10788), .A(n11153), .ZN(
        n10605) );
  INV_X1 U13263 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15867) );
  XNOR2_X1 U13264 ( .A(n10683), .B(n15867), .ZN(n13141) );
  NAND2_X1 U13265 ( .A1(n11233), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n13156) );
  INV_X1 U13266 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15871) );
  XNOR2_X1 U13267 ( .A(n10687), .B(n15871), .ZN(n13155) );
  XNOR2_X1 U13268 ( .A(n11869), .B(P3_REG1_REG_10__SCAN_IN), .ZN(n11863) );
  AOI21_X1 U13269 ( .B1(n11864), .B2(n6489), .A(n11863), .ZN(n11866) );
  INV_X1 U13270 ( .A(n10658), .ZN(n13175) );
  NOR2_X1 U13271 ( .A1(n10608), .A2(n10658), .ZN(n13194) );
  INV_X1 U13272 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n13701) );
  XNOR2_X1 U13273 ( .A(n13190), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13192) );
  INV_X1 U13274 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12202) );
  INV_X1 U13275 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13748) );
  INV_X1 U13276 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13742) );
  OR2_X1 U13277 ( .A1(n13230), .A2(n13742), .ZN(n10665) );
  NAND2_X1 U13278 ( .A1(n13230), .A2(n13742), .ZN(n10612) );
  AND2_X1 U13279 ( .A1(n10665), .A2(n10612), .ZN(n13232) );
  NOR3_X1 U13280 ( .A1(n13235), .A2(n7247), .A3(n6997), .ZN(n10613) );
  INV_X1 U13281 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13734) );
  NOR2_X1 U13282 ( .A1(n10699), .A2(n13734), .ZN(n10615) );
  AOI21_X1 U13283 ( .B1(n10699), .B2(n13734), .A(n10615), .ZN(n13272) );
  INV_X1 U13284 ( .A(n10976), .ZN(n13287) );
  INV_X1 U13285 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13730) );
  INV_X1 U13286 ( .A(n13303), .ZN(n11119) );
  NAND2_X1 U13287 ( .A1(n11119), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13298) );
  INV_X1 U13288 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13289 ( .A1(n13303), .A2(n10616), .ZN(n10617) );
  NAND2_X1 U13290 ( .A1(n13298), .A2(n10617), .ZN(n10618) );
  NAND3_X1 U13291 ( .A1(n13276), .A2(n10619), .A3(n10618), .ZN(n10625) );
  NAND2_X1 U13292 ( .A1(n10620), .A2(n11783), .ZN(n10713) );
  NAND2_X1 U13293 ( .A1(n6417), .A2(n10621), .ZN(n10623) );
  NAND2_X1 U13294 ( .A1(n10623), .A2(n10622), .ZN(n10712) );
  INV_X1 U13295 ( .A(n10712), .ZN(n10624) );
  AOI21_X1 U13296 ( .B1(n6538), .B2(n10625), .A(n13293), .ZN(n10717) );
  MUX2_X1 U13297 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13831), .Z(n10672) );
  MUX2_X1 U13298 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13831), .Z(n10670) );
  MUX2_X1 U13299 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13831), .Z(n10669) );
  INV_X1 U13300 ( .A(n10699), .ZN(n13266) );
  INV_X1 U13301 ( .A(n10893), .ZN(n13215) );
  MUX2_X1 U13302 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13831), .Z(n10661) );
  INV_X1 U13303 ( .A(n10661), .ZN(n10662) );
  MUX2_X1 U13304 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13831), .Z(n10659) );
  INV_X1 U13305 ( .A(n10659), .ZN(n10660) );
  MUX2_X1 U13306 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13831), .Z(n10653) );
  INV_X1 U13307 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15815) );
  INV_X1 U13308 ( .A(n10676), .ZN(n11017) );
  NAND2_X1 U13309 ( .A1(n10627), .A2(n11017), .ZN(n10628) );
  INV_X1 U13310 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11320) );
  MUX2_X1 U13311 ( .A(n11320), .B(n9460), .S(n13831), .Z(n11276) );
  NAND2_X1 U13312 ( .A1(n11276), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11008) );
  INV_X1 U13313 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10673) );
  MUX2_X1 U13314 ( .A(n10673), .B(n9487), .S(n13831), .Z(n10630) );
  INV_X1 U13315 ( .A(n10999), .ZN(n10629) );
  NAND2_X1 U13316 ( .A1(n10630), .A2(n10629), .ZN(n10633) );
  INV_X1 U13317 ( .A(n10630), .ZN(n10631) );
  NAND2_X1 U13318 ( .A1(n10631), .A2(n10999), .ZN(n10632) );
  NAND2_X1 U13319 ( .A1(n10633), .A2(n10632), .ZN(n10985) );
  INV_X1 U13320 ( .A(n10633), .ZN(n11027) );
  MUX2_X1 U13321 ( .A(n7134), .B(n15864), .S(n13831), .Z(n10634) );
  NAND2_X1 U13322 ( .A1(n10634), .A2(n7206), .ZN(n11163) );
  INV_X1 U13323 ( .A(n10634), .ZN(n10635) );
  NAND2_X1 U13324 ( .A1(n10635), .A2(n11033), .ZN(n10636) );
  AND2_X1 U13325 ( .A1(n11163), .A2(n10636), .ZN(n11026) );
  INV_X1 U13326 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11508) );
  MUX2_X1 U13327 ( .A(n11508), .B(n9505), .S(n13831), .Z(n10637) );
  INV_X1 U13328 ( .A(n10788), .ZN(n11169) );
  NAND2_X1 U13329 ( .A1(n10637), .A2(n11169), .ZN(n10640) );
  INV_X1 U13330 ( .A(n10637), .ZN(n10638) );
  NAND2_X1 U13331 ( .A1(n10638), .A2(n10788), .ZN(n10639) );
  NAND2_X1 U13332 ( .A1(n10640), .A2(n10639), .ZN(n11162) );
  INV_X1 U13333 ( .A(n10640), .ZN(n11344) );
  INV_X1 U13334 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11517) );
  INV_X1 U13335 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11545) );
  MUX2_X1 U13336 ( .A(n11517), .B(n11545), .S(n13831), .Z(n10641) );
  NAND2_X1 U13337 ( .A1(n10641), .A2(n11349), .ZN(n13129) );
  INV_X1 U13338 ( .A(n10641), .ZN(n10642) );
  NAND2_X1 U13339 ( .A1(n10642), .A2(n10791), .ZN(n10643) );
  AND2_X1 U13340 ( .A1(n13129), .A2(n10643), .ZN(n11343) );
  INV_X1 U13341 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11620) );
  MUX2_X1 U13342 ( .A(n11620), .B(n15867), .S(n13831), .Z(n10644) );
  NAND2_X1 U13343 ( .A1(n10644), .A2(n10683), .ZN(n11229) );
  INV_X1 U13344 ( .A(n10644), .ZN(n10645) );
  NAND2_X1 U13345 ( .A1(n10645), .A2(n13134), .ZN(n10646) );
  NAND2_X1 U13346 ( .A1(n11229), .A2(n10646), .ZN(n13128) );
  INV_X1 U13347 ( .A(n11229), .ZN(n10651) );
  INV_X1 U13348 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11606) );
  MUX2_X1 U13349 ( .A(n11606), .B(n15869), .S(n13831), .Z(n10647) );
  NAND2_X1 U13350 ( .A1(n10647), .A2(n10684), .ZN(n10652) );
  INV_X1 U13351 ( .A(n10647), .ZN(n10648) );
  NAND2_X1 U13352 ( .A1(n10648), .A2(n11238), .ZN(n10649) );
  NAND2_X1 U13353 ( .A1(n10652), .A2(n10649), .ZN(n11228) );
  INV_X1 U13354 ( .A(n11228), .ZN(n10650) );
  OAI21_X1 U13355 ( .B1(n13132), .B2(n10651), .A(n10650), .ZN(n11232) );
  NAND2_X1 U13356 ( .A1(n11232), .A2(n10652), .ZN(n13163) );
  XNOR2_X1 U13357 ( .A(n10653), .B(n10687), .ZN(n13162) );
  MUX2_X1 U13358 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13831), .Z(n10654) );
  NAND2_X1 U13359 ( .A1(n11490), .A2(n10654), .ZN(n11484) );
  MUX2_X1 U13360 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13831), .Z(n10655) );
  XNOR2_X1 U13361 ( .A(n11869), .B(n10655), .ZN(n11856) );
  MUX2_X1 U13362 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13831), .Z(n10656) );
  XNOR2_X1 U13363 ( .A(n10658), .B(n10656), .ZN(n13171) );
  INV_X1 U13364 ( .A(n10656), .ZN(n10657) );
  AOI22_X1 U13365 ( .A1(n13172), .A2(n13171), .B1(n10658), .B2(n10657), .ZN(
        n13199) );
  XNOR2_X1 U13366 ( .A(n13190), .B(n10659), .ZN(n13198) );
  XNOR2_X1 U13367 ( .A(n10893), .B(n10661), .ZN(n13211) );
  INV_X1 U13368 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n10663) );
  OR2_X1 U13369 ( .A1(n13230), .A2(n10663), .ZN(n10696) );
  NAND2_X1 U13370 ( .A1(n13230), .A2(n10663), .ZN(n10664) );
  AND2_X1 U13371 ( .A1(n10696), .A2(n10664), .ZN(n13221) );
  MUX2_X1 U13372 ( .A(n13232), .B(n13221), .S(n13305), .Z(n13237) );
  MUX2_X1 U13373 ( .A(n10665), .B(n10696), .S(n13305), .Z(n10666) );
  NAND2_X1 U13374 ( .A1(n13236), .A2(n10666), .ZN(n10668) );
  INV_X1 U13375 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n10667) );
  INV_X1 U13376 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13738) );
  MUX2_X1 U13377 ( .A(n10667), .B(n13738), .S(n13831), .Z(n13246) );
  XOR2_X1 U13378 ( .A(n10699), .B(n10669), .Z(n13262) );
  XOR2_X1 U13379 ( .A(n10670), .B(n10976), .Z(n13283) );
  AOI21_X1 U13380 ( .B1(n10670), .B2(n13287), .A(n13281), .ZN(n13304) );
  XNOR2_X1 U13381 ( .A(n13304), .B(n13303), .ZN(n10671) );
  NOR2_X1 U13382 ( .A1(n10671), .A2(n10672), .ZN(n13302) );
  AND2_X1 U13383 ( .A1(n12915), .A2(P3_U3897), .ZN(n13315) );
  INV_X1 U13384 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10693) );
  INV_X1 U13385 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10690) );
  XNOR2_X1 U13386 ( .A(n10999), .B(n10673), .ZN(n10984) );
  NAND2_X1 U13387 ( .A1(n10674), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10675) );
  NAND2_X1 U13388 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13389 ( .A1(n6516), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13390 ( .A1(n10677), .A2(n10678), .ZN(n11005) );
  OR2_X1 U13391 ( .A1(n11005), .A2(n15815), .ZN(n11003) );
  NAND2_X1 U13392 ( .A1(n11003), .A2(n10678), .ZN(n10983) );
  NAND2_X1 U13393 ( .A1(n10984), .A2(n10983), .ZN(n10982) );
  NAND2_X1 U13394 ( .A1(n10999), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13395 ( .A1(n10982), .A2(n10679), .ZN(n10680) );
  OR2_X1 U13396 ( .A1(n10680), .A2(n11033), .ZN(n10681) );
  NAND2_X1 U13397 ( .A1(n10680), .A2(n11033), .ZN(n11154) );
  XNOR2_X1 U13398 ( .A(n10788), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11155) );
  XNOR2_X1 U13399 ( .A(n10683), .B(n11620), .ZN(n13137) );
  AOI21_X1 U13400 ( .B1(n13138), .B2(n6661), .A(n13137), .ZN(n13140) );
  AOI21_X1 U13401 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n13134), .A(n13140), .ZN(
        n10685) );
  NOR2_X1 U13402 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  AOI21_X1 U13403 ( .B1(n10685), .B2(n10684), .A(n10686), .ZN(n11227) );
  NAND2_X1 U13404 ( .A1(n11227), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n13151) );
  INV_X1 U13405 ( .A(n10686), .ZN(n13149) );
  INV_X1 U13406 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11774) );
  XNOR2_X1 U13407 ( .A(n10687), .B(n11774), .ZN(n13150) );
  AOI21_X1 U13408 ( .B1(n13151), .B2(n13149), .A(n13150), .ZN(n13153) );
  AOI21_X1 U13409 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13158), .A(n13153), .ZN(
        n10689) );
  NOR2_X1 U13410 ( .A1(n10689), .A2(n10688), .ZN(n11859) );
  XNOR2_X1 U13411 ( .A(n11869), .B(n10690), .ZN(n11858) );
  NAND2_X1 U13412 ( .A1(n10691), .A2(n13175), .ZN(n10692) );
  INV_X1 U13413 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13170) );
  INV_X1 U13414 ( .A(n10692), .ZN(n13185) );
  XNOR2_X1 U13415 ( .A(n13190), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n13184) );
  INV_X1 U13416 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12214) );
  INV_X1 U13417 ( .A(n10694), .ZN(n13220) );
  NAND2_X1 U13418 ( .A1(n13219), .A2(n10696), .ZN(n10695) );
  INV_X1 U13419 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n10698) );
  NOR2_X1 U13420 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  AOI21_X1 U13421 ( .B1(n10699), .B2(n10698), .A(n10700), .ZN(n13260) );
  INV_X1 U13422 ( .A(n10700), .ZN(n10701) );
  NAND2_X1 U13423 ( .A1(n13279), .A2(n10707), .ZN(n10704) );
  NAND2_X1 U13424 ( .A1(n11119), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13295) );
  NAND2_X1 U13425 ( .A1(n13303), .A2(n10702), .ZN(n10703) );
  AND2_X1 U13426 ( .A1(n13295), .A2(n10703), .ZN(n10705) );
  NAND2_X1 U13427 ( .A1(n10704), .A2(n10705), .ZN(n13296) );
  INV_X1 U13428 ( .A(n10705), .ZN(n10706) );
  NAND3_X1 U13429 ( .A1(n13279), .A2(n10707), .A3(n10706), .ZN(n10710) );
  INV_X1 U13430 ( .A(n10708), .ZN(n10711) );
  AOI21_X1 U13431 ( .B1(n13296), .B2(n10710), .A(n13319), .ZN(n10716) );
  INV_X1 U13432 ( .A(P3_U3897), .ZN(n13114) );
  MUX2_X1 U13433 ( .A(n13114), .B(n10711), .S(n12915), .Z(n13313) );
  NAND2_X1 U13434 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13077)
         );
  NAND2_X1 U13435 ( .A1(n15779), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n10714) );
  OAI211_X1 U13436 ( .C1(n13313), .C2(n11119), .A(n13077), .B(n10714), .ZN(
        n10715) );
  NAND2_X1 U13437 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n11176) );
  MUX2_X1 U13438 ( .A(n8213), .B(P1_REG2_REG_1__SCAN_IN), .S(n10730), .Z(
        n10724) );
  NOR2_X1 U13439 ( .A1(n10724), .A2(n11176), .ZN(n14756) );
  INV_X1 U13440 ( .A(n10719), .ZN(n10718) );
  NAND2_X1 U13441 ( .A1(n10718), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12881) );
  INV_X1 U13442 ( .A(n12881), .ZN(n12101) );
  OR2_X1 U13443 ( .A1(n10756), .A2(n12101), .ZN(n10732) );
  NAND2_X1 U13444 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  NAND2_X1 U13445 ( .A1(n10721), .A2(n8235), .ZN(n10731) );
  INV_X1 U13446 ( .A(n10731), .ZN(n10722) );
  NAND2_X1 U13447 ( .A1(n10732), .A2(n10722), .ZN(n10887) );
  INV_X1 U13448 ( .A(n10101), .ZN(n11175) );
  NAND2_X1 U13449 ( .A1(n10881), .A2(n11175), .ZN(n10723) );
  AOI211_X1 U13450 ( .C1(n11176), .C2(n10724), .A(n14756), .B(n14805), .ZN(
        n10736) );
  NAND2_X1 U13451 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10729) );
  MUX2_X1 U13452 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10839), .S(n10730), .Z(
        n10725) );
  INV_X1 U13453 ( .A(n10725), .ZN(n10728) );
  INV_X1 U13454 ( .A(n10838), .ZN(n10727) );
  INV_X1 U13455 ( .A(n10887), .ZN(n10726) );
  NAND2_X1 U13456 ( .A1(n10726), .A2(n10101), .ZN(n14817) );
  AOI211_X1 U13457 ( .C1(n10729), .C2(n10728), .A(n10727), .B(n14817), .ZN(
        n10735) );
  INV_X1 U13458 ( .A(n10730), .ZN(n10848) );
  NOR2_X1 U13459 ( .A1(n14765), .A2(n10848), .ZN(n10734) );
  NAND2_X1 U13460 ( .A1(n10732), .A2(n10731), .ZN(n15483) );
  OAI22_X1 U13461 ( .A1(n15483), .A2(n7877), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15115), .ZN(n10733) );
  OR4_X1 U13462 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        P1_U3244) );
  AND2_X1 U13463 ( .A1(n10769), .A2(P2_U3088), .ZN(n14565) );
  INV_X2 U13464 ( .A(n14565), .ZN(n14562) );
  NAND2_X1 U13465 ( .A1(n10071), .A2(P2_U3088), .ZN(n14569) );
  OAI222_X1 U13466 ( .A1(n14562), .A2(n13590), .B1(n14569), .B2(n10778), .C1(
        P2_U3088), .C2(n15639), .ZN(P2_U3325) );
  NAND2_X1 U13467 ( .A1(n10737), .A2(n13816), .ZN(n10738) );
  OAI21_X1 U13468 ( .B1(n10739), .B2(n13816), .A(n10738), .ZN(P3_U3377) );
  INV_X1 U13469 ( .A(n10740), .ZN(n10785) );
  OAI222_X1 U13470 ( .A1(n14562), .A2(n10741), .B1(n14569), .B2(n10785), .C1(
        P2_U3088), .C2(n14031), .ZN(P2_U3324) );
  INV_X1 U13471 ( .A(n10742), .ZN(n10781) );
  OAI222_X1 U13472 ( .A1(n14562), .A2(n10743), .B1(n14569), .B2(n10781), .C1(
        P2_U3088), .C2(n11088), .ZN(P2_U3323) );
  NAND2_X1 U13473 ( .A1(n10071), .A2(P1_U3086), .ZN(n15307) );
  INV_X1 U13474 ( .A(n10744), .ZN(n10750) );
  INV_X1 U13475 ( .A(n10920), .ZN(n10905) );
  OAI222_X1 U13476 ( .A1(n15307), .A2(n10745), .B1(n15305), .B2(n10750), .C1(
        P1_U3086), .C2(n10905), .ZN(P1_U3348) );
  INV_X1 U13477 ( .A(n10746), .ZN(n10783) );
  OAI222_X1 U13478 ( .A1(n14058), .A2(P2_U3088), .B1(n14569), .B2(n10783), 
        .C1(n10747), .C2(n14562), .ZN(P2_U3321) );
  OAI222_X1 U13479 ( .A1(n15619), .A2(P2_U3088), .B1(n12913), .B2(n10777), 
        .C1(n10748), .C2(n14562), .ZN(P2_U3326) );
  INV_X1 U13480 ( .A(n14074), .ZN(n10751) );
  INV_X1 U13481 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10749) );
  OAI222_X1 U13482 ( .A1(n10751), .A2(P2_U3088), .B1(n12913), .B2(n10750), 
        .C1(n10749), .C2(n14562), .ZN(P2_U3320) );
  INV_X1 U13483 ( .A(n10752), .ZN(n10779) );
  OAI222_X1 U13484 ( .A1(n14562), .A2(n10753), .B1(n12913), .B2(n10779), .C1(
        P2_U3088), .C2(n14045), .ZN(P2_U3322) );
  INV_X1 U13485 ( .A(n10754), .ZN(n10755) );
  INV_X1 U13486 ( .A(n10757), .ZN(n10758) );
  AOI22_X1 U13487 ( .A1(n15541), .A2(n10759), .B1(n10758), .B2(n10761), .ZN(
        P1_U3446) );
  INV_X1 U13488 ( .A(n10760), .ZN(n10762) );
  AOI22_X1 U13489 ( .A1(n15541), .A2(n10763), .B1(n10762), .B2(n10761), .ZN(
        P1_U3445) );
  INV_X1 U13490 ( .A(n10764), .ZN(n10767) );
  OAI222_X1 U13491 ( .A1(n15307), .A2(n10765), .B1(n15305), .B2(n10767), .C1(
        P1_U3086), .C2(n6706), .ZN(P1_U3347) );
  INV_X1 U13492 ( .A(n14084), .ZN(n14080) );
  INV_X1 U13493 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10766) );
  OAI222_X1 U13494 ( .A1(n14080), .A2(P2_U3088), .B1(n12913), .B2(n10767), 
        .C1(n10766), .C2(n14562), .ZN(P2_U3319) );
  NAND2_X1 U13495 ( .A1(n10071), .A2(P3_U3151), .ZN(n12918) );
  INV_X1 U13496 ( .A(SI_6_), .ZN(n10772) );
  NAND2_X1 U13497 ( .A1(n10769), .A2(P3_U3151), .ZN(n12160) );
  INV_X1 U13498 ( .A(n10770), .ZN(n10771) );
  OAI222_X1 U13499 ( .A1(n12918), .A2(n10772), .B1(n12160), .B2(n10771), .C1(
        P3_U3151), .C2(n13134), .ZN(P3_U3289) );
  INV_X1 U13500 ( .A(n10773), .ZN(n10774) );
  OAI222_X1 U13501 ( .A1(n12918), .A2(n10775), .B1(n12160), .B2(n10774), .C1(
        n11017), .C2(P3_U3151), .ZN(P3_U3294) );
  INV_X1 U13502 ( .A(n15307), .ZN(n15299) );
  INV_X1 U13503 ( .A(n15299), .ZN(n12946) );
  OAI222_X1 U13504 ( .A1(n10848), .A2(P1_U3086), .B1(n15305), .B2(n10777), 
        .C1(n10776), .C2(n12946), .ZN(P1_U3354) );
  OAI222_X1 U13505 ( .A1(n8254), .A2(P1_U3086), .B1(n15305), .B2(n10778), .C1(
        n9472), .C2(n12946), .ZN(P1_U3353) );
  OAI222_X1 U13506 ( .A1(n10895), .A2(P1_U3086), .B1(n15305), .B2(n10779), 
        .C1(n7399), .C2(n12946), .ZN(P1_U3350) );
  INV_X1 U13507 ( .A(n10852), .ZN(n11183) );
  OAI222_X1 U13508 ( .A1(n11183), .A2(P1_U3086), .B1(n15305), .B2(n10781), 
        .C1(n10780), .C2(n12946), .ZN(P1_U3351) );
  INV_X1 U13509 ( .A(n10899), .ZN(n10932) );
  OAI222_X1 U13510 ( .A1(n10932), .A2(P1_U3086), .B1(n15305), .B2(n10783), 
        .C1(n10782), .C2(n12946), .ZN(P1_U3349) );
  OAI222_X1 U13511 ( .A1(n7034), .A2(P1_U3086), .B1(n15305), .B2(n10785), .C1(
        n10784), .C2(n12946), .ZN(P1_U3352) );
  INV_X1 U13512 ( .A(n15483), .ZN(n14768) );
  NOR2_X1 U13513 ( .A1(n14768), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13514 ( .A(SI_4_), .ZN(n10786) );
  OAI222_X1 U13515 ( .A1(P3_U3151), .A2(n10788), .B1(n12160), .B2(n10787), 
        .C1(n10786), .C2(n12918), .ZN(P3_U3291) );
  INV_X1 U13516 ( .A(SI_5_), .ZN(n10789) );
  OAI222_X1 U13517 ( .A1(P3_U3151), .A2(n10791), .B1(n12160), .B2(n10790), 
        .C1(n10789), .C2(n12918), .ZN(P3_U3290) );
  OAI222_X1 U13518 ( .A1(P3_U3151), .A2(n11033), .B1(n12160), .B2(n10793), 
        .C1(n10792), .C2(n12918), .ZN(P3_U3292) );
  INV_X1 U13519 ( .A(SI_2_), .ZN(n10794) );
  OAI222_X1 U13520 ( .A1(P3_U3151), .A2(n10999), .B1(n12160), .B2(n10795), 
        .C1(n10794), .C2(n12918), .ZN(P3_U3293) );
  INV_X1 U13521 ( .A(n10796), .ZN(n10798) );
  OAI222_X1 U13522 ( .A1(n15675), .A2(P2_U3088), .B1(n14569), .B2(n10798), 
        .C1(n10797), .C2(n14562), .ZN(P2_U3318) );
  INV_X1 U13523 ( .A(n10949), .ZN(n10961) );
  OAI222_X1 U13524 ( .A1(n15307), .A2(n10799), .B1(n15305), .B2(n10798), .C1(
        P1_U3086), .C2(n10961), .ZN(P1_U3346) );
  INV_X1 U13525 ( .A(n13816), .ZN(n10801) );
  NOR2_X1 U13526 ( .A1(n10801), .A2(n10800), .ZN(n10803) );
  INV_X1 U13527 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10802) );
  NOR2_X1 U13528 ( .A1(n10803), .A2(n10802), .ZN(P3_U3258) );
  CLKBUF_X1 U13529 ( .A(n10803), .Z(n10827) );
  INV_X1 U13530 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10804) );
  NOR2_X1 U13531 ( .A1(n10827), .A2(n10804), .ZN(P3_U3251) );
  INV_X1 U13532 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10805) );
  NOR2_X1 U13533 ( .A1(n10827), .A2(n10805), .ZN(P3_U3254) );
  INV_X1 U13534 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10806) );
  NOR2_X1 U13535 ( .A1(n10827), .A2(n10806), .ZN(P3_U3257) );
  INV_X1 U13536 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10807) );
  NOR2_X1 U13537 ( .A1(n10827), .A2(n10807), .ZN(P3_U3252) );
  INV_X1 U13538 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10808) );
  NOR2_X1 U13539 ( .A1(n10827), .A2(n10808), .ZN(P3_U3253) );
  INV_X1 U13540 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10809) );
  NOR2_X1 U13541 ( .A1(n10827), .A2(n10809), .ZN(P3_U3255) );
  INV_X1 U13542 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U13543 ( .A1(n10827), .A2(n10810), .ZN(P3_U3256) );
  INV_X1 U13544 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10811) );
  NOR2_X1 U13545 ( .A1(n10803), .A2(n10811), .ZN(P3_U3260) );
  INV_X1 U13546 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10812) );
  NOR2_X1 U13547 ( .A1(n10827), .A2(n10812), .ZN(P3_U3259) );
  INV_X1 U13548 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10813) );
  NOR2_X1 U13549 ( .A1(n10827), .A2(n10813), .ZN(P3_U3263) );
  INV_X1 U13550 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n13633) );
  NOR2_X1 U13551 ( .A1(n10803), .A2(n13633), .ZN(P3_U3262) );
  INV_X1 U13552 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10814) );
  NOR2_X1 U13553 ( .A1(n10803), .A2(n10814), .ZN(P3_U3235) );
  INV_X1 U13554 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10815) );
  NOR2_X1 U13555 ( .A1(n10803), .A2(n10815), .ZN(P3_U3238) );
  INV_X1 U13556 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10816) );
  NOR2_X1 U13557 ( .A1(n10803), .A2(n10816), .ZN(P3_U3239) );
  INV_X1 U13558 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10817) );
  NOR2_X1 U13559 ( .A1(n10827), .A2(n10817), .ZN(P3_U3247) );
  INV_X1 U13560 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10818) );
  NOR2_X1 U13561 ( .A1(n10803), .A2(n10818), .ZN(P3_U3234) );
  INV_X1 U13562 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10819) );
  NOR2_X1 U13563 ( .A1(n10827), .A2(n10819), .ZN(P3_U3246) );
  INV_X1 U13564 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10820) );
  NOR2_X1 U13565 ( .A1(n10827), .A2(n10820), .ZN(P3_U3261) );
  INV_X1 U13566 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10821) );
  NOR2_X1 U13567 ( .A1(n10803), .A2(n10821), .ZN(P3_U3236) );
  INV_X1 U13568 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10822) );
  NOR2_X1 U13569 ( .A1(n10803), .A2(n10822), .ZN(P3_U3245) );
  INV_X1 U13570 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10823) );
  NOR2_X1 U13571 ( .A1(n10803), .A2(n10823), .ZN(P3_U3237) );
  INV_X1 U13572 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10824) );
  NOR2_X1 U13573 ( .A1(n10827), .A2(n10824), .ZN(P3_U3250) );
  INV_X1 U13574 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10825) );
  NOR2_X1 U13575 ( .A1(n10827), .A2(n10825), .ZN(P3_U3249) );
  INV_X1 U13576 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10826) );
  NOR2_X1 U13577 ( .A1(n10827), .A2(n10826), .ZN(P3_U3248) );
  INV_X1 U13578 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10828) );
  NOR2_X1 U13579 ( .A1(n10803), .A2(n10828), .ZN(P3_U3240) );
  INV_X1 U13580 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10829) );
  NOR2_X1 U13581 ( .A1(n10827), .A2(n10829), .ZN(P3_U3241) );
  INV_X1 U13582 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10830) );
  NOR2_X1 U13583 ( .A1(n10827), .A2(n10830), .ZN(P3_U3243) );
  INV_X1 U13584 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13585 ( .A1(n10827), .A2(n10831), .ZN(P3_U3244) );
  INV_X1 U13586 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10832) );
  NOR2_X1 U13587 ( .A1(n10827), .A2(n10832), .ZN(P3_U3242) );
  INV_X1 U13588 ( .A(n11267), .ZN(n10835) );
  INV_X1 U13589 ( .A(n10833), .ZN(n10836) );
  INV_X1 U13590 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10834) );
  OAI222_X1 U13591 ( .A1(n10835), .A2(P2_U3088), .B1(n12913), .B2(n10836), 
        .C1(n10834), .C2(n14562), .ZN(P2_U3317) );
  INV_X1 U13592 ( .A(n11139), .ZN(n11135) );
  OAI222_X1 U13593 ( .A1(n15307), .A2(n10837), .B1(n15305), .B2(n10836), .C1(
        P1_U3086), .C2(n11135), .ZN(P1_U3345) );
  MUX2_X1 U13594 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10896), .S(n10895), .Z(
        n10844) );
  INV_X1 U13595 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10841) );
  INV_X1 U13596 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10840) );
  XOR2_X1 U13597 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10851), .Z(n14771) );
  NAND2_X1 U13598 ( .A1(n14770), .A2(n14771), .ZN(n14769) );
  OAI21_X1 U13599 ( .B1(n7034), .B2(n10841), .A(n14769), .ZN(n11187) );
  XOR2_X1 U13600 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10852), .Z(n11188) );
  AOI21_X1 U13601 ( .B1(n10844), .B2(n10843), .A(n10894), .ZN(n10858) );
  INV_X1 U13602 ( .A(n10895), .ZN(n10898) );
  INV_X1 U13603 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U13604 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11417) );
  OAI21_X1 U13605 ( .B1(n15483), .B2(n10845), .A(n11417), .ZN(n10846) );
  AOI21_X1 U13606 ( .B1(n15475), .B2(n10898), .A(n10846), .ZN(n10857) );
  MUX2_X1 U13607 ( .A(n10847), .B(P1_REG2_REG_5__SCAN_IN), .S(n10895), .Z(
        n10855) );
  NOR2_X1 U13608 ( .A1(n10848), .A2(n8213), .ZN(n14752) );
  MUX2_X1 U13609 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10849), .S(n14751), .Z(
        n10850) );
  NAND2_X1 U13610 ( .A1(n14751), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14773) );
  MUX2_X1 U13611 ( .A(n15512), .B(P1_REG2_REG_3__SCAN_IN), .S(n10851), .Z(
        n14772) );
  MUX2_X1 U13612 ( .A(n10853), .B(P1_REG2_REG_4__SCAN_IN), .S(n10852), .Z(
        n11184) );
  NAND2_X1 U13613 ( .A1(n10854), .A2(n10855), .ZN(n10938) );
  OAI211_X1 U13614 ( .C1(n10855), .C2(n10854), .A(n15479), .B(n10938), .ZN(
        n10856) );
  OAI211_X1 U13615 ( .C1(n10858), .C2(n14817), .A(n10857), .B(n10856), .ZN(
        P1_U3248) );
  INV_X1 U13616 ( .A(n13190), .ZN(n10862) );
  INV_X1 U13617 ( .A(n10859), .ZN(n10861) );
  INV_X1 U13618 ( .A(n12918), .ZN(n13822) );
  OAI222_X1 U13619 ( .A1(P3_U3151), .A2(n10862), .B1(n12160), .B2(n10861), 
        .C1(n10860), .C2(n13838), .ZN(P3_U3283) );
  OAI222_X1 U13620 ( .A1(n13175), .A2(P3_U3151), .B1(n12160), .B2(n10864), 
        .C1(n10863), .C2(n13838), .ZN(P3_U3284) );
  INV_X1 U13621 ( .A(n10865), .ZN(n10868) );
  OAI222_X1 U13622 ( .A1(n12946), .A2(n10866), .B1(n15305), .B2(n10868), .C1(
        P1_U3086), .C2(n7019), .ZN(P1_U3344) );
  INV_X1 U13623 ( .A(n11798), .ZN(n10869) );
  OAI222_X1 U13624 ( .A1(n10869), .A2(P2_U3088), .B1(n12913), .B2(n10868), 
        .C1(n10867), .C2(n14562), .ZN(P2_U3316) );
  INV_X1 U13625 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U13626 ( .A1(n11365), .A2(P3_U3897), .ZN(n10870) );
  OAI21_X1 U13627 ( .B1(P3_U3897), .B2(n13621), .A(n10870), .ZN(P3_U3495) );
  INV_X1 U13628 ( .A(n11781), .ZN(n13836) );
  OAI222_X1 U13629 ( .A1(n11869), .A2(P3_U3151), .B1(n13836), .B2(n10872), 
        .C1(n10871), .C2(n12918), .ZN(P3_U3285) );
  INV_X1 U13630 ( .A(n10873), .ZN(n10875) );
  INV_X1 U13631 ( .A(SI_8_), .ZN(n10874) );
  OAI222_X1 U13632 ( .A1(P3_U3151), .A2(n13158), .B1(n13836), .B2(n10875), 
        .C1(n10874), .C2(n12918), .ZN(P3_U3287) );
  OAI222_X1 U13633 ( .A1(n11238), .A2(P3_U3151), .B1(n13836), .B2(n10876), 
        .C1(n13591), .C2(n13838), .ZN(P3_U3288) );
  OAI222_X1 U13634 ( .A1(n11490), .A2(P3_U3151), .B1(n13836), .B2(n10878), 
        .C1(n10877), .C2(n12918), .ZN(P3_U3286) );
  NAND2_X1 U13635 ( .A1(n11175), .A2(n10879), .ZN(n10880) );
  NAND2_X1 U13636 ( .A1(n10881), .A2(n10880), .ZN(n11180) );
  INV_X1 U13637 ( .A(n11180), .ZN(n10883) );
  NAND2_X1 U13638 ( .A1(n10101), .A2(n8240), .ZN(n10882) );
  NAND2_X1 U13639 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  MUX2_X1 U13640 ( .A(n10884), .B(n10883), .S(P1_IR_REG_0__SCAN_IN), .Z(n10886) );
  OAI22_X1 U13641 ( .A1(n10887), .A2(n10886), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10885), .ZN(n10888) );
  AOI21_X1 U13642 ( .B1(n14768), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n10888), .ZN(
        n10890) );
  NAND3_X1 U13643 ( .A1(n15478), .A2(P1_IR_REG_0__SCAN_IN), .A3(n8240), .ZN(
        n10889) );
  NAND2_X1 U13644 ( .A1(n10890), .A2(n10889), .ZN(P1_U3243) );
  OAI222_X1 U13645 ( .A1(n10893), .A2(P3_U3151), .B1(n12160), .B2(n10892), 
        .C1(n10891), .C2(n13838), .ZN(P3_U3282) );
  INV_X1 U13646 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15613) );
  MUX2_X1 U13647 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15613), .S(n10899), .Z(
        n10931) );
  XNOR2_X1 U13648 ( .A(n10920), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10897) );
  AOI211_X1 U13649 ( .C1(n6642), .C2(n10897), .A(n14817), .B(n10919), .ZN(
        n10908) );
  NAND2_X1 U13650 ( .A1(n10898), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10937) );
  MUX2_X1 U13651 ( .A(n11955), .B(P1_REG2_REG_6__SCAN_IN), .S(n10899), .Z(
        n10936) );
  AOI21_X1 U13652 ( .B1(n10938), .B2(n10937), .A(n10936), .ZN(n10935) );
  NOR2_X1 U13653 ( .A1(n10932), .A2(n11955), .ZN(n10901) );
  MUX2_X1 U13654 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11942), .S(n10920), .Z(
        n10900) );
  INV_X1 U13655 ( .A(n10917), .ZN(n10903) );
  NOR3_X1 U13656 ( .A1(n10935), .A2(n10901), .A3(n10900), .ZN(n10902) );
  NOR3_X1 U13657 ( .A1(n10903), .A2(n10902), .A3(n14805), .ZN(n10907) );
  NAND2_X1 U13658 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U13659 ( .A1(n14768), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10904) );
  OAI211_X1 U13660 ( .C1(n14765), .C2(n10905), .A(n11712), .B(n10904), .ZN(
        n10906) );
  OR3_X1 U13661 ( .A1(n10908), .A2(n10907), .A3(n10906), .ZN(P1_U3250) );
  INV_X1 U13662 ( .A(n10909), .ZN(n10910) );
  OAI222_X1 U13663 ( .A1(P3_U3151), .A2(n6997), .B1(n12160), .B2(n10910), .C1(
        n13693), .C2(n13838), .ZN(P3_U3280) );
  INV_X1 U13664 ( .A(n10911), .ZN(n10913) );
  OAI222_X1 U13665 ( .A1(n15695), .A2(P2_U3088), .B1(n12913), .B2(n10913), 
        .C1(n10912), .C2(n14562), .ZN(P2_U3315) );
  INV_X1 U13666 ( .A(n11460), .ZN(n11289) );
  OAI222_X1 U13667 ( .A1(n15307), .A2(n10914), .B1(n15305), .B2(n10913), .C1(
        P1_U3086), .C2(n11289), .ZN(P1_U3343) );
  NAND2_X1 U13668 ( .A1(n10920), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10916) );
  MUX2_X1 U13669 ( .A(n12010), .B(P1_REG2_REG_8__SCAN_IN), .S(n10946), .Z(
        n10915) );
  NAND3_X1 U13670 ( .A1(n10917), .A2(n10916), .A3(n10915), .ZN(n10918) );
  NAND2_X1 U13671 ( .A1(n10918), .A2(n15479), .ZN(n10929) );
  AOI21_X1 U13672 ( .B1(n10920), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10919), .ZN(
        n10923) );
  MUX2_X1 U13673 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10921), .S(n10946), .Z(
        n10922) );
  OAI21_X1 U13674 ( .B1(n10923), .B2(n10922), .A(n10945), .ZN(n10924) );
  NAND2_X1 U13675 ( .A1(n10924), .A2(n15478), .ZN(n10928) );
  NAND2_X1 U13676 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11909) );
  INV_X1 U13677 ( .A(n11909), .ZN(n10926) );
  NOR2_X1 U13678 ( .A1(n14765), .A2(n6706), .ZN(n10925) );
  AOI211_X1 U13679 ( .C1(n14768), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10926), .B(
        n10925), .ZN(n10927) );
  OAI211_X1 U13680 ( .C1(n10952), .C2(n10929), .A(n10928), .B(n10927), .ZN(
        P1_U3251) );
  OAI21_X1 U13681 ( .B1(n10931), .B2(n10930), .A(n15478), .ZN(n10943) );
  AND2_X1 U13682 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10934) );
  NOR2_X1 U13683 ( .A1(n14765), .A2(n10932), .ZN(n10933) );
  AOI211_X1 U13684 ( .C1(n14768), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10934), .B(
        n10933), .ZN(n10942) );
  INV_X1 U13685 ( .A(n10935), .ZN(n10940) );
  NAND3_X1 U13686 ( .A1(n10938), .A2(n10937), .A3(n10936), .ZN(n10939) );
  NAND3_X1 U13687 ( .A1(n10940), .A2(n15479), .A3(n10939), .ZN(n10941) );
  OAI211_X1 U13688 ( .C1(n10944), .C2(n10943), .A(n10942), .B(n10941), .ZN(
        P1_U3249) );
  XNOR2_X1 U13689 ( .A(n10949), .B(n13696), .ZN(n10962) );
  XOR2_X1 U13690 ( .A(n10962), .B(n10963), .Z(n10955) );
  NOR2_X1 U13691 ( .A1(n13694), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12062) );
  NOR2_X1 U13692 ( .A1(n14765), .A2(n10961), .ZN(n10947) );
  AOI211_X1 U13693 ( .C1(n14768), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n12062), .B(
        n10947), .ZN(n10954) );
  MUX2_X1 U13694 ( .A(n8410), .B(P1_REG2_REG_9__SCAN_IN), .S(n10949), .Z(
        n10948) );
  NAND2_X1 U13695 ( .A1(n6659), .A2(n10948), .ZN(n10951) );
  NAND2_X1 U13696 ( .A1(n10949), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13697 ( .A1(n10961), .A2(n8410), .ZN(n10950) );
  OAI211_X1 U13698 ( .C1(n10952), .C2(n10951), .A(n10960), .B(n15479), .ZN(
        n10953) );
  OAI211_X1 U13699 ( .C1(n10955), .C2(n14817), .A(n10954), .B(n10953), .ZN(
        P1_U3252) );
  INV_X1 U13700 ( .A(n10956), .ZN(n10958) );
  OAI222_X1 U13701 ( .A1(P3_U3151), .A2(n13266), .B1(n12160), .B2(n10958), 
        .C1(n10957), .C2(n13838), .ZN(P3_U3279) );
  XNOR2_X1 U13702 ( .A(n11139), .B(n12183), .ZN(n11140) );
  XNOR2_X1 U13703 ( .A(n11141), .B(n11140), .ZN(n10970) );
  XOR2_X1 U13704 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11139), .Z(n10964) );
  OAI211_X1 U13705 ( .C1(n10965), .C2(n10964), .A(n11134), .B(n15478), .ZN(
        n10969) );
  NOR2_X1 U13706 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8448), .ZN(n10967) );
  NOR2_X1 U13707 ( .A1(n14765), .A2(n11135), .ZN(n10966) );
  AOI211_X1 U13708 ( .C1(n14768), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n10967), 
        .B(n10966), .ZN(n10968) );
  OAI211_X1 U13709 ( .C1(n10970), .C2(n14805), .A(n10969), .B(n10968), .ZN(
        P1_U3253) );
  INV_X1 U13710 ( .A(n13230), .ZN(n10974) );
  INV_X1 U13711 ( .A(n10971), .ZN(n10973) );
  OAI222_X1 U13712 ( .A1(P3_U3151), .A2(n10974), .B1(n12160), .B2(n10973), 
        .C1(n10972), .C2(n13838), .ZN(P3_U3281) );
  INV_X1 U13713 ( .A(n10975), .ZN(n10978) );
  OAI22_X1 U13714 ( .A1(n10976), .A2(P3_U3151), .B1(SI_17_), .B2(n13838), .ZN(
        n10977) );
  AOI21_X1 U13715 ( .B1(n10978), .B2(n11781), .A(n10977), .ZN(P3_U3278) );
  INV_X1 U13716 ( .A(n10979), .ZN(n10981) );
  OAI222_X1 U13717 ( .A1(P1_U3086), .A2(n11469), .B1(n15307), .B2(n10980), 
        .C1(n15305), .C2(n10981), .ZN(P1_U3342) );
  OAI222_X1 U13718 ( .A1(P2_U3088), .A2(n11803), .B1(n14562), .B2(n13593), 
        .C1(n12913), .C2(n10981), .ZN(P2_U3314) );
  OAI21_X1 U13719 ( .B1(n10984), .B2(n10983), .A(n10982), .ZN(n10997) );
  INV_X1 U13720 ( .A(n11028), .ZN(n10988) );
  NAND3_X1 U13721 ( .A1(n11006), .A2(n10986), .A3(n10985), .ZN(n10987) );
  AOI21_X1 U13722 ( .B1(n10988), .B2(n10987), .A(n13282), .ZN(n10996) );
  OAI21_X1 U13723 ( .B1(n10991), .B2(n10990), .A(n10989), .ZN(n10992) );
  NAND2_X1 U13724 ( .A1(n13300), .A2(n10992), .ZN(n10994) );
  AOI22_X1 U13725 ( .A1(n15779), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10993) );
  NAND2_X1 U13726 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  AOI211_X1 U13727 ( .C1(n13290), .C2(n10997), .A(n10996), .B(n10995), .ZN(
        n10998) );
  OAI21_X1 U13728 ( .B1(n10999), .B2(n13313), .A(n10998), .ZN(P3_U3184) );
  INV_X1 U13729 ( .A(n11000), .ZN(n11002) );
  OAI21_X1 U13730 ( .B1(n11002), .B2(P3_REG1_REG_1__SCAN_IN), .A(n11001), .ZN(
        n11015) );
  INV_X1 U13731 ( .A(n11003), .ZN(n11004) );
  AOI21_X1 U13732 ( .B1(n15815), .B2(n11005), .A(n11004), .ZN(n11011) );
  INV_X1 U13733 ( .A(n11006), .ZN(n11007) );
  AOI21_X1 U13734 ( .B1(n11009), .B2(n11008), .A(n11007), .ZN(n11010) );
  OAI22_X1 U13735 ( .A1(n13319), .A2(n11011), .B1(n13282), .B2(n11010), .ZN(
        n11014) );
  INV_X1 U13736 ( .A(n15779), .ZN(n13227) );
  INV_X1 U13737 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n11012) );
  INV_X1 U13738 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11115) );
  OAI22_X1 U13739 ( .A1(n13227), .A2(n11012), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11115), .ZN(n11013) );
  AOI211_X1 U13740 ( .C1(n13300), .C2(n11015), .A(n11014), .B(n11013), .ZN(
        n11016) );
  OAI21_X1 U13741 ( .B1(n11017), .B2(n13313), .A(n11016), .ZN(P3_U3183) );
  OAI21_X1 U13742 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11018), .A(n11156), .ZN(
        n11025) );
  INV_X1 U13743 ( .A(n11019), .ZN(n11021) );
  INV_X1 U13744 ( .A(n11151), .ZN(n11020) );
  AOI21_X1 U13745 ( .B1(n15864), .B2(n11021), .A(n11020), .ZN(n11023) );
  AOI22_X1 U13746 ( .A1(n15779), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11022) );
  OAI21_X1 U13747 ( .B1(n13293), .B2(n11023), .A(n11022), .ZN(n11024) );
  AOI21_X1 U13748 ( .B1(n13290), .B2(n11025), .A(n11024), .ZN(n11032) );
  INV_X1 U13749 ( .A(n11164), .ZN(n11030) );
  NOR3_X1 U13750 ( .A1(n11028), .A2(n11027), .A3(n11026), .ZN(n11029) );
  OAI21_X1 U13751 ( .B1(n11030), .B2(n11029), .A(n13315), .ZN(n11031) );
  OAI211_X1 U13752 ( .C1(n13313), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        P3_U3185) );
  OAI21_X1 U13753 ( .B1(n12595), .B2(n11035), .A(n11034), .ZN(n11036) );
  NAND2_X1 U13754 ( .A1(n11036), .A2(n14379), .ZN(n11038) );
  AOI22_X1 U13755 ( .A1(n14376), .A2(n14024), .B1(n14374), .B2(n14022), .ZN(
        n11037) );
  NAND2_X1 U13756 ( .A1(n11038), .A2(n11037), .ZN(n14395) );
  INV_X1 U13757 ( .A(n14395), .ZN(n11044) );
  OAI21_X1 U13758 ( .B1(n11572), .B2(n11039), .A(n14273), .ZN(n11040) );
  NOR2_X1 U13759 ( .A1(n11040), .A2(n11643), .ZN(n14398) );
  AND2_X1 U13760 ( .A1(n15750), .A2(n6421), .ZN(n11041) );
  NOR2_X1 U13761 ( .A1(n14398), .A2(n11041), .ZN(n11043) );
  INV_X1 U13762 ( .A(n12595), .ZN(n11639) );
  XNOR2_X1 U13763 ( .A(n11640), .B(n11639), .ZN(n14402) );
  NAND2_X1 U13764 ( .A1(n14402), .A2(n15764), .ZN(n11042) );
  AND3_X1 U13765 ( .A1(n11044), .A2(n11043), .A3(n11042), .ZN(n15739) );
  NAND2_X1 U13766 ( .A1(n15775), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11045) );
  OAI21_X1 U13767 ( .B1(n15775), .B2(n15739), .A(n11045), .ZN(P2_U3501) );
  NOR2_X1 U13768 ( .A1(n13094), .A2(P3_U3151), .ZN(n11226) );
  INV_X1 U13769 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11048) );
  OAI22_X1 U13770 ( .A1(n13079), .A2(n6837), .B1(n11358), .B2(n13083), .ZN(
        n11046) );
  AOI21_X1 U13771 ( .B1(n13074), .B2(n11254), .A(n11046), .ZN(n11047) );
  OAI21_X1 U13772 ( .B1(n11226), .B2(n11048), .A(n11047), .ZN(P3_U3172) );
  AOI21_X1 U13773 ( .B1(n11051), .B2(n11050), .A(n11049), .ZN(n11052) );
  OR2_X1 U13774 ( .A1(n11053), .A2(n11052), .ZN(n11076) );
  NOR2_X1 U13775 ( .A1(n11054), .A2(P2_U3088), .ZN(n14564) );
  AND2_X1 U13776 ( .A1(n11076), .A2(n14564), .ZN(n11101) );
  INV_X1 U13777 ( .A(n12942), .ZN(n12642) );
  NAND2_X1 U13778 ( .A1(n11101), .A2(n12642), .ZN(n14161) );
  INV_X1 U13779 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11583) );
  MUX2_X1 U13780 ( .A(n11583), .B(P2_REG2_REG_1__SCAN_IN), .S(n15619), .Z(
        n15628) );
  AND2_X1 U13781 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n15629) );
  NAND2_X1 U13782 ( .A1(n15628), .A2(n15629), .ZN(n15627) );
  NAND2_X1 U13783 ( .A1(n11082), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U13784 ( .A1(n15627), .A2(n11055), .ZN(n15642) );
  INV_X1 U13785 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11056) );
  MUX2_X1 U13786 ( .A(n11056), .B(P2_REG2_REG_2__SCAN_IN), .S(n15639), .Z(
        n15643) );
  NAND2_X1 U13787 ( .A1(n11084), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U13788 ( .A1(n15641), .A2(n14033), .ZN(n11058) );
  INV_X1 U13789 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11654) );
  MUX2_X1 U13790 ( .A(n11654), .B(P2_REG2_REG_3__SCAN_IN), .S(n14031), .Z(
        n11057) );
  NAND2_X1 U13791 ( .A1(n11058), .A2(n11057), .ZN(n14035) );
  INV_X1 U13792 ( .A(n14031), .ZN(n11086) );
  NAND2_X1 U13793 ( .A1(n11086), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n11059) );
  NAND2_X1 U13794 ( .A1(n14035), .A2(n11059), .ZN(n15656) );
  INV_X1 U13795 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11060) );
  MUX2_X1 U13796 ( .A(n11060), .B(P2_REG2_REG_4__SCAN_IN), .S(n11088), .Z(
        n15657) );
  INV_X1 U13797 ( .A(n11088), .ZN(n15654) );
  NAND2_X1 U13798 ( .A1(n15654), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14047) );
  INV_X1 U13799 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11635) );
  MUX2_X1 U13800 ( .A(n11635), .B(P2_REG2_REG_5__SCAN_IN), .S(n14045), .Z(
        n11061) );
  INV_X1 U13801 ( .A(n14045), .ZN(n11090) );
  NAND2_X1 U13802 ( .A1(n11090), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14060) );
  INV_X1 U13803 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11549) );
  MUX2_X1 U13804 ( .A(n11549), .B(P2_REG2_REG_6__SCAN_IN), .S(n14058), .Z(
        n11062) );
  OR2_X1 U13805 ( .A1(n14058), .A2(n11549), .ZN(n14067) );
  NAND2_X1 U13806 ( .A1(n14068), .A2(n14067), .ZN(n11065) );
  INV_X1 U13807 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11561) );
  MUX2_X1 U13808 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11561), .S(n14074), .Z(
        n11064) );
  NAND2_X1 U13809 ( .A1(n14074), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14086) );
  INV_X1 U13810 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11737) );
  MUX2_X1 U13811 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11737), .S(n14084), .Z(
        n11066) );
  NAND2_X1 U13812 ( .A1(n14084), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11067) );
  INV_X1 U13813 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11068) );
  MUX2_X1 U13814 ( .A(n11068), .B(P2_REG2_REG_9__SCAN_IN), .S(n15675), .Z(
        n15662) );
  NAND2_X1 U13815 ( .A1(n15663), .A2(n15662), .ZN(n15661) );
  NAND2_X1 U13816 ( .A1(n15675), .A2(n11068), .ZN(n11069) );
  NAND2_X1 U13817 ( .A1(n15661), .A2(n11069), .ZN(n11266) );
  INV_X1 U13818 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11070) );
  MUX2_X1 U13819 ( .A(n11070), .B(P2_REG2_REG_10__SCAN_IN), .S(n11267), .Z(
        n11265) );
  NAND2_X1 U13820 ( .A1(n11267), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11071) );
  INV_X1 U13821 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13667) );
  MUX2_X1 U13822 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13667), .S(n11798), .Z(
        n11072) );
  OAI21_X1 U13823 ( .B1(n11073), .B2(n11072), .A(n15682), .ZN(n11079) );
  NOR2_X2 U13824 ( .A1(n11076), .A2(P2_U3088), .ZN(n15634) );
  INV_X1 U13825 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U13826 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12293)
         );
  NOR2_X1 U13827 ( .A1(n11074), .A2(P2_U3088), .ZN(n11075) );
  NAND2_X1 U13828 ( .A1(n15707), .A2(n11798), .ZN(n11077) );
  OAI211_X1 U13829 ( .C1(n15715), .C2(n15449), .A(n12293), .B(n11077), .ZN(
        n11078) );
  AOI21_X1 U13830 ( .B1(n15708), .B2(n11079), .A(n11078), .ZN(n11105) );
  INV_X1 U13831 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11080) );
  XNOR2_X1 U13832 ( .A(n11798), .B(n11080), .ZN(n11103) );
  XNOR2_X1 U13833 ( .A(n15619), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n15620) );
  NAND2_X1 U13834 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15624) );
  INV_X1 U13835 ( .A(n15624), .ZN(n11081) );
  NAND2_X1 U13836 ( .A1(n15620), .A2(n11081), .ZN(n15621) );
  NAND2_X1 U13837 ( .A1(n11082), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U13838 ( .A1(n15621), .A2(n11083), .ZN(n15636) );
  XNOR2_X1 U13839 ( .A(n15639), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n15637) );
  NAND2_X1 U13840 ( .A1(n15636), .A2(n15637), .ZN(n15635) );
  NAND2_X1 U13841 ( .A1(n11084), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U13842 ( .A1(n15635), .A2(n11085), .ZN(n14029) );
  XNOR2_X1 U13843 ( .A(n14031), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n14030) );
  NAND2_X1 U13844 ( .A1(n14029), .A2(n14030), .ZN(n14028) );
  NAND2_X1 U13845 ( .A1(n11086), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U13846 ( .A1(n14028), .A2(n11087), .ZN(n15649) );
  XNOR2_X1 U13847 ( .A(n11088), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n15650) );
  NAND2_X1 U13848 ( .A1(n15649), .A2(n15650), .ZN(n15648) );
  NAND2_X1 U13849 ( .A1(n15654), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11089) );
  NAND2_X1 U13850 ( .A1(n15648), .A2(n11089), .ZN(n14043) );
  XNOR2_X1 U13851 ( .A(n14045), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U13852 ( .A1(n14043), .A2(n14044), .ZN(n14042) );
  NAND2_X1 U13853 ( .A1(n11090), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U13854 ( .A1(n14042), .A2(n11091), .ZN(n14056) );
  INV_X1 U13855 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11092) );
  MUX2_X1 U13856 ( .A(n11092), .B(P2_REG1_REG_6__SCAN_IN), .S(n14058), .Z(
        n14057) );
  NAND2_X1 U13857 ( .A1(n14056), .A2(n14057), .ZN(n14055) );
  OR2_X1 U13858 ( .A1(n14058), .A2(n11092), .ZN(n11093) );
  NAND2_X1 U13859 ( .A1(n14055), .A2(n11093), .ZN(n14071) );
  INV_X1 U13860 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11094) );
  XNOR2_X1 U13861 ( .A(n14074), .B(n11094), .ZN(n14072) );
  NAND2_X1 U13862 ( .A1(n14071), .A2(n14072), .ZN(n14070) );
  NAND2_X1 U13863 ( .A1(n14074), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13864 ( .A1(n14070), .A2(n11095), .ZN(n14082) );
  INV_X1 U13865 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11096) );
  XNOR2_X1 U13866 ( .A(n14084), .B(n11096), .ZN(n14083) );
  NAND2_X1 U13867 ( .A1(n14082), .A2(n14083), .ZN(n15670) );
  INV_X1 U13868 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11098) );
  XNOR2_X1 U13869 ( .A(n15675), .B(n11098), .ZN(n15667) );
  AND2_X1 U13870 ( .A1(n14084), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n15666) );
  NOR2_X1 U13871 ( .A1(n15667), .A2(n15666), .ZN(n11097) );
  NAND2_X1 U13872 ( .A1(n15670), .A2(n11097), .ZN(n15665) );
  NAND2_X1 U13873 ( .A1(n15675), .A2(n11098), .ZN(n11099) );
  NAND2_X1 U13874 ( .A1(n15665), .A2(n11099), .ZN(n11261) );
  XNOR2_X1 U13875 ( .A(n11267), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11262) );
  OR2_X1 U13876 ( .A1(n11261), .A2(n11262), .ZN(n11259) );
  NAND2_X1 U13877 ( .A1(n11267), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U13878 ( .A1(n11259), .A2(n11100), .ZN(n11102) );
  NAND2_X1 U13879 ( .A1(n11102), .A2(n11103), .ZN(n15689) );
  OAI211_X1 U13880 ( .C1(n11103), .C2(n11102), .A(n15690), .B(n15689), .ZN(
        n11104) );
  NAND2_X1 U13881 ( .A1(n11105), .A2(n11104), .ZN(P2_U3225) );
  OAI22_X1 U13882 ( .A1(n13079), .A2(n11441), .B1(n15807), .B2(n13083), .ZN(
        n11106) );
  AOI21_X1 U13883 ( .B1(n13076), .B2(n15798), .A(n11106), .ZN(n11114) );
  INV_X1 U13884 ( .A(n11107), .ZN(n11108) );
  NAND2_X1 U13885 ( .A1(n11108), .A2(n11218), .ZN(n11217) );
  NAND3_X1 U13886 ( .A1(n10442), .A2(n11110), .A3(n12895), .ZN(n11111) );
  OAI211_X1 U13887 ( .C1(n11218), .C2(n15800), .A(n11217), .B(n11111), .ZN(
        n11112) );
  NAND2_X1 U13888 ( .A1(n11112), .A2(n13074), .ZN(n11113) );
  OAI211_X1 U13889 ( .C1(n11226), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        P3_U3162) );
  INV_X1 U13890 ( .A(n11116), .ZN(n11118) );
  INV_X1 U13891 ( .A(SI_18_), .ZN(n11117) );
  OAI222_X1 U13892 ( .A1(P3_U3151), .A2(n11119), .B1(n12160), .B2(n11118), 
        .C1(n11117), .C2(n13838), .ZN(P3_U3277) );
  INV_X1 U13893 ( .A(n11120), .ZN(n11131) );
  INV_X1 U13894 ( .A(n12078), .ZN(n14781) );
  OAI222_X1 U13895 ( .A1(n12946), .A2(n11121), .B1(n15305), .B2(n11131), .C1(
        n14781), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13896 ( .A(n11123), .ZN(n11124) );
  AOI21_X1 U13897 ( .B1(n11125), .B2(n11122), .A(n11124), .ZN(n11130) );
  NAND2_X1 U13898 ( .A1(n14689), .A2(n11126), .ZN(n11201) );
  INV_X1 U13899 ( .A(n14700), .ZN(n14710) );
  INV_X1 U13900 ( .A(n15105), .ZN(n15108) );
  NAND2_X1 U13901 ( .A1(n14746), .A2(n14697), .ZN(n15113) );
  OAI21_X1 U13902 ( .B1(n15108), .B2(n14675), .A(n15113), .ZN(n11127) );
  AOI22_X1 U13903 ( .A1(n11201), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14710), 
        .B2(n11127), .ZN(n11129) );
  NAND2_X1 U13904 ( .A1(n14714), .A2(n15117), .ZN(n11128) );
  OAI211_X1 U13905 ( .C1(n11130), .C2(n14717), .A(n11129), .B(n11128), .ZN(
        P1_U3222) );
  INV_X1 U13906 ( .A(n14143), .ZN(n11133) );
  OAI222_X1 U13907 ( .A1(P2_U3088), .A2(n11133), .B1(n14562), .B2(n11132), 
        .C1(n12913), .C2(n11131), .ZN(P2_U3311) );
  XNOR2_X1 U13908 ( .A(n11285), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11138) );
  INV_X1 U13909 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11136) );
  AOI21_X1 U13910 ( .B1(n11138), .B2(n11137), .A(n11282), .ZN(n11147) );
  NAND2_X1 U13911 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12222)
         );
  OAI21_X1 U13912 ( .B1(n15483), .B2(n6955), .A(n12222), .ZN(n11145) );
  AOI22_X1 U13913 ( .A1(n11141), .A2(n11140), .B1(n11139), .B2(
        P1_REG2_REG_10__SCAN_IN), .ZN(n11143) );
  MUX2_X1 U13914 ( .A(n12276), .B(P1_REG2_REG_11__SCAN_IN), .S(n11285), .Z(
        n11142) );
  AOI211_X1 U13915 ( .C1(n11143), .C2(n11142), .A(n14805), .B(n11284), .ZN(
        n11144) );
  AOI211_X1 U13916 ( .C1(n15475), .C2(n11285), .A(n11145), .B(n11144), .ZN(
        n11146) );
  OAI21_X1 U13917 ( .B1(n11147), .B2(n14817), .A(n11146), .ZN(P1_U3254) );
  INV_X1 U13918 ( .A(P1_U4016), .ZN(n14733) );
  NAND2_X1 U13919 ( .A1(n14733), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n11148) );
  OAI21_X1 U13920 ( .B1(n14612), .B2(n14733), .A(n11148), .ZN(P1_U3582) );
  INV_X1 U13921 ( .A(n13313), .ZN(n13229) );
  AND3_X1 U13922 ( .A1(n11151), .A2(n11150), .A3(n11149), .ZN(n11152) );
  OAI21_X1 U13923 ( .B1(n11153), .B2(n11152), .A(n13300), .ZN(n11161) );
  AND3_X1 U13924 ( .A1(n11156), .A2(n11155), .A3(n11154), .ZN(n11157) );
  OAI21_X1 U13925 ( .B1(n11158), .B2(n11157), .A(n13290), .ZN(n11160) );
  AND2_X1 U13926 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11245) );
  AOI21_X1 U13927 ( .B1(n15779), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11245), .ZN(
        n11159) );
  NAND3_X1 U13928 ( .A1(n11161), .A2(n11160), .A3(n11159), .ZN(n11168) );
  INV_X1 U13929 ( .A(n11345), .ZN(n11166) );
  NAND3_X1 U13930 ( .A1(n11164), .A2(n11163), .A3(n11162), .ZN(n11165) );
  AOI21_X1 U13931 ( .B1(n11166), .B2(n11165), .A(n13282), .ZN(n11167) );
  AOI211_X1 U13932 ( .C1(n13229), .C2(n11169), .A(n11168), .B(n11167), .ZN(
        n11170) );
  INV_X1 U13933 ( .A(n11170), .ZN(P3_U3186) );
  INV_X1 U13934 ( .A(n14714), .ZN(n14681) );
  XOR2_X1 U13935 ( .A(n11172), .B(n11171), .Z(n11177) );
  NAND2_X1 U13936 ( .A1(n11177), .A2(n14685), .ZN(n11174) );
  NOR2_X1 U13937 ( .A1(n10301), .A2(n14706), .ZN(n15544) );
  AOI22_X1 U13938 ( .A1(n11201), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n15544), 
        .B2(n14710), .ZN(n11173) );
  OAI211_X1 U13939 ( .C1(n14681), .C2(n15525), .A(n11174), .B(n11173), .ZN(
        P1_U3232) );
  MUX2_X1 U13940 ( .A(n11177), .B(n11176), .S(n11175), .Z(n11178) );
  NOR2_X1 U13941 ( .A1(n11178), .A2(n8811), .ZN(n11179) );
  AOI211_X1 U13942 ( .C1(n11181), .C2(n11180), .A(n14733), .B(n11179), .ZN(
        n14748) );
  NAND2_X1 U13943 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U13944 ( .A1(n14768), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n11182) );
  OAI211_X1 U13945 ( .C1(n14765), .C2(n11183), .A(n11378), .B(n11182), .ZN(
        n11192) );
  XNOR2_X1 U13946 ( .A(n11185), .B(n11184), .ZN(n11190) );
  OAI211_X1 U13947 ( .C1(n11188), .C2(n11187), .A(n15478), .B(n11186), .ZN(
        n11189) );
  OAI21_X1 U13948 ( .B1(n14805), .B2(n11190), .A(n11189), .ZN(n11191) );
  OR3_X1 U13949 ( .A1(n14748), .A2(n11192), .A3(n11191), .ZN(P1_U3247) );
  OAI222_X1 U13950 ( .A1(n13836), .A2(n11194), .B1(P3_U3151), .B2(n13312), 
        .C1(n11193), .C2(n13838), .ZN(P3_U3276) );
  OAI21_X1 U13951 ( .B1(n11197), .B2(n11195), .A(n11196), .ZN(n11198) );
  NAND2_X1 U13952 ( .A1(n11198), .A2(n14685), .ZN(n11203) );
  NAND2_X1 U13953 ( .A1(n14747), .A2(n15111), .ZN(n11200) );
  NAND2_X1 U13954 ( .A1(n14745), .A2(n14697), .ZN(n11199) );
  NAND2_X1 U13955 ( .A1(n11200), .A2(n11199), .ZN(n15554) );
  AOI22_X1 U13956 ( .A1(n11201), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14710), 
        .B2(n15554), .ZN(n11202) );
  OAI211_X1 U13957 ( .C1(n11204), .C2(n14681), .A(n11203), .B(n11202), .ZN(
        P1_U3237) );
  INV_X1 U13958 ( .A(n11205), .ZN(n11207) );
  OAI222_X1 U13959 ( .A1(P2_U3088), .A2(n11806), .B1(n14562), .B2(n11206), 
        .C1(n12913), .C2(n11207), .ZN(P2_U3313) );
  INV_X1 U13960 ( .A(n12076), .ZN(n11688) );
  OAI222_X1 U13961 ( .A1(P1_U3086), .A2(n11688), .B1(n15307), .B2(n11208), 
        .C1(n15305), .C2(n11207), .ZN(P1_U3341) );
  OAI211_X1 U13962 ( .C1(n11210), .C2(n11209), .A(n8317), .B(n14685), .ZN(
        n11215) );
  INV_X1 U13963 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U13964 ( .A1(n14746), .A2(n15111), .ZN(n11212) );
  NAND2_X1 U13965 ( .A1(n14744), .A2(n14697), .ZN(n11211) );
  AND2_X1 U13966 ( .A1(n11212), .A2(n11211), .ZN(n15505) );
  OAI22_X1 U13967 ( .A1(n15505), .A2(n14700), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14764), .ZN(n11213) );
  AOI21_X1 U13968 ( .B1(n14698), .B2(n14764), .A(n11213), .ZN(n11214) );
  OAI211_X1 U13969 ( .C1(n12685), .C2(n14681), .A(n11215), .B(n11214), .ZN(
        P1_U3218) );
  INV_X1 U13970 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11225) );
  XNOR2_X1 U13971 ( .A(n11216), .B(n15797), .ZN(n11220) );
  OAI21_X1 U13972 ( .B1(n11218), .B2(n13127), .A(n11217), .ZN(n11219) );
  NAND2_X1 U13973 ( .A1(n11219), .A2(n11220), .ZN(n11297) );
  OAI21_X1 U13974 ( .B1(n11220), .B2(n11219), .A(n11297), .ZN(n11221) );
  NAND2_X1 U13975 ( .A1(n11221), .A2(n13074), .ZN(n11224) );
  OAI22_X1 U13976 ( .A1(n13079), .A2(n15784), .B1(n15790), .B2(n13083), .ZN(
        n11222) );
  AOI21_X1 U13977 ( .B1(n13076), .B2(n13127), .A(n11222), .ZN(n11223) );
  OAI211_X1 U13978 ( .C1(n11226), .C2(n11225), .A(n11224), .B(n11223), .ZN(
        P3_U3177) );
  OAI21_X1 U13979 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11227), .A(n13151), .ZN(
        n11241) );
  INV_X1 U13980 ( .A(n13132), .ZN(n11230) );
  NAND3_X1 U13981 ( .A1(n11230), .A2(n11229), .A3(n11228), .ZN(n11231) );
  AOI21_X1 U13982 ( .B1(n11232), .B2(n11231), .A(n13282), .ZN(n11240) );
  OAI21_X1 U13983 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11233), .A(n13156), .ZN(
        n11234) );
  NAND2_X1 U13984 ( .A1(n11234), .A2(n13300), .ZN(n11237) );
  NOR2_X1 U13985 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7300), .ZN(n11235) );
  AOI21_X1 U13986 ( .B1(n15779), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11235), .ZN(
        n11236) );
  OAI211_X1 U13987 ( .C1(n13313), .C2(n11238), .A(n11237), .B(n11236), .ZN(
        n11239) );
  AOI211_X1 U13988 ( .C1(n13290), .C2(n11241), .A(n11240), .B(n11239), .ZN(
        n11242) );
  INV_X1 U13989 ( .A(n11242), .ZN(P3_U3189) );
  INV_X1 U13990 ( .A(n13076), .ZN(n13030) );
  OAI22_X1 U13991 ( .A1(n15784), .A2(n13030), .B1(n13079), .B2(n11243), .ZN(
        n11244) );
  AOI211_X1 U13992 ( .C1(n13098), .C2(n11509), .A(n11245), .B(n11244), .ZN(
        n11250) );
  NAND2_X1 U13993 ( .A1(n11248), .A2(n13074), .ZN(n11249) );
  OAI211_X1 U13994 ( .C1(n11510), .C2(n13088), .A(n11250), .B(n11249), .ZN(
        P3_U3170) );
  INV_X1 U13995 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11255) );
  AND2_X1 U13996 ( .A1(n11251), .A2(n15806), .ZN(n11253) );
  AND2_X1 U13997 ( .A1(n13127), .A2(n15796), .ZN(n11252) );
  AOI21_X1 U13998 ( .B1(n11254), .B2(n11253), .A(n11252), .ZN(n11356) );
  MUX2_X1 U13999 ( .A(n11255), .B(n11356), .S(n15860), .Z(n11256) );
  OAI21_X1 U14000 ( .B1(n13815), .B2(n11358), .A(n11256), .ZN(P3_U3390) );
  INV_X1 U14001 ( .A(n11257), .ZN(n11307) );
  INV_X1 U14002 ( .A(n15476), .ZN(n12077) );
  OAI222_X1 U14003 ( .A1(n15307), .A2(n11258), .B1(n15305), .B2(n11307), .C1(
        n12077), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U14004 ( .A(n11259), .ZN(n11260) );
  AOI211_X1 U14005 ( .C1(n11262), .C2(n11261), .A(n11260), .B(n15701), .ZN(
        n11272) );
  INV_X1 U14006 ( .A(n11263), .ZN(n11264) );
  AOI211_X1 U14007 ( .C1(n11266), .C2(n11265), .A(n14161), .B(n11264), .ZN(
        n11271) );
  NAND2_X1 U14008 ( .A1(n15634), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14009 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11995)
         );
  NAND2_X1 U14010 ( .A1(n15707), .A2(n11267), .ZN(n11268) );
  NAND3_X1 U14011 ( .A1(n11269), .A2(n11995), .A3(n11268), .ZN(n11270) );
  OR3_X1 U14012 ( .A1(n11272), .A2(n11271), .A3(n11270), .ZN(P2_U3224) );
  NAND2_X1 U14013 ( .A1(n13290), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11274) );
  NAND2_X1 U14014 ( .A1(n13300), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11273) );
  OAI211_X1 U14015 ( .C1(n13282), .C2(n11276), .A(n11274), .B(n11273), .ZN(
        n11275) );
  INV_X1 U14016 ( .A(n11275), .ZN(n11279) );
  NAND3_X1 U14017 ( .A1(n13293), .A2(n13282), .A3(n13319), .ZN(n11277) );
  AOI21_X1 U14018 ( .B1(n11277), .B2(n11276), .A(n13229), .ZN(n11278) );
  MUX2_X1 U14019 ( .A(n11279), .B(n11278), .S(P3_IR_REG_0__SCAN_IN), .Z(n11281) );
  AOI22_X1 U14020 ( .A1(n15779), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11280) );
  NAND2_X1 U14021 ( .A1(n11281), .A2(n11280), .ZN(P3_U3182) );
  XNOR2_X1 U14022 ( .A(n11460), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n11456) );
  AOI21_X1 U14023 ( .B1(n11283), .B2(n7019), .A(n11282), .ZN(n11457) );
  XOR2_X1 U14024 ( .A(n11456), .B(n11457), .Z(n11293) );
  MUX2_X1 U14025 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12312), .S(n11460), .Z(
        n11287) );
  OAI21_X1 U14026 ( .B1(n11287), .B2(n11286), .A(n11466), .ZN(n11291) );
  NAND2_X1 U14027 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12258)
         );
  NAND2_X1 U14028 ( .A1(n14768), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11288) );
  OAI211_X1 U14029 ( .C1(n14765), .C2(n11289), .A(n12258), .B(n11288), .ZN(
        n11290) );
  AOI21_X1 U14030 ( .B1(n11291), .B2(n15479), .A(n11290), .ZN(n11292) );
  OAI21_X1 U14031 ( .B1(n11293), .B2(n14817), .A(n11292), .ZN(P1_U3255) );
  XNOR2_X1 U14032 ( .A(n11294), .B(n13126), .ZN(n11296) );
  AOI21_X1 U14033 ( .B1(n11297), .B2(n11295), .A(n11296), .ZN(n11304) );
  NAND3_X1 U14034 ( .A1(n11297), .A2(n11296), .A3(n11295), .ZN(n11298) );
  NAND2_X1 U14035 ( .A1(n11298), .A2(n13074), .ZN(n11303) );
  OAI22_X1 U14036 ( .A1(n13079), .A2(n11440), .B1(n13083), .B2(n11299), .ZN(
        n11301) );
  MUX2_X1 U14037 ( .A(n13094), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11300) );
  AOI211_X1 U14038 ( .C1(n13076), .C2(n15797), .A(n11301), .B(n11300), .ZN(
        n11302) );
  OAI21_X1 U14039 ( .B1(n11304), .B2(n11303), .A(n11302), .ZN(P3_U3158) );
  INV_X1 U14040 ( .A(n11305), .ZN(n11322) );
  INV_X1 U14041 ( .A(n14787), .ZN(n14797) );
  OAI222_X1 U14042 ( .A1(n12946), .A2(n11306), .B1(n15305), .B2(n11322), .C1(
        n14797), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U14043 ( .A1(P2_U3088), .A2(n11808), .B1(n14562), .B2(n11308), 
        .C1(n12913), .C2(n11307), .ZN(P2_U3312) );
  INV_X1 U14044 ( .A(n11309), .ZN(n11359) );
  AOI22_X1 U14045 ( .A1(n14809), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15299), .ZN(n11310) );
  OAI21_X1 U14046 ( .B1(n11359), .B2(n15305), .A(n11310), .ZN(P1_U3337) );
  NAND2_X1 U14047 ( .A1(n11311), .A2(n13817), .ZN(n11313) );
  INV_X1 U14048 ( .A(n11356), .ZN(n11317) );
  AOI21_X1 U14049 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15812), .A(n11317), .ZN(
        n11319) );
  MUX2_X1 U14050 ( .A(n11320), .B(n11319), .S(n15813), .Z(n11321) );
  OAI21_X1 U14051 ( .B1(n11358), .B2(n13534), .A(n11321), .ZN(P3_U3233) );
  INV_X1 U14052 ( .A(n15706), .ZN(n11324) );
  OAI222_X1 U14053 ( .A1(P2_U3088), .A2(n11324), .B1(n14562), .B2(n11323), 
        .C1(n12913), .C2(n11322), .ZN(P2_U3310) );
  OAI21_X1 U14054 ( .B1(n11327), .B2(n11326), .A(n11325), .ZN(n11333) );
  NAND2_X1 U14055 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15647) );
  NAND2_X1 U14056 ( .A1(n13998), .A2(n12396), .ZN(n11328) );
  OAI211_X1 U14057 ( .C1(n13993), .C2(n11595), .A(n15647), .B(n11328), .ZN(
        n11332) );
  INV_X1 U14058 ( .A(n13952), .ZN(n13890) );
  NAND2_X1 U14059 ( .A1(n13890), .A2(n14376), .ZN(n13995) );
  OAI22_X1 U14060 ( .A1(n13995), .A2(n11330), .B1(n13991), .B2(n11329), .ZN(
        n11331) );
  AOI211_X1 U14061 ( .C1(n13986), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        n11334) );
  INV_X1 U14062 ( .A(n11334), .ZN(P2_U3202) );
  AOI22_X1 U14063 ( .A1(n15690), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15708), .ZN(n11337) );
  INV_X1 U14064 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11669) );
  INV_X1 U14065 ( .A(n15707), .ZN(n15696) );
  OAI21_X1 U14066 ( .B1(n15701), .B2(P2_REG1_REG_0__SCAN_IN), .A(n15696), .ZN(
        n11335) );
  AOI21_X1 U14067 ( .B1(n15708), .B2(n11669), .A(n11335), .ZN(n11336) );
  MUX2_X1 U14068 ( .A(n11337), .B(n11336), .S(P2_IR_REG_0__SCAN_IN), .Z(n11339) );
  AOI22_X1 U14069 ( .A1(n15634), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11338) );
  NAND2_X1 U14070 ( .A1(n11339), .A2(n11338), .ZN(P2_U3214) );
  INV_X1 U14071 ( .A(n11340), .ZN(n11342) );
  INV_X1 U14072 ( .A(n13142), .ZN(n11341) );
  AOI21_X1 U14073 ( .B1(n11545), .B2(n11342), .A(n11341), .ZN(n11355) );
  INV_X1 U14074 ( .A(n13130), .ZN(n11347) );
  NOR3_X1 U14075 ( .A1(n11345), .A2(n11344), .A3(n11343), .ZN(n11346) );
  OAI21_X1 U14076 ( .B1(n11347), .B2(n11346), .A(n13315), .ZN(n11354) );
  OAI21_X1 U14077 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11348), .A(n13138), .ZN(
        n11352) );
  NAND2_X1 U14078 ( .A1(n13229), .A2(n11349), .ZN(n11350) );
  NAND2_X1 U14079 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n11366) );
  OAI211_X1 U14080 ( .C1(n7363), .C2(n13227), .A(n11350), .B(n11366), .ZN(
        n11351) );
  AOI21_X1 U14081 ( .B1(n11352), .B2(n13290), .A(n11351), .ZN(n11353) );
  OAI211_X1 U14082 ( .C1(n11355), .C2(n13293), .A(n11354), .B(n11353), .ZN(
        P3_U3187) );
  MUX2_X1 U14083 ( .A(n9460), .B(n11356), .S(n15873), .Z(n11357) );
  OAI21_X1 U14084 ( .B1(n13750), .B2(n11358), .A(n11357), .ZN(P3_U3459) );
  INV_X1 U14085 ( .A(n14147), .ZN(n14144) );
  OAI222_X1 U14086 ( .A1(P2_U3088), .A2(n14144), .B1(n14562), .B2(n11360), 
        .C1(n12913), .C2(n11359), .ZN(P2_U3309) );
  INV_X1 U14087 ( .A(n11518), .ZN(n11370) );
  OAI21_X1 U14088 ( .B1(n11363), .B2(n11362), .A(n11361), .ZN(n11364) );
  NAND2_X1 U14089 ( .A1(n11364), .A2(n13074), .ZN(n11369) );
  AOI22_X1 U14090 ( .A1(n11365), .A2(n15799), .B1(n15796), .B2(n13124), .ZN(
        n11404) );
  INV_X1 U14091 ( .A(n13086), .ZN(n13096) );
  OAI21_X1 U14092 ( .B1(n11404), .B2(n13096), .A(n11366), .ZN(n11367) );
  AOI21_X1 U14093 ( .B1(n11519), .B2(n13098), .A(n11367), .ZN(n11368) );
  OAI211_X1 U14094 ( .C1(n11370), .C2(n13088), .A(n11369), .B(n11368), .ZN(
        P3_U3167) );
  NAND2_X1 U14095 ( .A1(n11371), .A2(n11372), .ZN(n11374) );
  XNOR2_X1 U14096 ( .A(n11374), .B(n11373), .ZN(n11381) );
  NAND2_X1 U14097 ( .A1(n14745), .A2(n15111), .ZN(n11376) );
  NAND2_X1 U14098 ( .A1(n14743), .A2(n14697), .ZN(n11375) );
  NAND2_X1 U14099 ( .A1(n11376), .A2(n11375), .ZN(n11963) );
  NAND2_X1 U14100 ( .A1(n14710), .A2(n11963), .ZN(n11377) );
  OAI211_X1 U14101 ( .C1(n14712), .C2(n11965), .A(n11378), .B(n11377), .ZN(
        n11379) );
  AOI21_X1 U14102 ( .B1(n14714), .B2(n15569), .A(n11379), .ZN(n11380) );
  OAI21_X1 U14103 ( .B1(n11381), .B2(n14717), .A(n11380), .ZN(P1_U3230) );
  INV_X1 U14104 ( .A(n11382), .ZN(n11629) );
  OAI21_X1 U14105 ( .B1(n11385), .B2(n11384), .A(n11383), .ZN(n11386) );
  NAND2_X1 U14106 ( .A1(n11386), .A2(n13986), .ZN(n11389) );
  AOI22_X1 U14107 ( .A1(n14376), .A2(n14021), .B1(n14374), .B2(n14019), .ZN(
        n11632) );
  NAND2_X1 U14108 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14039) );
  OAI21_X1 U14109 ( .B1(n13952), .B2(n11632), .A(n14039), .ZN(n11387) );
  AOI21_X1 U14110 ( .B1(n12404), .B2(n13998), .A(n11387), .ZN(n11388) );
  OAI211_X1 U14111 ( .C1(n13993), .C2(n11629), .A(n11389), .B(n11388), .ZN(
        P2_U3199) );
  INV_X1 U14112 ( .A(n11390), .ZN(n11391) );
  OAI21_X1 U14113 ( .B1(n11391), .B2(n13984), .A(n13973), .ZN(n11393) );
  OR2_X1 U14114 ( .A1(n11392), .A2(P2_U3088), .ZN(n13957) );
  AOI22_X1 U14115 ( .A1(n11393), .A2(n11663), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13957), .ZN(n11395) );
  NAND4_X1 U14116 ( .A1(n13986), .A2(n14025), .A3(n11662), .A4(n9166), .ZN(
        n11394) );
  OAI211_X1 U14117 ( .C1(n12380), .C2(n13991), .A(n11395), .B(n11394), .ZN(
        P2_U3204) );
  XOR2_X1 U14118 ( .A(n11396), .B(n11399), .Z(n11513) );
  NAND2_X1 U14119 ( .A1(n11442), .A2(n11437), .ZN(n11443) );
  INV_X1 U14120 ( .A(n11397), .ZN(n11398) );
  NAND2_X1 U14121 ( .A1(n11443), .A2(n11398), .ZN(n11504) );
  NAND2_X1 U14122 ( .A1(n11504), .A2(n11503), .ZN(n11502) );
  AOI21_X1 U14123 ( .B1(n11502), .B2(n11400), .A(n11399), .ZN(n11403) );
  INV_X1 U14124 ( .A(n11401), .ZN(n11402) );
  OAI21_X1 U14125 ( .B1(n11403), .B2(n11402), .A(n15801), .ZN(n11405) );
  NAND2_X1 U14126 ( .A1(n11405), .A2(n11404), .ZN(n11515) );
  AOI21_X1 U14127 ( .B1(n11513), .B2(n15851), .A(n11515), .ZN(n11544) );
  AOI22_X1 U14128 ( .A1(n13759), .A2(n11519), .B1(n15858), .B2(
        P3_REG0_REG_5__SCAN_IN), .ZN(n11406) );
  OAI21_X1 U14129 ( .B1(n11544), .B2(n15858), .A(n11406), .ZN(P3_U3405) );
  INV_X1 U14130 ( .A(n11407), .ZN(n11409) );
  OAI222_X1 U14131 ( .A1(n12630), .A2(P2_U3088), .B1(n12913), .B2(n11409), 
        .C1(n11408), .C2(n14562), .ZN(P2_U3308) );
  OAI222_X1 U14132 ( .A1(n12946), .A2(n11410), .B1(n15305), .B2(n11409), .C1(
        n11828), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U14133 ( .A1(n6648), .A2(n11411), .ZN(n11412) );
  XNOR2_X1 U14134 ( .A(n11413), .B(n11412), .ZN(n11420) );
  OR2_X1 U14135 ( .A1(n12699), .A2(n14706), .ZN(n11415) );
  NAND2_X1 U14136 ( .A1(n14744), .A2(n15111), .ZN(n11414) );
  NAND2_X1 U14137 ( .A1(n11415), .A2(n11414), .ZN(n15491) );
  NAND2_X1 U14138 ( .A1(n14710), .A2(n15491), .ZN(n11416) );
  OAI211_X1 U14139 ( .C1(n14712), .C2(n15493), .A(n11417), .B(n11416), .ZN(
        n11418) );
  AOI21_X1 U14140 ( .B1(n14714), .B2(n15495), .A(n11418), .ZN(n11419) );
  OAI21_X1 U14141 ( .B1(n11420), .B2(n14717), .A(n11419), .ZN(P1_U3227) );
  AOI21_X1 U14142 ( .B1(n11422), .B2(n11421), .A(n6647), .ZN(n11426) );
  OAI22_X1 U14143 ( .A1(n13973), .A2(n11574), .B1(n13991), .B2(n11578), .ZN(
        n11423) );
  AOI21_X1 U14144 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n13957), .A(n11423), .ZN(
        n11425) );
  INV_X1 U14145 ( .A(n13995), .ZN(n13958) );
  NAND2_X1 U14146 ( .A1(n13958), .A2(n14025), .ZN(n11424) );
  OAI211_X1 U14147 ( .C1(n11426), .C2(n13984), .A(n11425), .B(n11424), .ZN(
        P2_U3194) );
  XNOR2_X1 U14148 ( .A(n11428), .B(n11427), .ZN(n11434) );
  NAND2_X1 U14149 ( .A1(n14374), .A2(n14018), .ZN(n11430) );
  NAND2_X1 U14150 ( .A1(n14376), .A2(n14020), .ZN(n11429) );
  AND2_X1 U14151 ( .A1(n11430), .A2(n11429), .ZN(n11476) );
  NAND2_X1 U14152 ( .A1(n13998), .A2(n12420), .ZN(n11431) );
  NAND2_X1 U14153 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14052) );
  OAI211_X1 U14154 ( .C1(n11476), .C2(n13952), .A(n11431), .B(n14052), .ZN(
        n11432) );
  AOI21_X1 U14155 ( .B1(n11550), .B2(n13873), .A(n11432), .ZN(n11433) );
  OAI21_X1 U14156 ( .B1(n11434), .B2(n13984), .A(n11433), .ZN(P2_U3211) );
  NAND2_X1 U14157 ( .A1(n11435), .A2(n11436), .ZN(n11500) );
  INV_X1 U14158 ( .A(n11437), .ZN(n11499) );
  XNOR2_X1 U14159 ( .A(n11500), .B(n11499), .ZN(n15829) );
  INV_X1 U14160 ( .A(n15829), .ZN(n11451) );
  OR2_X1 U14161 ( .A1(n11438), .A2(n11660), .ZN(n15810) );
  INV_X1 U14162 ( .A(n15810), .ZN(n11439) );
  NAND2_X1 U14163 ( .A1(n15813), .A2(n11439), .ZN(n13414) );
  OAI22_X1 U14164 ( .A1(n11441), .A2(n15785), .B1(n11440), .B2(n15783), .ZN(
        n11447) );
  INV_X1 U14165 ( .A(n11442), .ZN(n11445) );
  INV_X1 U14166 ( .A(n11443), .ZN(n11444) );
  AOI211_X1 U14167 ( .C1(n11499), .C2(n11445), .A(n15789), .B(n11444), .ZN(
        n11446) );
  AOI211_X1 U14168 ( .C1(n15829), .C2(n15843), .A(n11447), .B(n11446), .ZN(
        n15826) );
  MUX2_X1 U14169 ( .A(n7134), .B(n15826), .S(n15813), .Z(n11450) );
  AND2_X1 U14170 ( .A1(n11448), .A2(n15836), .ZN(n15828) );
  AOI22_X1 U14171 ( .A1(n11777), .A2(n15828), .B1(n15812), .B2(n7745), .ZN(
        n11449) );
  OAI211_X1 U14172 ( .C1(n11451), .C2(n13414), .A(n11450), .B(n11449), .ZN(
        P3_U3230) );
  INV_X1 U14173 ( .A(SI_20_), .ZN(n11455) );
  INV_X1 U14174 ( .A(n11452), .ZN(n11453) );
  OAI222_X1 U14175 ( .A1(n12918), .A2(n11455), .B1(P3_U3151), .B2(n11454), 
        .C1(n13836), .C2(n11453), .ZN(P3_U3275) );
  XNOR2_X1 U14176 ( .A(n11684), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11459) );
  OAI22_X1 U14177 ( .A1(n11457), .A2(n11456), .B1(n11460), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11458) );
  NOR2_X1 U14178 ( .A1(n11458), .A2(n11459), .ZN(n11683) );
  AOI211_X1 U14179 ( .C1(n11459), .C2(n11458), .A(n14817), .B(n11683), .ZN(
        n11472) );
  INV_X1 U14180 ( .A(n11466), .ZN(n11462) );
  NOR2_X1 U14181 ( .A1(n11460), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11464) );
  MUX2_X1 U14182 ( .A(n11463), .B(P1_REG2_REG_13__SCAN_IN), .S(n11684), .Z(
        n11461) );
  OAI21_X1 U14183 ( .B1(n11462), .B2(n11464), .A(n11461), .ZN(n11467) );
  NOR2_X1 U14184 ( .A1(n11469), .A2(n11463), .ZN(n11679) );
  AOI211_X1 U14185 ( .C1(n11463), .C2(n11469), .A(n11679), .B(n11464), .ZN(
        n11465) );
  AND3_X1 U14186 ( .A1(n11467), .A2(n15479), .A3(n11681), .ZN(n11471) );
  NAND2_X1 U14187 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12301)
         );
  NAND2_X1 U14188 ( .A1(n14768), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11468) );
  OAI211_X1 U14189 ( .C1(n14765), .C2(n11469), .A(n12301), .B(n11468), .ZN(
        n11470) );
  OR3_X1 U14190 ( .A1(n11472), .A2(n11471), .A3(n11470), .ZN(P1_U3256) );
  XOR2_X1 U14191 ( .A(n12599), .B(n11473), .Z(n11557) );
  INV_X1 U14192 ( .A(n11557), .ZN(n11480) );
  INV_X1 U14193 ( .A(n11533), .ZN(n11474) );
  AOI211_X1 U14194 ( .C1(n12420), .C2(n6639), .A(n14380), .B(n11474), .ZN(
        n11554) );
  XNOR2_X1 U14195 ( .A(n11475), .B(n12599), .ZN(n11478) );
  INV_X1 U14196 ( .A(n11476), .ZN(n11477) );
  AOI21_X1 U14197 ( .B1(n11478), .B2(n14379), .A(n11477), .ZN(n11548) );
  INV_X1 U14198 ( .A(n11548), .ZN(n11479) );
  AOI211_X1 U14199 ( .C1(n15764), .C2(n11480), .A(n11554), .B(n11479), .ZN(
        n11483) );
  AOI22_X1 U14200 ( .A1(n12108), .A2(n12420), .B1(n15775), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11481) );
  OAI21_X1 U14201 ( .B1(n11483), .B2(n15775), .A(n11481), .ZN(P2_U3505) );
  AOI22_X1 U14202 ( .A1(n12114), .A2(n12420), .B1(n15765), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n11482) );
  OAI21_X1 U14203 ( .B1(n11483), .B2(n15765), .A(n11482), .ZN(P2_U3448) );
  NAND2_X1 U14204 ( .A1(n6658), .A2(n11484), .ZN(n11485) );
  XNOR2_X1 U14205 ( .A(n11486), .B(n11485), .ZN(n11497) );
  OAI21_X1 U14206 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n11487), .A(n11864), .ZN(
        n11492) );
  NOR2_X1 U14207 ( .A1(n11488), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12044) );
  AOI21_X1 U14208 ( .B1(n15779), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12044), .ZN(
        n11489) );
  OAI21_X1 U14209 ( .B1(n13313), .B2(n11490), .A(n11489), .ZN(n11491) );
  AOI21_X1 U14210 ( .B1(n11492), .B2(n13300), .A(n11491), .ZN(n11496) );
  NOR2_X1 U14211 ( .A1(n11493), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11494) );
  OAI21_X1 U14212 ( .B1(n11494), .B2(n11860), .A(n13290), .ZN(n11495) );
  OAI211_X1 U14213 ( .C1(n11497), .C2(n13282), .A(n11496), .B(n11495), .ZN(
        P3_U3191) );
  AOI21_X1 U14214 ( .B1(n11500), .B2(n11499), .A(n11498), .ZN(n11501) );
  XOR2_X1 U14215 ( .A(n11503), .B(n11501), .Z(n15831) );
  AOI22_X1 U14216 ( .A1(n13126), .A2(n15799), .B1(n15796), .B2(n13125), .ZN(
        n11506) );
  OAI211_X1 U14217 ( .C1(n11504), .C2(n11503), .A(n11502), .B(n15801), .ZN(
        n11505) );
  OAI211_X1 U14218 ( .C1(n15831), .C2(n15805), .A(n11506), .B(n11505), .ZN(
        n15832) );
  INV_X1 U14219 ( .A(n15832), .ZN(n11507) );
  MUX2_X1 U14220 ( .A(n11508), .B(n11507), .S(n15813), .Z(n11512) );
  AND2_X1 U14221 ( .A1(n11509), .A2(n15836), .ZN(n15833) );
  AOI22_X1 U14222 ( .A1(n11777), .A2(n15833), .B1(n15812), .B2(n9510), .ZN(
        n11511) );
  OAI211_X1 U14223 ( .C1(n15831), .C2(n13414), .A(n11512), .B(n11511), .ZN(
        P3_U3229) );
  INV_X1 U14224 ( .A(n11513), .ZN(n11522) );
  NAND2_X1 U14225 ( .A1(n15805), .A2(n15810), .ZN(n11514) );
  INV_X1 U14226 ( .A(n11515), .ZN(n11516) );
  MUX2_X1 U14227 ( .A(n11517), .B(n11516), .S(n15813), .Z(n11521) );
  INV_X1 U14228 ( .A(n13534), .ZN(n13410) );
  AOI22_X1 U14229 ( .A1(n13410), .A2(n11519), .B1(n15812), .B2(n11518), .ZN(
        n11520) );
  OAI211_X1 U14230 ( .C1(n11522), .C2(n13528), .A(n11521), .B(n11520), .ZN(
        P3_U3228) );
  INV_X1 U14231 ( .A(n11621), .ZN(n11529) );
  OAI211_X1 U14232 ( .C1(n11525), .C2(n11524), .A(n11523), .B(n13074), .ZN(
        n11528) );
  AOI22_X1 U14233 ( .A1(n13123), .A2(n15796), .B1(n15799), .B2(n13125), .ZN(
        n11617) );
  NAND2_X1 U14234 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n13133) );
  OAI21_X1 U14235 ( .B1(n13096), .B2(n11617), .A(n13133), .ZN(n11526) );
  AOI21_X1 U14236 ( .B1(n13098), .B2(n15837), .A(n11526), .ZN(n11527) );
  OAI211_X1 U14237 ( .C1(n11529), .C2(n13088), .A(n11528), .B(n11527), .ZN(
        P3_U3179) );
  OAI21_X1 U14238 ( .B1(n11531), .B2(n11534), .A(n11530), .ZN(n11558) );
  INV_X1 U14239 ( .A(n11738), .ZN(n11532) );
  AOI211_X1 U14240 ( .C1(n12428), .C2(n11533), .A(n14380), .B(n11532), .ZN(
        n11565) );
  XNOR2_X1 U14241 ( .A(n11535), .B(n11534), .ZN(n11536) );
  AOI22_X1 U14242 ( .A1(n14376), .A2(n14019), .B1(n14374), .B2(n14017), .ZN(
        n11695) );
  OAI21_X1 U14243 ( .B1(n11536), .B2(n14302), .A(n11695), .ZN(n11559) );
  AOI211_X1 U14244 ( .C1(n15764), .C2(n11558), .A(n11565), .B(n11559), .ZN(
        n11539) );
  AOI22_X1 U14245 ( .A1(n12108), .A2(n12428), .B1(n15775), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11537) );
  OAI21_X1 U14246 ( .B1(n11539), .B2(n15775), .A(n11537), .ZN(P2_U3506) );
  AOI22_X1 U14247 ( .A1(n12114), .A2(n12428), .B1(n15765), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n11538) );
  OAI21_X1 U14248 ( .B1(n11539), .B2(n15765), .A(n11538), .ZN(P2_U3451) );
  INV_X1 U14249 ( .A(n11540), .ZN(n11542) );
  OAI222_X1 U14250 ( .A1(P2_U3088), .A2(n12626), .B1(n14562), .B2(n11541), 
        .C1(n12913), .C2(n11542), .ZN(P2_U3307) );
  OAI222_X1 U14251 ( .A1(n12946), .A2(n11543), .B1(P1_U3086), .B2(n15526), 
        .C1(n15305), .C2(n11542), .ZN(P1_U3335) );
  MUX2_X1 U14252 ( .A(n11545), .B(n11544), .S(n15873), .Z(n11546) );
  OAI21_X1 U14253 ( .B1(n13750), .B2(n11547), .A(n11546), .ZN(P3_U3464) );
  MUX2_X1 U14254 ( .A(n11549), .B(n11548), .S(n14396), .Z(n11556) );
  INV_X1 U14255 ( .A(n11550), .ZN(n11551) );
  OAI22_X1 U14256 ( .A1(n14368), .A2(n11552), .B1(n14385), .B2(n11551), .ZN(
        n11553) );
  AOI21_X1 U14257 ( .B1(n14399), .B2(n11554), .A(n11553), .ZN(n11555) );
  OAI211_X1 U14258 ( .C1(n11557), .C2(n14371), .A(n11556), .B(n11555), .ZN(
        P2_U3259) );
  INV_X1 U14259 ( .A(n11558), .ZN(n11568) );
  INV_X1 U14260 ( .A(n11559), .ZN(n11560) );
  MUX2_X1 U14261 ( .A(n11561), .B(n11560), .S(n14396), .Z(n11567) );
  INV_X1 U14262 ( .A(n12428), .ZN(n11563) );
  INV_X1 U14263 ( .A(n11697), .ZN(n11562) );
  OAI22_X1 U14264 ( .A1(n14368), .A2(n11563), .B1(n11562), .B2(n14385), .ZN(
        n11564) );
  AOI21_X1 U14265 ( .B1(n11565), .B2(n14399), .A(n11564), .ZN(n11566) );
  OAI211_X1 U14266 ( .C1(n11568), .C2(n14371), .A(n11567), .B(n11566), .ZN(
        P2_U3258) );
  NAND2_X1 U14267 ( .A1(n11570), .A2(n14273), .ZN(n11571) );
  NOR2_X1 U14268 ( .A1(n11572), .A2(n11571), .ZN(n15733) );
  AOI22_X1 U14269 ( .A1(n14399), .A2(n15733), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14397), .ZN(n11573) );
  OAI21_X1 U14270 ( .B1(n11574), .B2(n14368), .A(n11573), .ZN(n11575) );
  INV_X1 U14271 ( .A(n11575), .ZN(n11585) );
  INV_X1 U14272 ( .A(n14025), .ZN(n11579) );
  OAI22_X1 U14273 ( .A1(n11579), .A2(n14329), .B1(n14331), .B2(n11578), .ZN(
        n11581) );
  NOR2_X1 U14274 ( .A1(n15736), .A2(n14337), .ZN(n11580) );
  AOI211_X1 U14275 ( .C1(n14379), .C2(n11582), .A(n11581), .B(n11580), .ZN(
        n15735) );
  MUX2_X1 U14276 ( .A(n15735), .B(n11583), .S(n14352), .Z(n11584) );
  OAI211_X1 U14277 ( .C1(n15736), .C2(n14348), .A(n11585), .B(n11584), .ZN(
        P2_U3264) );
  XNOR2_X1 U14278 ( .A(n11586), .B(n12596), .ZN(n15749) );
  NAND3_X1 U14279 ( .A1(n11587), .A2(n11589), .A3(n11588), .ZN(n11590) );
  NAND2_X1 U14280 ( .A1(n11591), .A2(n14379), .ZN(n11593) );
  AOI22_X1 U14281 ( .A1(n14376), .A2(n14022), .B1(n14374), .B2(n14020), .ZN(
        n11592) );
  NAND2_X1 U14282 ( .A1(n11593), .A2(n11592), .ZN(n15753) );
  INV_X1 U14283 ( .A(n14399), .ZN(n14274) );
  AOI21_X1 U14284 ( .B1(n11644), .B2(n12396), .A(n14380), .ZN(n11594) );
  NAND2_X1 U14285 ( .A1(n11594), .A2(n11627), .ZN(n15751) );
  OAI22_X1 U14286 ( .A1(n14274), .A2(n15751), .B1(n11595), .B2(n14385), .ZN(
        n11596) );
  AOI21_X1 U14287 ( .B1(n14352), .B2(P2_REG2_REG_4__SCAN_IN), .A(n11596), .ZN(
        n11597) );
  OAI21_X1 U14288 ( .B1(n7888), .B2(n14368), .A(n11597), .ZN(n11598) );
  AOI21_X1 U14289 ( .B1(n14396), .B2(n15753), .A(n11598), .ZN(n11599) );
  OAI21_X1 U14290 ( .B1(n14371), .B2(n15749), .A(n11599), .ZN(P2_U3261) );
  NOR2_X1 U14291 ( .A1(n7366), .A2(n11616), .ZN(n11614) );
  NOR2_X1 U14292 ( .A1(n11614), .A2(n11601), .ZN(n11603) );
  XNOR2_X1 U14293 ( .A(n11603), .B(n11602), .ZN(n11605) );
  OAI22_X1 U14294 ( .A1(n11673), .A2(n15785), .B1(n12042), .B2(n15783), .ZN(
        n11604) );
  AOI21_X1 U14295 ( .B1(n11605), .B2(n15801), .A(n11604), .ZN(n15847) );
  MUX2_X1 U14296 ( .A(n11606), .B(n15847), .S(n15813), .Z(n11610) );
  AND2_X1 U14297 ( .A1(n11607), .A2(n15836), .ZN(n15849) );
  INV_X1 U14298 ( .A(n11608), .ZN(n11676) );
  AOI22_X1 U14299 ( .A1(n11777), .A2(n15849), .B1(n15812), .B2(n11676), .ZN(
        n11609) );
  OAI211_X1 U14300 ( .C1(n15846), .C2(n13528), .A(n11610), .B(n11609), .ZN(
        P3_U3226) );
  NAND2_X1 U14301 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  XOR2_X1 U14302 ( .A(n11616), .B(n11613), .Z(n15840) );
  AOI211_X1 U14303 ( .C1(n11616), .C2(n7366), .A(n15789), .B(n11614), .ZN(
        n11619) );
  INV_X1 U14304 ( .A(n11617), .ZN(n11618) );
  NOR2_X1 U14305 ( .A1(n11619), .A2(n11618), .ZN(n15839) );
  MUX2_X1 U14306 ( .A(n11620), .B(n15839), .S(n15813), .Z(n11623) );
  AOI22_X1 U14307 ( .A1(n13410), .A2(n15837), .B1(n15812), .B2(n11621), .ZN(
        n11622) );
  OAI211_X1 U14308 ( .C1(n13528), .C2(n15840), .A(n11623), .B(n11622), .ZN(
        P3_U3227) );
  AND2_X1 U14309 ( .A1(n11625), .A2(n11624), .ZN(n12597) );
  XNOR2_X1 U14310 ( .A(n11626), .B(n12597), .ZN(n15756) );
  INV_X1 U14311 ( .A(n11627), .ZN(n11628) );
  OAI211_X1 U14312 ( .C1(n15759), .C2(n11628), .A(n6639), .B(n14273), .ZN(
        n15757) );
  OAI22_X1 U14313 ( .A1(n14274), .A2(n15757), .B1(n11629), .B2(n14385), .ZN(
        n11630) );
  AOI21_X1 U14314 ( .B1(n14401), .B2(n12404), .A(n11630), .ZN(n11637) );
  XNOR2_X1 U14315 ( .A(n11631), .B(n12597), .ZN(n11634) );
  INV_X1 U14316 ( .A(n11632), .ZN(n11633) );
  AOI21_X1 U14317 ( .B1(n11634), .B2(n14379), .A(n11633), .ZN(n15760) );
  MUX2_X1 U14318 ( .A(n11635), .B(n15760), .S(n14396), .Z(n11636) );
  OAI211_X1 U14319 ( .C1(n15756), .C2(n14371), .A(n11637), .B(n11636), .ZN(
        P2_U3260) );
  AOI21_X1 U14320 ( .B1(n11640), .B2(n11639), .A(n11638), .ZN(n11642) );
  XNOR2_X1 U14321 ( .A(n11642), .B(n11641), .ZN(n15745) );
  INV_X1 U14322 ( .A(n11643), .ZN(n11646) );
  INV_X1 U14323 ( .A(n11644), .ZN(n11645) );
  AOI211_X1 U14324 ( .C1(n15742), .C2(n11646), .A(n14380), .B(n11645), .ZN(
        n15740) );
  AOI22_X1 U14325 ( .A1(n14401), .A2(n15742), .B1(n15740), .B2(n14399), .ZN(
        n11657) );
  OR2_X1 U14326 ( .A1(n11647), .A2(n12598), .ZN(n11648) );
  NAND2_X1 U14327 ( .A1(n11587), .A2(n11648), .ZN(n11649) );
  NAND2_X1 U14328 ( .A1(n11649), .A2(n14379), .ZN(n15743) );
  NAND2_X1 U14329 ( .A1(n14374), .A2(n14021), .ZN(n11651) );
  NAND2_X1 U14330 ( .A1(n14376), .A2(n14023), .ZN(n11650) );
  NAND2_X1 U14331 ( .A1(n11651), .A2(n11650), .ZN(n15741) );
  AOI21_X1 U14332 ( .B1(n14397), .B2(n11652), .A(n15741), .ZN(n11653) );
  AND2_X1 U14333 ( .A1(n15743), .A2(n11653), .ZN(n11655) );
  MUX2_X1 U14334 ( .A(n11655), .B(n11654), .S(n14352), .Z(n11656) );
  OAI211_X1 U14335 ( .C1(n15745), .C2(n14371), .A(n11657), .B(n11656), .ZN(
        P2_U3262) );
  INV_X1 U14336 ( .A(SI_21_), .ZN(n11661) );
  INV_X1 U14337 ( .A(n11658), .ZN(n11659) );
  OAI222_X1 U14338 ( .A1(n12918), .A2(n11661), .B1(P3_U3151), .B2(n11660), 
        .C1(n13836), .C2(n11659), .ZN(P3_U3274) );
  INV_X1 U14339 ( .A(n14348), .ZN(n11664) );
  OAI21_X1 U14340 ( .B1(n14025), .B2(n11663), .A(n11662), .ZN(n12594) );
  INV_X1 U14341 ( .A(n12594), .ZN(n15731) );
  AOI22_X1 U14342 ( .A1(n11664), .A2(n15731), .B1(n14401), .B2(n11663), .ZN(
        n11668) );
  AOI21_X1 U14343 ( .B1(n14302), .B2(n14337), .A(n12594), .ZN(n11665) );
  AOI21_X1 U14344 ( .B1(n14374), .B2(n14024), .A(n11665), .ZN(n15728) );
  OAI21_X1 U14345 ( .B1(n15727), .B2(n9166), .A(n15728), .ZN(n11666) );
  AOI22_X1 U14346 ( .A1(n14396), .A2(n11666), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14397), .ZN(n11667) );
  OAI211_X1 U14347 ( .C1(n11669), .C2(n14396), .A(n11668), .B(n11667), .ZN(
        P2_U3265) );
  XNOR2_X1 U14348 ( .A(n11671), .B(n11670), .ZN(n11678) );
  OAI22_X1 U14349 ( .A1(n13083), .A2(n11672), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7300), .ZN(n11675) );
  OAI22_X1 U14350 ( .A1(n11673), .A2(n13030), .B1(n13079), .B2(n12042), .ZN(
        n11674) );
  AOI211_X1 U14351 ( .C1(n11676), .C2(n13094), .A(n11675), .B(n11674), .ZN(
        n11677) );
  OAI21_X1 U14352 ( .B1(n11678), .B2(n13100), .A(n11677), .ZN(P3_U3153) );
  INV_X1 U14353 ( .A(n11679), .ZN(n11680) );
  NAND2_X1 U14354 ( .A1(n11681), .A2(n11680), .ZN(n12067) );
  XOR2_X1 U14355 ( .A(n12076), .B(P1_REG2_REG_14__SCAN_IN), .Z(n12066) );
  XNOR2_X1 U14356 ( .A(n12067), .B(n12066), .ZN(n11692) );
  XNOR2_X1 U14357 ( .A(n12076), .B(n11682), .ZN(n11686) );
  AOI21_X1 U14358 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n11684), .A(n11683), 
        .ZN(n11685) );
  NAND2_X1 U14359 ( .A1(n11685), .A2(n11686), .ZN(n12075) );
  OAI21_X1 U14360 ( .B1(n11686), .B2(n11685), .A(n12075), .ZN(n11687) );
  NAND2_X1 U14361 ( .A1(n11687), .A2(n15478), .ZN(n11691) );
  NOR2_X1 U14362 ( .A1(n13679), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14588) );
  NOR2_X1 U14363 ( .A1(n14765), .A2(n11688), .ZN(n11689) );
  AOI211_X1 U14364 ( .C1(n14768), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14588), 
        .B(n11689), .ZN(n11690) );
  OAI211_X1 U14365 ( .C1(n11692), .C2(n14805), .A(n11691), .B(n11690), .ZN(
        P1_U3257) );
  XNOR2_X1 U14366 ( .A(n11693), .B(n11694), .ZN(n11700) );
  OAI22_X1 U14367 ( .A1(n13952), .A2(n11695), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8997), .ZN(n11696) );
  AOI21_X1 U14368 ( .B1(n12428), .B2(n13998), .A(n11696), .ZN(n11699) );
  NAND2_X1 U14369 ( .A1(n13873), .A2(n11697), .ZN(n11698) );
  OAI211_X1 U14370 ( .C1(n11700), .C2(n13984), .A(n11699), .B(n11698), .ZN(
        P2_U3185) );
  INV_X1 U14371 ( .A(n11701), .ZN(n11704) );
  OAI22_X1 U14372 ( .A1(n11702), .A2(P3_U3151), .B1(SI_22_), .B2(n13838), .ZN(
        n11703) );
  AOI21_X1 U14373 ( .B1(n11704), .B2(n11781), .A(n11703), .ZN(P3_U3273) );
  INV_X1 U14374 ( .A(n11705), .ZN(n12909) );
  OAI222_X1 U14375 ( .A1(n12946), .A2(n11706), .B1(n15305), .B2(n12909), .C1(
        n12822), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U14376 ( .A(n11708), .B(n11707), .ZN(n11715) );
  OR2_X1 U14377 ( .A1(n12699), .A2(n14675), .ZN(n11710) );
  NAND2_X1 U14378 ( .A1(n14740), .A2(n14697), .ZN(n11709) );
  NAND2_X1 U14379 ( .A1(n11710), .A2(n11709), .ZN(n15596) );
  NAND2_X1 U14380 ( .A1(n14710), .A2(n15596), .ZN(n11711) );
  OAI211_X1 U14381 ( .C1(n14712), .C2(n11944), .A(n11712), .B(n11711), .ZN(
        n11713) );
  AOI21_X1 U14382 ( .B1(n14714), .B2(n15597), .A(n11713), .ZN(n11714) );
  OAI21_X1 U14383 ( .B1(n11715), .B2(n14717), .A(n11714), .ZN(P1_U3213) );
  NAND2_X1 U14384 ( .A1(n11717), .A2(n11718), .ZN(n12016) );
  NAND3_X1 U14385 ( .A1(n11716), .A2(n12016), .A3(n15604), .ZN(n11724) );
  XNOR2_X1 U14386 ( .A(n11719), .B(n11718), .ZN(n12008) );
  NAND2_X1 U14387 ( .A1(n12008), .A2(n15572), .ZN(n11723) );
  NAND2_X1 U14388 ( .A1(n14739), .A2(n14697), .ZN(n11721) );
  NAND2_X1 U14389 ( .A1(n14741), .A2(n15111), .ZN(n11720) );
  AND2_X1 U14390 ( .A1(n11721), .A2(n11720), .ZN(n12009) );
  OAI211_X1 U14391 ( .C1(n11939), .C2(n11914), .A(n15500), .B(n11722), .ZN(
        n12013) );
  NAND4_X1 U14392 ( .A1(n11724), .A2(n11723), .A3(n12009), .A4(n12013), .ZN(
        n11729) );
  OAI22_X1 U14393 ( .A1(n15228), .A2(n11914), .B1(n15618), .B2(n10921), .ZN(
        n11725) );
  AOI21_X1 U14394 ( .B1(n11729), .B2(n15618), .A(n11725), .ZN(n11726) );
  INV_X1 U14395 ( .A(n11726), .ZN(P1_U3536) );
  INV_X1 U14396 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11727) );
  OAI22_X1 U14397 ( .A1(n15288), .A2(n11914), .B1(n15606), .B2(n11727), .ZN(
        n11728) );
  AOI21_X1 U14398 ( .B1(n11729), .B2(n15606), .A(n11728), .ZN(n11730) );
  INV_X1 U14399 ( .A(n11730), .ZN(P1_U3483) );
  OAI21_X1 U14400 ( .B1(n11732), .B2(n10013), .A(n11731), .ZN(n14512) );
  XNOR2_X1 U14401 ( .A(n11733), .B(n12601), .ZN(n11736) );
  AOI22_X1 U14402 ( .A1(n14376), .A2(n14018), .B1(n14015), .B2(n14374), .ZN(
        n11734) );
  OAI21_X1 U14403 ( .B1(n14512), .B2(n14337), .A(n11734), .ZN(n11735) );
  AOI21_X1 U14404 ( .B1(n14379), .B2(n11736), .A(n11735), .ZN(n14511) );
  MUX2_X1 U14405 ( .A(n11737), .B(n14511), .S(n14396), .Z(n11744) );
  NAND2_X1 U14406 ( .A1(n11738), .A2(n14509), .ZN(n11739) );
  NAND2_X1 U14407 ( .A1(n11739), .A2(n14273), .ZN(n11740) );
  NOR2_X1 U14408 ( .A1(n11762), .A2(n11740), .ZN(n14508) );
  INV_X1 U14409 ( .A(n14509), .ZN(n11851) );
  INV_X1 U14410 ( .A(n11849), .ZN(n11741) );
  OAI22_X1 U14411 ( .A1(n14368), .A2(n11851), .B1(n11741), .B2(n14385), .ZN(
        n11742) );
  AOI21_X1 U14412 ( .B1(n14399), .B2(n14508), .A(n11742), .ZN(n11743) );
  OAI211_X1 U14413 ( .C1(n14512), .C2(n14348), .A(n11744), .B(n11743), .ZN(
        P2_U3257) );
  XNOR2_X1 U14414 ( .A(n11745), .B(n11746), .ZN(n11753) );
  NOR2_X1 U14415 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11747), .ZN(n13160) );
  OAI22_X1 U14416 ( .A1(n13030), .A2(n11749), .B1(n11748), .B2(n13083), .ZN(
        n11750) );
  AOI211_X1 U14417 ( .C1(n13027), .C2(n13121), .A(n13160), .B(n11750), .ZN(
        n11752) );
  NAND2_X1 U14418 ( .A1(n13094), .A2(n11776), .ZN(n11751) );
  OAI211_X1 U14419 ( .C1(n11753), .C2(n13100), .A(n11752), .B(n11751), .ZN(
        P3_U3161) );
  XOR2_X1 U14420 ( .A(n11754), .B(n12604), .Z(n11840) );
  INV_X1 U14421 ( .A(n11840), .ZN(n11769) );
  INV_X1 U14422 ( .A(n11755), .ZN(n11757) );
  INV_X1 U14423 ( .A(n12604), .ZN(n11756) );
  OAI21_X1 U14424 ( .B1(n11757), .B2(n11756), .A(n14379), .ZN(n11760) );
  NOR2_X1 U14425 ( .A1(n11755), .A2(n12604), .ZN(n12024) );
  NAND2_X1 U14426 ( .A1(n14374), .A2(n14014), .ZN(n11759) );
  NAND2_X1 U14427 ( .A1(n14376), .A2(n14017), .ZN(n11758) );
  AND2_X1 U14428 ( .A1(n11759), .A2(n11758), .ZN(n11899) );
  OAI21_X1 U14429 ( .B1(n11760), .B2(n12024), .A(n11899), .ZN(n11838) );
  INV_X1 U14430 ( .A(n11838), .ZN(n11761) );
  MUX2_X1 U14431 ( .A(n11068), .B(n11761), .S(n14396), .Z(n11768) );
  OAI21_X1 U14432 ( .B1(n11762), .B2(n11896), .A(n14273), .ZN(n11764) );
  NOR2_X1 U14433 ( .A1(n11764), .A2(n11763), .ZN(n11839) );
  INV_X1 U14434 ( .A(n11897), .ZN(n11765) );
  OAI22_X1 U14435 ( .A1(n14368), .A2(n11896), .B1(n11765), .B2(n14385), .ZN(
        n11766) );
  AOI21_X1 U14436 ( .B1(n11839), .B2(n14399), .A(n11766), .ZN(n11767) );
  OAI211_X1 U14437 ( .C1(n14371), .C2(n11769), .A(n11768), .B(n11767), .ZN(
        P2_U3256) );
  XNOR2_X1 U14438 ( .A(n11878), .B(n11770), .ZN(n15857) );
  INV_X1 U14439 ( .A(n15857), .ZN(n11780) );
  AOI22_X1 U14440 ( .A1(n15796), .A2(n13121), .B1(n13123), .B2(n15799), .ZN(
        n11771) );
  OAI21_X1 U14441 ( .B1(n11772), .B2(n15789), .A(n11771), .ZN(n11773) );
  AOI21_X1 U14442 ( .B1(n15857), .B2(n15843), .A(n11773), .ZN(n15853) );
  MUX2_X1 U14443 ( .A(n11774), .B(n15853), .S(n15813), .Z(n11779) );
  AND2_X1 U14444 ( .A1(n11775), .A2(n15836), .ZN(n15855) );
  AOI22_X1 U14445 ( .A1(n11777), .A2(n15855), .B1(n11776), .B2(n15812), .ZN(
        n11778) );
  OAI211_X1 U14446 ( .C1(n11780), .C2(n13414), .A(n11779), .B(n11778), .ZN(
        P3_U3225) );
  NAND2_X1 U14447 ( .A1(n11782), .A2(n11781), .ZN(n11784) );
  OAI211_X1 U14448 ( .C1(n11785), .C2(n12918), .A(n11784), .B(n11783), .ZN(
        P3_U3272) );
  INV_X1 U14449 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11786) );
  XNOR2_X1 U14450 ( .A(n14143), .B(n11786), .ZN(n14131) );
  OR2_X1 U14451 ( .A1(n11798), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15680) );
  MUX2_X1 U14452 ( .A(n11788), .B(P2_REG2_REG_12__SCAN_IN), .S(n15695), .Z(
        n15679) );
  NAND2_X1 U14453 ( .A1(n11787), .A2(n15679), .ZN(n15684) );
  NAND2_X1 U14454 ( .A1(n15695), .A2(n11788), .ZN(n11789) );
  INV_X1 U14455 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11790) );
  MUX2_X1 U14456 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11790), .S(n11803), .Z(
        n14093) );
  OR2_X1 U14457 ( .A1(n11803), .A2(n11790), .ZN(n11791) );
  NAND2_X1 U14458 ( .A1(n14108), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11794) );
  INV_X1 U14459 ( .A(n11806), .ZN(n14112) );
  NAND2_X1 U14460 ( .A1(n11792), .A2(n14112), .ZN(n11793) );
  NAND2_X1 U14461 ( .A1(n11794), .A2(n11793), .ZN(n11795) );
  XNOR2_X1 U14462 ( .A(n11795), .B(n11808), .ZN(n14120) );
  NAND2_X1 U14463 ( .A1(n14120), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11797) );
  INV_X1 U14464 ( .A(n11808), .ZN(n14124) );
  NAND2_X1 U14465 ( .A1(n11795), .A2(n14124), .ZN(n11796) );
  XOR2_X1 U14466 ( .A(n14131), .B(n14132), .Z(n11819) );
  NAND2_X1 U14467 ( .A1(n11798), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n15688) );
  XNOR2_X1 U14468 ( .A(n15695), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n15687) );
  AND2_X1 U14469 ( .A1(n15688), .A2(n15687), .ZN(n11799) );
  NAND2_X1 U14470 ( .A1(n15689), .A2(n11799), .ZN(n15686) );
  NAND2_X1 U14471 ( .A1(n15695), .A2(n11800), .ZN(n11801) );
  NAND2_X1 U14472 ( .A1(n15686), .A2(n11801), .ZN(n14101) );
  INV_X1 U14473 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11802) );
  XNOR2_X1 U14474 ( .A(n11803), .B(n11802), .ZN(n14100) );
  INV_X1 U14475 ( .A(n11803), .ZN(n14099) );
  NAND2_X1 U14476 ( .A1(n14099), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U14477 ( .A1(n14103), .A2(n11804), .ZN(n14115) );
  XNOR2_X1 U14478 ( .A(n11806), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U14479 ( .A1(n14115), .A2(n14114), .ZN(n14113) );
  OR2_X1 U14480 ( .A1(n11806), .A2(n11805), .ZN(n11807) );
  NAND2_X1 U14481 ( .A1(n14113), .A2(n11807), .ZN(n11809) );
  XNOR2_X1 U14482 ( .A(n11809), .B(n11808), .ZN(n14126) );
  NAND2_X1 U14483 ( .A1(n14126), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U14484 ( .A1(n11809), .A2(n14124), .ZN(n11810) );
  NAND2_X1 U14485 ( .A1(n14125), .A2(n11810), .ZN(n11813) );
  XNOR2_X1 U14486 ( .A(n14143), .B(n11811), .ZN(n11812) );
  OAI21_X1 U14487 ( .B1(n11813), .B2(n11812), .A(n15690), .ZN(n11817) );
  NAND2_X1 U14488 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13901)
         );
  INV_X1 U14489 ( .A(n13901), .ZN(n11814) );
  AOI21_X1 U14490 ( .B1(n15707), .B2(n14143), .A(n11814), .ZN(n11816) );
  NAND2_X1 U14491 ( .A1(n15634), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n11815) );
  OAI211_X1 U14492 ( .C1(n11817), .C2(n14142), .A(n11816), .B(n11815), .ZN(
        n11818) );
  AOI21_X1 U14493 ( .B1(n11819), .B2(n15708), .A(n11818), .ZN(n11820) );
  INV_X1 U14494 ( .A(n11820), .ZN(P2_U3230) );
  INV_X1 U14495 ( .A(n11821), .ZN(n11822) );
  AOI21_X1 U14496 ( .B1(n11824), .B2(n11823), .A(n11822), .ZN(n15557) );
  NAND2_X1 U14497 ( .A1(n11826), .A2(n11825), .ZN(n14842) );
  NAND2_X1 U14498 ( .A1(n15513), .A2(n15604), .ZN(n15528) );
  INV_X1 U14499 ( .A(n15518), .ZN(n11827) );
  AOI211_X1 U14500 ( .C1(n10303), .C2(n15107), .A(n15517), .B(n11827), .ZN(
        n15553) );
  NOR2_X1 U14501 ( .A1(n15524), .A2(n15526), .ZN(n11829) );
  NAND2_X1 U14502 ( .A1(n15515), .A2(n10303), .ZN(n11831) );
  AOI22_X1 U14503 ( .A1(n15513), .A2(n15554), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15531), .ZN(n11830) );
  OAI211_X1 U14504 ( .C1(n10849), .C2(n15513), .A(n11831), .B(n11830), .ZN(
        n11832) );
  AOI21_X1 U14505 ( .B1(n15553), .B2(n15519), .A(n11832), .ZN(n11837) );
  XNOR2_X1 U14506 ( .A(n14747), .B(n15117), .ZN(n15106) );
  INV_X1 U14507 ( .A(n15106), .ZN(n11834) );
  NOR2_X1 U14508 ( .A1(n14747), .A2(n15117), .ZN(n12679) );
  AOI21_X1 U14509 ( .B1(n11834), .B2(n15104), .A(n12679), .ZN(n11835) );
  XNOR2_X1 U14510 ( .A(n11835), .B(n12829), .ZN(n15560) );
  NAND2_X1 U14511 ( .A1(n15100), .A2(n15560), .ZN(n11836) );
  OAI211_X1 U14512 ( .C1(n15557), .C2(n15528), .A(n11837), .B(n11836), .ZN(
        P1_U3291) );
  AOI211_X1 U14513 ( .C1(n15764), .C2(n11840), .A(n11839), .B(n11838), .ZN(
        n11843) );
  AOI22_X1 U14514 ( .A1(n12114), .A2(n12455), .B1(n15765), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n11841) );
  OAI21_X1 U14515 ( .B1(n11843), .B2(n15765), .A(n11841), .ZN(P2_U3457) );
  AOI22_X1 U14516 ( .A1(n12108), .A2(n12455), .B1(n15775), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11842) );
  OAI21_X1 U14517 ( .B1(n11843), .B2(n15775), .A(n11842), .ZN(P2_U3508) );
  OAI21_X1 U14518 ( .B1(n11846), .B2(n11845), .A(n11844), .ZN(n11854) );
  OAI22_X1 U14519 ( .A1(n13995), .A2(n11848), .B1(n13991), .B2(n11847), .ZN(
        n11853) );
  NAND2_X1 U14520 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14079) );
  NAND2_X1 U14521 ( .A1(n13873), .A2(n11849), .ZN(n11850) );
  OAI211_X1 U14522 ( .C1(n13973), .C2(n11851), .A(n14079), .B(n11850), .ZN(
        n11852) );
  AOI211_X1 U14523 ( .C1(n11854), .C2(n13986), .A(n11853), .B(n11852), .ZN(
        n11855) );
  INV_X1 U14524 ( .A(n11855), .ZN(P2_U3193) );
  XNOR2_X1 U14525 ( .A(n11857), .B(n11856), .ZN(n11872) );
  OR3_X1 U14526 ( .A1(n11860), .A2(n11859), .A3(n11858), .ZN(n11861) );
  AOI21_X1 U14527 ( .B1(n11862), .B2(n11861), .A(n13319), .ZN(n11871) );
  AND3_X1 U14528 ( .A1(n11864), .A2(n11863), .A3(n6489), .ZN(n11865) );
  OAI21_X1 U14529 ( .B1(n11866), .B2(n11865), .A(n13300), .ZN(n11868) );
  AND2_X1 U14530 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11986) );
  AOI21_X1 U14531 ( .B1(n15779), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11986), 
        .ZN(n11867) );
  OAI211_X1 U14532 ( .C1(n13313), .C2(n11869), .A(n11868), .B(n11867), .ZN(
        n11870) );
  AOI211_X1 U14533 ( .C1(n13315), .C2(n11872), .A(n11871), .B(n11870), .ZN(
        n11873) );
  INV_X1 U14534 ( .A(n11873), .ZN(P3_U3192) );
  INV_X1 U14535 ( .A(n11874), .ZN(n11876) );
  OAI222_X1 U14536 ( .A1(P2_U3088), .A2(n12625), .B1(n12913), .B2(n11876), 
        .C1(n11875), .C2(n14562), .ZN(P2_U3305) );
  OR2_X1 U14537 ( .A1(n11878), .A2(n11877), .ZN(n11880) );
  NAND2_X1 U14538 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14539 ( .A(n11881), .B(n6895), .ZN(n11890) );
  INV_X1 U14540 ( .A(n11890), .ZN(n11919) );
  OR2_X1 U14541 ( .A1(n11884), .A2(n11883), .ZN(n11973) );
  NAND2_X1 U14542 ( .A1(n11884), .A2(n11883), .ZN(n11885) );
  NAND2_X1 U14543 ( .A1(n11973), .A2(n11885), .ZN(n11886) );
  NAND2_X1 U14544 ( .A1(n11886), .A2(n15801), .ZN(n11888) );
  AOI22_X1 U14545 ( .A1(n15799), .A2(n13122), .B1(n13120), .B2(n15796), .ZN(
        n11887) );
  NAND2_X1 U14546 ( .A1(n11888), .A2(n11887), .ZN(n11889) );
  AOI21_X1 U14547 ( .B1(n15843), .B2(n11890), .A(n11889), .ZN(n11915) );
  OAI21_X1 U14548 ( .B1(n11919), .B2(n15841), .A(n11915), .ZN(n11891) );
  INV_X1 U14549 ( .A(n11891), .ZN(n12104) );
  INV_X1 U14550 ( .A(n12107), .ZN(n12048) );
  AOI22_X1 U14551 ( .A1(n13759), .A2(n12048), .B1(n15858), .B2(
        P3_REG0_REG_9__SCAN_IN), .ZN(n11892) );
  OAI21_X1 U14552 ( .B1(n12104), .B2(n15858), .A(n11892), .ZN(P3_U3417) );
  OAI21_X1 U14553 ( .B1(n11895), .B2(n11894), .A(n11893), .ZN(n11902) );
  NOR2_X1 U14554 ( .A1(n13973), .A2(n11896), .ZN(n11901) );
  NAND2_X1 U14555 ( .A1(n13873), .A2(n11897), .ZN(n11898) );
  NAND2_X1 U14556 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n15677) );
  OAI211_X1 U14557 ( .C1(n11899), .C2(n13952), .A(n11898), .B(n15677), .ZN(
        n11900) );
  AOI211_X1 U14558 ( .C1(n11902), .C2(n13986), .A(n11901), .B(n11900), .ZN(
        n11903) );
  INV_X1 U14559 ( .A(n11903), .ZN(P2_U3203) );
  XOR2_X1 U14560 ( .A(n11905), .B(n11904), .Z(n11906) );
  NAND2_X1 U14561 ( .A1(n11907), .A2(n11906), .ZN(n12056) );
  OAI21_X1 U14562 ( .B1(n11907), .B2(n11906), .A(n12056), .ZN(n11908) );
  NAND2_X1 U14563 ( .A1(n11908), .A2(n14685), .ZN(n11913) );
  INV_X1 U14564 ( .A(n12012), .ZN(n11911) );
  OAI21_X1 U14565 ( .B1(n12009), .B2(n14700), .A(n11909), .ZN(n11910) );
  AOI21_X1 U14566 ( .B1(n11911), .B2(n14698), .A(n11910), .ZN(n11912) );
  OAI211_X1 U14567 ( .C1(n11914), .C2(n14681), .A(n11913), .B(n11912), .ZN(
        P1_U3221) );
  MUX2_X1 U14568 ( .A(n7706), .B(n11915), .S(n15813), .Z(n11918) );
  INV_X1 U14569 ( .A(n12046), .ZN(n11916) );
  AOI22_X1 U14570 ( .A1(n13410), .A2(n12048), .B1(n15812), .B2(n11916), .ZN(
        n11917) );
  OAI211_X1 U14571 ( .C1(n11919), .C2(n13414), .A(n11918), .B(n11917), .ZN(
        P3_U3224) );
  OAI21_X1 U14572 ( .B1(n11921), .B2(n10020), .A(n11920), .ZN(n14502) );
  NAND2_X1 U14573 ( .A1(n12125), .A2(n14500), .ZN(n11922) );
  NAND2_X1 U14574 ( .A1(n11922), .A2(n14273), .ZN(n11923) );
  NOR2_X1 U14575 ( .A1(n6857), .A2(n11923), .ZN(n14499) );
  OAI22_X1 U14576 ( .A1(n14368), .A2(n7885), .B1(n12325), .B2(n14385), .ZN(
        n11924) );
  AOI21_X1 U14577 ( .B1(n14499), .B2(n14399), .A(n11924), .ZN(n11937) );
  OR2_X1 U14578 ( .A1(n11755), .A2(n7400), .ZN(n11927) );
  NAND2_X1 U14579 ( .A1(n11927), .A2(n11926), .ZN(n12121) );
  NAND2_X1 U14580 ( .A1(n12121), .A2(n11928), .ZN(n11929) );
  NAND2_X1 U14581 ( .A1(n11929), .A2(n10020), .ZN(n11931) );
  NAND3_X1 U14582 ( .A1(n11931), .A2(n14379), .A3(n11930), .ZN(n11934) );
  NAND2_X1 U14583 ( .A1(n14376), .A2(n14013), .ZN(n11933) );
  NAND2_X1 U14584 ( .A1(n14374), .A2(n14011), .ZN(n11932) );
  AND2_X1 U14585 ( .A1(n11933), .A2(n11932), .ZN(n12328) );
  NAND2_X1 U14586 ( .A1(n11934), .A2(n12328), .ZN(n14498) );
  MUX2_X1 U14587 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n14498), .S(n14396), .Z(
        n11935) );
  INV_X1 U14588 ( .A(n11935), .ZN(n11936) );
  OAI211_X1 U14589 ( .C1(n14502), .C2(n14371), .A(n11937), .B(n11936), .ZN(
        P2_U3253) );
  XNOR2_X1 U14590 ( .A(n11938), .B(n12834), .ZN(n15600) );
  AOI211_X1 U14591 ( .C1(n15597), .C2(n7631), .A(n15517), .B(n11939), .ZN(
        n15595) );
  NOR2_X1 U14592 ( .A1(n15096), .A2(n11940), .ZN(n11946) );
  INV_X1 U14593 ( .A(n15596), .ZN(n11941) );
  MUX2_X1 U14594 ( .A(n11942), .B(n11941), .S(n15513), .Z(n11943) );
  OAI21_X1 U14595 ( .B1(n15511), .B2(n11944), .A(n11943), .ZN(n11945) );
  AOI211_X1 U14596 ( .C1(n15595), .C2(n15519), .A(n11946), .B(n11945), .ZN(
        n11949) );
  XNOR2_X1 U14597 ( .A(n11947), .B(n12834), .ZN(n15603) );
  INV_X1 U14598 ( .A(n15528), .ZN(n15075) );
  NAND2_X1 U14599 ( .A1(n15603), .A2(n15075), .ZN(n11948) );
  OAI211_X1 U14600 ( .C1(n15529), .C2(n15600), .A(n11949), .B(n11948), .ZN(
        P1_U3286) );
  XNOR2_X1 U14601 ( .A(n11950), .B(n12833), .ZN(n15590) );
  XNOR2_X1 U14602 ( .A(n11951), .B(n12833), .ZN(n11954) );
  NAND2_X1 U14603 ( .A1(n14741), .A2(n14697), .ZN(n11953) );
  NAND2_X1 U14604 ( .A1(n14743), .A2(n15111), .ZN(n11952) );
  NAND2_X1 U14605 ( .A1(n11953), .A2(n11952), .ZN(n14687) );
  AOI21_X1 U14606 ( .B1(n11954), .B2(n15604), .A(n14687), .ZN(n15587) );
  MUX2_X1 U14607 ( .A(n11955), .B(n15587), .S(n15513), .Z(n11959) );
  AOI211_X1 U14608 ( .C1(n12700), .C2(n15499), .A(n15517), .B(n11956), .ZN(
        n15591) );
  OAI22_X1 U14609 ( .A1(n15096), .A2(n14688), .B1(n14690), .B2(n15511), .ZN(
        n11957) );
  AOI21_X1 U14610 ( .B1(n15591), .B2(n15519), .A(n11957), .ZN(n11958) );
  OAI211_X1 U14611 ( .C1(n15529), .C2(n15590), .A(n11959), .B(n11958), .ZN(
        P1_U3287) );
  NAND3_X1 U14612 ( .A1(n11960), .A2(n7177), .A3(n11961), .ZN(n11962) );
  AOI21_X1 U14613 ( .B1(n11964), .B2(n15604), .A(n11963), .ZN(n15576) );
  INV_X2 U14614 ( .A(n15513), .ZN(n15534) );
  OAI22_X1 U14615 ( .A1(n15513), .A2(n10853), .B1(n11965), .B2(n15511), .ZN(
        n11967) );
  OAI211_X1 U14616 ( .C1(n15516), .C2(n12689), .A(n15500), .B(n15498), .ZN(
        n15571) );
  NOR2_X1 U14617 ( .A1(n15571), .A2(n15015), .ZN(n11966) );
  AOI211_X1 U14618 ( .C1(n15515), .C2(n15569), .A(n11967), .B(n11966), .ZN(
        n11970) );
  XNOR2_X1 U14619 ( .A(n11968), .B(n7177), .ZN(n15573) );
  NAND2_X1 U14620 ( .A1(n15573), .A2(n15100), .ZN(n11969) );
  OAI211_X1 U14621 ( .C1(n15576), .C2(n15534), .A(n11970), .B(n11969), .ZN(
        P1_U3289) );
  XNOR2_X1 U14622 ( .A(n11971), .B(n11974), .ZN(n12133) );
  NAND2_X1 U14623 ( .A1(n12133), .A2(n15843), .ZN(n11981) );
  NAND2_X1 U14624 ( .A1(n11973), .A2(n11972), .ZN(n11976) );
  INV_X1 U14625 ( .A(n11976), .ZN(n11975) );
  NAND2_X1 U14626 ( .A1(n11975), .A2(n11974), .ZN(n12085) );
  AOI21_X1 U14627 ( .B1(n11976), .B2(n7503), .A(n15789), .ZN(n11979) );
  NAND2_X1 U14628 ( .A1(n13119), .A2(n15796), .ZN(n11977) );
  AOI21_X1 U14629 ( .B1(n12085), .B2(n11979), .A(n11978), .ZN(n11980) );
  NAND2_X1 U14630 ( .A1(n11981), .A2(n11980), .ZN(n12134) );
  AOI21_X1 U14631 ( .B1(n15856), .B2(n12133), .A(n12134), .ZN(n12141) );
  AOI22_X1 U14632 ( .A1(n13759), .A2(n12137), .B1(n15858), .B2(
        P3_REG0_REG_10__SCAN_IN), .ZN(n11982) );
  OAI21_X1 U14633 ( .B1(n12141), .B2(n15858), .A(n11982), .ZN(P3_U3420) );
  NAND2_X1 U14634 ( .A1(n11983), .A2(n13074), .ZN(n11992) );
  AOI21_X1 U14635 ( .B1(n12038), .B2(n11985), .A(n11984), .ZN(n11991) );
  NAND2_X1 U14636 ( .A1(n13094), .A2(n12136), .ZN(n11988) );
  AOI21_X1 U14637 ( .B1(n13027), .B2(n13119), .A(n11986), .ZN(n11987) );
  AOI21_X1 U14638 ( .B1(n12137), .B2(n13098), .A(n11989), .ZN(n11990) );
  OAI21_X1 U14639 ( .B1(n11992), .B2(n11991), .A(n11990), .ZN(P3_U3157) );
  XNOR2_X1 U14640 ( .A(n11994), .B(n11993), .ZN(n11999) );
  AOI22_X1 U14641 ( .A1(n14374), .A2(n14013), .B1(n14376), .B2(n14015), .ZN(
        n12027) );
  NAND2_X1 U14642 ( .A1(n13873), .A2(n12032), .ZN(n11996) );
  OAI211_X1 U14643 ( .C1(n12027), .C2(n13952), .A(n11996), .B(n11995), .ZN(
        n11997) );
  AOI21_X1 U14644 ( .B1(n12460), .B2(n13998), .A(n11997), .ZN(n11998) );
  OAI21_X1 U14645 ( .B1(n11999), .B2(n13984), .A(n11998), .ZN(P2_U3189) );
  OAI21_X1 U14646 ( .B1(n6636), .B2(n10235), .A(n12000), .ZN(n13538) );
  XNOR2_X1 U14647 ( .A(n12002), .B(n12001), .ZN(n12003) );
  NAND2_X1 U14648 ( .A1(n12003), .A2(n15801), .ZN(n12006) );
  NAND2_X1 U14649 ( .A1(n13117), .A2(n15796), .ZN(n12005) );
  NAND2_X1 U14650 ( .A1(n13119), .A2(n15799), .ZN(n12004) );
  AND2_X1 U14651 ( .A1(n12005), .A2(n12004), .ZN(n12999) );
  NAND2_X1 U14652 ( .A1(n12006), .A2(n12999), .ZN(n13530) );
  AOI21_X1 U14653 ( .B1(n13538), .B2(n15851), .A(n13530), .ZN(n12203) );
  AOI22_X1 U14654 ( .A1(n12201), .A2(n13759), .B1(n15858), .B2(
        P3_REG0_REG_12__SCAN_IN), .ZN(n12007) );
  OAI21_X1 U14655 ( .B1(n12203), .B2(n15858), .A(n12007), .ZN(P3_U3426) );
  INV_X1 U14656 ( .A(n12008), .ZN(n12019) );
  MUX2_X1 U14657 ( .A(n12010), .B(n12009), .S(n15513), .Z(n12011) );
  OAI21_X1 U14658 ( .B1(n15511), .B2(n12012), .A(n12011), .ZN(n12015) );
  NOR2_X1 U14659 ( .A1(n12013), .A2(n15015), .ZN(n12014) );
  AOI211_X1 U14660 ( .C1(n15515), .C2(n12706), .A(n12015), .B(n12014), .ZN(
        n12018) );
  NAND3_X1 U14661 ( .A1(n11716), .A2(n12016), .A3(n15075), .ZN(n12017) );
  OAI211_X1 U14662 ( .C1(n12019), .C2(n15529), .A(n12018), .B(n12017), .ZN(
        P1_U3285) );
  OAI21_X1 U14663 ( .B1(n12021), .B2(n10015), .A(n12020), .ZN(n12111) );
  INV_X1 U14664 ( .A(n12111), .ZN(n12037) );
  INV_X1 U14665 ( .A(n12022), .ZN(n12023) );
  NOR2_X1 U14666 ( .A1(n12024), .A2(n12023), .ZN(n12026) );
  INV_X1 U14667 ( .A(n12026), .ZN(n12025) );
  OAI21_X1 U14668 ( .B1(n12025), .B2(n12606), .A(n14379), .ZN(n12028) );
  NOR2_X1 U14669 ( .A1(n12026), .A2(n10015), .ZN(n12119) );
  OAI21_X1 U14670 ( .B1(n12028), .B2(n12119), .A(n12027), .ZN(n12109) );
  INV_X1 U14671 ( .A(n12109), .ZN(n12029) );
  MUX2_X1 U14672 ( .A(n11070), .B(n12029), .S(n14396), .Z(n12036) );
  INV_X1 U14673 ( .A(n11763), .ZN(n12031) );
  INV_X1 U14674 ( .A(n12127), .ZN(n12030) );
  AOI211_X1 U14675 ( .C1(n12460), .C2(n12031), .A(n14380), .B(n12030), .ZN(
        n12110) );
  INV_X1 U14676 ( .A(n12032), .ZN(n12033) );
  OAI22_X1 U14677 ( .A1(n14368), .A2(n12120), .B1(n12033), .B2(n14385), .ZN(
        n12034) );
  AOI21_X1 U14678 ( .B1(n12110), .B2(n14399), .A(n12034), .ZN(n12035) );
  OAI211_X1 U14679 ( .C1(n14371), .C2(n12037), .A(n12036), .B(n12035), .ZN(
        P2_U3255) );
  INV_X1 U14680 ( .A(n12038), .ZN(n12039) );
  AOI21_X1 U14681 ( .B1(n12041), .B2(n12040), .A(n12039), .ZN(n12050) );
  NOR2_X1 U14682 ( .A1(n13030), .A2(n12042), .ZN(n12043) );
  AOI211_X1 U14683 ( .C1(n13027), .C2(n13120), .A(n12044), .B(n12043), .ZN(
        n12045) );
  OAI21_X1 U14684 ( .B1(n12046), .B2(n13088), .A(n12045), .ZN(n12047) );
  AOI21_X1 U14685 ( .B1(n12048), .B2(n13098), .A(n12047), .ZN(n12049) );
  OAI21_X1 U14686 ( .B1(n12050), .B2(n13100), .A(n12049), .ZN(P3_U3171) );
  INV_X1 U14687 ( .A(n15242), .ZN(n12172) );
  INV_X1 U14688 ( .A(n12056), .ZN(n12052) );
  NOR2_X1 U14689 ( .A1(n12052), .A2(n12051), .ZN(n12058) );
  XNOR2_X1 U14690 ( .A(n12054), .B(n12053), .ZN(n12057) );
  NAND3_X1 U14691 ( .A1(n12056), .A2(n12057), .A3(n12055), .ZN(n12191) );
  OAI211_X1 U14692 ( .C1(n12058), .C2(n12057), .A(n14685), .B(n12191), .ZN(
        n12064) );
  NAND2_X1 U14693 ( .A1(n14738), .A2(n14697), .ZN(n12060) );
  NAND2_X1 U14694 ( .A1(n14740), .A2(n15111), .ZN(n12059) );
  NAND2_X1 U14695 ( .A1(n12060), .A2(n12059), .ZN(n12166) );
  NOR2_X1 U14696 ( .A1(n14712), .A2(n12169), .ZN(n12061) );
  AOI211_X1 U14697 ( .C1(n14710), .C2(n12166), .A(n12062), .B(n12061), .ZN(
        n12063) );
  OAI211_X1 U14698 ( .C1(n12172), .C2(n14681), .A(n12064), .B(n12063), .ZN(
        P1_U3231) );
  INV_X1 U14699 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n12065) );
  NAND2_X1 U14700 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14632)
         );
  OAI21_X1 U14701 ( .B1(n15483), .B2(n12065), .A(n14632), .ZN(n12074) );
  INV_X1 U14702 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12070) );
  MUX2_X1 U14703 ( .A(n12070), .B(P1_REG2_REG_16__SCAN_IN), .S(n12078), .Z(
        n12072) );
  AOI22_X1 U14704 ( .A1(n12067), .A2(n12066), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n12076), .ZN(n12068) );
  NAND2_X1 U14705 ( .A1(n12068), .A2(n12077), .ZN(n12069) );
  OAI21_X1 U14706 ( .B1(n12068), .B2(n12077), .A(n12069), .ZN(n15469) );
  OR2_X1 U14707 ( .A1(n15469), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n15470) );
  NOR2_X1 U14708 ( .A1(n14781), .A2(n12070), .ZN(n14789) );
  AOI211_X1 U14709 ( .C1(n12072), .C2(n12071), .A(n14805), .B(n14790), .ZN(
        n12073) );
  AOI211_X1 U14710 ( .C1(n15475), .C2(n12078), .A(n12074), .B(n12073), .ZN(
        n12082) );
  XOR2_X1 U14711 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12078), .Z(n12079) );
  OAI211_X1 U14712 ( .C1(n12080), .C2(n12079), .A(n14779), .B(n15478), .ZN(
        n12081) );
  NAND2_X1 U14713 ( .A1(n12082), .A2(n12081), .ZN(P1_U3259) );
  INV_X1 U14714 ( .A(n12083), .ZN(n12084) );
  NAND2_X1 U14715 ( .A1(n12085), .A2(n12084), .ZN(n12087) );
  XNOR2_X1 U14716 ( .A(n12087), .B(n12086), .ZN(n12090) );
  NAND2_X1 U14717 ( .A1(n13120), .A2(n15799), .ZN(n12089) );
  NAND2_X1 U14718 ( .A1(n13118), .A2(n15796), .ZN(n12088) );
  NAND2_X1 U14719 ( .A1(n12089), .A2(n12088), .ZN(n13066) );
  AOI21_X1 U14720 ( .B1(n12090), .B2(n15801), .A(n13066), .ZN(n12144) );
  NAND2_X1 U14721 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  NAND2_X1 U14722 ( .A1(n12094), .A2(n12093), .ZN(n12147) );
  OR2_X1 U14723 ( .A1(n12147), .A2(n13745), .ZN(n12095) );
  NAND2_X1 U14724 ( .A1(n12144), .A2(n12095), .ZN(n13751) );
  INV_X1 U14725 ( .A(n13751), .ZN(n12097) );
  AOI22_X1 U14726 ( .A1(n13759), .A2(n13753), .B1(n15858), .B2(
        P3_REG0_REG_11__SCAN_IN), .ZN(n12096) );
  OAI21_X1 U14727 ( .B1(n12097), .B2(n15858), .A(n12096), .ZN(P3_U3423) );
  INV_X1 U14728 ( .A(n12098), .ZN(n12103) );
  NAND2_X1 U14729 ( .A1(n12099), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12644) );
  INV_X1 U14730 ( .A(n12644), .ZN(n12631) );
  AOI21_X1 U14731 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14565), .A(n12631), 
        .ZN(n12100) );
  OAI21_X1 U14732 ( .B1(n12103), .B2(n14569), .A(n12100), .ZN(P2_U3304) );
  AOI21_X1 U14733 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15299), .A(n12101), 
        .ZN(n12102) );
  OAI21_X1 U14734 ( .B1(n12103), .B2(n15305), .A(n12102), .ZN(P1_U3332) );
  INV_X1 U14735 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12105) );
  MUX2_X1 U14736 ( .A(n12105), .B(n12104), .S(n15873), .Z(n12106) );
  OAI21_X1 U14737 ( .B1(n13750), .B2(n12107), .A(n12106), .ZN(P3_U3468) );
  INV_X1 U14738 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n12112) );
  AOI211_X1 U14739 ( .C1(n15764), .C2(n12111), .A(n12110), .B(n12109), .ZN(
        n12115) );
  MUX2_X1 U14740 ( .A(n12112), .B(n12115), .S(n15778), .Z(n12113) );
  OAI21_X1 U14741 ( .B1(n12120), .B2(n14487), .A(n12113), .ZN(P2_U3509) );
  INV_X1 U14742 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12116) );
  MUX2_X1 U14743 ( .A(n12116), .B(n12115), .S(n15767), .Z(n12117) );
  OAI21_X1 U14744 ( .B1(n12120), .B2(n14551), .A(n12117), .ZN(P2_U3460) );
  XNOR2_X1 U14745 ( .A(n12118), .B(n12605), .ZN(n14507) );
  AOI21_X1 U14746 ( .B1(n12120), .B2(n14014), .A(n12119), .ZN(n12122) );
  OAI21_X1 U14747 ( .B1(n12122), .B2(n12605), .A(n12121), .ZN(n12124) );
  AOI22_X1 U14748 ( .A1(n14374), .A2(n14012), .B1(n14376), .B2(n14014), .ZN(
        n12295) );
  INV_X1 U14749 ( .A(n12295), .ZN(n12123) );
  AOI21_X1 U14750 ( .B1(n12124), .B2(n14379), .A(n12123), .ZN(n14506) );
  MUX2_X1 U14751 ( .A(n13667), .B(n14506), .S(n14396), .Z(n12132) );
  INV_X1 U14752 ( .A(n12125), .ZN(n12126) );
  AOI211_X1 U14753 ( .C1(n14504), .C2(n12127), .A(n14380), .B(n12126), .ZN(
        n14503) );
  INV_X1 U14754 ( .A(n14504), .ZN(n12129) );
  INV_X1 U14755 ( .A(n12292), .ZN(n12128) );
  OAI22_X1 U14756 ( .A1(n14368), .A2(n12129), .B1(n12128), .B2(n14385), .ZN(
        n12130) );
  AOI21_X1 U14757 ( .B1(n14503), .B2(n14399), .A(n12130), .ZN(n12131) );
  OAI211_X1 U14758 ( .C1(n14507), .C2(n14371), .A(n12132), .B(n12131), .ZN(
        P2_U3254) );
  INV_X1 U14759 ( .A(n12133), .ZN(n12140) );
  MUX2_X1 U14760 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n12134), .S(n15813), .Z(
        n12135) );
  INV_X1 U14761 ( .A(n12135), .ZN(n12139) );
  AOI22_X1 U14762 ( .A1(n13410), .A2(n12137), .B1(n15812), .B2(n12136), .ZN(
        n12138) );
  OAI211_X1 U14763 ( .C1(n12140), .C2(n13414), .A(n12139), .B(n12138), .ZN(
        P3_U3223) );
  INV_X1 U14764 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n13684) );
  MUX2_X1 U14765 ( .A(n13684), .B(n12141), .S(n15873), .Z(n12142) );
  OAI21_X1 U14766 ( .B1(n13750), .B2(n12143), .A(n12142), .ZN(P3_U3469) );
  MUX2_X1 U14767 ( .A(n12144), .B(n13170), .S(n15816), .Z(n12146) );
  AOI22_X1 U14768 ( .A1(n13410), .A2(n13753), .B1(n15812), .B2(n13065), .ZN(
        n12145) );
  OAI211_X1 U14769 ( .C1(n12147), .C2(n13528), .A(n12146), .B(n12145), .ZN(
        P3_U3222) );
  XNOR2_X1 U14770 ( .A(n12148), .B(n12610), .ZN(n14497) );
  OAI211_X1 U14771 ( .C1(n12151), .C2(n12150), .A(n12149), .B(n14379), .ZN(
        n12152) );
  AOI22_X1 U14772 ( .A1(n14374), .A2(n14010), .B1(n14376), .B2(n14012), .ZN(
        n12363) );
  NAND2_X1 U14773 ( .A1(n12152), .A2(n12363), .ZN(n14493) );
  AOI211_X1 U14774 ( .C1(n14495), .C2(n7887), .A(n14380), .B(n12153), .ZN(
        n14494) );
  NAND2_X1 U14775 ( .A1(n14494), .A2(n14399), .ZN(n12155) );
  AOI22_X1 U14776 ( .A1(n14352), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12365), 
        .B2(n14397), .ZN(n12154) );
  OAI211_X1 U14777 ( .C1(n12368), .C2(n14368), .A(n12155), .B(n12154), .ZN(
        n12156) );
  AOI21_X1 U14778 ( .B1(n14396), .B2(n14493), .A(n12156), .ZN(n12157) );
  OAI21_X1 U14779 ( .B1(n14497), .B2(n14371), .A(n12157), .ZN(P2_U3252) );
  INV_X1 U14780 ( .A(SI_24_), .ZN(n12161) );
  INV_X1 U14781 ( .A(n12158), .ZN(n12159) );
  OAI222_X1 U14782 ( .A1(n12918), .A2(n12161), .B1(n12160), .B2(n12159), .C1(
        P3_U3151), .C2(n9442), .ZN(P3_U3271) );
  INV_X1 U14783 ( .A(n12162), .ZN(n12165) );
  INV_X1 U14784 ( .A(n12163), .ZN(n12164) );
  OAI21_X1 U14785 ( .B1(n12165), .B2(n7011), .A(n12164), .ZN(n12167) );
  AOI21_X1 U14786 ( .B1(n12167), .B2(n15604), .A(n12166), .ZN(n15244) );
  AOI211_X1 U14787 ( .C1(n15242), .C2(n11722), .A(n15517), .B(n12168), .ZN(
        n15241) );
  INV_X1 U14788 ( .A(n12169), .ZN(n12170) );
  AOI22_X1 U14789 ( .A1(n15534), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12170), 
        .B2(n15531), .ZN(n12171) );
  OAI21_X1 U14790 ( .B1(n12172), .B2(n15096), .A(n12171), .ZN(n12175) );
  XOR2_X1 U14791 ( .A(n12173), .B(n12837), .Z(n15245) );
  NOR2_X1 U14792 ( .A1(n15245), .A2(n15529), .ZN(n12174) );
  AOI211_X1 U14793 ( .C1(n15241), .C2(n15519), .A(n12175), .B(n12174), .ZN(
        n12176) );
  OAI21_X1 U14794 ( .B1(n15534), .B2(n15244), .A(n12176), .ZN(P1_U3284) );
  NAND2_X1 U14795 ( .A1(n12178), .A2(n12177), .ZN(n12263) );
  XNOR2_X1 U14796 ( .A(n12263), .B(n12181), .ZN(n15240) );
  OAI211_X1 U14797 ( .C1(n12181), .C2(n12180), .A(n12179), .B(n15604), .ZN(
        n15238) );
  NAND2_X1 U14798 ( .A1(n14739), .A2(n15111), .ZN(n12195) );
  AOI21_X1 U14799 ( .B1(n15238), .B2(n12195), .A(n15534), .ZN(n12182) );
  INV_X1 U14800 ( .A(n12182), .ZN(n12189) );
  OAI22_X1 U14801 ( .A1(n15513), .A2(n12183), .B1(n12196), .B2(n15511), .ZN(
        n12187) );
  AOI21_X1 U14802 ( .B1(n12184), .B2(n15234), .A(n15517), .ZN(n12185) );
  NAND2_X1 U14803 ( .A1(n12185), .A2(n12272), .ZN(n15236) );
  NAND2_X1 U14804 ( .A1(n14737), .A2(n14697), .ZN(n12194) );
  AOI21_X1 U14805 ( .B1(n15236), .B2(n12194), .A(n15015), .ZN(n12186) );
  AOI211_X1 U14806 ( .C1(n15515), .C2(n15234), .A(n12187), .B(n12186), .ZN(
        n12188) );
  OAI211_X1 U14807 ( .C1(n15240), .C2(n15529), .A(n12189), .B(n12188), .ZN(
        P1_U3283) );
  NAND2_X1 U14808 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  XOR2_X1 U14809 ( .A(n12193), .B(n12192), .Z(n12200) );
  AND2_X1 U14810 ( .A1(n12195), .A2(n12194), .ZN(n15237) );
  OAI22_X1 U14811 ( .A1(n15237), .A2(n14700), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8448), .ZN(n12198) );
  NOR2_X1 U14812 ( .A1(n14712), .A2(n12196), .ZN(n12197) );
  AOI211_X1 U14813 ( .C1(n14714), .C2(n15234), .A(n12198), .B(n12197), .ZN(
        n12199) );
  OAI21_X1 U14814 ( .B1(n12200), .B2(n14717), .A(n12199), .ZN(P1_U3217) );
  MUX2_X1 U14815 ( .A(n12203), .B(n12202), .S(n10255), .Z(n12204) );
  OAI21_X1 U14816 ( .B1(n7110), .B2(n13750), .A(n12204), .ZN(P3_U3471) );
  XNOR2_X1 U14817 ( .A(n12206), .B(n12205), .ZN(n13746) );
  INV_X1 U14818 ( .A(n13048), .ZN(n12207) );
  OAI22_X1 U14819 ( .A1(n13814), .A2(n13534), .B1(n12207), .B2(n13532), .ZN(
        n12208) );
  INV_X1 U14820 ( .A(n12208), .ZN(n12216) );
  XNOR2_X1 U14821 ( .A(n12210), .B(n12209), .ZN(n12213) );
  OAI22_X1 U14822 ( .A1(n13045), .A2(n15783), .B1(n12211), .B2(n15785), .ZN(
        n12212) );
  AOI21_X1 U14823 ( .B1(n12213), .B2(n15801), .A(n12212), .ZN(n13744) );
  MUX2_X1 U14824 ( .A(n13744), .B(n12214), .S(n15816), .Z(n12215) );
  OAI211_X1 U14825 ( .C1(n13746), .C2(n13528), .A(n12216), .B(n12215), .ZN(
        P3_U3220) );
  INV_X1 U14826 ( .A(n15291), .ZN(n12227) );
  OAI21_X1 U14827 ( .B1(n12218), .B2(n12217), .A(n12252), .ZN(n12219) );
  NAND2_X1 U14828 ( .A1(n12219), .A2(n14685), .ZN(n12226) );
  INV_X1 U14829 ( .A(n12275), .ZN(n12224) );
  NAND2_X1 U14830 ( .A1(n14738), .A2(n15111), .ZN(n12221) );
  NAND2_X1 U14831 ( .A1(n14736), .A2(n14697), .ZN(n12220) );
  AND2_X1 U14832 ( .A1(n12221), .A2(n12220), .ZN(n12270) );
  OAI21_X1 U14833 ( .B1(n12270), .B2(n14700), .A(n12222), .ZN(n12223) );
  AOI21_X1 U14834 ( .B1(n12224), .B2(n14698), .A(n12223), .ZN(n12225) );
  OAI211_X1 U14835 ( .C1(n12227), .C2(n14681), .A(n12226), .B(n12225), .ZN(
        P1_U3236) );
  INV_X1 U14836 ( .A(n12228), .ZN(n12232) );
  OAI222_X1 U14837 ( .A1(n12946), .A2(n12230), .B1(n15305), .B2(n12232), .C1(
        P1_U3086), .C2(n12229), .ZN(P1_U3331) );
  OAI222_X1 U14838 ( .A1(n12233), .A2(P2_U3088), .B1(n12913), .B2(n12232), 
        .C1(n12231), .C2(n14562), .ZN(P2_U3303) );
  INV_X1 U14839 ( .A(n12234), .ZN(n12236) );
  OAI222_X1 U14840 ( .A1(P3_U3151), .A2(n12237), .B1(n13836), .B2(n12236), 
        .C1(n12235), .C2(n13838), .ZN(P3_U3270) );
  NAND2_X1 U14841 ( .A1(n12240), .A2(n12239), .ZN(n12611) );
  XOR2_X1 U14842 ( .A(n12238), .B(n12611), .Z(n14492) );
  XNOR2_X1 U14843 ( .A(n12241), .B(n12611), .ZN(n12242) );
  OAI222_X1 U14844 ( .A1(n14331), .A2(n13902), .B1(n14329), .B2(n13845), .C1(
        n12242), .C2(n14302), .ZN(n14488) );
  INV_X1 U14845 ( .A(n12153), .ZN(n12244) );
  INV_X1 U14846 ( .A(n12337), .ZN(n12243) );
  AOI211_X1 U14847 ( .C1(n14490), .C2(n12244), .A(n14380), .B(n12243), .ZN(
        n14489) );
  NAND2_X1 U14848 ( .A1(n14489), .A2(n14399), .ZN(n12247) );
  INV_X1 U14849 ( .A(n13844), .ZN(n12245) );
  AOI22_X1 U14850 ( .A1(n14352), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12245), 
        .B2(n14397), .ZN(n12246) );
  OAI211_X1 U14851 ( .C1(n12248), .C2(n14368), .A(n12247), .B(n12246), .ZN(
        n12249) );
  AOI21_X1 U14852 ( .B1(n14488), .B2(n14396), .A(n12249), .ZN(n12250) );
  OAI21_X1 U14853 ( .B1(n14492), .B2(n14371), .A(n12250), .ZN(P2_U3251) );
  AND2_X1 U14854 ( .A1(n12252), .A2(n12251), .ZN(n12255) );
  OAI211_X1 U14855 ( .C1(n12255), .C2(n12254), .A(n14685), .B(n12253), .ZN(
        n12262) );
  INV_X1 U14856 ( .A(n12311), .ZN(n12260) );
  OR2_X1 U14857 ( .A1(n14584), .A2(n14706), .ZN(n12257) );
  NAND2_X1 U14858 ( .A1(n14737), .A2(n15111), .ZN(n12256) );
  AND2_X1 U14859 ( .A1(n12257), .A2(n12256), .ZN(n12309) );
  OAI21_X1 U14860 ( .B1(n12309), .B2(n14700), .A(n12258), .ZN(n12259) );
  AOI21_X1 U14861 ( .B1(n12260), .B2(n14698), .A(n12259), .ZN(n12261) );
  OAI211_X1 U14862 ( .C1(n15225), .C2(n14681), .A(n12262), .B(n12261), .ZN(
        P1_U3224) );
  NAND2_X1 U14863 ( .A1(n12263), .A2(n12839), .ZN(n12265) );
  NAND2_X1 U14864 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  XNOR2_X1 U14865 ( .A(n12266), .B(n12840), .ZN(n15231) );
  NAND3_X1 U14866 ( .A1(n12179), .A2(n7010), .A3(n12267), .ZN(n12268) );
  NAND3_X1 U14867 ( .A1(n12269), .A2(n15604), .A3(n12268), .ZN(n12271) );
  AND2_X1 U14868 ( .A1(n12271), .A2(n12270), .ZN(n15230) );
  INV_X1 U14869 ( .A(n15230), .ZN(n12280) );
  INV_X1 U14870 ( .A(n12314), .ZN(n12274) );
  AOI21_X1 U14871 ( .B1(n12272), .B2(n15291), .A(n15517), .ZN(n12273) );
  NAND2_X1 U14872 ( .A1(n12274), .A2(n12273), .ZN(n15229) );
  OAI22_X1 U14873 ( .A1(n15513), .A2(n12276), .B1(n12275), .B2(n15511), .ZN(
        n12277) );
  AOI21_X1 U14874 ( .B1(n15291), .B2(n15515), .A(n12277), .ZN(n12278) );
  OAI21_X1 U14875 ( .B1(n15229), .B2(n15015), .A(n12278), .ZN(n12279) );
  AOI21_X1 U14876 ( .B1(n12280), .B2(n15513), .A(n12279), .ZN(n12281) );
  OAI21_X1 U14877 ( .B1(n15529), .B2(n15231), .A(n12281), .ZN(P1_U3282) );
  INV_X1 U14878 ( .A(n12282), .ZN(n12286) );
  OAI222_X1 U14879 ( .A1(n12284), .A2(P1_U3086), .B1(n15305), .B2(n12286), 
        .C1(n12283), .C2(n12946), .ZN(P1_U3330) );
  OAI222_X1 U14880 ( .A1(n12287), .A2(P2_U3088), .B1(n12913), .B2(n12286), 
        .C1(n12285), .C2(n14562), .ZN(P2_U3302) );
  INV_X1 U14881 ( .A(n12288), .ZN(n12289) );
  AOI21_X1 U14882 ( .B1(n12291), .B2(n12290), .A(n12289), .ZN(n12298) );
  NAND2_X1 U14883 ( .A1(n13873), .A2(n12292), .ZN(n12294) );
  OAI211_X1 U14884 ( .C1(n12295), .C2(n13952), .A(n12294), .B(n12293), .ZN(
        n12296) );
  AOI21_X1 U14885 ( .B1(n14504), .B2(n13998), .A(n12296), .ZN(n12297) );
  OAI21_X1 U14886 ( .B1(n12298), .B2(n13984), .A(n12297), .ZN(P2_U3208) );
  XNOR2_X1 U14887 ( .A(n12300), .B(n12299), .ZN(n12305) );
  NOR2_X1 U14888 ( .A1(n14712), .A2(n12353), .ZN(n12303) );
  AOI22_X1 U14889 ( .A1(n14734), .A2(n14697), .B1(n15111), .B2(n14736), .ZN(
        n12347) );
  OAI21_X1 U14890 ( .B1(n12347), .B2(n14700), .A(n12301), .ZN(n12302) );
  AOI211_X1 U14891 ( .C1(n12738), .C2(n14714), .A(n12303), .B(n12302), .ZN(
        n12304) );
  OAI21_X1 U14892 ( .B1(n12305), .B2(n14717), .A(n12304), .ZN(P1_U3234) );
  XNOR2_X1 U14893 ( .A(n12306), .B(n7008), .ZN(n15222) );
  INV_X1 U14894 ( .A(n15222), .ZN(n12319) );
  OAI211_X1 U14895 ( .C1(n12308), .C2(n12842), .A(n12307), .B(n15604), .ZN(
        n12310) );
  NAND2_X1 U14896 ( .A1(n12310), .A2(n12309), .ZN(n15227) );
  NAND2_X1 U14897 ( .A1(n15227), .A2(n15513), .ZN(n12318) );
  OAI22_X1 U14898 ( .A1(n15513), .A2(n12312), .B1(n12311), .B2(n15511), .ZN(
        n12316) );
  OAI211_X1 U14899 ( .C1(n12314), .C2(n15225), .A(n15500), .B(n12313), .ZN(
        n15223) );
  NOR2_X1 U14900 ( .A1(n15223), .A2(n15015), .ZN(n12315) );
  AOI211_X1 U14901 ( .C1(n15515), .C2(n12724), .A(n12316), .B(n12315), .ZN(
        n12317) );
  OAI211_X1 U14902 ( .C1(n15529), .C2(n12319), .A(n12318), .B(n12317), .ZN(
        P1_U3281) );
  INV_X1 U14903 ( .A(n12320), .ZN(n12322) );
  NAND2_X1 U14904 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  XNOR2_X1 U14905 ( .A(n12324), .B(n12323), .ZN(n12331) );
  INV_X1 U14906 ( .A(n12325), .ZN(n12326) );
  NAND2_X1 U14907 ( .A1(n13873), .A2(n12326), .ZN(n12327) );
  NAND2_X1 U14908 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15698)
         );
  OAI211_X1 U14909 ( .C1(n12328), .C2(n13952), .A(n12327), .B(n15698), .ZN(
        n12329) );
  AOI21_X1 U14910 ( .B1(n14500), .B2(n13998), .A(n12329), .ZN(n12330) );
  OAI21_X1 U14911 ( .B1(n12331), .B2(n13984), .A(n12330), .ZN(P2_U3196) );
  XNOR2_X1 U14912 ( .A(n12332), .B(n12333), .ZN(n14484) );
  INV_X1 U14913 ( .A(n14484), .ZN(n12343) );
  XNOR2_X1 U14914 ( .A(n12334), .B(n12333), .ZN(n12335) );
  OAI222_X1 U14915 ( .A1(n14331), .A2(n13990), .B1(n14329), .B2(n13994), .C1(
        n12335), .C2(n14302), .ZN(n14482) );
  INV_X1 U14916 ( .A(n14381), .ZN(n12336) );
  AOI211_X1 U14917 ( .C1(n13999), .C2(n12337), .A(n14380), .B(n12336), .ZN(
        n14483) );
  NAND2_X1 U14918 ( .A1(n14483), .A2(n14399), .ZN(n12340) );
  INV_X1 U14919 ( .A(n13992), .ZN(n12338) );
  AOI22_X1 U14920 ( .A1(n14352), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12338), 
        .B2(n14397), .ZN(n12339) );
  OAI211_X1 U14921 ( .C1(n6858), .C2(n14368), .A(n12340), .B(n12339), .ZN(
        n12341) );
  AOI21_X1 U14922 ( .B1(n14482), .B2(n14396), .A(n12341), .ZN(n12342) );
  OAI21_X1 U14923 ( .B1(n12343), .B2(n14371), .A(n12342), .ZN(P2_U3250) );
  OAI211_X1 U14924 ( .C1(n12346), .C2(n12345), .A(n12344), .B(n15604), .ZN(
        n12348) );
  NAND2_X1 U14925 ( .A1(n12348), .A2(n12347), .ZN(n15217) );
  INV_X1 U14926 ( .A(n15217), .ZN(n12359) );
  NAND2_X1 U14927 ( .A1(n12350), .A2(n12349), .ZN(n12351) );
  XNOR2_X1 U14928 ( .A(n12351), .B(n12844), .ZN(n15219) );
  INV_X1 U14929 ( .A(n15091), .ZN(n12352) );
  AOI211_X1 U14930 ( .C1(n12738), .C2(n12313), .A(n15517), .B(n12352), .ZN(
        n15218) );
  NAND2_X1 U14931 ( .A1(n15218), .A2(n15519), .ZN(n12356) );
  INV_X1 U14932 ( .A(n12353), .ZN(n12354) );
  AOI22_X1 U14933 ( .A1(n15534), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n12354), 
        .B2(n15531), .ZN(n12355) );
  OAI211_X1 U14934 ( .C1(n15286), .C2(n15096), .A(n12356), .B(n12355), .ZN(
        n12357) );
  AOI21_X1 U14935 ( .B1(n15100), .B2(n15219), .A(n12357), .ZN(n12358) );
  OAI21_X1 U14936 ( .B1(n12359), .B2(n15534), .A(n12358), .ZN(P1_U3280) );
  OAI211_X1 U14937 ( .C1(n12362), .C2(n12361), .A(n12360), .B(n13986), .ZN(
        n12367) );
  OAI22_X1 U14938 ( .A1(n13952), .A2(n12363), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14097), .ZN(n12364) );
  AOI21_X1 U14939 ( .B1(n12365), .B2(n13873), .A(n12364), .ZN(n12366) );
  OAI211_X1 U14940 ( .C1(n12368), .C2(n13973), .A(n12367), .B(n12366), .ZN(
        P2_U3206) );
  INV_X1 U14941 ( .A(n12369), .ZN(n12372) );
  OAI222_X1 U14942 ( .A1(n13836), .A2(n12372), .B1(P3_U3151), .B2(n12371), 
        .C1(n12370), .C2(n12918), .ZN(P3_U3265) );
  NOR2_X1 U14943 ( .A1(n12381), .A2(n15727), .ZN(n12379) );
  OAI21_X1 U14944 ( .B1(n14025), .B2(n11663), .A(n12374), .ZN(n12378) );
  NAND2_X1 U14945 ( .A1(n14025), .A2(n15727), .ZN(n12376) );
  NAND2_X1 U14946 ( .A1(n12625), .A2(n14386), .ZN(n12375) );
  NAND3_X1 U14947 ( .A1(n12376), .A2(n12582), .A3(n12375), .ZN(n12377) );
  OAI21_X1 U14948 ( .B1(n12379), .B2(n12378), .A(n12377), .ZN(n12390) );
  NAND2_X1 U14949 ( .A1(n12383), .A2(n12382), .ZN(n12389) );
  NAND2_X1 U14950 ( .A1(n6617), .A2(n6421), .ZN(n12385) );
  NAND2_X1 U14951 ( .A1(n14023), .A2(n12381), .ZN(n12384) );
  AND2_X1 U14952 ( .A1(n12385), .A2(n12384), .ZN(n12394) );
  NAND2_X1 U14953 ( .A1(n12547), .A2(n14023), .ZN(n12387) );
  NAND2_X1 U14954 ( .A1(n12556), .A2(n6421), .ZN(n12386) );
  NAND2_X1 U14955 ( .A1(n12387), .A2(n12386), .ZN(n12393) );
  OAI22_X1 U14956 ( .A1(n12390), .A2(n12389), .B1(n12394), .B2(n12393), .ZN(
        n12392) );
  AOI22_X1 U14957 ( .A1(n12547), .A2(n10044), .B1(n14024), .B2(n12381), .ZN(
        n12388) );
  AOI21_X1 U14958 ( .B1(n12390), .B2(n12389), .A(n12388), .ZN(n12391) );
  NOR2_X1 U14959 ( .A1(n12392), .A2(n12391), .ZN(n12407) );
  NAND2_X1 U14960 ( .A1(n14021), .A2(n12381), .ZN(n12395) );
  NAND2_X1 U14961 ( .A1(n12547), .A2(n14021), .ZN(n12398) );
  NAND2_X1 U14962 ( .A1(n12556), .A2(n12396), .ZN(n12397) );
  NAND2_X1 U14963 ( .A1(n12398), .A2(n12397), .ZN(n12408) );
  NAND2_X1 U14964 ( .A1(n12547), .A2(n14022), .ZN(n12400) );
  NAND2_X1 U14965 ( .A1(n12381), .A2(n15742), .ZN(n12399) );
  AND2_X1 U14966 ( .A1(n12400), .A2(n12399), .ZN(n12413) );
  NAND2_X1 U14967 ( .A1(n6617), .A2(n15742), .ZN(n12402) );
  NAND2_X1 U14968 ( .A1(n14022), .A2(n12556), .ZN(n12401) );
  NAND2_X1 U14969 ( .A1(n12402), .A2(n12401), .ZN(n12412) );
  NAND2_X1 U14970 ( .A1(n12404), .A2(n12381), .ZN(n12406) );
  NAND2_X1 U14971 ( .A1(n12547), .A2(n14020), .ZN(n12405) );
  NAND2_X1 U14972 ( .A1(n12406), .A2(n12405), .ZN(n12416) );
  INV_X1 U14973 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14974 ( .A(n12409), .ZN(n12410) );
  AOI22_X1 U14975 ( .A1(n12413), .A2(n12412), .B1(n12411), .B2(n12410), .ZN(
        n12427) );
  NAND2_X1 U14976 ( .A1(n12415), .A2(n12414), .ZN(n12426) );
  INV_X1 U14977 ( .A(n12416), .ZN(n12424) );
  INV_X1 U14978 ( .A(n12417), .ZN(n12423) );
  NAND2_X1 U14979 ( .A1(n12420), .A2(n12381), .ZN(n12419) );
  NAND2_X1 U14980 ( .A1(n12547), .A2(n14019), .ZN(n12418) );
  AND2_X1 U14981 ( .A1(n12419), .A2(n12418), .ZN(n12432) );
  NAND2_X1 U14982 ( .A1(n12420), .A2(n6617), .ZN(n12422) );
  NAND2_X1 U14983 ( .A1(n14019), .A2(n12381), .ZN(n12421) );
  NAND2_X1 U14984 ( .A1(n12422), .A2(n12421), .ZN(n12431) );
  AOI22_X1 U14985 ( .A1(n12424), .A2(n12423), .B1(n12432), .B2(n12431), .ZN(
        n12425) );
  OAI21_X1 U14986 ( .B1(n12427), .B2(n12426), .A(n12425), .ZN(n12436) );
  INV_X1 U14987 ( .A(n6617), .ZN(n12556) );
  AOI22_X1 U14988 ( .A1(n12428), .A2(n12547), .B1(n14018), .B2(n12556), .ZN(
        n12439) );
  NAND2_X1 U14989 ( .A1(n12428), .A2(n12381), .ZN(n12430) );
  NAND2_X1 U14990 ( .A1(n12547), .A2(n14018), .ZN(n12429) );
  NAND2_X1 U14991 ( .A1(n12430), .A2(n12429), .ZN(n12438) );
  INV_X1 U14992 ( .A(n12431), .ZN(n12434) );
  INV_X1 U14993 ( .A(n12432), .ZN(n12433) );
  AOI22_X1 U14994 ( .A1(n12439), .A2(n12438), .B1(n12434), .B2(n12433), .ZN(
        n12435) );
  INV_X1 U14995 ( .A(n12437), .ZN(n12452) );
  INV_X1 U14996 ( .A(n12438), .ZN(n12441) );
  INV_X1 U14997 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14998 ( .A1(n12441), .A2(n12440), .ZN(n12447) );
  AOI22_X1 U14999 ( .A1(n14509), .A2(n6617), .B1(n14017), .B2(n12381), .ZN(
        n12449) );
  INV_X1 U15000 ( .A(n12449), .ZN(n12445) );
  NAND2_X1 U15001 ( .A1(n14509), .A2(n12556), .ZN(n12443) );
  NAND2_X1 U15002 ( .A1(n6617), .A2(n14017), .ZN(n12442) );
  NAND2_X1 U15003 ( .A1(n12443), .A2(n12442), .ZN(n12448) );
  NAND2_X1 U15004 ( .A1(n12447), .A2(n12446), .ZN(n12451) );
  NAND2_X1 U15005 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  NAND2_X1 U15006 ( .A1(n12455), .A2(n12556), .ZN(n12454) );
  NAND2_X1 U15007 ( .A1(n12547), .A2(n14015), .ZN(n12453) );
  NAND2_X1 U15008 ( .A1(n12454), .A2(n12453), .ZN(n12457) );
  AOI22_X1 U15009 ( .A1(n12455), .A2(n12547), .B1(n14015), .B2(n12556), .ZN(
        n12456) );
  NAND2_X1 U15010 ( .A1(n12460), .A2(n6617), .ZN(n12459) );
  NAND2_X1 U15011 ( .A1(n14014), .A2(n12556), .ZN(n12458) );
  NAND2_X1 U15012 ( .A1(n12460), .A2(n12381), .ZN(n12461) );
  OAI21_X1 U15013 ( .B1(n12462), .B2(n12381), .A(n12461), .ZN(n12463) );
  AOI22_X1 U15014 ( .A1(n14504), .A2(n12547), .B1(n14013), .B2(n12381), .ZN(
        n12468) );
  NAND2_X1 U15015 ( .A1(n14504), .A2(n12381), .ZN(n12465) );
  NAND2_X1 U15016 ( .A1(n12547), .A2(n14013), .ZN(n12464) );
  NAND2_X1 U15017 ( .A1(n12465), .A2(n12464), .ZN(n12467) );
  NAND2_X1 U15018 ( .A1(n12468), .A2(n12467), .ZN(n12466) );
  INV_X1 U15019 ( .A(n12467), .ZN(n12470) );
  INV_X1 U15020 ( .A(n12468), .ZN(n12469) );
  NAND2_X1 U15021 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  NAND2_X1 U15022 ( .A1(n12472), .A2(n12471), .ZN(n12477) );
  NAND2_X1 U15023 ( .A1(n14500), .A2(n6617), .ZN(n12474) );
  NAND2_X1 U15024 ( .A1(n14012), .A2(n12556), .ZN(n12473) );
  NAND2_X1 U15025 ( .A1(n12474), .A2(n12473), .ZN(n12476) );
  AOI22_X1 U15026 ( .A1(n14500), .A2(n12556), .B1(n6617), .B2(n14012), .ZN(
        n12475) );
  NAND2_X1 U15027 ( .A1(n14495), .A2(n12556), .ZN(n12479) );
  NAND2_X1 U15028 ( .A1(n6617), .A2(n14011), .ZN(n12478) );
  NAND2_X1 U15029 ( .A1(n12479), .A2(n12478), .ZN(n12483) );
  NAND2_X1 U15030 ( .A1(n14495), .A2(n6617), .ZN(n12480) );
  OAI21_X1 U15031 ( .B1(n13845), .B2(n12547), .A(n12480), .ZN(n12481) );
  NAND2_X1 U15032 ( .A1(n12482), .A2(n12481), .ZN(n12485) );
  NAND2_X1 U15033 ( .A1(n14490), .A2(n6617), .ZN(n12487) );
  NAND2_X1 U15034 ( .A1(n14010), .A2(n12556), .ZN(n12486) );
  NAND2_X1 U15035 ( .A1(n12487), .A2(n12486), .ZN(n12489) );
  AOI22_X1 U15036 ( .A1(n14490), .A2(n12556), .B1(n6617), .B2(n14010), .ZN(
        n12488) );
  NAND2_X1 U15037 ( .A1(n13999), .A2(n12556), .ZN(n12491) );
  NAND2_X1 U15038 ( .A1(n14377), .A2(n6617), .ZN(n12490) );
  NAND2_X1 U15039 ( .A1(n12491), .A2(n12490), .ZN(n12493) );
  AOI22_X1 U15040 ( .A1(n13999), .A2(n12547), .B1(n14377), .B2(n12381), .ZN(
        n12492) );
  AOI22_X1 U15041 ( .A1(n14477), .A2(n12547), .B1(n14359), .B2(n12381), .ZN(
        n12497) );
  INV_X1 U15042 ( .A(n14477), .ZN(n12495) );
  OAI22_X1 U15043 ( .A1(n12495), .A2(n12547), .B1(n13990), .B2(n12556), .ZN(
        n12496) );
  OAI22_X1 U15044 ( .A1(n14546), .A2(n12547), .B1(n14330), .B2(n12381), .ZN(
        n12501) );
  OAI22_X1 U15045 ( .A1(n14546), .A2(n12381), .B1(n14330), .B2(n12547), .ZN(
        n12503) );
  INV_X1 U15046 ( .A(n12501), .ZN(n12502) );
  AOI22_X1 U15047 ( .A1(n14466), .A2(n12547), .B1(n14360), .B2(n12381), .ZN(
        n12505) );
  OAI22_X1 U15048 ( .A1(n14347), .A2(n12547), .B1(n14314), .B2(n12381), .ZN(
        n12504) );
  AOI22_X1 U15049 ( .A1(n14321), .A2(n12556), .B1(n6617), .B2(n14009), .ZN(
        n12508) );
  OAI22_X1 U15050 ( .A1(n7890), .A2(n12381), .B1(n14332), .B2(n12547), .ZN(
        n12506) );
  OAI22_X1 U15051 ( .A1(n14308), .A2(n12556), .B1(n14315), .B2(n12547), .ZN(
        n12510) );
  NAND2_X1 U15052 ( .A1(n12509), .A2(n12510), .ZN(n12514) );
  OAI22_X1 U15053 ( .A1(n14308), .A2(n12547), .B1(n14315), .B2(n12381), .ZN(
        n12513) );
  INV_X1 U15054 ( .A(n12510), .ZN(n12511) );
  OAI22_X1 U15055 ( .A1(n14537), .A2(n12547), .B1(n14303), .B2(n12381), .ZN(
        n12517) );
  INV_X1 U15056 ( .A(n12517), .ZN(n12516) );
  OAI22_X1 U15057 ( .A1(n14537), .A2(n12381), .B1(n14303), .B2(n12547), .ZN(
        n12515) );
  AOI22_X1 U15058 ( .A1(n14277), .A2(n12547), .B1(n14285), .B2(n12381), .ZN(
        n12520) );
  OAI22_X1 U15059 ( .A1(n14533), .A2(n12547), .B1(n14255), .B2(n12556), .ZN(
        n12519) );
  AOI22_X1 U15060 ( .A1(n14440), .A2(n12381), .B1(n6617), .B2(n14227), .ZN(
        n12524) );
  INV_X1 U15061 ( .A(n12524), .ZN(n12522) );
  AOI22_X1 U15062 ( .A1(n14440), .A2(n6617), .B1(n14227), .B2(n12381), .ZN(
        n12521) );
  OAI22_X1 U15063 ( .A1(n14233), .A2(n12381), .B1(n14256), .B2(n12547), .ZN(
        n12527) );
  OAI22_X1 U15064 ( .A1(n14233), .A2(n12547), .B1(n14256), .B2(n12381), .ZN(
        n12526) );
  OAI22_X1 U15065 ( .A1(n14527), .A2(n12547), .B1(n13980), .B2(n12381), .ZN(
        n12528) );
  OAI22_X1 U15066 ( .A1(n14527), .A2(n12381), .B1(n13980), .B2(n12547), .ZN(
        n12529) );
  AOI22_X1 U15067 ( .A1(n14425), .A2(n12547), .B1(n14006), .B2(n12381), .ZN(
        n12530) );
  AOI22_X1 U15068 ( .A1(n14425), .A2(n12381), .B1(n6617), .B2(n14006), .ZN(
        n12531) );
  AOI22_X1 U15069 ( .A1(n14420), .A2(n12381), .B1(n6617), .B2(n14196), .ZN(
        n12560) );
  OAI22_X1 U15070 ( .A1(n14190), .A2(n12381), .B1(n13979), .B2(n12547), .ZN(
        n12561) );
  NAND2_X1 U15071 ( .A1(n12910), .A2(n9302), .ZN(n12533) );
  NAND2_X1 U15072 ( .A1(n12550), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12532) );
  NAND2_X1 U15073 ( .A1(n12640), .A2(n12534), .ZN(n12535) );
  AOI21_X1 U15074 ( .B1(n12536), .B2(n12626), .A(n12535), .ZN(n12541) );
  INV_X1 U15075 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U15076 ( .A1(n6474), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15077 ( .A1(n9375), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12537) );
  OAI211_X1 U15078 ( .C1(n12539), .C2(n14514), .A(n12538), .B(n12537), .ZN(
        n14002) );
  NAND2_X1 U15079 ( .A1(n14002), .A2(n12381), .ZN(n12540) );
  AOI21_X1 U15080 ( .B1(n12541), .B2(n12540), .A(n12543), .ZN(n12542) );
  AOI21_X1 U15081 ( .B1(n14169), .B2(n12547), .A(n12542), .ZN(n12573) );
  NAND2_X1 U15082 ( .A1(n14169), .A2(n12556), .ZN(n12545) );
  INV_X1 U15083 ( .A(n12543), .ZN(n14003) );
  NAND2_X1 U15084 ( .A1(n12547), .A2(n14003), .ZN(n12544) );
  NAND2_X1 U15085 ( .A1(n12545), .A2(n12544), .ZN(n12572) );
  AND2_X1 U15086 ( .A1(n14004), .A2(n12556), .ZN(n12546) );
  AOI21_X1 U15087 ( .B1(n14415), .B2(n12547), .A(n12546), .ZN(n12565) );
  NAND2_X1 U15088 ( .A1(n14415), .A2(n12556), .ZN(n12549) );
  NAND2_X1 U15089 ( .A1(n14004), .A2(n6617), .ZN(n12548) );
  NAND2_X1 U15090 ( .A1(n12549), .A2(n12548), .ZN(n12564) );
  OAI22_X1 U15091 ( .A1(n12573), .A2(n12572), .B1(n12565), .B2(n12564), .ZN(
        n12554) );
  NAND2_X1 U15092 ( .A1(n12550), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15093 ( .A1(n14516), .A2(n14002), .ZN(n12553) );
  INV_X1 U15094 ( .A(n14002), .ZN(n14171) );
  NAND2_X1 U15095 ( .A1(n12552), .A2(n14171), .ZN(n12581) );
  NAND2_X1 U15096 ( .A1(n12554), .A2(n12624), .ZN(n12575) );
  AND2_X1 U15097 ( .A1(n14005), .A2(n6617), .ZN(n12555) );
  AOI21_X1 U15098 ( .B1(n12934), .B2(n12556), .A(n12555), .ZN(n12567) );
  NAND2_X1 U15099 ( .A1(n12934), .A2(n6617), .ZN(n12558) );
  NAND2_X1 U15100 ( .A1(n14005), .A2(n12556), .ZN(n12557) );
  NAND2_X1 U15101 ( .A1(n12558), .A2(n12557), .ZN(n12566) );
  NAND2_X1 U15102 ( .A1(n12567), .A2(n12566), .ZN(n12559) );
  NAND2_X1 U15103 ( .A1(n12575), .A2(n12559), .ZN(n12578) );
  AOI21_X1 U15104 ( .B1(n12560), .B2(n12561), .A(n12578), .ZN(n12580) );
  INV_X1 U15105 ( .A(n12560), .ZN(n12563) );
  INV_X1 U15106 ( .A(n12561), .ZN(n12562) );
  NAND2_X1 U15107 ( .A1(n12563), .A2(n12562), .ZN(n12577) );
  INV_X1 U15108 ( .A(n12564), .ZN(n12571) );
  INV_X1 U15109 ( .A(n12565), .ZN(n12570) );
  INV_X1 U15110 ( .A(n12566), .ZN(n12569) );
  INV_X1 U15111 ( .A(n12567), .ZN(n12568) );
  AOI22_X1 U15112 ( .A1(n12575), .A2(n12574), .B1(n12573), .B2(n12572), .ZN(
        n12576) );
  OAI21_X1 U15113 ( .B1(n12578), .B2(n12577), .A(n12576), .ZN(n12579) );
  NOR2_X1 U15114 ( .A1(n12581), .A2(n6617), .ZN(n12639) );
  INV_X1 U15115 ( .A(n12639), .ZN(n12586) );
  NAND3_X1 U15116 ( .A1(n14516), .A2(n12547), .A3(n14002), .ZN(n12585) );
  NAND2_X1 U15117 ( .A1(n12582), .A2(n12625), .ZN(n12583) );
  OAI211_X1 U15118 ( .C1(n14386), .C2(n8895), .A(n12583), .B(n12640), .ZN(
        n12584) );
  NAND4_X1 U15119 ( .A1(n12586), .A2(n12631), .A3(n12585), .A4(n12584), .ZN(
        n12650) );
  XNOR2_X1 U15120 ( .A(n14169), .B(n14003), .ZN(n12623) );
  XNOR2_X1 U15121 ( .A(n14425), .B(n12587), .ZN(n14203) );
  NAND2_X1 U15122 ( .A1(n12589), .A2(n12588), .ZN(n14253) );
  NAND2_X1 U15123 ( .A1(n12591), .A2(n12590), .ZN(n14312) );
  AND4_X1 U15124 ( .A1(n6590), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12602) );
  NAND4_X1 U15125 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12603) );
  NOR2_X1 U15126 ( .A1(n12604), .A2(n12603), .ZN(n12607) );
  NAND4_X1 U15127 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        n12609) );
  NOR2_X1 U15128 ( .A1(n12610), .A2(n12609), .ZN(n12612) );
  NAND4_X1 U15129 ( .A1(n14353), .A2(n12612), .A3(n14389), .A4(n12611), .ZN(
        n12613) );
  NOR2_X1 U15130 ( .A1(n12614), .A2(n12613), .ZN(n12615) );
  NAND3_X1 U15131 ( .A1(n14312), .A2(n12615), .A3(n14336), .ZN(n12616) );
  NOR2_X1 U15132 ( .A1(n14300), .A2(n12616), .ZN(n12617) );
  NAND4_X1 U15133 ( .A1(n14253), .A2(n14266), .A3(n12617), .A4(n14281), .ZN(
        n12618) );
  AND3_X1 U15134 ( .A1(n12620), .A2(n6504), .A3(n14180), .ZN(n12622) );
  NAND4_X1 U15135 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12635) );
  INV_X1 U15136 ( .A(n12635), .ZN(n12632) );
  NAND3_X1 U15137 ( .A1(n12631), .A2(n14386), .A3(n8895), .ZN(n12633) );
  INV_X1 U15138 ( .A(n12625), .ZN(n15726) );
  MUX2_X1 U15139 ( .A(n12534), .B(n15726), .S(n12626), .Z(n12628) );
  NOR2_X1 U15140 ( .A1(n12644), .A2(n12630), .ZN(n12627) );
  NAND2_X1 U15141 ( .A1(n12628), .A2(n12627), .ZN(n12637) );
  OAI21_X1 U15142 ( .B1(n12632), .B2(n12633), .A(n12637), .ZN(n12629) );
  NAND4_X1 U15143 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n8895), .ZN(
        n12648) );
  INV_X1 U15144 ( .A(n12633), .ZN(n12634) );
  OAI211_X1 U15145 ( .C1(n12636), .C2(n12639), .A(n12635), .B(n12634), .ZN(
        n12647) );
  INV_X1 U15146 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U15147 ( .A1(n12639), .A2(n12638), .ZN(n12646) );
  INV_X1 U15148 ( .A(n12640), .ZN(n12641) );
  NAND4_X1 U15149 ( .A1(n15722), .A2(n12642), .A3(n14376), .A4(n12641), .ZN(
        n12643) );
  OAI211_X1 U15150 ( .C1(n15726), .C2(n12644), .A(n12643), .B(P2_B_REG_SCAN_IN), .ZN(n12645) );
  INV_X2 U15151 ( .A(n12737), .ZN(n12823) );
  MUX2_X1 U15152 ( .A(n12653), .B(n15131), .S(n12823), .Z(n12807) );
  MUX2_X1 U15153 ( .A(n14720), .B(n14834), .S(n12691), .Z(n12806) );
  NAND2_X1 U15154 ( .A1(n12807), .A2(n12806), .ZN(n12665) );
  INV_X1 U15155 ( .A(n12665), .ZN(n12813) );
  NAND2_X1 U15156 ( .A1(n14719), .A2(n12823), .ZN(n12654) );
  OAI21_X1 U15157 ( .B1(n8801), .B2(n12655), .A(n12654), .ZN(n12661) );
  INV_X1 U15158 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15126) );
  NAND2_X1 U15159 ( .A1(n12656), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12659) );
  NAND2_X1 U15160 ( .A1(n12657), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12658) );
  OAI211_X1 U15161 ( .C1(n12660), .C2(n15126), .A(n12659), .B(n12658), .ZN(
        n14841) );
  AND2_X1 U15162 ( .A1(n12661), .A2(n14841), .ZN(n12662) );
  AOI21_X1 U15163 ( .B1(n14826), .B2(n12691), .A(n12662), .ZN(n12809) );
  INV_X1 U15164 ( .A(n12809), .ZN(n12812) );
  OAI21_X1 U15165 ( .B1(n14719), .B2(n15526), .A(n14841), .ZN(n12663) );
  INV_X1 U15166 ( .A(n12663), .ZN(n12664) );
  MUX2_X1 U15167 ( .A(n12664), .B(n14826), .S(n12823), .Z(n12810) );
  AOI21_X1 U15168 ( .B1(n12809), .B2(n12665), .A(n12810), .ZN(n12811) );
  INV_X1 U15169 ( .A(n14743), .ZN(n12666) );
  AOI21_X1 U15170 ( .B1(n12666), .B2(n12803), .A(n15580), .ZN(n12698) );
  AOI21_X1 U15171 ( .B1(n14743), .B2(n12823), .A(n15495), .ZN(n12697) );
  INV_X1 U15172 ( .A(n12667), .ZN(n12669) );
  OAI21_X1 U15173 ( .B1(n15525), .B2(n12670), .A(n15105), .ZN(n12671) );
  NAND2_X1 U15174 ( .A1(n14747), .A2(n12768), .ZN(n12681) );
  NAND2_X1 U15175 ( .A1(n15117), .A2(n12691), .ZN(n12680) );
  NAND2_X1 U15176 ( .A1(n12684), .A2(n12691), .ZN(n12687) );
  NAND3_X1 U15177 ( .A1(n14745), .A2(n12685), .A3(n12768), .ZN(n12686) );
  NAND2_X1 U15178 ( .A1(n12688), .A2(n8053), .ZN(n12696) );
  INV_X1 U15179 ( .A(n14744), .ZN(n12690) );
  AOI21_X1 U15180 ( .B1(n12690), .B2(n12768), .A(n12689), .ZN(n12693) );
  AOI21_X1 U15181 ( .B1(n14744), .B2(n12691), .A(n15569), .ZN(n12692) );
  MUX2_X1 U15182 ( .A(n14688), .B(n12699), .S(n12737), .Z(n12702) );
  MUX2_X1 U15183 ( .A(n12700), .B(n14742), .S(n12768), .Z(n12701) );
  MUX2_X1 U15184 ( .A(n15597), .B(n14741), .S(n12823), .Z(n12704) );
  MUX2_X1 U15185 ( .A(n14741), .B(n15597), .S(n12823), .Z(n12703) );
  INV_X1 U15186 ( .A(n12704), .ZN(n12705) );
  MUX2_X1 U15187 ( .A(n14740), .B(n12706), .S(n12768), .Z(n12709) );
  MUX2_X1 U15188 ( .A(n14740), .B(n12706), .S(n12691), .Z(n12707) );
  MUX2_X1 U15189 ( .A(n14739), .B(n15242), .S(n12737), .Z(n12711) );
  MUX2_X1 U15190 ( .A(n14739), .B(n15242), .S(n12768), .Z(n12710) );
  MUX2_X1 U15191 ( .A(n14738), .B(n15234), .S(n12768), .Z(n12715) );
  NAND2_X1 U15192 ( .A1(n12714), .A2(n12715), .ZN(n12713) );
  MUX2_X1 U15193 ( .A(n14738), .B(n15234), .S(n12691), .Z(n12712) );
  NAND2_X1 U15194 ( .A1(n12713), .A2(n12712), .ZN(n12719) );
  INV_X1 U15195 ( .A(n12714), .ZN(n12717) );
  INV_X1 U15196 ( .A(n12715), .ZN(n12716) );
  NAND2_X1 U15197 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  NAND2_X1 U15198 ( .A1(n12719), .A2(n12718), .ZN(n12721) );
  MUX2_X1 U15199 ( .A(n14737), .B(n15291), .S(n12691), .Z(n12722) );
  MUX2_X1 U15200 ( .A(n14737), .B(n15291), .S(n12823), .Z(n12720) );
  INV_X1 U15201 ( .A(n12722), .ZN(n12723) );
  MUX2_X1 U15202 ( .A(n12724), .B(n14736), .S(n12737), .Z(n12728) );
  MUX2_X1 U15203 ( .A(n12724), .B(n14736), .S(n12823), .Z(n12725) );
  NAND2_X1 U15204 ( .A1(n12726), .A2(n12725), .ZN(n12732) );
  INV_X1 U15205 ( .A(n12727), .ZN(n12730) );
  INV_X1 U15206 ( .A(n12728), .ZN(n12729) );
  NAND2_X1 U15207 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  NAND2_X1 U15208 ( .A1(n10372), .A2(n12733), .ZN(n12734) );
  NAND2_X1 U15209 ( .A1(n12734), .A2(n12803), .ZN(n12742) );
  NAND2_X1 U15210 ( .A1(n12747), .A2(n12735), .ZN(n12736) );
  NAND2_X1 U15211 ( .A1(n12736), .A2(n12823), .ZN(n12741) );
  MUX2_X1 U15212 ( .A(n14584), .B(n15286), .S(n12803), .Z(n12743) );
  INV_X1 U15213 ( .A(n14584), .ZN(n14735) );
  MUX2_X1 U15214 ( .A(n14735), .B(n12738), .S(n12823), .Z(n12739) );
  NAND3_X1 U15215 ( .A1(n15099), .A2(n12743), .A3(n12739), .ZN(n12740) );
  INV_X1 U15216 ( .A(n12743), .ZN(n12745) );
  NAND2_X1 U15217 ( .A1(n14735), .A2(n12803), .ZN(n12744) );
  OAI211_X1 U15218 ( .C1(n15286), .C2(n12803), .A(n12745), .B(n12744), .ZN(
        n12746) );
  AND2_X1 U15219 ( .A1(n15099), .A2(n12746), .ZN(n12752) );
  MUX2_X1 U15220 ( .A(n12747), .B(n10372), .S(n12823), .Z(n12749) );
  MUX2_X1 U15221 ( .A(n14707), .B(n15064), .S(n12823), .Z(n12757) );
  MUX2_X1 U15222 ( .A(n14731), .B(n15200), .S(n12803), .Z(n12756) );
  NAND2_X1 U15223 ( .A1(n12757), .A2(n12756), .ZN(n12748) );
  AND2_X1 U15224 ( .A1(n12749), .A2(n12748), .ZN(n12751) );
  XNOR2_X1 U15225 ( .A(n15188), .B(n14729), .ZN(n12750) );
  OAI211_X1 U15226 ( .C1(n6608), .C2(n12752), .A(n12751), .B(n12755), .ZN(
        n12753) );
  NOR2_X1 U15227 ( .A1(n12753), .A2(n15006), .ZN(n12754) );
  INV_X1 U15228 ( .A(n12756), .ZN(n12759) );
  INV_X1 U15229 ( .A(n12757), .ZN(n12758) );
  MUX2_X1 U15230 ( .A(n14730), .B(n15045), .S(n12803), .Z(n12764) );
  NAND2_X1 U15231 ( .A1(n12762), .A2(n14729), .ZN(n12760) );
  OAI22_X1 U15232 ( .A1(n12764), .A2(n12760), .B1(n14729), .B2(n12803), .ZN(
        n12761) );
  NAND2_X1 U15233 ( .A1(n12761), .A2(n15188), .ZN(n12767) );
  NAND2_X1 U15234 ( .A1(n12762), .A2(n14599), .ZN(n12763) );
  OAI22_X1 U15235 ( .A1(n12764), .A2(n12763), .B1(n14599), .B2(n12823), .ZN(
        n12765) );
  NAND2_X1 U15236 ( .A1(n12765), .A2(n15032), .ZN(n12766) );
  AND2_X1 U15237 ( .A1(n15012), .A2(n12768), .ZN(n12770) );
  NOR2_X1 U15238 ( .A1(n15012), .A2(n12823), .ZN(n12769) );
  MUX2_X1 U15239 ( .A(n12770), .B(n12769), .S(n14728), .Z(n12771) );
  MUX2_X1 U15240 ( .A(n14611), .B(n15271), .S(n12803), .Z(n12774) );
  MUX2_X1 U15241 ( .A(n14727), .B(n14994), .S(n12823), .Z(n12773) );
  MUX2_X1 U15242 ( .A(n14726), .B(n14974), .S(n12823), .Z(n12776) );
  MUX2_X1 U15243 ( .A(n14726), .B(n14974), .S(n12803), .Z(n12775) );
  INV_X1 U15244 ( .A(n12776), .ZN(n12777) );
  MUX2_X1 U15245 ( .A(n15263), .B(n14612), .S(n12823), .Z(n12778) );
  INV_X1 U15246 ( .A(n12778), .ZN(n12780) );
  MUX2_X1 U15247 ( .A(n15263), .B(n14612), .S(n12803), .Z(n12779) );
  MUX2_X1 U15248 ( .A(n14725), .B(n14940), .S(n12823), .Z(n12785) );
  MUX2_X1 U15249 ( .A(n14725), .B(n14940), .S(n12803), .Z(n12784) );
  MUX2_X1 U15250 ( .A(n14724), .B(n14921), .S(n12803), .Z(n12789) );
  MUX2_X1 U15251 ( .A(n14724), .B(n14921), .S(n12823), .Z(n12786) );
  NAND2_X1 U15252 ( .A1(n12787), .A2(n12786), .ZN(n12794) );
  INV_X1 U15253 ( .A(n12789), .ZN(n12790) );
  AND2_X1 U15254 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  NAND2_X1 U15255 ( .A1(n12788), .A2(n12792), .ZN(n12793) );
  MUX2_X1 U15256 ( .A(n14723), .B(n14903), .S(n12823), .Z(n12796) );
  MUX2_X1 U15257 ( .A(n14723), .B(n14903), .S(n12691), .Z(n12795) );
  MUX2_X1 U15258 ( .A(n14722), .B(n14890), .S(n12691), .Z(n12798) );
  MUX2_X1 U15259 ( .A(n14722), .B(n14890), .S(n12823), .Z(n12797) );
  INV_X1 U15260 ( .A(n12798), .ZN(n12799) );
  MUX2_X1 U15261 ( .A(n14721), .B(n14880), .S(n12823), .Z(n12801) );
  MUX2_X1 U15262 ( .A(n14721), .B(n14880), .S(n12803), .Z(n12800) );
  INV_X1 U15263 ( .A(n12801), .ZN(n12802) );
  MUX2_X1 U15264 ( .A(n14839), .B(n12804), .S(n12803), .Z(n12808) );
  MUX2_X1 U15265 ( .A(n14851), .B(n14861), .S(n12823), .Z(n12805) );
  INV_X1 U15266 ( .A(n12875), .ZN(n12819) );
  XNOR2_X1 U15267 ( .A(n12862), .B(n14719), .ZN(n12825) );
  NAND2_X1 U15268 ( .A1(n12815), .A2(n12814), .ZN(n12817) );
  NAND2_X1 U15269 ( .A1(n12652), .A2(n12816), .ZN(n14866) );
  AND2_X1 U15270 ( .A1(n12817), .A2(n14866), .ZN(n12820) );
  NAND2_X1 U15271 ( .A1(n12819), .A2(n12818), .ZN(n12877) );
  NOR2_X1 U15272 ( .A1(n12862), .A2(n12823), .ZN(n12861) );
  INV_X1 U15273 ( .A(n12820), .ZN(n12860) );
  AND2_X1 U15274 ( .A1(n12822), .A2(n12821), .ZN(n12863) );
  INV_X1 U15275 ( .A(n12863), .ZN(n12871) );
  NAND2_X1 U15276 ( .A1(n12860), .A2(n12871), .ZN(n12859) );
  NAND2_X1 U15277 ( .A1(n12862), .A2(n12823), .ZN(n12868) );
  NOR2_X1 U15278 ( .A1(n12868), .A2(n14719), .ZN(n12824) );
  AOI211_X1 U15279 ( .C1(n12861), .C2(n14719), .A(n12859), .B(n12824), .ZN(
        n12874) );
  INV_X1 U15280 ( .A(n12825), .ZN(n12855) );
  NAND2_X1 U15281 ( .A1(n15105), .A2(n15525), .ZN(n12827) );
  AND2_X1 U15282 ( .A1(n7957), .A2(n12827), .ZN(n15542) );
  NAND4_X1 U15283 ( .A1(n12829), .A2(n15542), .A3(n12828), .A4(n15106), .ZN(
        n12832) );
  NOR3_X1 U15284 ( .A1(n12832), .A2(n12831), .A3(n12830), .ZN(n12836) );
  NAND4_X1 U15285 ( .A1(n12836), .A2(n12835), .A3(n12834), .A4(n12833), .ZN(
        n12838) );
  NOR3_X1 U15286 ( .A1(n12839), .A2(n12838), .A3(n12837), .ZN(n12841) );
  NAND3_X1 U15287 ( .A1(n12842), .A2(n12841), .A3(n12840), .ZN(n12843) );
  NOR2_X1 U15288 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  AND3_X1 U15289 ( .A1(n15041), .A2(n15099), .A3(n12845), .ZN(n12846) );
  XNOR2_X1 U15290 ( .A(n15200), .B(n14731), .ZN(n15055) );
  NAND4_X1 U15291 ( .A1(n12846), .A2(n15070), .A3(n15033), .A4(n15055), .ZN(
        n12847) );
  NOR2_X1 U15292 ( .A1(n14987), .A2(n12847), .ZN(n12848) );
  NAND4_X1 U15293 ( .A1(n12849), .A2(n12848), .A3(n15001), .A4(n14967), .ZN(
        n12850) );
  NOR2_X1 U15294 ( .A1(n14934), .A2(n12850), .ZN(n12852) );
  NAND4_X1 U15295 ( .A1(n14891), .A2(n12852), .A3(n14902), .A4(n12851), .ZN(
        n12853) );
  XNOR2_X1 U15296 ( .A(n14826), .B(n14841), .ZN(n12856) );
  NAND3_X1 U15297 ( .A1(n12857), .A2(n14852), .A3(n12856), .ZN(n12858) );
  XOR2_X1 U15298 ( .A(n12652), .B(n12858), .Z(n12872) );
  NOR3_X1 U15299 ( .A1(n14825), .A2(n14719), .A3(n12859), .ZN(n12869) );
  NOR3_X1 U15300 ( .A1(n12868), .A2(n14719), .A3(n12860), .ZN(n12867) );
  XNOR2_X1 U15301 ( .A(n12861), .B(n12860), .ZN(n12865) );
  INV_X1 U15302 ( .A(n14719), .ZN(n12864) );
  NOR4_X1 U15303 ( .A1(n12865), .A2(n12864), .A3(n12863), .A4(n12862), .ZN(
        n12866) );
  AOI211_X1 U15304 ( .C1(n12869), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        n12870) );
  AOI21_X1 U15305 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12876) );
  AND2_X1 U15306 ( .A1(n12877), .A2(n12876), .ZN(n12882) );
  NOR3_X1 U15307 ( .A1(n12878), .A2(n10101), .A3(n14675), .ZN(n12880) );
  OAI21_X1 U15308 ( .B1(n12881), .B2(n12651), .A(P1_B_REG_SCAN_IN), .ZN(n12879) );
  OAI22_X1 U15309 ( .A1(n12882), .A2(n12881), .B1(n12880), .B2(n12879), .ZN(
        P1_U3242) );
  INV_X1 U15310 ( .A(n12885), .ZN(n12887) );
  OAI21_X1 U15311 ( .B1(n12885), .B2(n12884), .A(n13003), .ZN(n12886) );
  XNOR2_X1 U15312 ( .A(n10160), .B(n12895), .ZN(n12889) );
  NAND2_X1 U15313 ( .A1(n12889), .A2(n13389), .ZN(n12891) );
  OAI21_X1 U15314 ( .B1(n12889), .B2(n13389), .A(n12891), .ZN(n13004) );
  INV_X1 U15315 ( .A(n12891), .ZN(n12892) );
  XNOR2_X1 U15316 ( .A(n13553), .B(n12895), .ZN(n12893) );
  NAND2_X1 U15317 ( .A1(n12893), .A2(n13010), .ZN(n12894) );
  OAI21_X1 U15318 ( .B1(n12893), .B2(n13010), .A(n12894), .ZN(n13084) );
  XNOR2_X1 U15319 ( .A(n13549), .B(n12895), .ZN(n12901) );
  NAND2_X1 U15320 ( .A1(n12901), .A2(n7457), .ZN(n12897) );
  OAI21_X1 U15321 ( .B1(n12901), .B2(n7457), .A(n12897), .ZN(n12949) );
  XNOR2_X1 U15322 ( .A(n13332), .B(n12896), .ZN(n12898) );
  INV_X1 U15323 ( .A(n12898), .ZN(n12903) );
  NAND3_X1 U15324 ( .A1(n12903), .A2(n13074), .A3(n12897), .ZN(n12907) );
  OAI22_X1 U15325 ( .A1(n13030), .A2(n7457), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13665), .ZN(n12899) );
  AOI21_X1 U15326 ( .B1(n13027), .B2(n13103), .A(n12899), .ZN(n12900) );
  OAI21_X1 U15327 ( .B1(n13341), .B2(n13088), .A(n12900), .ZN(n12905) );
  INV_X1 U15328 ( .A(n12901), .ZN(n12902) );
  NOR4_X1 U15329 ( .A1(n12903), .A2(n12902), .A3(n13100), .A4(n13334), .ZN(
        n12904) );
  AOI211_X1 U15330 ( .C1(n13098), .C2(n13340), .A(n12905), .B(n12904), .ZN(
        n12906) );
  INV_X1 U15331 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12908) );
  OAI222_X1 U15332 ( .A1(n8895), .A2(P2_U3088), .B1(n12913), .B2(n12909), .C1(
        n12908), .C2(n14562), .ZN(P2_U3306) );
  INV_X1 U15333 ( .A(n12910), .ZN(n12943) );
  OAI222_X1 U15334 ( .A1(n12913), .A2(n12943), .B1(P2_U3088), .B2(n12912), 
        .C1(n12911), .C2(n14562), .ZN(P2_U3297) );
  INV_X1 U15335 ( .A(n12914), .ZN(n12916) );
  OAI222_X1 U15336 ( .A1(n12918), .A2(n12917), .B1(n13836), .B2(n12916), .C1(
        n12915), .C2(P3_U3151), .ZN(P3_U3267) );
  INV_X1 U15337 ( .A(n12920), .ZN(n12924) );
  NAND2_X1 U15338 ( .A1(n15816), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12923) );
  INV_X1 U15339 ( .A(n12921), .ZN(n12922) );
  NAND2_X1 U15340 ( .A1(n15812), .A2(n12922), .ZN(n13323) );
  OAI211_X1 U15341 ( .C1(n12924), .C2(n13534), .A(n12923), .B(n13323), .ZN(
        n12925) );
  AOI21_X1 U15342 ( .B1(n12926), .B2(n13537), .A(n12925), .ZN(n12927) );
  OAI21_X1 U15343 ( .B1(n12919), .B2(n15816), .A(n12927), .ZN(P3_U3204) );
  INV_X1 U15344 ( .A(n12928), .ZN(n14560) );
  OAI222_X1 U15345 ( .A1(n15307), .A2(n12930), .B1(P1_U3086), .B2(n12929), 
        .C1(n15305), .C2(n14560), .ZN(P1_U3326) );
  INV_X1 U15346 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n12931) );
  OAI22_X1 U15347 ( .A1(n12932), .A2(n14385), .B1(n12931), .B2(n14396), .ZN(
        n12933) );
  AOI21_X1 U15348 ( .B1(n12934), .B2(n14401), .A(n12933), .ZN(n12939) );
  OAI21_X1 U15349 ( .B1(n14386), .B2(n12936), .A(n12935), .ZN(n12937) );
  NAND2_X1 U15350 ( .A1(n12937), .A2(n14396), .ZN(n12938) );
  OAI211_X1 U15351 ( .C1(n12940), .C2(n14371), .A(n12939), .B(n12938), .ZN(
        P2_U3237) );
  INV_X1 U15352 ( .A(n12941), .ZN(n15303) );
  OAI222_X1 U15353 ( .A1(P2_U3088), .A2(n12942), .B1(n14562), .B2(n13654), 
        .C1(n14569), .C2(n15303), .ZN(P2_U3300) );
  OAI222_X1 U15354 ( .A1(n8172), .A2(P1_U3086), .B1(n15307), .B2(n12944), .C1(
        n15305), .C2(n12943), .ZN(P1_U3325) );
  INV_X1 U15355 ( .A(n12945), .ZN(n14567) );
  OAI222_X1 U15356 ( .A1(P1_U3086), .A2(n8811), .B1(n15305), .B2(n14567), .C1(
        n12947), .C2(n12946), .ZN(P1_U3327) );
  NAND2_X1 U15357 ( .A1(n13094), .A2(n13359), .ZN(n12952) );
  AOI22_X1 U15358 ( .A1(n13027), .A2(n13349), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12951) );
  OAI211_X1 U15359 ( .C1(n13010), .C2(n13030), .A(n12952), .B(n12951), .ZN(
        n12953) );
  AOI21_X1 U15360 ( .B1(n13549), .B2(n13098), .A(n12953), .ZN(n12954) );
  OAI21_X1 U15361 ( .B1(n12955), .B2(n13100), .A(n12954), .ZN(P3_U3154) );
  OAI21_X1 U15362 ( .B1(n6917), .B2(n13521), .A(n12956), .ZN(n12957) );
  OAI21_X1 U15363 ( .B1(n12958), .B2(n13117), .A(n12957), .ZN(n12961) );
  XNOR2_X1 U15364 ( .A(n12959), .B(n13116), .ZN(n12960) );
  XNOR2_X1 U15365 ( .A(n12961), .B(n12960), .ZN(n12966) );
  NAND2_X1 U15366 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13225)
         );
  NAND2_X1 U15367 ( .A1(n13076), .A2(n13117), .ZN(n12962) );
  OAI211_X1 U15368 ( .C1(n13079), .C2(n13522), .A(n13225), .B(n12962), .ZN(
        n12963) );
  AOI21_X1 U15369 ( .B1(n13524), .B2(n13094), .A(n12963), .ZN(n12965) );
  NAND2_X1 U15370 ( .A1(n13523), .A2(n13098), .ZN(n12964) );
  OAI211_X1 U15371 ( .C1(n12966), .C2(n13100), .A(n12965), .B(n12964), .ZN(
        P3_U3155) );
  AOI22_X1 U15372 ( .A1(n13107), .A2(n13076), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12969) );
  NAND2_X1 U15373 ( .A1(n13406), .A2(n13094), .ZN(n12968) );
  OAI211_X1 U15374 ( .C1(n13402), .C2(n13079), .A(n12969), .B(n12968), .ZN(
        n12970) );
  AOI21_X1 U15375 ( .B1(n13411), .B2(n13098), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15376 ( .B1(n12972), .B2(n13100), .A(n12971), .ZN(P3_U3156) );
  AND2_X1 U15377 ( .A1(n12973), .A2(n12974), .ZN(n12977) );
  OAI211_X1 U15378 ( .C1(n12977), .C2(n12976), .A(n13074), .B(n12975), .ZN(
        n12981) );
  NAND2_X1 U15379 ( .A1(n13111), .A2(n13076), .ZN(n12978) );
  NAND2_X1 U15380 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13311)
         );
  OAI211_X1 U15381 ( .C1(n13457), .C2(n13079), .A(n12978), .B(n13311), .ZN(
        n12979) );
  AOI21_X1 U15382 ( .B1(n13458), .B2(n13094), .A(n12979), .ZN(n12980) );
  OAI211_X1 U15383 ( .C1(n13083), .C2(n13794), .A(n12981), .B(n12980), .ZN(
        P3_U3159) );
  INV_X1 U15384 ( .A(n12982), .ZN(n12983) );
  AOI21_X1 U15385 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(n12992) );
  OAI22_X1 U15386 ( .A1(n13401), .A2(n15783), .B1(n13457), .B2(n15785), .ZN(
        n13432) );
  INV_X1 U15387 ( .A(n13435), .ZN(n12987) );
  OAI22_X1 U15388 ( .A1(n12987), .A2(n13088), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12986), .ZN(n12990) );
  INV_X1 U15389 ( .A(n12988), .ZN(n13786) );
  NOR2_X1 U15390 ( .A1(n13786), .A2(n13083), .ZN(n12989) );
  AOI211_X1 U15391 ( .C1(n13086), .C2(n13432), .A(n12990), .B(n12989), .ZN(
        n12991) );
  OAI21_X1 U15392 ( .B1(n12992), .B2(n13100), .A(n12991), .ZN(P3_U3163) );
  INV_X1 U15393 ( .A(n12993), .ZN(n13064) );
  INV_X1 U15394 ( .A(n13063), .ZN(n12995) );
  NOR3_X1 U15395 ( .A1(n13064), .A2(n12995), .A3(n12994), .ZN(n12998) );
  INV_X1 U15396 ( .A(n12996), .ZN(n12997) );
  OAI21_X1 U15397 ( .B1(n12998), .B2(n12997), .A(n13074), .ZN(n13002) );
  NAND2_X1 U15398 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13188)
         );
  OAI21_X1 U15399 ( .B1(n13096), .B2(n12999), .A(n13188), .ZN(n13000) );
  AOI21_X1 U15400 ( .B1(n13531), .B2(n13094), .A(n13000), .ZN(n13001) );
  OAI211_X1 U15401 ( .C1(n7110), .C2(n13083), .A(n13002), .B(n13001), .ZN(
        P3_U3164) );
  INV_X1 U15402 ( .A(n10160), .ZN(n13015) );
  INV_X1 U15403 ( .A(n13003), .ZN(n13006) );
  INV_X1 U15404 ( .A(n13004), .ZN(n13005) );
  NOR3_X1 U15405 ( .A1(n13007), .A2(n13006), .A3(n13005), .ZN(n13009) );
  OAI21_X1 U15406 ( .B1(n13009), .B2(n13008), .A(n13074), .ZN(n13014) );
  OAI22_X1 U15407 ( .A1(n13402), .A2(n15785), .B1(n13010), .B2(n15783), .ZN(
        n13381) );
  INV_X1 U15408 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13011) );
  OAI22_X1 U15409 ( .A1(n13088), .A2(n13377), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13011), .ZN(n13012) );
  AOI21_X1 U15410 ( .B1(n13381), .B2(n13086), .A(n13012), .ZN(n13013) );
  OAI211_X1 U15411 ( .C1(n13015), .C2(n13083), .A(n13014), .B(n13013), .ZN(
        P3_U3165) );
  NAND2_X1 U15412 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  XNOR2_X1 U15413 ( .A(n13016), .B(n13019), .ZN(n13024) );
  INV_X1 U15414 ( .A(n13498), .ZN(n13021) );
  OAI22_X1 U15415 ( .A1(n13469), .A2(n15783), .B1(n13522), .B2(n15785), .ZN(
        n13491) );
  AND2_X1 U15416 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13264) );
  AOI21_X1 U15417 ( .B1(n13491), .B2(n13086), .A(n13264), .ZN(n13020) );
  OAI21_X1 U15418 ( .B1(n13021), .B2(n13088), .A(n13020), .ZN(n13022) );
  AOI21_X1 U15419 ( .B1(n13497), .B2(n13098), .A(n13022), .ZN(n13023) );
  OAI21_X1 U15420 ( .B1(n13024), .B2(n13100), .A(n13023), .ZN(P3_U3166) );
  XNOR2_X1 U15421 ( .A(n13026), .B(n13025), .ZN(n13033) );
  AND2_X1 U15422 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13285) );
  AOI21_X1 U15423 ( .B1(n13111), .B2(n13027), .A(n13285), .ZN(n13029) );
  NAND2_X1 U15424 ( .A1(n13094), .A2(n13485), .ZN(n13028) );
  OAI211_X1 U15425 ( .C1(n13479), .C2(n13030), .A(n13029), .B(n13028), .ZN(
        n13031) );
  AOI21_X1 U15426 ( .B1(n13484), .B2(n13098), .A(n13031), .ZN(n13032) );
  OAI21_X1 U15427 ( .B1(n13033), .B2(n13100), .A(n13032), .ZN(P3_U3168) );
  XNOR2_X1 U15428 ( .A(n13034), .B(n13035), .ZN(n13041) );
  AOI22_X1 U15429 ( .A1(n13108), .A2(n15796), .B1(n15799), .B2(n13110), .ZN(
        n13444) );
  OAI22_X1 U15430 ( .A1(n13444), .A2(n13096), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13036), .ZN(n13039) );
  INV_X1 U15431 ( .A(n13037), .ZN(n13790) );
  NOR2_X1 U15432 ( .A1(n13790), .A2(n13083), .ZN(n13038) );
  AOI211_X1 U15433 ( .C1(n13446), .C2(n13094), .A(n13039), .B(n13038), .ZN(
        n13040) );
  OAI21_X1 U15434 ( .B1(n13041), .B2(n13100), .A(n13040), .ZN(P3_U3173) );
  XNOR2_X1 U15435 ( .A(n13042), .B(n13117), .ZN(n13043) );
  XNOR2_X1 U15436 ( .A(n6917), .B(n13043), .ZN(n13050) );
  NAND2_X1 U15437 ( .A1(n13076), .A2(n13118), .ZN(n13044) );
  NAND2_X1 U15438 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13208)
         );
  OAI211_X1 U15439 ( .C1(n13079), .C2(n13045), .A(n13044), .B(n13208), .ZN(
        n13047) );
  NOR2_X1 U15440 ( .A1(n13814), .A2(n13083), .ZN(n13046) );
  AOI211_X1 U15441 ( .C1(n13048), .C2(n13094), .A(n13047), .B(n13046), .ZN(
        n13049) );
  OAI21_X1 U15442 ( .B1(n13050), .B2(n13100), .A(n13049), .ZN(P3_U3174) );
  INV_X1 U15443 ( .A(n13051), .ZN(n13052) );
  AOI21_X1 U15444 ( .B1(n13107), .B2(n13053), .A(n13052), .ZN(n13059) );
  AOI22_X1 U15445 ( .A1(n13108), .A2(n13076), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13055) );
  NAND2_X1 U15446 ( .A1(n13422), .A2(n13094), .ZN(n13054) );
  OAI211_X1 U15447 ( .C1(n13419), .C2(n13079), .A(n13055), .B(n13054), .ZN(
        n13056) );
  AOI21_X1 U15448 ( .B1(n13057), .B2(n13098), .A(n13056), .ZN(n13058) );
  OAI21_X1 U15449 ( .B1(n13059), .B2(n13100), .A(n13058), .ZN(P3_U3175) );
  AOI21_X1 U15450 ( .B1(n13061), .B2(n13063), .A(n13060), .ZN(n13062) );
  AOI21_X1 U15451 ( .B1(n13064), .B2(n13063), .A(n13062), .ZN(n13071) );
  INV_X1 U15452 ( .A(n13065), .ZN(n13068) );
  AOI22_X1 U15453 ( .A1(n13086), .A2(n13066), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13067) );
  OAI21_X1 U15454 ( .B1(n13088), .B2(n13068), .A(n13067), .ZN(n13069) );
  AOI21_X1 U15455 ( .B1(n13753), .B2(n13098), .A(n13069), .ZN(n13070) );
  OAI21_X1 U15456 ( .B1(n13071), .B2(n13100), .A(n13070), .ZN(P3_U3176) );
  INV_X1 U15457 ( .A(n13587), .ZN(n13473) );
  OAI21_X1 U15458 ( .B1(n13073), .B2(n13072), .A(n12973), .ZN(n13075) );
  NAND2_X1 U15459 ( .A1(n13075), .A2(n13074), .ZN(n13082) );
  NAND2_X1 U15460 ( .A1(n13112), .A2(n13076), .ZN(n13078) );
  OAI211_X1 U15461 ( .C1(n13470), .C2(n13079), .A(n13078), .B(n13077), .ZN(
        n13080) );
  AOI21_X1 U15462 ( .B1(n13471), .B2(n13094), .A(n13080), .ZN(n13081) );
  OAI211_X1 U15463 ( .C1(n13473), .C2(n13083), .A(n13082), .B(n13081), .ZN(
        P3_U3178) );
  OAI22_X1 U15464 ( .A1(n7457), .A2(n15783), .B1(n13389), .B2(n15785), .ZN(
        n13366) );
  AOI22_X1 U15465 ( .A1(n13366), .A2(n13086), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13087) );
  OAI21_X1 U15466 ( .B1(n13088), .B2(n13370), .A(n13087), .ZN(n13089) );
  AOI21_X1 U15467 ( .B1(n13553), .B2(n13098), .A(n13089), .ZN(n13090) );
  OAI21_X1 U15468 ( .B1(n13091), .B2(n13100), .A(n13090), .ZN(P3_U3180) );
  AOI21_X1 U15469 ( .B1(n13093), .B2(n13092), .A(n6626), .ZN(n13101) );
  AOI22_X1 U15470 ( .A1(n13113), .A2(n15796), .B1(n15799), .B2(n13116), .ZN(
        n13505) );
  NAND2_X1 U15471 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13249)
         );
  NAND2_X1 U15472 ( .A1(n13094), .A2(n13511), .ZN(n13095) );
  OAI211_X1 U15473 ( .C1(n13505), .C2(n13096), .A(n13249), .B(n13095), .ZN(
        n13097) );
  AOI21_X1 U15474 ( .B1(n13510), .B2(n13098), .A(n13097), .ZN(n13099) );
  OAI21_X1 U15475 ( .B1(n13101), .B2(n13100), .A(n13099), .ZN(P3_U3181) );
  MUX2_X1 U15476 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13322), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15477 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13102), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15478 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13103), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15479 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13349), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15480 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13334), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15481 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13350), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15482 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13104), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15483 ( .A(n13105), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13114), .Z(
        P3_U3515) );
  MUX2_X1 U15484 ( .A(n13106), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13114), .Z(
        P3_U3514) );
  MUX2_X1 U15485 ( .A(n13107), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13114), .Z(
        P3_U3513) );
  MUX2_X1 U15486 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13108), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15487 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13109), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15488 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13110), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15489 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13111), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15490 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13112), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15491 ( .A(n13113), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13114), .Z(
        P3_U3507) );
  MUX2_X1 U15492 ( .A(n13115), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13114), .Z(
        P3_U3506) );
  MUX2_X1 U15493 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13116), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15494 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13117), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15495 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13118), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15496 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13119), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15497 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13120), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15498 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13121), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15499 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13122), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15500 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13123), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15501 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13124), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15502 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13125), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15503 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13126), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15504 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15797), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15505 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13127), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15506 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15798), .S(P3_U3897), .Z(
        P3_U3491) );
  AND3_X1 U15507 ( .A1(n13130), .A2(n13129), .A3(n13128), .ZN(n13131) );
  OAI21_X1 U15508 ( .B1(n13132), .B2(n13131), .A(n13315), .ZN(n13148) );
  INV_X1 U15509 ( .A(n13133), .ZN(n13136) );
  NOR2_X1 U15510 ( .A1(n13313), .A2(n13134), .ZN(n13135) );
  AOI211_X1 U15511 ( .C1(n15779), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n13136), .B(
        n13135), .ZN(n13147) );
  AND3_X1 U15512 ( .A1(n13138), .A2(n13137), .A3(n6661), .ZN(n13139) );
  OAI21_X1 U15513 ( .B1(n13140), .B2(n13139), .A(n13290), .ZN(n13146) );
  AND3_X1 U15514 ( .A1(n13142), .A2(n13141), .A3(n7563), .ZN(n13143) );
  OAI21_X1 U15515 ( .B1(n13144), .B2(n13143), .A(n13300), .ZN(n13145) );
  NAND4_X1 U15516 ( .A1(n13148), .A2(n13147), .A3(n13146), .A4(n13145), .ZN(
        P3_U3188) );
  AND3_X1 U15517 ( .A1(n13151), .A2(n13150), .A3(n13149), .ZN(n13152) );
  OAI21_X1 U15518 ( .B1(n13153), .B2(n13152), .A(n13290), .ZN(n13168) );
  AND3_X1 U15519 ( .A1(n13156), .A2(n13155), .A3(n13154), .ZN(n13157) );
  OAI21_X1 U15520 ( .B1(n6657), .B2(n13157), .A(n13300), .ZN(n13167) );
  NOR2_X1 U15521 ( .A1(n13313), .A2(n13158), .ZN(n13159) );
  AOI211_X1 U15522 ( .C1(n15779), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n13160), .B(
        n13159), .ZN(n13166) );
  OAI21_X1 U15523 ( .B1(n13163), .B2(n13162), .A(n13161), .ZN(n13164) );
  NAND2_X1 U15524 ( .A1(n13164), .A2(n13315), .ZN(n13165) );
  NAND4_X1 U15525 ( .A1(n13168), .A2(n13167), .A3(n13166), .A4(n13165), .ZN(
        P3_U3190) );
  AOI21_X1 U15526 ( .B1(n13170), .B2(n13169), .A(n6619), .ZN(n13182) );
  XNOR2_X1 U15527 ( .A(n13172), .B(n13171), .ZN(n13180) );
  AND2_X1 U15528 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13173) );
  AOI21_X1 U15529 ( .B1(n15779), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n13173), 
        .ZN(n13174) );
  OAI21_X1 U15530 ( .B1(n13313), .B2(n13175), .A(n13174), .ZN(n13179) );
  AOI21_X1 U15531 ( .B1(n13701), .B2(n13176), .A(n13193), .ZN(n13177) );
  NOR2_X1 U15532 ( .A1(n13177), .A2(n13293), .ZN(n13178) );
  AOI211_X1 U15533 ( .C1(n13315), .C2(n13180), .A(n13179), .B(n13178), .ZN(
        n13181) );
  OAI21_X1 U15534 ( .B1(n13182), .B2(n13319), .A(n13181), .ZN(P3_U3193) );
  INV_X1 U15535 ( .A(n13183), .ZN(n13187) );
  NOR3_X1 U15536 ( .A1(n6619), .A2(n13185), .A3(n13184), .ZN(n13186) );
  OAI21_X1 U15537 ( .B1(n13187), .B2(n13186), .A(n13290), .ZN(n13203) );
  OAI21_X1 U15538 ( .B1(n13227), .B2(n15339), .A(n13188), .ZN(n13189) );
  AOI21_X1 U15539 ( .B1(n13190), .B2(n13229), .A(n13189), .ZN(n13202) );
  INV_X1 U15540 ( .A(n13191), .ZN(n13196) );
  NOR3_X1 U15541 ( .A1(n13194), .A2(n13193), .A3(n13192), .ZN(n13195) );
  OAI21_X1 U15542 ( .B1(n13196), .B2(n13195), .A(n13300), .ZN(n13201) );
  OAI211_X1 U15543 ( .C1(n13199), .C2(n13198), .A(n13197), .B(n13315), .ZN(
        n13200) );
  NAND4_X1 U15544 ( .A1(n13203), .A2(n13202), .A3(n13201), .A4(n13200), .ZN(
        P3_U3194) );
  AOI21_X1 U15545 ( .B1(n13748), .B2(n13204), .A(n13233), .ZN(n13218) );
  INV_X1 U15546 ( .A(n13205), .ZN(n13206) );
  NOR2_X1 U15547 ( .A1(n13206), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13207) );
  OAI21_X1 U15548 ( .B1(n13207), .B2(n13222), .A(n13290), .ZN(n13217) );
  INV_X1 U15549 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15402) );
  OAI21_X1 U15550 ( .B1(n13227), .B2(n15402), .A(n13208), .ZN(n13214) );
  AOI21_X1 U15551 ( .B1(n13211), .B2(n13210), .A(n13209), .ZN(n13212) );
  NOR2_X1 U15552 ( .A1(n13212), .A2(n13282), .ZN(n13213) );
  AOI211_X1 U15553 ( .C1(n13229), .C2(n13215), .A(n13214), .B(n13213), .ZN(
        n13216) );
  OAI211_X1 U15554 ( .C1(n13218), .C2(n13293), .A(n13217), .B(n13216), .ZN(
        P3_U3195) );
  INV_X1 U15555 ( .A(n13219), .ZN(n13224) );
  NOR3_X1 U15556 ( .A1(n13222), .A2(n13221), .A3(n13220), .ZN(n13223) );
  OAI21_X1 U15557 ( .B1(n13224), .B2(n13223), .A(n13290), .ZN(n13242) );
  INV_X1 U15558 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13226) );
  OAI21_X1 U15559 ( .B1(n13227), .B2(n13226), .A(n13225), .ZN(n13228) );
  AOI21_X1 U15560 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(n13241) );
  NOR3_X1 U15561 ( .A1(n13233), .A2(n13232), .A3(n13231), .ZN(n13234) );
  OAI21_X1 U15562 ( .B1(n13235), .B2(n13234), .A(n13300), .ZN(n13240) );
  OAI211_X1 U15563 ( .C1(n13238), .C2(n13237), .A(n13236), .B(n13315), .ZN(
        n13239) );
  NAND4_X1 U15564 ( .A1(n13242), .A2(n13241), .A3(n13240), .A4(n13239), .ZN(
        P3_U3196) );
  OAI21_X1 U15565 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n13244), .A(n13243), 
        .ZN(n13252) );
  AOI211_X1 U15566 ( .C1(n13247), .C2(n13246), .A(n13282), .B(n13245), .ZN(
        n13251) );
  NAND2_X1 U15567 ( .A1(n15779), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n13248) );
  OAI211_X1 U15568 ( .C1(n6997), .C2(n13313), .A(n13249), .B(n13248), .ZN(
        n13250) );
  AOI211_X1 U15569 ( .C1(n13252), .C2(n13290), .A(n13251), .B(n13250), .ZN(
        n13257) );
  OAI21_X1 U15570 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13254), .A(n13253), 
        .ZN(n13255) );
  NAND2_X1 U15571 ( .A1(n13255), .A2(n13300), .ZN(n13256) );
  NAND2_X1 U15572 ( .A1(n13257), .A2(n13256), .ZN(P3_U3197) );
  OAI21_X1 U15573 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n13269) );
  AOI211_X1 U15574 ( .C1(n13263), .C2(n13262), .A(n13282), .B(n13261), .ZN(
        n13268) );
  AOI21_X1 U15575 ( .B1(n15779), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13264), 
        .ZN(n13265) );
  OAI21_X1 U15576 ( .B1(n13313), .B2(n13266), .A(n13265), .ZN(n13267) );
  AOI211_X1 U15577 ( .C1(n13269), .C2(n13290), .A(n13268), .B(n13267), .ZN(
        n13275) );
  OAI21_X1 U15578 ( .B1(n13272), .B2(n13271), .A(n13270), .ZN(n13273) );
  NAND2_X1 U15579 ( .A1(n13273), .A2(n13300), .ZN(n13274) );
  NAND2_X1 U15580 ( .A1(n13275), .A2(n13274), .ZN(P3_U3198) );
  INV_X1 U15581 ( .A(n13276), .ZN(n13277) );
  AOI21_X1 U15582 ( .B1(n13730), .B2(n13278), .A(n13277), .ZN(n13294) );
  OAI21_X1 U15583 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13280), .A(n13279), 
        .ZN(n13291) );
  AOI211_X1 U15584 ( .C1(n13284), .C2(n13283), .A(n13282), .B(n13281), .ZN(
        n13289) );
  AOI21_X1 U15585 ( .B1(n15779), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13285), 
        .ZN(n13286) );
  OAI21_X1 U15586 ( .B1(n13313), .B2(n13287), .A(n13286), .ZN(n13288) );
  AOI211_X1 U15587 ( .C1(n13291), .C2(n13290), .A(n13289), .B(n13288), .ZN(
        n13292) );
  OAI21_X1 U15588 ( .B1(n13294), .B2(n13293), .A(n13292), .ZN(P3_U3199) );
  NAND2_X1 U15589 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  XNOR2_X1 U15590 ( .A(n13312), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13306) );
  XNOR2_X1 U15591 ( .A(n13297), .B(n13306), .ZN(n13320) );
  INV_X1 U15592 ( .A(n13298), .ZN(n13299) );
  XNOR2_X1 U15593 ( .A(n13312), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U15594 ( .A1(n13301), .A2(n13300), .ZN(n13318) );
  AOI21_X1 U15595 ( .B1(n13304), .B2(n13303), .A(n13302), .ZN(n13309) );
  MUX2_X1 U15596 ( .A(n13307), .B(n13306), .S(n13305), .Z(n13308) );
  XNOR2_X1 U15597 ( .A(n13309), .B(n13308), .ZN(n13316) );
  NAND2_X1 U15598 ( .A1(n15779), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13310) );
  OAI211_X1 U15599 ( .C1(n13313), .C2(n13312), .A(n13311), .B(n13310), .ZN(
        n13314) );
  AOI21_X1 U15600 ( .B1(n13316), .B2(n13315), .A(n13314), .ZN(n13317) );
  OAI211_X1 U15601 ( .C1(n13320), .C2(n13319), .A(n13318), .B(n13317), .ZN(
        P3_U3201) );
  NAND2_X1 U15602 ( .A1(n13322), .A2(n13321), .ZN(n13756) );
  OAI21_X1 U15603 ( .B1(n15816), .B2(n13756), .A(n13323), .ZN(n13325) );
  AOI21_X1 U15604 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15816), .A(n13325), 
        .ZN(n13324) );
  OAI21_X1 U15605 ( .B1(n13758), .B2(n13534), .A(n13324), .ZN(P3_U3202) );
  AOI21_X1 U15606 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15816), .A(n13325), 
        .ZN(n13326) );
  OAI21_X1 U15607 ( .B1(n13327), .B2(n13534), .A(n13326), .ZN(P3_U3203) );
  INV_X1 U15608 ( .A(n13546), .ZN(n13346) );
  NAND2_X1 U15609 ( .A1(n13334), .A2(n15799), .ZN(n13335) );
  OAI21_X1 U15610 ( .B1(n13336), .B2(n15783), .A(n13335), .ZN(n13337) );
  INV_X1 U15611 ( .A(n13341), .ZN(n13342) );
  AOI22_X1 U15612 ( .A1(n15816), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15812), 
        .B2(n13342), .ZN(n13343) );
  OAI21_X1 U15613 ( .B1(n13767), .B2(n13534), .A(n13343), .ZN(n13344) );
  AOI21_X1 U15614 ( .B1(n13545), .B2(n15813), .A(n13344), .ZN(n13345) );
  OAI21_X1 U15615 ( .B1(n13346), .B2(n13528), .A(n13345), .ZN(P3_U3205) );
  INV_X1 U15616 ( .A(n13355), .ZN(n13356) );
  AOI21_X1 U15617 ( .B1(n13358), .B2(n13357), .A(n13356), .ZN(n13552) );
  INV_X1 U15618 ( .A(n13552), .ZN(n13363) );
  INV_X1 U15619 ( .A(n13549), .ZN(n13361) );
  AOI22_X1 U15620 ( .A1(n15816), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15812), 
        .B2(n13359), .ZN(n13360) );
  OAI21_X1 U15621 ( .B1(n13361), .B2(n13534), .A(n13360), .ZN(n13362) );
  AOI21_X1 U15622 ( .B1(n13363), .B2(n13537), .A(n13362), .ZN(n13364) );
  OAI21_X1 U15623 ( .B1(n15816), .B2(n13551), .A(n13364), .ZN(P3_U3206) );
  XNOR2_X1 U15624 ( .A(n13365), .B(n13368), .ZN(n13367) );
  AOI21_X1 U15625 ( .B1(n13367), .B2(n15801), .A(n13366), .ZN(n13555) );
  XOR2_X1 U15626 ( .A(n13369), .B(n13368), .Z(n13554) );
  INV_X1 U15627 ( .A(n13370), .ZN(n13371) );
  AOI22_X1 U15628 ( .A1(n15816), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15812), 
        .B2(n13371), .ZN(n13372) );
  OAI21_X1 U15629 ( .B1(n7369), .B2(n13534), .A(n13372), .ZN(n13373) );
  AOI21_X1 U15630 ( .B1(n13554), .B2(n13537), .A(n13373), .ZN(n13374) );
  OAI21_X1 U15631 ( .B1(n15816), .B2(n13555), .A(n13374), .ZN(P3_U3207) );
  XNOR2_X1 U15632 ( .A(n13376), .B(n13375), .ZN(n13559) );
  INV_X1 U15633 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13378) );
  OAI22_X1 U15634 ( .A1(n15813), .A2(n13378), .B1(n13377), .B2(n13532), .ZN(
        n13385) );
  AOI21_X1 U15635 ( .B1(n13380), .B2(n13379), .A(n15789), .ZN(n13383) );
  AOI21_X1 U15636 ( .B1(n13383), .B2(n13382), .A(n13381), .ZN(n13558) );
  NOR2_X1 U15637 ( .A1(n13558), .A2(n15816), .ZN(n13384) );
  OAI21_X1 U15638 ( .B1(n13528), .B2(n13559), .A(n13386), .ZN(P3_U3208) );
  XNOR2_X1 U15639 ( .A(n13387), .B(n6586), .ZN(n13560) );
  XNOR2_X1 U15640 ( .A(n13388), .B(n6586), .ZN(n13391) );
  OAI22_X1 U15641 ( .A1(n13419), .A2(n15785), .B1(n13389), .B2(n15783), .ZN(
        n13390) );
  AOI21_X1 U15642 ( .B1(n13391), .B2(n15801), .A(n13390), .ZN(n13392) );
  OAI21_X1 U15643 ( .B1(n13560), .B2(n15805), .A(n13392), .ZN(n13561) );
  NAND2_X1 U15644 ( .A1(n13561), .A2(n15813), .ZN(n13397) );
  OAI22_X1 U15645 ( .A1(n13394), .A2(n13532), .B1(n15813), .B2(n13393), .ZN(
        n13395) );
  AOI21_X1 U15646 ( .B1(n10238), .B2(n13410), .A(n13395), .ZN(n13396) );
  OAI211_X1 U15647 ( .C1(n13560), .C2(n13414), .A(n13397), .B(n13396), .ZN(
        P3_U3209) );
  XNOR2_X1 U15648 ( .A(n13398), .B(n13399), .ZN(n13565) );
  XNOR2_X1 U15649 ( .A(n13400), .B(n13399), .ZN(n13404) );
  OAI22_X1 U15650 ( .A1(n13402), .A2(n15783), .B1(n13401), .B2(n15785), .ZN(
        n13403) );
  AOI21_X1 U15651 ( .B1(n13404), .B2(n15801), .A(n13403), .ZN(n13405) );
  OAI21_X1 U15652 ( .B1(n13565), .B2(n15805), .A(n13405), .ZN(n13566) );
  NAND2_X1 U15653 ( .A1(n13566), .A2(n15813), .ZN(n13413) );
  INV_X1 U15654 ( .A(n13406), .ZN(n13408) );
  OAI22_X1 U15655 ( .A1(n13408), .A2(n13532), .B1(n15813), .B2(n13407), .ZN(
        n13409) );
  AOI21_X1 U15656 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13412) );
  OAI211_X1 U15657 ( .C1(n13565), .C2(n13414), .A(n13413), .B(n13412), .ZN(
        P3_U3210) );
  XNOR2_X1 U15658 ( .A(n13416), .B(n13415), .ZN(n13417) );
  OAI222_X1 U15659 ( .A1(n15783), .A2(n13419), .B1(n15785), .B2(n13418), .C1(
        n15789), .C2(n13417), .ZN(n13570) );
  INV_X1 U15660 ( .A(n13570), .ZN(n13426) );
  XNOR2_X1 U15661 ( .A(n13420), .B(n13421), .ZN(n13571) );
  AOI22_X1 U15662 ( .A1(n13422), .A2(n15812), .B1(n15816), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U15663 ( .B1(n13782), .B2(n13534), .A(n13423), .ZN(n13424) );
  AOI21_X1 U15664 ( .B1(n13571), .B2(n13537), .A(n13424), .ZN(n13425) );
  OAI21_X1 U15665 ( .B1(n13426), .B2(n15816), .A(n13425), .ZN(P3_U3211) );
  XNOR2_X1 U15666 ( .A(n13427), .B(n13430), .ZN(n13575) );
  INV_X1 U15667 ( .A(n13575), .ZN(n13439) );
  AND2_X1 U15668 ( .A1(n13441), .A2(n13428), .ZN(n13431) );
  OAI21_X1 U15669 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13433) );
  AOI21_X1 U15670 ( .B1(n13433), .B2(n15801), .A(n13432), .ZN(n13434) );
  INV_X1 U15671 ( .A(n13434), .ZN(n13574) );
  AOI22_X1 U15672 ( .A1(n13435), .A2(n15812), .B1(n15816), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U15673 ( .B1(n13786), .B2(n13534), .A(n13436), .ZN(n13437) );
  AOI21_X1 U15674 ( .B1(n13574), .B2(n15813), .A(n13437), .ZN(n13438) );
  OAI21_X1 U15675 ( .B1(n13439), .B2(n13528), .A(n13438), .ZN(P3_U3212) );
  XOR2_X1 U15676 ( .A(n13440), .B(n13442), .Z(n13579) );
  INV_X1 U15677 ( .A(n13579), .ZN(n13450) );
  OAI211_X1 U15678 ( .C1(n13443), .C2(n13442), .A(n13441), .B(n15801), .ZN(
        n13445) );
  NAND2_X1 U15679 ( .A1(n13445), .A2(n13444), .ZN(n13578) );
  AOI22_X1 U15680 ( .A1(n13446), .A2(n15812), .B1(n15816), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n13447) );
  OAI21_X1 U15681 ( .B1(n13790), .B2(n13534), .A(n13447), .ZN(n13448) );
  AOI21_X1 U15682 ( .B1(n13578), .B2(n15813), .A(n13448), .ZN(n13449) );
  OAI21_X1 U15683 ( .B1(n13450), .B2(n13528), .A(n13449), .ZN(P3_U3213) );
  NAND2_X1 U15684 ( .A1(n13451), .A2(n13452), .ZN(n13453) );
  XOR2_X1 U15685 ( .A(n13454), .B(n13453), .Z(n13583) );
  INV_X1 U15686 ( .A(n13583), .ZN(n13462) );
  XNOR2_X1 U15687 ( .A(n13455), .B(n13454), .ZN(n13456) );
  OAI222_X1 U15688 ( .A1(n15783), .A2(n13457), .B1(n15785), .B2(n13480), .C1(
        n13456), .C2(n15789), .ZN(n13582) );
  AOI22_X1 U15689 ( .A1(n15816), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13458), 
        .B2(n15812), .ZN(n13459) );
  OAI21_X1 U15690 ( .B1(n13794), .B2(n13534), .A(n13459), .ZN(n13460) );
  AOI21_X1 U15691 ( .B1(n13582), .B2(n15813), .A(n13460), .ZN(n13461) );
  OAI21_X1 U15692 ( .B1(n13462), .B2(n13528), .A(n13461), .ZN(P3_U3214) );
  XOR2_X1 U15693 ( .A(n13463), .B(n13467), .Z(n13589) );
  INV_X1 U15694 ( .A(n13464), .ZN(n13465) );
  AOI21_X1 U15695 ( .B1(n13467), .B2(n13466), .A(n13465), .ZN(n13468) );
  OAI222_X1 U15696 ( .A1(n15783), .A2(n13470), .B1(n15785), .B2(n13469), .C1(
        n15789), .C2(n13468), .ZN(n13586) );
  AOI22_X1 U15697 ( .A1(n15816), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15812), 
        .B2(n13471), .ZN(n13472) );
  OAI21_X1 U15698 ( .B1(n13473), .B2(n13534), .A(n13472), .ZN(n13474) );
  AOI21_X1 U15699 ( .B1(n13586), .B2(n15813), .A(n13474), .ZN(n13475) );
  OAI21_X1 U15700 ( .B1(n13589), .B2(n13528), .A(n13475), .ZN(P3_U3215) );
  XNOR2_X1 U15701 ( .A(n13476), .B(n13477), .ZN(n13478) );
  OAI222_X1 U15702 ( .A1(n15783), .A2(n13480), .B1(n15785), .B2(n13479), .C1(
        n13478), .C2(n15789), .ZN(n13728) );
  INV_X1 U15703 ( .A(n13728), .ZN(n13489) );
  OAI21_X1 U15704 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(n13729) );
  INV_X1 U15705 ( .A(n13484), .ZN(n13799) );
  AOI22_X1 U15706 ( .A1(n15816), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15812), 
        .B2(n13485), .ZN(n13486) );
  OAI21_X1 U15707 ( .B1(n13799), .B2(n13534), .A(n13486), .ZN(n13487) );
  AOI21_X1 U15708 ( .B1(n13729), .B2(n13537), .A(n13487), .ZN(n13488) );
  OAI21_X1 U15709 ( .B1(n15816), .B2(n13489), .A(n13488), .ZN(P3_U3216) );
  XNOR2_X1 U15710 ( .A(n13490), .B(n13495), .ZN(n13493) );
  INV_X1 U15711 ( .A(n13491), .ZN(n13492) );
  OAI21_X1 U15712 ( .B1(n13493), .B2(n15789), .A(n13492), .ZN(n13732) );
  INV_X1 U15713 ( .A(n13732), .ZN(n13502) );
  OAI21_X1 U15714 ( .B1(n13496), .B2(n13495), .A(n13494), .ZN(n13733) );
  INV_X1 U15715 ( .A(n13497), .ZN(n13803) );
  AOI22_X1 U15716 ( .A1(n15816), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15812), 
        .B2(n13498), .ZN(n13499) );
  OAI21_X1 U15717 ( .B1(n13803), .B2(n13534), .A(n13499), .ZN(n13500) );
  AOI21_X1 U15718 ( .B1(n13733), .B2(n13537), .A(n13500), .ZN(n13501) );
  OAI21_X1 U15719 ( .B1(n15816), .B2(n13502), .A(n13501), .ZN(P3_U3217) );
  XNOR2_X1 U15720 ( .A(n13503), .B(n13504), .ZN(n13506) );
  OAI21_X1 U15721 ( .B1(n13506), .B2(n15789), .A(n13505), .ZN(n13736) );
  INV_X1 U15722 ( .A(n13736), .ZN(n13515) );
  OAI21_X1 U15723 ( .B1(n13509), .B2(n13508), .A(n13507), .ZN(n13737) );
  AOI22_X1 U15724 ( .A1(n15816), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15812), 
        .B2(n13511), .ZN(n13512) );
  OAI21_X1 U15725 ( .B1(n7713), .B2(n13534), .A(n13512), .ZN(n13513) );
  AOI21_X1 U15726 ( .B1(n13737), .B2(n13537), .A(n13513), .ZN(n13514) );
  OAI21_X1 U15727 ( .B1(n15816), .B2(n13515), .A(n13514), .ZN(P3_U3218) );
  XNOR2_X1 U15728 ( .A(n13516), .B(n13517), .ZN(n13741) );
  INV_X1 U15729 ( .A(n13741), .ZN(n13529) );
  XNOR2_X1 U15730 ( .A(n13518), .B(n13519), .ZN(n13520) );
  OAI222_X1 U15731 ( .A1(n15783), .A2(n13522), .B1(n15785), .B2(n13521), .C1(
        n13520), .C2(n15789), .ZN(n13740) );
  INV_X1 U15732 ( .A(n13523), .ZN(n13810) );
  AOI22_X1 U15733 ( .A1(n15816), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15812), 
        .B2(n13524), .ZN(n13525) );
  OAI21_X1 U15734 ( .B1(n13810), .B2(n13534), .A(n13525), .ZN(n13526) );
  AOI21_X1 U15735 ( .B1(n13740), .B2(n15813), .A(n13526), .ZN(n13527) );
  OAI21_X1 U15736 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(P3_U3219) );
  MUX2_X1 U15737 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n13530), .S(n15813), .Z(
        n13536) );
  INV_X1 U15738 ( .A(n13531), .ZN(n13533) );
  OAI22_X1 U15739 ( .A1(n7110), .A2(n13534), .B1(n13533), .B2(n13532), .ZN(
        n13535) );
  AOI211_X1 U15740 ( .C1(n13538), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13539) );
  INV_X1 U15741 ( .A(n13539), .ZN(P3_U3221) );
  NOR2_X1 U15742 ( .A1(n10255), .A2(n13756), .ZN(n13541) );
  AOI21_X1 U15743 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n10255), .A(n13541), 
        .ZN(n13540) );
  OAI21_X1 U15744 ( .B1(n13758), .B2(n13750), .A(n13540), .ZN(P3_U3490) );
  INV_X1 U15745 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13544) );
  NAND2_X1 U15746 ( .A1(n13760), .A2(n13754), .ZN(n13543) );
  INV_X1 U15747 ( .A(n13541), .ZN(n13542) );
  OAI211_X1 U15748 ( .C1(n15873), .C2(n13544), .A(n13543), .B(n13542), .ZN(
        P3_U3489) );
  INV_X1 U15749 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13547) );
  MUX2_X1 U15750 ( .A(n13766), .B(n13547), .S(n10255), .Z(n13548) );
  NAND2_X1 U15751 ( .A1(n13549), .A2(n15836), .ZN(n13550) );
  OAI211_X1 U15752 ( .C1(n13552), .C2(n13745), .A(n13551), .B(n13550), .ZN(
        n13768) );
  MUX2_X1 U15753 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13768), .S(n15873), .Z(
        P3_U3486) );
  AOI22_X1 U15754 ( .A1(n13554), .A2(n15851), .B1(n15836), .B2(n13553), .ZN(
        n13556) );
  NAND2_X1 U15755 ( .A1(n13556), .A2(n13555), .ZN(n13769) );
  MUX2_X1 U15756 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13769), .S(n15873), .Z(
        P3_U3485) );
  NAND2_X1 U15757 ( .A1(n10160), .A2(n15836), .ZN(n13557) );
  OAI211_X1 U15758 ( .C1(n13559), .C2(n13745), .A(n13558), .B(n13557), .ZN(
        n13770) );
  MUX2_X1 U15759 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13770), .S(n15873), .Z(
        P3_U3484) );
  INV_X1 U15760 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13563) );
  INV_X1 U15761 ( .A(n13560), .ZN(n13562) );
  AOI21_X1 U15762 ( .B1(n15856), .B2(n13562), .A(n13561), .ZN(n13771) );
  MUX2_X1 U15763 ( .A(n13563), .B(n13771), .S(n15873), .Z(n13564) );
  OAI21_X1 U15764 ( .B1(n13774), .B2(n13750), .A(n13564), .ZN(P3_U3483) );
  INV_X1 U15765 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13568) );
  INV_X1 U15766 ( .A(n13565), .ZN(n13567) );
  AOI21_X1 U15767 ( .B1(n15856), .B2(n13567), .A(n13566), .ZN(n13775) );
  MUX2_X1 U15768 ( .A(n13568), .B(n13775), .S(n15873), .Z(n13569) );
  OAI21_X1 U15769 ( .B1(n13778), .B2(n13750), .A(n13569), .ZN(P3_U3482) );
  INV_X1 U15770 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13572) );
  AOI21_X1 U15771 ( .B1(n15851), .B2(n13571), .A(n13570), .ZN(n13779) );
  MUX2_X1 U15772 ( .A(n13572), .B(n13779), .S(n15873), .Z(n13573) );
  OAI21_X1 U15773 ( .B1(n13782), .B2(n13750), .A(n13573), .ZN(P3_U3481) );
  INV_X1 U15774 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13576) );
  AOI21_X1 U15775 ( .B1(n13575), .B2(n15851), .A(n13574), .ZN(n13783) );
  MUX2_X1 U15776 ( .A(n13576), .B(n13783), .S(n15873), .Z(n13577) );
  OAI21_X1 U15777 ( .B1(n13786), .B2(n13750), .A(n13577), .ZN(P3_U3480) );
  INV_X1 U15778 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13580) );
  AOI21_X1 U15779 ( .B1(n13579), .B2(n15851), .A(n13578), .ZN(n13787) );
  MUX2_X1 U15780 ( .A(n13580), .B(n13787), .S(n15873), .Z(n13581) );
  OAI21_X1 U15781 ( .B1(n13790), .B2(n13750), .A(n13581), .ZN(P3_U3479) );
  INV_X1 U15782 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13584) );
  AOI21_X1 U15783 ( .B1(n13583), .B2(n15851), .A(n13582), .ZN(n13791) );
  MUX2_X1 U15784 ( .A(n13584), .B(n13791), .S(n15873), .Z(n13585) );
  OAI21_X1 U15785 ( .B1(n13750), .B2(n13794), .A(n13585), .ZN(P3_U3478) );
  AOI21_X1 U15786 ( .B1(n15836), .B2(n13587), .A(n13586), .ZN(n13588) );
  OAI21_X1 U15787 ( .B1(n13745), .B2(n13589), .A(n13588), .ZN(n13795) );
  MUX2_X1 U15788 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13795), .S(n15873), .Z(
        n13727) );
  XNOR2_X1 U15789 ( .A(n13590), .B(keyinput14), .ZN(n13597) );
  XNOR2_X1 U15790 ( .A(n13591), .B(keyinput47), .ZN(n13596) );
  XNOR2_X1 U15791 ( .A(n13592), .B(keyinput1), .ZN(n13595) );
  XNOR2_X1 U15792 ( .A(n13593), .B(keyinput25), .ZN(n13594) );
  NOR4_X1 U15793 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13619) );
  XOR2_X1 U15794 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput37), .Z(n13602) );
  XNOR2_X1 U15795 ( .A(n13797), .B(keyinput48), .ZN(n13601) );
  XNOR2_X1 U15796 ( .A(n13598), .B(keyinput34), .ZN(n13600) );
  XNOR2_X1 U15797 ( .A(n14122), .B(keyinput0), .ZN(n13599) );
  NOR4_X1 U15798 ( .A1(n13602), .A2(n13601), .A3(n13600), .A4(n13599), .ZN(
        n13618) );
  XOR2_X1 U15799 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput40), .Z(n13608) );
  XOR2_X1 U15800 ( .A(P3_REG1_REG_11__SCAN_IN), .B(keyinput20), .Z(n13607) );
  XNOR2_X1 U15801 ( .A(n13603), .B(keyinput3), .ZN(n13606) );
  XNOR2_X1 U15802 ( .A(n13604), .B(keyinput41), .ZN(n13605) );
  NOR4_X1 U15803 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13617) );
  XNOR2_X1 U15804 ( .A(n13609), .B(keyinput51), .ZN(n13615) );
  XNOR2_X1 U15805 ( .A(n13610), .B(keyinput33), .ZN(n13614) );
  XNOR2_X1 U15806 ( .A(n13695), .B(keyinput26), .ZN(n13613) );
  XNOR2_X1 U15807 ( .A(n13611), .B(keyinput29), .ZN(n13612) );
  NOR4_X1 U15808 ( .A1(n13615), .A2(n13614), .A3(n13613), .A4(n13612), .ZN(
        n13616) );
  NAND4_X1 U15809 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13629) );
  AOI22_X1 U15810 ( .A1(n15335), .A2(keyinput7), .B1(n13857), .B2(keyinput19), 
        .ZN(n13620) );
  OAI221_X1 U15811 ( .B1(n15335), .B2(keyinput7), .C1(n13857), .C2(keyinput19), 
        .A(n13620), .ZN(n13628) );
  XOR2_X1 U15812 ( .A(n15536), .B(keyinput24), .Z(n13625) );
  XOR2_X1 U15813 ( .A(n13621), .B(keyinput54), .Z(n13624) );
  XNOR2_X1 U15814 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput6), .ZN(n13623)
         );
  XNOR2_X1 U15815 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput22), .ZN(n13622) );
  NAND4_X1 U15816 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13627) );
  XNOR2_X1 U15817 ( .A(n15535), .B(keyinput32), .ZN(n13626) );
  OR4_X1 U15818 ( .A1(n13629), .A2(n13628), .A3(n13627), .A4(n13626), .ZN(
        n13663) );
  INV_X1 U15819 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15845) );
  INV_X1 U15820 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U15821 ( .A1(n15845), .A2(keyinput17), .B1(n15755), .B2(keyinput13), 
        .ZN(n13630) );
  OAI221_X1 U15822 ( .B1(n15845), .B2(keyinput17), .C1(n15755), .C2(keyinput13), .A(n13630), .ZN(n13640) );
  INV_X1 U15823 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15738) );
  INV_X1 U15824 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15717) );
  AOI22_X1 U15825 ( .A1(n15738), .A2(keyinput43), .B1(n15717), .B2(keyinput31), 
        .ZN(n13631) );
  OAI221_X1 U15826 ( .B1(n15738), .B2(keyinput43), .C1(n15717), .C2(keyinput31), .A(n13631), .ZN(n13639) );
  AOI22_X1 U15827 ( .A1(n15537), .A2(keyinput42), .B1(n13633), .B2(keyinput62), 
        .ZN(n13632) );
  OAI221_X1 U15828 ( .B1(n15537), .B2(keyinput42), .C1(n13633), .C2(keyinput62), .A(n13632), .ZN(n13638) );
  INV_X1 U15829 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13635) );
  AOI22_X1 U15830 ( .A1(n13636), .A2(keyinput53), .B1(n13635), .B2(keyinput30), 
        .ZN(n13634) );
  OAI221_X1 U15831 ( .B1(n13636), .B2(keyinput53), .C1(n13635), .C2(keyinput30), .A(n13634), .ZN(n13637) );
  OR4_X1 U15832 ( .A1(n13640), .A2(n13639), .A3(n13638), .A4(n13637), .ZN(
        n13662) );
  INV_X1 U15833 ( .A(P1_WR_REG_SCAN_IN), .ZN(n13642) );
  AOI22_X1 U15834 ( .A1(n13696), .A2(keyinput50), .B1(keyinput49), .B2(n13642), 
        .ZN(n13641) );
  OAI221_X1 U15835 ( .B1(n13696), .B2(keyinput50), .C1(n13642), .C2(keyinput49), .A(n13641), .ZN(n13645) );
  AOI22_X1 U15836 ( .A1(n7363), .A2(keyinput23), .B1(n10879), .B2(keyinput46), 
        .ZN(n13643) );
  OAI221_X1 U15837 ( .B1(n7363), .B2(keyinput23), .C1(n10879), .C2(keyinput46), 
        .A(n13643), .ZN(n13644) );
  NOR2_X1 U15838 ( .A1(n13645), .A2(n13644), .ZN(n13660) );
  XNOR2_X1 U15839 ( .A(keyinput45), .B(n12010), .ZN(n13647) );
  XNOR2_X1 U15840 ( .A(keyinput15), .B(n14874), .ZN(n13646) );
  NOR2_X1 U15841 ( .A1(n13647), .A2(n13646), .ZN(n13659) );
  AOI22_X1 U15842 ( .A1(n14808), .A2(keyinput60), .B1(n13649), .B2(keyinput36), 
        .ZN(n13648) );
  OAI221_X1 U15843 ( .B1(n14808), .B2(keyinput60), .C1(n13649), .C2(keyinput36), .A(n13648), .ZN(n13652) );
  AOI22_X1 U15844 ( .A1(n14799), .A2(keyinput61), .B1(n13788), .B2(keyinput5), 
        .ZN(n13650) );
  OAI221_X1 U15845 ( .B1(n14799), .B2(keyinput61), .C1(n13788), .C2(keyinput5), 
        .A(n13650), .ZN(n13651) );
  NOR2_X1 U15846 ( .A1(n13652), .A2(n13651), .ZN(n13658) );
  AOI22_X1 U15847 ( .A1(n13655), .A2(keyinput28), .B1(n13654), .B2(keyinput35), 
        .ZN(n13653) );
  OAI221_X1 U15848 ( .B1(n13655), .B2(keyinput28), .C1(n13654), .C2(keyinput35), .A(n13653), .ZN(n13656) );
  INV_X1 U15849 ( .A(n13656), .ZN(n13657) );
  NAND4_X1 U15850 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  NOR3_X1 U15851 ( .A1(n13663), .A2(n13662), .A3(n13661), .ZN(n13725) );
  AOI22_X1 U15852 ( .A1(n13665), .A2(keyinput39), .B1(n14134), .B2(keyinput2), 
        .ZN(n13664) );
  OAI221_X1 U15853 ( .B1(n13665), .B2(keyinput39), .C1(n14134), .C2(keyinput2), 
        .A(n13664), .ZN(n13674) );
  INV_X1 U15854 ( .A(P2_WR_REG_SCAN_IN), .ZN(n13668) );
  AOI22_X1 U15855 ( .A1(n13668), .A2(keyinput56), .B1(n13667), .B2(keyinput52), 
        .ZN(n13666) );
  OAI221_X1 U15856 ( .B1(n13668), .B2(keyinput56), .C1(n13667), .C2(keyinput52), .A(n13666), .ZN(n13673) );
  AOI22_X1 U15857 ( .A1(n15339), .A2(keyinput38), .B1(n11060), .B2(keyinput55), 
        .ZN(n13669) );
  OAI221_X1 U15858 ( .B1(n15339), .B2(keyinput38), .C1(n11060), .C2(keyinput55), .A(n13669), .ZN(n13672) );
  AOI22_X1 U15859 ( .A1(n15261), .A2(keyinput11), .B1(n15539), .B2(keyinput10), 
        .ZN(n13670) );
  OAI221_X1 U15860 ( .B1(n15261), .B2(keyinput11), .C1(n15539), .C2(keyinput10), .A(n13670), .ZN(n13671) );
  NOR4_X1 U15861 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13724) );
  INV_X1 U15862 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15821) );
  AOI22_X1 U15863 ( .A1(n15821), .A2(keyinput8), .B1(keyinput21), .B2(n15316), 
        .ZN(n13675) );
  OAI221_X1 U15864 ( .B1(n15821), .B2(keyinput8), .C1(n15316), .C2(keyinput21), 
        .A(n13675), .ZN(n13692) );
  AOI22_X1 U15865 ( .A1(n13784), .A2(keyinput12), .B1(keyinput59), .B2(n15313), 
        .ZN(n13676) );
  OAI221_X1 U15866 ( .B1(n13784), .B2(keyinput12), .C1(n15313), .C2(keyinput59), .A(n13676), .ZN(n13682) );
  INV_X1 U15867 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U15868 ( .A1(n15538), .A2(keyinput18), .B1(n13693), .B2(keyinput27), 
        .ZN(n13677) );
  OAI221_X1 U15869 ( .B1(n15538), .B2(keyinput18), .C1(n13693), .C2(keyinput27), .A(n13677), .ZN(n13681) );
  AOI22_X1 U15870 ( .A1(n13679), .A2(keyinput63), .B1(P2_U3088), .B2(keyinput4), .ZN(n13678) );
  OAI221_X1 U15871 ( .B1(n13679), .B2(keyinput63), .C1(P2_U3088), .C2(
        keyinput4), .A(n13678), .ZN(n13680) );
  OR3_X1 U15872 ( .A1(n13682), .A2(n13681), .A3(n13680), .ZN(n13691) );
  INV_X1 U15873 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U15874 ( .A1(n13685), .A2(keyinput44), .B1(keyinput16), .B2(n13684), 
        .ZN(n13683) );
  OAI221_X1 U15875 ( .B1(n13685), .B2(keyinput44), .C1(n13684), .C2(keyinput16), .A(n13683), .ZN(n13690) );
  INV_X1 U15876 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n13688) );
  INV_X1 U15877 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13687) );
  AOI22_X1 U15878 ( .A1(n13688), .A2(keyinput58), .B1(keyinput9), .B2(n13687), 
        .ZN(n13686) );
  OAI221_X1 U15879 ( .B1(n13688), .B2(keyinput58), .C1(n13687), .C2(keyinput9), 
        .A(n13686), .ZN(n13689) );
  NOR4_X1 U15880 ( .A1(n13692), .A2(n13691), .A3(n13690), .A4(n13689), .ZN(
        n13723) );
  NAND3_X1 U15881 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_WR_REG_SCAN_IN), .A3(
        n13693), .ZN(n13700) );
  NAND4_X1 U15882 ( .A1(n13695), .A2(n13694), .A3(P1_REG3_REG_12__SCAN_IN), 
        .A4(P2_REG2_REG_26__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U15883 ( .A1(n13609), .A2(P3_REG0_REG_1__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .A4(P2_REG3_REG_10__SCAN_IN), .ZN(n13698) );
  NAND4_X1 U15884 ( .A1(n13696), .A2(P1_REG3_REG_23__SCAN_IN), .A3(
        P1_REG2_REG_8__SCAN_IN), .A4(P1_REG1_REG_19__SCAN_IN), .ZN(n13697) );
  NOR4_X1 U15885 ( .A1(n13700), .A2(n13699), .A3(n13698), .A4(n13697), .ZN(
        n13714) );
  NOR4_X1 U15886 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P1_DATAO_REG_27__SCAN_IN), 
        .A3(P1_REG0_REG_14__SCAN_IN), .A4(n15738), .ZN(n13713) );
  NAND4_X1 U15887 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .A3(P3_ADDR_REG_12__SCAN_IN), .A4(n15313), .ZN(n13708) );
  NAND4_X1 U15888 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(P1_REG0_REG_28__SCAN_IN), .A4(n14122), .ZN(n13704) );
  NAND4_X1 U15889 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(P3_REG0_REG_20__SCAN_IN), 
        .A3(P1_REG1_REG_18__SCAN_IN), .A4(n11060), .ZN(n13703) );
  OR4_X1 U15890 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P3_REG3_REG_28__SCAN_IN), .A4(n13701), .ZN(n13702) );
  NOR4_X1 U15891 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n13704), .A3(n13703), 
        .A4(n13702), .ZN(n13705) );
  NAND4_X1 U15892 ( .A1(n13705), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P3_DATAO_REG_4__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n13707) );
  NAND4_X1 U15893 ( .A1(SI_7_), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_REG0_REG_22__SCAN_IN), .ZN(n13706) );
  NOR3_X1 U15894 ( .A1(n13708), .A2(n13707), .A3(n13706), .ZN(n13712) );
  NOR3_X1 U15895 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_REG0_REG_21__SCAN_IN), 
        .A3(P3_REG0_REG_17__SCAN_IN), .ZN(n13710) );
  NOR4_X1 U15896 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(P2_DATAO_REG_5__SCAN_IN), 
        .A3(P2_REG0_REG_13__SCAN_IN), .A4(P3_REG1_REG_10__SCAN_IN), .ZN(n13709) );
  AND3_X1 U15897 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n13710), .A3(n13709), .ZN(
        n13711) );
  AND4_X1 U15898 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        n13719) );
  NAND4_X1 U15899 ( .A1(P2_STATE_REG_SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(n13857), .A4(n15335), .ZN(n13717) );
  NAND4_X1 U15900 ( .A1(P3_REG0_REG_10__SCAN_IN), .A2(P3_REG2_REG_31__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .A4(P2_WR_REG_SCAN_IN), .ZN(n13716) );
  NAND3_X1 U15901 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(P3_REG0_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .ZN(n13715) );
  NOR4_X1 U15902 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(n13717), .A3(n13716), .A4(
        n13715), .ZN(n13718) );
  AOI21_X1 U15903 ( .B1(n13719), .B2(n13718), .A(keyinput57), .ZN(n13721) );
  MUX2_X1 U15904 ( .A(keyinput57), .B(n13721), .S(n13720), .Z(n13722) );
  NAND4_X1 U15905 ( .A1(n13725), .A2(n13724), .A3(n13723), .A4(n13722), .ZN(
        n13726) );
  XNOR2_X1 U15906 ( .A(n13727), .B(n13726), .ZN(P3_U3477) );
  AOI21_X1 U15907 ( .B1(n13729), .B2(n15851), .A(n13728), .ZN(n13796) );
  MUX2_X1 U15908 ( .A(n13730), .B(n13796), .S(n15873), .Z(n13731) );
  OAI21_X1 U15909 ( .B1(n13799), .B2(n13750), .A(n13731), .ZN(P3_U3476) );
  AOI21_X1 U15910 ( .B1(n13733), .B2(n15851), .A(n13732), .ZN(n13800) );
  MUX2_X1 U15911 ( .A(n13734), .B(n13800), .S(n15873), .Z(n13735) );
  OAI21_X1 U15912 ( .B1(n13803), .B2(n13750), .A(n13735), .ZN(P3_U3475) );
  AOI21_X1 U15913 ( .B1(n13737), .B2(n15851), .A(n13736), .ZN(n13804) );
  MUX2_X1 U15914 ( .A(n13738), .B(n13804), .S(n15873), .Z(n13739) );
  OAI21_X1 U15915 ( .B1(n7713), .B2(n13750), .A(n13739), .ZN(P3_U3474) );
  AOI21_X1 U15916 ( .B1(n13741), .B2(n15851), .A(n13740), .ZN(n13808) );
  MUX2_X1 U15917 ( .A(n13808), .B(n13742), .S(n10255), .Z(n13743) );
  OAI21_X1 U15918 ( .B1(n13810), .B2(n13750), .A(n13743), .ZN(P3_U3473) );
  OAI21_X1 U15919 ( .B1(n13746), .B2(n13745), .A(n13744), .ZN(n13747) );
  INV_X1 U15920 ( .A(n13747), .ZN(n13811) );
  MUX2_X1 U15921 ( .A(n13748), .B(n13811), .S(n15873), .Z(n13749) );
  OAI21_X1 U15922 ( .B1(n13750), .B2(n13814), .A(n13749), .ZN(P3_U3472) );
  MUX2_X1 U15923 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n13751), .S(n15873), .Z(
        n13752) );
  AOI21_X1 U15924 ( .B1(n13754), .B2(n13753), .A(n13752), .ZN(n13755) );
  INV_X1 U15925 ( .A(n13755), .ZN(P3_U3470) );
  NOR2_X1 U15926 ( .A1(n15858), .A2(n13756), .ZN(n13761) );
  AOI21_X1 U15927 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15858), .A(n13761), 
        .ZN(n13757) );
  OAI21_X1 U15928 ( .B1(n13758), .B2(n13815), .A(n13757), .ZN(P3_U3458) );
  INV_X1 U15929 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U15930 ( .A1(n13760), .A2(n13759), .ZN(n13763) );
  INV_X1 U15931 ( .A(n13761), .ZN(n13762) );
  OAI211_X1 U15932 ( .C1(n15860), .C2(n13764), .A(n13763), .B(n13762), .ZN(
        P3_U3457) );
  INV_X1 U15933 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13765) );
  MUX2_X1 U15934 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13768), .S(n15860), .Z(
        P3_U3454) );
  MUX2_X1 U15935 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13769), .S(n15860), .Z(
        P3_U3453) );
  MUX2_X1 U15936 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13770), .S(n15860), .Z(
        P3_U3452) );
  INV_X1 U15937 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13772) );
  MUX2_X1 U15938 ( .A(n13772), .B(n13771), .S(n15860), .Z(n13773) );
  OAI21_X1 U15939 ( .B1(n13774), .B2(n13815), .A(n13773), .ZN(P3_U3451) );
  INV_X1 U15940 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13776) );
  MUX2_X1 U15941 ( .A(n13776), .B(n13775), .S(n15860), .Z(n13777) );
  OAI21_X1 U15942 ( .B1(n13778), .B2(n13815), .A(n13777), .ZN(P3_U3450) );
  INV_X1 U15943 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13780) );
  MUX2_X1 U15944 ( .A(n13780), .B(n13779), .S(n15860), .Z(n13781) );
  OAI21_X1 U15945 ( .B1(n13782), .B2(n13815), .A(n13781), .ZN(P3_U3449) );
  MUX2_X1 U15946 ( .A(n13784), .B(n13783), .S(n15860), .Z(n13785) );
  OAI21_X1 U15947 ( .B1(n13786), .B2(n13815), .A(n13785), .ZN(P3_U3448) );
  MUX2_X1 U15948 ( .A(n13788), .B(n13787), .S(n15860), .Z(n13789) );
  OAI21_X1 U15949 ( .B1(n13790), .B2(n13815), .A(n13789), .ZN(P3_U3447) );
  INV_X1 U15950 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13792) );
  MUX2_X1 U15951 ( .A(n13792), .B(n13791), .S(n15860), .Z(n13793) );
  OAI21_X1 U15952 ( .B1(n13815), .B2(n13794), .A(n13793), .ZN(P3_U3446) );
  MUX2_X1 U15953 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13795), .S(n15860), .Z(
        P3_U3444) );
  MUX2_X1 U15954 ( .A(n13797), .B(n13796), .S(n15860), .Z(n13798) );
  OAI21_X1 U15955 ( .B1(n13799), .B2(n13815), .A(n13798), .ZN(P3_U3441) );
  MUX2_X1 U15956 ( .A(n13801), .B(n13800), .S(n15860), .Z(n13802) );
  OAI21_X1 U15957 ( .B1(n13803), .B2(n13815), .A(n13802), .ZN(P3_U3438) );
  MUX2_X1 U15958 ( .A(n13805), .B(n13804), .S(n15860), .Z(n13806) );
  OAI21_X1 U15959 ( .B1(n7713), .B2(n13815), .A(n13806), .ZN(P3_U3435) );
  INV_X1 U15960 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13807) );
  MUX2_X1 U15961 ( .A(n13808), .B(n13807), .S(n15858), .Z(n13809) );
  OAI21_X1 U15962 ( .B1(n13810), .B2(n13815), .A(n13809), .ZN(P3_U3432) );
  INV_X1 U15963 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13812) );
  MUX2_X1 U15964 ( .A(n13812), .B(n13811), .S(n15860), .Z(n13813) );
  OAI21_X1 U15965 ( .B1(n13815), .B2(n13814), .A(n13813), .ZN(P3_U3429) );
  MUX2_X1 U15966 ( .A(P3_D_REG_0__SCAN_IN), .B(n13817), .S(n13816), .Z(
        P3_U3376) );
  INV_X1 U15967 ( .A(n13818), .ZN(n13824) );
  INV_X1 U15968 ( .A(n13819), .ZN(n13820) );
  NOR4_X1 U15969 ( .A1(n13820), .A2(P3_IR_REG_30__SCAN_IN), .A3(n9411), .A4(
        P3_U3151), .ZN(n13821) );
  AOI21_X1 U15970 ( .B1(n13822), .B2(SI_31_), .A(n13821), .ZN(n13823) );
  OAI21_X1 U15971 ( .B1(n13824), .B2(n13836), .A(n13823), .ZN(P3_U3264) );
  INV_X1 U15972 ( .A(n13825), .ZN(n13826) );
  OAI222_X1 U15973 ( .A1(n13838), .A2(n13828), .B1(P3_U3151), .B2(n13827), 
        .C1(n13836), .C2(n13826), .ZN(P3_U3266) );
  INV_X1 U15974 ( .A(SI_27_), .ZN(n13832) );
  INV_X1 U15975 ( .A(n13829), .ZN(n13830) );
  OAI222_X1 U15976 ( .A1(n13838), .A2(n13832), .B1(P3_U3151), .B2(n13831), 
        .C1(n13836), .C2(n13830), .ZN(P3_U3268) );
  INV_X1 U15977 ( .A(n13833), .ZN(n13835) );
  OAI222_X1 U15978 ( .A1(n13838), .A2(n13837), .B1(n13836), .B2(n13835), .C1(
        P3_U3151), .C2(n13834), .ZN(P3_U3269) );
  MUX2_X1 U15979 ( .A(n13839), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15980 ( .A(n13840), .ZN(n13841) );
  AOI21_X1 U15981 ( .B1(n13843), .B2(n13842), .A(n13841), .ZN(n13849) );
  NAND2_X1 U15982 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n14110)
         );
  OAI21_X1 U15983 ( .B1(n13991), .B2(n13902), .A(n14110), .ZN(n13847) );
  OAI22_X1 U15984 ( .A1(n13995), .A2(n13845), .B1(n13993), .B2(n13844), .ZN(
        n13846) );
  AOI211_X1 U15985 ( .C1(n14490), .C2(n13998), .A(n13847), .B(n13846), .ZN(
        n13848) );
  OAI21_X1 U15986 ( .B1(n13849), .B2(n13984), .A(n13848), .ZN(P2_U3187) );
  INV_X1 U15987 ( .A(n13856), .ZN(n13853) );
  OAI21_X1 U15988 ( .B1(n13853), .B2(n13854), .A(n13986), .ZN(n13861) );
  INV_X1 U15989 ( .A(n13854), .ZN(n13855) );
  NOR2_X1 U15990 ( .A1(n13856), .A2(n13855), .ZN(n13922) );
  OAI22_X1 U15991 ( .A1(n14256), .A2(n13991), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13857), .ZN(n13859) );
  OAI22_X1 U15992 ( .A1(n13995), .A2(n14255), .B1(n13993), .B2(n14257), .ZN(
        n13858) );
  AOI211_X1 U15993 ( .C1(n14440), .C2(n13998), .A(n13859), .B(n13858), .ZN(
        n13860) );
  OAI21_X1 U15994 ( .B1(n13861), .B2(n13922), .A(n13860), .ZN(P2_U3188) );
  INV_X1 U15995 ( .A(n13991), .ZN(n13970) );
  AOI22_X1 U15996 ( .A1(n13958), .A2(n14023), .B1(n13970), .B2(n14021), .ZN(
        n13868) );
  AOI22_X1 U15997 ( .A1(n13998), .A2(n15742), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13867) );
  XOR2_X1 U15998 ( .A(n13863), .B(n13862), .Z(n13864) );
  NAND2_X1 U15999 ( .A1(n13864), .A2(n13986), .ZN(n13866) );
  NAND2_X1 U16000 ( .A1(n13873), .A2(n11652), .ZN(n13865) );
  NAND4_X1 U16001 ( .A1(n13868), .A2(n13867), .A3(n13866), .A4(n13865), .ZN(
        P2_U3190) );
  NAND2_X1 U16002 ( .A1(n13870), .A2(n13869), .ZN(n13872) );
  XOR2_X1 U16003 ( .A(n13872), .B(n13871), .Z(n13877) );
  AOI22_X1 U16004 ( .A1(n13970), .A2(n14284), .B1(n13873), .B2(n14322), .ZN(
        n13874) );
  NAND2_X1 U16005 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14167)
         );
  OAI211_X1 U16006 ( .C1(n14314), .C2(n13995), .A(n13874), .B(n14167), .ZN(
        n13875) );
  AOI21_X1 U16007 ( .B1(n14321), .B2(n13998), .A(n13875), .ZN(n13876) );
  OAI21_X1 U16008 ( .B1(n13877), .B2(n13984), .A(n13876), .ZN(P2_U3191) );
  INV_X1 U16009 ( .A(n13878), .ZN(n13880) );
  OAI211_X1 U16010 ( .C1(n13880), .C2(n6782), .A(n13986), .B(n13944), .ZN(
        n13884) );
  NOR2_X1 U16011 ( .A1(n13991), .A2(n14255), .ZN(n13882) );
  OAI22_X1 U16012 ( .A1(n13995), .A2(n14315), .B1(n13993), .B2(n14291), .ZN(
        n13881) );
  AOI211_X1 U16013 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n13882), 
        .B(n13881), .ZN(n13883) );
  OAI211_X1 U16014 ( .C1(n14537), .C2(n13973), .A(n13884), .B(n13883), .ZN(
        P2_U3195) );
  OAI211_X1 U16015 ( .C1(n13887), .C2(n13886), .A(n13885), .B(n13986), .ZN(
        n13893) );
  AOI22_X1 U16016 ( .A1(n14006), .A2(n14374), .B1(n14007), .B2(n14376), .ZN(
        n14212) );
  INV_X1 U16017 ( .A(n14212), .ZN(n13891) );
  OAI22_X1 U16018 ( .A1(n13993), .A2(n14218), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13888), .ZN(n13889) );
  AOI21_X1 U16019 ( .B1(n13891), .B2(n13890), .A(n13889), .ZN(n13892) );
  OAI211_X1 U16020 ( .C1(n14527), .C2(n13973), .A(n13893), .B(n13892), .ZN(
        P2_U3197) );
  XNOR2_X1 U16021 ( .A(n13895), .B(n13894), .ZN(n13900) );
  INV_X1 U16022 ( .A(n13896), .ZN(n13898) );
  XNOR2_X1 U16023 ( .A(n13897), .B(n13896), .ZN(n13989) );
  NAND2_X1 U16024 ( .A1(n13989), .A2(n13988), .ZN(n13987) );
  OAI21_X1 U16025 ( .B1(n13898), .B2(n13897), .A(n13987), .ZN(n13899) );
  NOR2_X1 U16026 ( .A1(n13899), .A2(n13900), .ZN(n13910) );
  AOI21_X1 U16027 ( .B1(n13900), .B2(n13899), .A(n13910), .ZN(n13906) );
  OAI21_X1 U16028 ( .B1(n13991), .B2(n14330), .A(n13901), .ZN(n13904) );
  OAI22_X1 U16029 ( .A1(n13995), .A2(n13902), .B1(n13993), .B2(n14384), .ZN(
        n13903) );
  AOI211_X1 U16030 ( .C1(n14477), .C2(n13998), .A(n13904), .B(n13903), .ZN(
        n13905) );
  OAI21_X1 U16031 ( .B1(n13906), .B2(n13984), .A(n13905), .ZN(P2_U3198) );
  INV_X1 U16032 ( .A(n13907), .ZN(n13909) );
  NOR3_X1 U16033 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(n13913) );
  INV_X1 U16034 ( .A(n13911), .ZN(n13912) );
  OAI21_X1 U16035 ( .B1(n13913), .B2(n13912), .A(n13986), .ZN(n13918) );
  NOR2_X1 U16036 ( .A1(n13914), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15705) );
  INV_X1 U16037 ( .A(n14365), .ZN(n13915) );
  OAI22_X1 U16038 ( .A1(n13995), .A2(n13990), .B1(n13993), .B2(n13915), .ZN(
        n13916) );
  AOI211_X1 U16039 ( .C1(n13970), .C2(n14360), .A(n15705), .B(n13916), .ZN(
        n13917) );
  OAI211_X1 U16040 ( .C1(n14546), .C2(n13973), .A(n13918), .B(n13917), .ZN(
        P2_U3200) );
  AND2_X1 U16041 ( .A1(n13920), .A2(n13919), .ZN(n13921) );
  NAND2_X1 U16042 ( .A1(n13924), .A2(n13923), .ZN(n13925) );
  XNOR2_X1 U16043 ( .A(n13926), .B(n13925), .ZN(n13933) );
  OAI22_X1 U16044 ( .A1(n13980), .A2(n13991), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13927), .ZN(n13931) );
  INV_X1 U16045 ( .A(n14231), .ZN(n13928) );
  OAI22_X1 U16046 ( .A1(n13995), .A2(n13929), .B1(n13993), .B2(n13928), .ZN(
        n13930) );
  AOI211_X1 U16047 ( .C1(n14434), .C2(n13998), .A(n13931), .B(n13930), .ZN(
        n13932) );
  OAI21_X1 U16048 ( .B1(n13933), .B2(n13984), .A(n13932), .ZN(P2_U3201) );
  XNOR2_X1 U16049 ( .A(n13935), .B(n13934), .ZN(n13936) );
  XNOR2_X1 U16050 ( .A(n13937), .B(n13936), .ZN(n13943) );
  OAI22_X1 U16051 ( .A1(n13995), .A2(n14332), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13938), .ZN(n13941) );
  INV_X1 U16052 ( .A(n14305), .ZN(n13939) );
  OAI22_X1 U16053 ( .A1(n13993), .A2(n13939), .B1(n13991), .B2(n14303), .ZN(
        n13940) );
  AOI211_X1 U16054 ( .C1(n14456), .C2(n13998), .A(n13941), .B(n13940), .ZN(
        n13942) );
  OAI21_X1 U16055 ( .B1(n13943), .B2(n13984), .A(n13942), .ZN(P2_U3205) );
  NOR2_X1 U16056 ( .A1(n13850), .A2(n13945), .ZN(n13949) );
  XNOR2_X1 U16057 ( .A(n13947), .B(n13946), .ZN(n13948) );
  XNOR2_X1 U16058 ( .A(n13949), .B(n13948), .ZN(n13956) );
  NOR2_X1 U16059 ( .A1(n13993), .A2(n14270), .ZN(n13954) );
  NOR2_X1 U16060 ( .A1(n14303), .A2(n14329), .ZN(n13950) );
  AOI21_X1 U16061 ( .B1(n14227), .B2(n14374), .A(n13950), .ZN(n14264) );
  OAI22_X1 U16062 ( .A1(n14264), .A2(n13952), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13951), .ZN(n13953) );
  AOI211_X1 U16063 ( .C1(n14277), .C2(n13998), .A(n13954), .B(n13953), .ZN(
        n13955) );
  OAI21_X1 U16064 ( .B1(n13956), .B2(n13984), .A(n13955), .ZN(P2_U3207) );
  AOI22_X1 U16065 ( .A1(n13958), .A2(n14024), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13957), .ZN(n13965) );
  AOI22_X1 U16066 ( .A1(n13970), .A2(n14022), .B1(n6421), .B2(n13998), .ZN(
        n13964) );
  OAI21_X1 U16067 ( .B1(n13961), .B2(n13959), .A(n13960), .ZN(n13962) );
  NAND2_X1 U16068 ( .A1(n13986), .A2(n13962), .ZN(n13963) );
  NAND3_X1 U16069 ( .A1(n13965), .A2(n13964), .A3(n13963), .ZN(P2_U3209) );
  OAI211_X1 U16070 ( .C1(n13968), .C2(n13967), .A(n13966), .B(n13986), .ZN(
        n13972) );
  AND2_X1 U16071 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14140) );
  OAI22_X1 U16072 ( .A1(n13995), .A2(n14330), .B1(n13993), .B2(n14344), .ZN(
        n13969) );
  AOI211_X1 U16073 ( .C1(n13970), .C2(n14009), .A(n14140), .B(n13969), .ZN(
        n13971) );
  OAI211_X1 U16074 ( .C1(n14347), .C2(n13973), .A(n13972), .B(n13971), .ZN(
        P2_U3210) );
  INV_X1 U16075 ( .A(n13974), .ZN(n13975) );
  AOI21_X1 U16076 ( .B1(n13977), .B2(n13976), .A(n13975), .ZN(n13985) );
  OAI22_X1 U16077 ( .A1(n13979), .A2(n13991), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13978), .ZN(n13982) );
  OAI22_X1 U16078 ( .A1(n13980), .A2(n13995), .B1(n14201), .B2(n13993), .ZN(
        n13981) );
  AOI211_X1 U16079 ( .C1(n14425), .C2(n13998), .A(n13982), .B(n13981), .ZN(
        n13983) );
  OAI21_X1 U16080 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(P2_U3212) );
  OAI211_X1 U16081 ( .C1(n13989), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n14001) );
  OAI22_X1 U16082 ( .A1(n13991), .A2(n13990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14122), .ZN(n13997) );
  OAI22_X1 U16083 ( .A1(n13995), .A2(n13994), .B1(n13993), .B2(n13992), .ZN(
        n13996) );
  AOI211_X1 U16084 ( .C1(n13999), .C2(n13998), .A(n13997), .B(n13996), .ZN(
        n14000) );
  NAND2_X1 U16085 ( .A1(n14001), .A2(n14000), .ZN(P2_U3213) );
  INV_X2 U16086 ( .A(P2_U3947), .ZN(n14016) );
  MUX2_X1 U16087 ( .A(n14002), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14016), .Z(
        P2_U3562) );
  MUX2_X1 U16088 ( .A(n14003), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14016), .Z(
        P2_U3561) );
  MUX2_X1 U16089 ( .A(n14004), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14016), .Z(
        P2_U3560) );
  MUX2_X1 U16090 ( .A(n14005), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14016), .Z(
        P2_U3559) );
  MUX2_X1 U16091 ( .A(n14196), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14016), .Z(
        P2_U3558) );
  MUX2_X1 U16092 ( .A(n14006), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14016), .Z(
        P2_U3557) );
  MUX2_X1 U16093 ( .A(n14226), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14016), .Z(
        P2_U3556) );
  MUX2_X1 U16094 ( .A(n14007), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14016), .Z(
        P2_U3555) );
  MUX2_X1 U16095 ( .A(n14227), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14016), .Z(
        P2_U3554) );
  MUX2_X1 U16096 ( .A(n14285), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14016), .Z(
        P2_U3553) );
  MUX2_X1 U16097 ( .A(n14008), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14016), .Z(
        P2_U3552) );
  MUX2_X1 U16098 ( .A(n14284), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14016), .Z(
        P2_U3551) );
  MUX2_X1 U16099 ( .A(n14009), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14016), .Z(
        P2_U3550) );
  MUX2_X1 U16100 ( .A(n14360), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14016), .Z(
        P2_U3549) );
  INV_X1 U16101 ( .A(n14330), .ZN(n14375) );
  MUX2_X1 U16102 ( .A(n14375), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14016), .Z(
        P2_U3548) );
  MUX2_X1 U16103 ( .A(n14359), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14016), .Z(
        P2_U3547) );
  MUX2_X1 U16104 ( .A(n14377), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14016), .Z(
        P2_U3546) );
  MUX2_X1 U16105 ( .A(n14010), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14016), .Z(
        P2_U3545) );
  MUX2_X1 U16106 ( .A(n14011), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14016), .Z(
        P2_U3544) );
  MUX2_X1 U16107 ( .A(n14012), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14016), .Z(
        P2_U3543) );
  MUX2_X1 U16108 ( .A(n14013), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14016), .Z(
        P2_U3542) );
  MUX2_X1 U16109 ( .A(n14014), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14016), .Z(
        P2_U3541) );
  MUX2_X1 U16110 ( .A(n14015), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14016), .Z(
        P2_U3540) );
  MUX2_X1 U16111 ( .A(n14017), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14016), .Z(
        P2_U3539) );
  MUX2_X1 U16112 ( .A(n14018), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14016), .Z(
        P2_U3538) );
  MUX2_X1 U16113 ( .A(n14019), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14016), .Z(
        P2_U3537) );
  MUX2_X1 U16114 ( .A(n14020), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14016), .Z(
        P2_U3536) );
  MUX2_X1 U16115 ( .A(n14021), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14016), .Z(
        P2_U3535) );
  MUX2_X1 U16116 ( .A(n14022), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14016), .Z(
        P2_U3534) );
  MUX2_X1 U16117 ( .A(n14023), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14016), .Z(
        P2_U3533) );
  MUX2_X1 U16118 ( .A(n14024), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14016), .Z(
        P2_U3532) );
  MUX2_X1 U16119 ( .A(n14025), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14016), .Z(
        P2_U3531) );
  NOR2_X1 U16120 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11652), .ZN(n14027) );
  NOR2_X1 U16121 ( .A1(n15696), .A2(n14031), .ZN(n14026) );
  AOI211_X1 U16122 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n15634), .A(n14027), .B(
        n14026), .ZN(n14038) );
  OAI211_X1 U16123 ( .C1(n14030), .C2(n14029), .A(n15690), .B(n14028), .ZN(
        n14037) );
  MUX2_X1 U16124 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11654), .S(n14031), .Z(
        n14032) );
  NAND3_X1 U16125 ( .A1(n15641), .A2(n14033), .A3(n14032), .ZN(n14034) );
  NAND3_X1 U16126 ( .A1(n15708), .A2(n14035), .A3(n14034), .ZN(n14036) );
  NAND3_X1 U16127 ( .A1(n14038), .A2(n14037), .A3(n14036), .ZN(P2_U3217) );
  INV_X1 U16128 ( .A(n14039), .ZN(n14041) );
  NOR2_X1 U16129 ( .A1(n15696), .A2(n14045), .ZN(n14040) );
  AOI211_X1 U16130 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n15634), .A(n14041), .B(
        n14040), .ZN(n14051) );
  OAI211_X1 U16131 ( .C1(n14044), .C2(n14043), .A(n15690), .B(n14042), .ZN(
        n14050) );
  MUX2_X1 U16132 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11635), .S(n14045), .Z(
        n14046) );
  NAND3_X1 U16133 ( .A1(n15655), .A2(n14047), .A3(n14046), .ZN(n14048) );
  NAND3_X1 U16134 ( .A1(n15708), .A2(n14061), .A3(n14048), .ZN(n14049) );
  NAND3_X1 U16135 ( .A1(n14051), .A2(n14050), .A3(n14049), .ZN(P2_U3219) );
  INV_X1 U16136 ( .A(n14052), .ZN(n14054) );
  NOR2_X1 U16137 ( .A1(n15696), .A2(n14058), .ZN(n14053) );
  AOI211_X1 U16138 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n15634), .A(n14054), .B(
        n14053), .ZN(n14065) );
  OAI211_X1 U16139 ( .C1(n14057), .C2(n14056), .A(n15690), .B(n14055), .ZN(
        n14064) );
  MUX2_X1 U16140 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11549), .S(n14058), .Z(
        n14059) );
  NAND3_X1 U16141 ( .A1(n14061), .A2(n14060), .A3(n14059), .ZN(n14062) );
  NAND3_X1 U16142 ( .A1(n15708), .A2(n14068), .A3(n14062), .ZN(n14063) );
  NAND3_X1 U16143 ( .A1(n14065), .A2(n14064), .A3(n14063), .ZN(P2_U3220) );
  MUX2_X1 U16144 ( .A(n11561), .B(P2_REG2_REG_7__SCAN_IN), .S(n14074), .Z(
        n14066) );
  NAND3_X1 U16145 ( .A1(n14068), .A2(n14067), .A3(n14066), .ZN(n14069) );
  NAND3_X1 U16146 ( .A1(n15708), .A2(n14087), .A3(n14069), .ZN(n14078) );
  OAI211_X1 U16147 ( .C1(n14072), .C2(n14071), .A(n15690), .B(n14070), .ZN(
        n14077) );
  NOR2_X1 U16148 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8997), .ZN(n14073) );
  AOI21_X1 U16149 ( .B1(n15707), .B2(n14074), .A(n14073), .ZN(n14076) );
  NAND2_X1 U16150 ( .A1(n15634), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n14075) );
  NAND4_X1 U16151 ( .A1(n14078), .A2(n14077), .A3(n14076), .A4(n14075), .ZN(
        P2_U3221) );
  OAI21_X1 U16152 ( .B1(n15696), .B2(n14080), .A(n14079), .ZN(n14081) );
  AOI21_X1 U16153 ( .B1(n15634), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n14081), .ZN(
        n14092) );
  OAI211_X1 U16154 ( .C1(n14083), .C2(n14082), .A(n15690), .B(n15670), .ZN(
        n14091) );
  MUX2_X1 U16155 ( .A(n11737), .B(P2_REG2_REG_8__SCAN_IN), .S(n14084), .Z(
        n14085) );
  NAND3_X1 U16156 ( .A1(n14087), .A2(n14086), .A3(n14085), .ZN(n14088) );
  NAND3_X1 U16157 ( .A1(n15708), .A2(n14089), .A3(n14088), .ZN(n14090) );
  NAND3_X1 U16158 ( .A1(n14092), .A2(n14091), .A3(n14090), .ZN(P2_U3222) );
  AOI21_X1 U16159 ( .B1(n14094), .B2(n14093), .A(n14161), .ZN(n14096) );
  NAND2_X1 U16160 ( .A1(n14096), .A2(n14095), .ZN(n14107) );
  NOR2_X1 U16161 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14097), .ZN(n14098) );
  AOI21_X1 U16162 ( .B1(n15707), .B2(n14099), .A(n14098), .ZN(n14106) );
  NAND2_X1 U16163 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  NAND3_X1 U16164 ( .A1(n14103), .A2(n15690), .A3(n14102), .ZN(n14105) );
  NAND2_X1 U16165 ( .A1(n15634), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n14104) );
  NAND4_X1 U16166 ( .A1(n14107), .A2(n14106), .A3(n14105), .A4(n14104), .ZN(
        P2_U3227) );
  XOR2_X1 U16167 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n14108), .Z(n14109) );
  NAND2_X1 U16168 ( .A1(n14109), .A2(n15708), .ZN(n14119) );
  INV_X1 U16169 ( .A(n14110), .ZN(n14111) );
  AOI21_X1 U16170 ( .B1(n15707), .B2(n14112), .A(n14111), .ZN(n14118) );
  OAI211_X1 U16171 ( .C1(n14115), .C2(n14114), .A(n14113), .B(n15690), .ZN(
        n14117) );
  NAND2_X1 U16172 ( .A1(n15634), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n14116) );
  NAND4_X1 U16173 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        P2_U3228) );
  XOR2_X1 U16174 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n14120), .Z(n14121) );
  NAND2_X1 U16175 ( .A1(n14121), .A2(n15708), .ZN(n14130) );
  NOR2_X1 U16176 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14122), .ZN(n14123) );
  AOI21_X1 U16177 ( .B1(n15707), .B2(n14124), .A(n14123), .ZN(n14129) );
  OAI211_X1 U16178 ( .C1(n14126), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14125), 
        .B(n15690), .ZN(n14128) );
  NAND2_X1 U16179 ( .A1(n15634), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n14127) );
  NAND4_X1 U16180 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14127), .ZN(
        P2_U3229) );
  NAND2_X1 U16181 ( .A1(n14143), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14133) );
  MUX2_X1 U16182 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14134), .S(n15706), .Z(
        n15710) );
  NAND2_X1 U16183 ( .A1(n15706), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14135) );
  NAND2_X1 U16184 ( .A1(n15709), .A2(n14135), .ZN(n14136) );
  OR2_X1 U16185 ( .A1(n14136), .A2(n14147), .ZN(n14158) );
  NAND2_X1 U16186 ( .A1(n14136), .A2(n14147), .ZN(n14137) );
  INV_X1 U16187 ( .A(n14159), .ZN(n14138) );
  AOI21_X1 U16188 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14139), .A(n14138), 
        .ZN(n14154) );
  INV_X1 U16189 ( .A(n14140), .ZN(n14141) );
  OAI21_X1 U16190 ( .B1(n15696), .B2(n14144), .A(n14141), .ZN(n14152) );
  AOI21_X1 U16191 ( .B1(n14143), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14142), 
        .ZN(n15703) );
  XNOR2_X1 U16192 ( .A(n15706), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15702) );
  NOR2_X1 U16193 ( .A1(n15703), .A2(n15702), .ZN(n15700) );
  AOI21_X1 U16194 ( .B1(n15706), .B2(P2_REG1_REG_17__SCAN_IN), .A(n15700), 
        .ZN(n14145) );
  INV_X1 U16195 ( .A(n14145), .ZN(n14148) );
  NOR2_X1 U16196 ( .A1(n14145), .A2(n14144), .ZN(n14156) );
  INV_X1 U16197 ( .A(n14156), .ZN(n14146) );
  OAI21_X1 U16198 ( .B1(n14148), .B2(n14147), .A(n14146), .ZN(n14149) );
  NOR2_X1 U16199 ( .A1(n14149), .A2(n14150), .ZN(n14155) );
  AOI211_X1 U16200 ( .C1(n14150), .C2(n14149), .A(n15701), .B(n14155), .ZN(
        n14151) );
  AOI211_X1 U16201 ( .C1(n15634), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14152), 
        .B(n14151), .ZN(n14153) );
  OAI21_X1 U16202 ( .B1(n14154), .B2(n14161), .A(n14153), .ZN(P2_U3232) );
  NOR2_X1 U16203 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  XNOR2_X1 U16204 ( .A(n14157), .B(n14463), .ZN(n14164) );
  INV_X1 U16205 ( .A(n14164), .ZN(n14160) );
  AOI22_X1 U16206 ( .A1(n14160), .A2(n15690), .B1(n14162), .B2(n15708), .ZN(
        n14166) );
  AOI211_X1 U16207 ( .C1(n15690), .C2(n14164), .A(n15707), .B(n14163), .ZN(
        n14165) );
  MUX2_X1 U16208 ( .A(n14166), .B(n14165), .S(n14386), .Z(n14168) );
  OAI211_X1 U16209 ( .C1(n8064), .C2(n15715), .A(n14168), .B(n14167), .ZN(
        P2_U3233) );
  XNOR2_X1 U16210 ( .A(n14175), .B(n14516), .ZN(n14170) );
  NAND2_X1 U16211 ( .A1(n14170), .A2(n14273), .ZN(n14407) );
  OR2_X1 U16212 ( .A1(n14172), .A2(n14171), .ZN(n14410) );
  NOR2_X1 U16213 ( .A1(n14352), .A2(n14410), .ZN(n14178) );
  NOR2_X1 U16214 ( .A1(n14516), .A2(n14368), .ZN(n14173) );
  AOI211_X1 U16215 ( .C1(n14352), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14178), 
        .B(n14173), .ZN(n14174) );
  OAI21_X1 U16216 ( .B1(n14407), .B2(n14274), .A(n14174), .ZN(P2_U3234) );
  OAI211_X1 U16217 ( .C1(n14520), .C2(n14176), .A(n14273), .B(n14175), .ZN(
        n14411) );
  NOR2_X1 U16218 ( .A1(n14520), .A2(n14368), .ZN(n14177) );
  AOI211_X1 U16219 ( .C1(n14352), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14178), 
        .B(n14177), .ZN(n14179) );
  OAI21_X1 U16220 ( .B1(n14274), .B2(n14411), .A(n14179), .ZN(P2_U3235) );
  XNOR2_X1 U16221 ( .A(n14181), .B(n14180), .ZN(n14184) );
  INV_X1 U16222 ( .A(n14182), .ZN(n14183) );
  AOI21_X1 U16223 ( .B1(n14184), .B2(n14379), .A(n14183), .ZN(n14423) );
  INV_X1 U16224 ( .A(n14371), .ZN(n14403) );
  NAND3_X1 U16225 ( .A1(n6498), .A2(n14403), .A3(n14419), .ZN(n14194) );
  OAI211_X1 U16226 ( .C1(n14190), .C2(n14197), .A(n14273), .B(n14187), .ZN(
        n14422) );
  INV_X1 U16227 ( .A(n14422), .ZN(n14192) );
  AOI22_X1 U16228 ( .A1(n14188), .A2(n14397), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14352), .ZN(n14189) );
  OAI21_X1 U16229 ( .B1(n14190), .B2(n14368), .A(n14189), .ZN(n14191) );
  AOI21_X1 U16230 ( .B1(n14192), .B2(n14399), .A(n14191), .ZN(n14193) );
  OAI211_X1 U16231 ( .C1(n14352), .C2(n14423), .A(n14194), .B(n14193), .ZN(
        P2_U3238) );
  AOI21_X1 U16232 ( .B1(n14425), .B2(n14214), .A(n14380), .ZN(n14198) );
  AND2_X1 U16233 ( .A1(n14198), .A2(n6861), .ZN(n14424) );
  NAND2_X1 U16234 ( .A1(n14425), .A2(n14401), .ZN(n14200) );
  NAND2_X1 U16235 ( .A1(n14352), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n14199) );
  OAI211_X1 U16236 ( .C1(n14385), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14205) );
  XNOR2_X1 U16237 ( .A(n14202), .B(n14203), .ZN(n14428) );
  NOR2_X1 U16238 ( .A1(n14428), .A2(n14371), .ZN(n14204) );
  AOI211_X1 U16239 ( .C1(n14424), .C2(n14399), .A(n14205), .B(n14204), .ZN(
        n14206) );
  OAI21_X1 U16240 ( .B1(n14352), .B2(n14427), .A(n14206), .ZN(P2_U3239) );
  XNOR2_X1 U16241 ( .A(n14207), .B(n14209), .ZN(n14431) );
  INV_X1 U16242 ( .A(n14431), .ZN(n14224) );
  OAI21_X1 U16243 ( .B1(n14210), .B2(n14209), .A(n14208), .ZN(n14211) );
  NAND2_X1 U16244 ( .A1(n14211), .A2(n14379), .ZN(n14213) );
  NAND2_X1 U16245 ( .A1(n14213), .A2(n14212), .ZN(n14429) );
  INV_X1 U16246 ( .A(n14229), .ZN(n14216) );
  INV_X1 U16247 ( .A(n14214), .ZN(n14215) );
  AOI211_X1 U16248 ( .C1(n14217), .C2(n14216), .A(n14380), .B(n14215), .ZN(
        n14430) );
  NAND2_X1 U16249 ( .A1(n14430), .A2(n14399), .ZN(n14221) );
  INV_X1 U16250 ( .A(n14218), .ZN(n14219) );
  AOI22_X1 U16251 ( .A1(n14219), .A2(n14397), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14352), .ZN(n14220) );
  OAI211_X1 U16252 ( .C1(n14527), .C2(n14368), .A(n14221), .B(n14220), .ZN(
        n14222) );
  AOI21_X1 U16253 ( .B1(n14429), .B2(n14396), .A(n14222), .ZN(n14223) );
  OAI21_X1 U16254 ( .B1(n14224), .B2(n14371), .A(n14223), .ZN(P2_U3240) );
  XNOR2_X1 U16255 ( .A(n14225), .B(n14236), .ZN(n14228) );
  AOI222_X1 U16256 ( .A1(n14379), .A2(n14228), .B1(n14227), .B2(n14376), .C1(
        n14226), .C2(n14374), .ZN(n14436) );
  NOR2_X1 U16257 ( .A1(n6475), .A2(n14233), .ZN(n14230) );
  AOI22_X1 U16258 ( .A1(n14231), .A2(n14397), .B1(n14352), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n14232) );
  OAI21_X1 U16259 ( .B1(n14233), .B2(n14368), .A(n14232), .ZN(n14238) );
  OAI21_X1 U16260 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14437) );
  NOR2_X1 U16261 ( .A1(n14437), .A2(n14371), .ZN(n14237) );
  AOI211_X1 U16262 ( .C1(n8061), .C2(n14399), .A(n14238), .B(n14237), .ZN(
        n14239) );
  OAI21_X1 U16263 ( .B1(n14352), .B2(n14436), .A(n14239), .ZN(P2_U3241) );
  INV_X1 U16264 ( .A(n14240), .ZN(n14241) );
  NAND2_X1 U16265 ( .A1(n14242), .A2(n14241), .ZN(n14280) );
  INV_X1 U16266 ( .A(n14243), .ZN(n14244) );
  OAI21_X1 U16267 ( .B1(n14280), .B2(n14281), .A(n14244), .ZN(n14267) );
  NAND2_X1 U16268 ( .A1(n14269), .A2(n14245), .ZN(n14246) );
  XOR2_X1 U16269 ( .A(n14253), .B(n14246), .Z(n14442) );
  NAND2_X1 U16270 ( .A1(n14272), .A2(n14440), .ZN(n14247) );
  NAND2_X1 U16271 ( .A1(n14247), .A2(n14273), .ZN(n14248) );
  NOR2_X1 U16272 ( .A1(n6475), .A2(n14248), .ZN(n14439) );
  INV_X1 U16273 ( .A(n14440), .ZN(n14250) );
  INV_X1 U16274 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14249) );
  OAI22_X1 U16275 ( .A1(n14250), .A2(n14368), .B1(n14249), .B2(n14396), .ZN(
        n14251) );
  AOI21_X1 U16276 ( .B1(n14439), .B2(n14399), .A(n14251), .ZN(n14260) );
  OAI222_X1 U16277 ( .A1(n14331), .A2(n14256), .B1(n14329), .B2(n14255), .C1(
        n14254), .C2(n14302), .ZN(n14438) );
  NOR2_X1 U16278 ( .A1(n14257), .A2(n14385), .ZN(n14258) );
  OAI21_X1 U16279 ( .B1(n14438), .B2(n14258), .A(n14396), .ZN(n14259) );
  OAI211_X1 U16280 ( .C1(n14442), .C2(n14371), .A(n14260), .B(n14259), .ZN(
        P2_U3242) );
  NAND2_X1 U16281 ( .A1(n14261), .A2(n7386), .ZN(n14262) );
  NAND3_X1 U16282 ( .A1(n14263), .A2(n14379), .A3(n14262), .ZN(n14265) );
  AND2_X1 U16283 ( .A1(n14265), .A2(n14264), .ZN(n14444) );
  NAND2_X1 U16284 ( .A1(n14267), .A2(n14266), .ZN(n14268) );
  AND2_X1 U16285 ( .A1(n14269), .A2(n14268), .ZN(n14446) );
  NAND2_X1 U16286 ( .A1(n14446), .A2(n14403), .ZN(n14279) );
  INV_X1 U16287 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14271) );
  OAI22_X1 U16288 ( .A1(n14396), .A2(n14271), .B1(n14270), .B2(n14385), .ZN(
        n14276) );
  OAI211_X1 U16289 ( .C1(n14288), .C2(n14533), .A(n14273), .B(n14272), .ZN(
        n14443) );
  NOR2_X1 U16290 ( .A1(n14443), .A2(n14274), .ZN(n14275) );
  AOI211_X1 U16291 ( .C1(n14401), .C2(n14277), .A(n14276), .B(n14275), .ZN(
        n14278) );
  OAI211_X1 U16292 ( .C1(n14352), .C2(n14444), .A(n14279), .B(n14278), .ZN(
        P2_U3243) );
  XNOR2_X1 U16293 ( .A(n14280), .B(n14281), .ZN(n14451) );
  INV_X1 U16294 ( .A(n14451), .ZN(n14297) );
  XNOR2_X1 U16295 ( .A(n14282), .B(n14281), .ZN(n14283) );
  NAND2_X1 U16296 ( .A1(n14283), .A2(n14379), .ZN(n14287) );
  AOI22_X1 U16297 ( .A1(n14285), .A2(n14374), .B1(n14284), .B2(n14376), .ZN(
        n14286) );
  NAND2_X1 U16298 ( .A1(n14287), .A2(n14286), .ZN(n14449) );
  INV_X1 U16299 ( .A(n14304), .ZN(n14289) );
  AOI211_X1 U16300 ( .C1(n14290), .C2(n14289), .A(n14380), .B(n14288), .ZN(
        n14450) );
  NAND2_X1 U16301 ( .A1(n14450), .A2(n14399), .ZN(n14294) );
  INV_X1 U16302 ( .A(n14291), .ZN(n14292) );
  AOI22_X1 U16303 ( .A1(n14352), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14292), 
        .B2(n14397), .ZN(n14293) );
  OAI211_X1 U16304 ( .C1(n14537), .C2(n14368), .A(n14294), .B(n14293), .ZN(
        n14295) );
  AOI21_X1 U16305 ( .B1(n14449), .B2(n14396), .A(n14295), .ZN(n14296) );
  OAI21_X1 U16306 ( .B1(n14297), .B2(n14371), .A(n14296), .ZN(P2_U3244) );
  XOR2_X1 U16307 ( .A(n14298), .B(n14300), .Z(n14458) );
  AOI21_X1 U16308 ( .B1(n14300), .B2(n14299), .A(n6529), .ZN(n14301) );
  OAI222_X1 U16309 ( .A1(n14329), .A2(n14332), .B1(n14331), .B2(n14303), .C1(
        n14302), .C2(n14301), .ZN(n14454) );
  AOI211_X1 U16310 ( .C1(n14456), .C2(n14319), .A(n14380), .B(n14304), .ZN(
        n14455) );
  NAND2_X1 U16311 ( .A1(n14455), .A2(n14399), .ZN(n14307) );
  AOI22_X1 U16312 ( .A1(n14352), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14305), 
        .B2(n14397), .ZN(n14306) );
  OAI211_X1 U16313 ( .C1(n14308), .C2(n14368), .A(n14307), .B(n14306), .ZN(
        n14309) );
  AOI21_X1 U16314 ( .B1(n14454), .B2(n14396), .A(n14309), .ZN(n14310) );
  OAI21_X1 U16315 ( .B1(n14458), .B2(n14371), .A(n14310), .ZN(P2_U3245) );
  XNOR2_X1 U16316 ( .A(n14311), .B(n14312), .ZN(n14459) );
  XNOR2_X1 U16317 ( .A(n14313), .B(n14312), .ZN(n14317) );
  OAI22_X1 U16318 ( .A1(n14315), .A2(n14331), .B1(n14314), .B2(n14329), .ZN(
        n14316) );
  AOI21_X1 U16319 ( .B1(n14317), .B2(n14379), .A(n14316), .ZN(n14318) );
  OAI21_X1 U16320 ( .B1(n14459), .B2(n14337), .A(n14318), .ZN(n14460) );
  NAND2_X1 U16321 ( .A1(n14460), .A2(n14396), .ZN(n14326) );
  INV_X1 U16322 ( .A(n14319), .ZN(n14320) );
  AOI211_X1 U16323 ( .C1(n14321), .C2(n14341), .A(n14380), .B(n14320), .ZN(
        n14461) );
  AOI22_X1 U16324 ( .A1(n14352), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14322), 
        .B2(n14397), .ZN(n14323) );
  OAI21_X1 U16325 ( .B1(n7890), .B2(n14368), .A(n14323), .ZN(n14324) );
  AOI21_X1 U16326 ( .B1(n14461), .B2(n14399), .A(n14324), .ZN(n14325) );
  OAI211_X1 U16327 ( .C1(n14459), .C2(n14348), .A(n14326), .B(n14325), .ZN(
        P2_U3246) );
  INV_X1 U16328 ( .A(n14353), .ZN(n14355) );
  NOR2_X1 U16329 ( .A1(n14356), .A2(n14355), .ZN(n14358) );
  NOR2_X1 U16330 ( .A1(n14358), .A2(n14327), .ZN(n14328) );
  XOR2_X1 U16331 ( .A(n14336), .B(n14328), .Z(n14340) );
  OAI22_X1 U16332 ( .A1(n14332), .A2(n14331), .B1(n14330), .B2(n14329), .ZN(
        n14339) );
  INV_X1 U16333 ( .A(n14333), .ZN(n14334) );
  AOI21_X1 U16334 ( .B1(n14336), .B2(n14335), .A(n14334), .ZN(n14469) );
  NOR2_X1 U16335 ( .A1(n14469), .A2(n14337), .ZN(n14338) );
  AOI211_X1 U16336 ( .C1(n14379), .C2(n14340), .A(n14339), .B(n14338), .ZN(
        n14468) );
  INV_X1 U16337 ( .A(n14363), .ZN(n14343) );
  INV_X1 U16338 ( .A(n14341), .ZN(n14342) );
  AOI211_X1 U16339 ( .C1(n14466), .C2(n14343), .A(n14380), .B(n14342), .ZN(
        n14465) );
  INV_X1 U16340 ( .A(n14344), .ZN(n14345) );
  AOI22_X1 U16341 ( .A1(n14352), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14345), 
        .B2(n14397), .ZN(n14346) );
  OAI21_X1 U16342 ( .B1(n14347), .B2(n14368), .A(n14346), .ZN(n14350) );
  NOR2_X1 U16343 ( .A1(n14469), .A2(n14348), .ZN(n14349) );
  AOI211_X1 U16344 ( .C1(n14465), .C2(n14399), .A(n14350), .B(n14349), .ZN(
        n14351) );
  OAI21_X1 U16345 ( .B1(n14468), .B2(n14352), .A(n14351), .ZN(P2_U3247) );
  XNOR2_X1 U16346 ( .A(n14354), .B(n14353), .ZN(n14472) );
  INV_X1 U16347 ( .A(n14472), .ZN(n14372) );
  AND2_X1 U16348 ( .A1(n14356), .A2(n14355), .ZN(n14357) );
  OAI21_X1 U16349 ( .B1(n14358), .B2(n14357), .A(n14379), .ZN(n14362) );
  AOI22_X1 U16350 ( .A1(n14360), .A2(n14374), .B1(n14376), .B2(n14359), .ZN(
        n14361) );
  NAND2_X1 U16351 ( .A1(n14362), .A2(n14361), .ZN(n14470) );
  AOI211_X1 U16352 ( .C1(n14364), .C2(n14382), .A(n14380), .B(n14363), .ZN(
        n14471) );
  NAND2_X1 U16353 ( .A1(n14471), .A2(n14399), .ZN(n14367) );
  AOI22_X1 U16354 ( .A1(n14352), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14365), 
        .B2(n14397), .ZN(n14366) );
  OAI211_X1 U16355 ( .C1(n14546), .C2(n14368), .A(n14367), .B(n14366), .ZN(
        n14369) );
  AOI21_X1 U16356 ( .B1(n14470), .B2(n14396), .A(n14369), .ZN(n14370) );
  OAI21_X1 U16357 ( .B1(n14372), .B2(n14371), .A(n14370), .ZN(P2_U3248) );
  XOR2_X1 U16358 ( .A(n14373), .B(n14389), .Z(n14378) );
  AOI222_X1 U16359 ( .A1(n14379), .A2(n14378), .B1(n14377), .B2(n14376), .C1(
        n14375), .C2(n14374), .ZN(n14480) );
  INV_X1 U16360 ( .A(n14480), .ZN(n14388) );
  AOI21_X1 U16361 ( .B1(n14381), .B2(n14477), .A(n14380), .ZN(n14383) );
  NAND2_X1 U16362 ( .A1(n14383), .A2(n14382), .ZN(n14478) );
  OAI22_X1 U16363 ( .A1(n14478), .A2(n14386), .B1(n14385), .B2(n14384), .ZN(
        n14387) );
  OAI21_X1 U16364 ( .B1(n14388), .B2(n14387), .A(n14396), .ZN(n14393) );
  AOI22_X1 U16365 ( .A1(n14477), .A2(n14401), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n14352), .ZN(n14392) );
  NAND2_X1 U16366 ( .A1(n14390), .A2(n14389), .ZN(n14475) );
  NAND3_X1 U16367 ( .A1(n14476), .A2(n14475), .A3(n14403), .ZN(n14391) );
  NAND3_X1 U16368 ( .A1(n14393), .A2(n14392), .A3(n14391), .ZN(P2_U3249) );
  NOR2_X1 U16369 ( .A1(n14396), .A2(n11056), .ZN(n14394) );
  AOI21_X1 U16370 ( .B1(n14396), .B2(n14395), .A(n14394), .ZN(n14406) );
  AOI22_X1 U16371 ( .A1(n14399), .A2(n14398), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14397), .ZN(n14405) );
  AOI22_X1 U16372 ( .A1(n14403), .A2(n14402), .B1(n14401), .B2(n6421), .ZN(
        n14404) );
  NAND3_X1 U16373 ( .A1(n14406), .A2(n14405), .A3(n14404), .ZN(P2_U3263) );
  INV_X1 U16374 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14408) );
  OAI21_X1 U16375 ( .B1(n14516), .B2(n14487), .A(n14409), .ZN(P2_U3530) );
  INV_X1 U16376 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14412) );
  AND2_X1 U16377 ( .A1(n14411), .A2(n14410), .ZN(n14517) );
  MUX2_X1 U16378 ( .A(n14412), .B(n14517), .S(n15778), .Z(n14413) );
  OAI21_X1 U16379 ( .B1(n14520), .B2(n14487), .A(n14413), .ZN(P2_U3529) );
  AOI21_X1 U16380 ( .B1(n15750), .B2(n14415), .A(n14414), .ZN(n14416) );
  MUX2_X1 U16381 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14521), .S(n15778), .Z(
        P2_U3528) );
  NAND2_X1 U16382 ( .A1(n14420), .A2(n15750), .ZN(n14421) );
  AOI21_X1 U16383 ( .B1(n15750), .B2(n14425), .A(n14424), .ZN(n14426) );
  OAI211_X1 U16384 ( .C1(n15748), .C2(n14428), .A(n14427), .B(n14426), .ZN(
        n14523) );
  MUX2_X1 U16385 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14523), .S(n15778), .Z(
        P2_U3525) );
  AOI211_X1 U16386 ( .C1(n14431), .C2(n15764), .A(n14430), .B(n14429), .ZN(
        n14524) );
  MUX2_X1 U16387 ( .A(n14432), .B(n14524), .S(n15778), .Z(n14433) );
  OAI21_X1 U16388 ( .B1(n14527), .B2(n14487), .A(n14433), .ZN(P2_U3524) );
  AOI21_X1 U16389 ( .B1(n15750), .B2(n14434), .A(n8061), .ZN(n14435) );
  OAI211_X1 U16390 ( .C1(n14437), .C2(n15748), .A(n14436), .B(n14435), .ZN(
        n14528) );
  MUX2_X1 U16391 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14528), .S(n15778), .Z(
        P2_U3523) );
  OAI21_X1 U16392 ( .B1(n14442), .B2(n15748), .A(n14441), .ZN(n14529) );
  MUX2_X1 U16393 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14529), .S(n15778), .Z(
        P2_U3522) );
  NAND2_X1 U16394 ( .A1(n14444), .A2(n14443), .ZN(n14445) );
  AOI21_X1 U16395 ( .B1(n14446), .B2(n15764), .A(n14445), .ZN(n14530) );
  MUX2_X1 U16396 ( .A(n14447), .B(n14530), .S(n15778), .Z(n14448) );
  OAI21_X1 U16397 ( .B1(n14533), .B2(n14487), .A(n14448), .ZN(P2_U3521) );
  AOI211_X1 U16398 ( .C1(n14451), .C2(n15764), .A(n14450), .B(n14449), .ZN(
        n14534) );
  MUX2_X1 U16399 ( .A(n14452), .B(n14534), .S(n15778), .Z(n14453) );
  OAI21_X1 U16400 ( .B1(n14537), .B2(n14487), .A(n14453), .ZN(P2_U3520) );
  AOI211_X1 U16401 ( .C1(n15750), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        n14457) );
  OAI21_X1 U16402 ( .B1(n14458), .B2(n15748), .A(n14457), .ZN(n14538) );
  MUX2_X1 U16403 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14538), .S(n15778), .Z(
        P2_U3519) );
  INV_X1 U16404 ( .A(n14459), .ZN(n14462) );
  AOI211_X1 U16405 ( .C1(n14462), .C2(n6951), .A(n14461), .B(n14460), .ZN(
        n14539) );
  MUX2_X1 U16406 ( .A(n14463), .B(n14539), .S(n15778), .Z(n14464) );
  OAI21_X1 U16407 ( .B1(n7890), .B2(n14487), .A(n14464), .ZN(P2_U3518) );
  AOI21_X1 U16408 ( .B1(n15750), .B2(n14466), .A(n14465), .ZN(n14467) );
  OAI211_X1 U16409 ( .C1(n14469), .C2(n12373), .A(n14468), .B(n14467), .ZN(
        n14542) );
  MUX2_X1 U16410 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14542), .S(n15778), .Z(
        P2_U3517) );
  INV_X1 U16411 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14473) );
  AOI211_X1 U16412 ( .C1(n14472), .C2(n15764), .A(n14471), .B(n14470), .ZN(
        n14543) );
  MUX2_X1 U16413 ( .A(n14473), .B(n14543), .S(n15778), .Z(n14474) );
  OAI21_X1 U16414 ( .B1(n14546), .B2(n14487), .A(n14474), .ZN(P2_U3516) );
  NAND3_X1 U16415 ( .A1(n14476), .A2(n15764), .A3(n14475), .ZN(n14481) );
  NAND2_X1 U16416 ( .A1(n14477), .A2(n15750), .ZN(n14479) );
  NAND4_X1 U16417 ( .A1(n14481), .A2(n14480), .A3(n14479), .A4(n14478), .ZN(
        n14547) );
  MUX2_X1 U16418 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14547), .S(n15778), .Z(
        P2_U3515) );
  AOI211_X1 U16419 ( .C1(n14484), .C2(n15764), .A(n14483), .B(n14482), .ZN(
        n14548) );
  MUX2_X1 U16420 ( .A(n14485), .B(n14548), .S(n15778), .Z(n14486) );
  OAI21_X1 U16421 ( .B1(n6858), .B2(n14487), .A(n14486), .ZN(P2_U3514) );
  AOI211_X1 U16422 ( .C1(n15750), .C2(n14490), .A(n14489), .B(n14488), .ZN(
        n14491) );
  OAI21_X1 U16423 ( .B1(n14492), .B2(n15748), .A(n14491), .ZN(n14552) );
  MUX2_X1 U16424 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14552), .S(n15778), .Z(
        P2_U3513) );
  AOI211_X1 U16425 ( .C1(n15750), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        n14496) );
  OAI21_X1 U16426 ( .B1(n14497), .B2(n15748), .A(n14496), .ZN(n14553) );
  MUX2_X1 U16427 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14553), .S(n15778), .Z(
        P2_U3512) );
  AOI211_X1 U16428 ( .C1(n15750), .C2(n14500), .A(n14499), .B(n14498), .ZN(
        n14501) );
  OAI21_X1 U16429 ( .B1(n14502), .B2(n15748), .A(n14501), .ZN(n14554) );
  MUX2_X1 U16430 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14554), .S(n15778), .Z(
        P2_U3511) );
  AOI21_X1 U16431 ( .B1(n15750), .B2(n14504), .A(n14503), .ZN(n14505) );
  OAI211_X1 U16432 ( .C1(n15748), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14555) );
  MUX2_X1 U16433 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14555), .S(n15778), .Z(
        P2_U3510) );
  AOI21_X1 U16434 ( .B1(n15750), .B2(n14509), .A(n14508), .ZN(n14510) );
  OAI211_X1 U16435 ( .C1(n12373), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14556) );
  MUX2_X1 U16436 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14556), .S(n15778), .Z(
        P2_U3507) );
  OAI21_X1 U16437 ( .B1(n14516), .B2(n14551), .A(n14515), .ZN(P2_U3498) );
  INV_X1 U16438 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14518) );
  MUX2_X1 U16439 ( .A(n14518), .B(n14517), .S(n15767), .Z(n14519) );
  OAI21_X1 U16440 ( .B1(n14520), .B2(n14551), .A(n14519), .ZN(P2_U3497) );
  MUX2_X1 U16441 ( .A(n14522), .B(P2_REG0_REG_27__SCAN_IN), .S(n15765), .Z(
        P2_U3494) );
  MUX2_X1 U16442 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14523), .S(n15767), .Z(
        P2_U3493) );
  INV_X1 U16443 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14525) );
  MUX2_X1 U16444 ( .A(n14525), .B(n14524), .S(n15767), .Z(n14526) );
  OAI21_X1 U16445 ( .B1(n14527), .B2(n14551), .A(n14526), .ZN(P2_U3492) );
  MUX2_X1 U16446 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14528), .S(n15767), .Z(
        P2_U3491) );
  MUX2_X1 U16447 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14529), .S(n15767), .Z(
        P2_U3490) );
  INV_X1 U16448 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14531) );
  MUX2_X1 U16449 ( .A(n14531), .B(n14530), .S(n15767), .Z(n14532) );
  OAI21_X1 U16450 ( .B1(n14533), .B2(n14551), .A(n14532), .ZN(P2_U3489) );
  INV_X1 U16451 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14535) );
  MUX2_X1 U16452 ( .A(n14535), .B(n14534), .S(n15767), .Z(n14536) );
  OAI21_X1 U16453 ( .B1(n14537), .B2(n14551), .A(n14536), .ZN(P2_U3488) );
  MUX2_X1 U16454 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14538), .S(n15767), .Z(
        P2_U3487) );
  INV_X1 U16455 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14540) );
  MUX2_X1 U16456 ( .A(n14540), .B(n14539), .S(n15767), .Z(n14541) );
  OAI21_X1 U16457 ( .B1(n7890), .B2(n14551), .A(n14541), .ZN(P2_U3486) );
  MUX2_X1 U16458 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14542), .S(n15767), .Z(
        P2_U3484) );
  INV_X1 U16459 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14544) );
  MUX2_X1 U16460 ( .A(n14544), .B(n14543), .S(n15767), .Z(n14545) );
  OAI21_X1 U16461 ( .B1(n14546), .B2(n14551), .A(n14545), .ZN(P2_U3481) );
  MUX2_X1 U16462 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14547), .S(n15767), .Z(
        P2_U3478) );
  INV_X1 U16463 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14549) );
  MUX2_X1 U16464 ( .A(n14549), .B(n14548), .S(n15767), .Z(n14550) );
  OAI21_X1 U16465 ( .B1(n6858), .B2(n14551), .A(n14550), .ZN(P2_U3475) );
  MUX2_X1 U16466 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14552), .S(n15767), .Z(
        P2_U3472) );
  MUX2_X1 U16467 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14553), .S(n15767), .Z(
        P2_U3469) );
  MUX2_X1 U16468 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14554), .S(n15767), .Z(
        P2_U3466) );
  MUX2_X1 U16469 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14555), .S(n15767), .Z(
        P2_U3463) );
  MUX2_X1 U16470 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14556), .S(n15767), .Z(
        P2_U3454) );
  INV_X1 U16471 ( .A(n14557), .ZN(n15301) );
  NOR4_X1 U16472 ( .A1(n8889), .A2(P2_IR_REG_30__SCAN_IN), .A3(n10274), .A4(
        P2_U3088), .ZN(n14558) );
  AOI21_X1 U16473 ( .B1(n14565), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14558), 
        .ZN(n14559) );
  OAI21_X1 U16474 ( .B1(n15301), .B2(n14569), .A(n14559), .ZN(P2_U3296) );
  OAI222_X1 U16475 ( .A1(P2_U3088), .A2(n14563), .B1(n14562), .B2(n14561), 
        .C1(n14569), .C2(n14560), .ZN(P2_U3298) );
  AOI21_X1 U16476 ( .B1(n14565), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14564), 
        .ZN(n14566) );
  OAI21_X1 U16477 ( .B1(n14567), .B2(n14569), .A(n14566), .ZN(P2_U3299) );
  INV_X1 U16478 ( .A(n14568), .ZN(n15304) );
  OAI222_X1 U16479 ( .A1(P2_U3088), .A2(n14571), .B1(n14562), .B2(n14570), 
        .C1(n14569), .C2(n15304), .ZN(P2_U3301) );
  INV_X1 U16480 ( .A(n14572), .ZN(n14573) );
  MUX2_X1 U16481 ( .A(n14573), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AND2_X1 U16482 ( .A1(n14722), .A2(n15111), .ZN(n14575) );
  AOI21_X1 U16483 ( .B1(n14839), .B2(n14697), .A(n14575), .ZN(n14872) );
  INV_X1 U16484 ( .A(n14875), .ZN(n14576) );
  AOI22_X1 U16485 ( .A1(n14576), .A2(n14698), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14577) );
  OAI21_X1 U16486 ( .B1(n14872), .B2(n14700), .A(n14577), .ZN(n14578) );
  AOI21_X1 U16487 ( .B1(n15135), .B2(n14689), .A(n14578), .ZN(n14579) );
  INV_X1 U16488 ( .A(n15212), .ZN(n15097) );
  OAI21_X1 U16489 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n14583) );
  NAND2_X1 U16490 ( .A1(n14583), .A2(n14685), .ZN(n14590) );
  OR2_X1 U16491 ( .A1(n14584), .A2(n14675), .ZN(n14585) );
  OAI21_X1 U16492 ( .B1(n14586), .B2(n14706), .A(n14585), .ZN(n15088) );
  NOR2_X1 U16493 ( .A1(n14712), .A2(n15093), .ZN(n14587) );
  AOI211_X1 U16494 ( .C1(n14710), .C2(n15088), .A(n14588), .B(n14587), .ZN(
        n14589) );
  OAI211_X1 U16495 ( .C1(n15097), .C2(n14681), .A(n14590), .B(n14589), .ZN(
        P1_U3215) );
  XOR2_X1 U16496 ( .A(n14592), .B(n14591), .Z(n14598) );
  NOR2_X1 U16497 ( .A1(n14944), .A2(n15579), .ZN(n15158) );
  NOR2_X1 U16498 ( .A1(n14612), .A2(n14675), .ZN(n14593) );
  AOI21_X1 U16499 ( .B1(n14724), .B2(n14697), .A(n14593), .ZN(n14930) );
  INV_X1 U16500 ( .A(n14594), .ZN(n14941) );
  AOI22_X1 U16501 ( .A1(n14941), .A2(n14698), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14595) );
  OAI21_X1 U16502 ( .B1(n14930), .B2(n14700), .A(n14595), .ZN(n14596) );
  AOI21_X1 U16503 ( .B1(n15158), .B2(n14689), .A(n14596), .ZN(n14597) );
  OAI21_X1 U16504 ( .B1(n14598), .B2(n14717), .A(n14597), .ZN(P1_U3216) );
  OAI22_X1 U16505 ( .A1(n14611), .A2(n14706), .B1(n14599), .B2(n14675), .ZN(
        n15179) );
  NAND2_X1 U16506 ( .A1(n15179), .A2(n14710), .ZN(n14600) );
  NAND2_X1 U16507 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14820)
         );
  OAI211_X1 U16508 ( .C1(n14712), .C2(n15010), .A(n14600), .B(n14820), .ZN(
        n14605) );
  AOI211_X1 U16509 ( .C1(n14603), .C2(n14602), .A(n14717), .B(n14601), .ZN(
        n14604) );
  AOI211_X1 U16510 ( .C1(n14714), .C2(n15012), .A(n14605), .B(n14604), .ZN(
        n14606) );
  INV_X1 U16511 ( .A(n14606), .ZN(P1_U3219) );
  INV_X1 U16512 ( .A(n14974), .ZN(n15267) );
  OAI21_X1 U16513 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14610) );
  NAND2_X1 U16514 ( .A1(n14610), .A2(n14685), .ZN(n14617) );
  OAI22_X1 U16515 ( .A1(n14612), .A2(n14706), .B1(n14611), .B2(n14675), .ZN(
        n14971) );
  INV_X1 U16516 ( .A(n14978), .ZN(n14614) );
  OAI22_X1 U16517 ( .A1(n14614), .A2(n14712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14613), .ZN(n14615) );
  AOI21_X1 U16518 ( .B1(n14971), .B2(n14710), .A(n14615), .ZN(n14616) );
  OAI211_X1 U16519 ( .C1(n15267), .C2(n14681), .A(n14617), .B(n14616), .ZN(
        P1_U3223) );
  XOR2_X1 U16520 ( .A(n14619), .B(n14618), .Z(n14624) );
  AOI22_X1 U16521 ( .A1(n14722), .A2(n14697), .B1(n15111), .B2(n14724), .ZN(
        n14898) );
  INV_X1 U16522 ( .A(n14620), .ZN(n14904) );
  AOI22_X1 U16523 ( .A1(n14904), .A2(n14698), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14621) );
  OAI21_X1 U16524 ( .B1(n14898), .B2(n14700), .A(n14621), .ZN(n14622) );
  AOI21_X1 U16525 ( .B1(n14903), .B2(n14714), .A(n14622), .ZN(n14623) );
  OAI21_X1 U16526 ( .B1(n14624), .B2(n14717), .A(n14623), .ZN(P1_U3225) );
  NAND2_X1 U16527 ( .A1(n14626), .A2(n14625), .ZN(n14630) );
  XNOR2_X1 U16528 ( .A(n14627), .B(n14628), .ZN(n14705) );
  OAI22_X1 U16529 ( .A1(n14705), .A2(n14704), .B1(n14628), .B2(n14627), .ZN(
        n14629) );
  XOR2_X1 U16530 ( .A(n14630), .B(n14629), .Z(n14635) );
  AOI22_X1 U16531 ( .A1(n14730), .A2(n14697), .B1(n15111), .B2(n14732), .ZN(
        n15060) );
  NAND2_X1 U16532 ( .A1(n14698), .A2(n15061), .ZN(n14631) );
  OAI211_X1 U16533 ( .C1(n15060), .C2(n14700), .A(n14632), .B(n14631), .ZN(
        n14633) );
  AOI21_X1 U16534 ( .B1(n15200), .B2(n14714), .A(n14633), .ZN(n14634) );
  OAI21_X1 U16535 ( .B1(n14635), .B2(n14717), .A(n14634), .ZN(P1_U3226) );
  INV_X1 U16536 ( .A(n14636), .ZN(n14641) );
  AOI21_X1 U16537 ( .B1(n14638), .B2(n14640), .A(n14637), .ZN(n14639) );
  AOI21_X1 U16538 ( .B1(n14641), .B2(n14640), .A(n14639), .ZN(n14645) );
  NOR2_X1 U16539 ( .A1(n14712), .A2(n15046), .ZN(n14643) );
  AOI22_X1 U16540 ( .A1(n14729), .A2(n14697), .B1(n14731), .B2(n15111), .ZN(
        n15042) );
  NAND2_X1 U16541 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14784)
         );
  OAI21_X1 U16542 ( .B1(n15042), .B2(n14700), .A(n14784), .ZN(n14642) );
  AOI211_X1 U16543 ( .C1(n15045), .C2(n14714), .A(n14643), .B(n14642), .ZN(
        n14644) );
  OAI21_X1 U16544 ( .B1(n14645), .B2(n14717), .A(n14644), .ZN(P1_U3228) );
  XOR2_X1 U16545 ( .A(n14647), .B(n14646), .Z(n14652) );
  AND2_X1 U16546 ( .A1(n14921), .A2(n15598), .ZN(n15154) );
  AND2_X1 U16547 ( .A1(n14725), .A2(n15111), .ZN(n14648) );
  AOI21_X1 U16548 ( .B1(n14723), .B2(n14697), .A(n14648), .ZN(n14918) );
  AOI22_X1 U16549 ( .A1(n14922), .A2(n14698), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14649) );
  OAI21_X1 U16550 ( .B1(n14918), .B2(n14700), .A(n14649), .ZN(n14650) );
  AOI21_X1 U16551 ( .B1(n15154), .B2(n14689), .A(n14650), .ZN(n14651) );
  OAI21_X1 U16552 ( .B1(n14652), .B2(n14717), .A(n14651), .ZN(P1_U3229) );
  AOI22_X1 U16553 ( .A1(n14726), .A2(n14697), .B1(n15111), .B2(n14728), .ZN(
        n14990) );
  AOI22_X1 U16554 ( .A1(n14653), .A2(n14698), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14654) );
  OAI21_X1 U16555 ( .B1(n14990), .B2(n14700), .A(n14654), .ZN(n14659) );
  AOI211_X1 U16556 ( .C1(n14657), .C2(n14656), .A(n14717), .B(n14655), .ZN(
        n14658) );
  AOI211_X1 U16557 ( .C1(n14714), .C2(n14994), .A(n14659), .B(n14658), .ZN(
        n14660) );
  INV_X1 U16558 ( .A(n14660), .ZN(P1_U3233) );
  OAI21_X1 U16559 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(n14664) );
  NAND2_X1 U16560 ( .A1(n14664), .A2(n14685), .ZN(n14670) );
  OAI22_X1 U16561 ( .A1(n14666), .A2(n14706), .B1(n14665), .B2(n14675), .ZN(
        n14950) );
  OAI22_X1 U16562 ( .A1(n14958), .A2(n14712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14667), .ZN(n14668) );
  AOI21_X1 U16563 ( .B1(n14950), .B2(n14710), .A(n14668), .ZN(n14669) );
  OAI211_X1 U16564 ( .C1(n14681), .C2(n15263), .A(n14670), .B(n14669), .ZN(
        P1_U3235) );
  OAI21_X1 U16565 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n14674) );
  NAND2_X1 U16566 ( .A1(n14674), .A2(n14685), .ZN(n14680) );
  OAI22_X1 U16567 ( .A1(n14677), .A2(n14706), .B1(n14676), .B2(n14675), .ZN(
        n15024) );
  NAND2_X1 U16568 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14800)
         );
  OAI21_X1 U16569 ( .B1(n14712), .B2(n15029), .A(n14800), .ZN(n14678) );
  AOI21_X1 U16570 ( .B1(n15024), .B2(n14710), .A(n14678), .ZN(n14679) );
  OAI211_X1 U16571 ( .C1(n15032), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        P1_U3238) );
  NAND2_X1 U16572 ( .A1(n6646), .A2(n14682), .ZN(n14683) );
  XNOR2_X1 U16573 ( .A(n14684), .B(n14683), .ZN(n14686) );
  NAND2_X1 U16574 ( .A1(n14686), .A2(n14685), .ZN(n14695) );
  AOI22_X1 U16575 ( .A1(n14710), .A2(n14687), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14694) );
  NOR2_X1 U16576 ( .A1(n14688), .A2(n15579), .ZN(n15593) );
  NAND2_X1 U16577 ( .A1(n14689), .A2(n15593), .ZN(n14693) );
  INV_X1 U16578 ( .A(n14690), .ZN(n14691) );
  NAND2_X1 U16579 ( .A1(n14698), .A2(n14691), .ZN(n14692) );
  NAND4_X1 U16580 ( .A1(n14695), .A2(n14694), .A3(n14693), .A4(n14692), .ZN(
        P1_U3239) );
  AOI22_X1 U16581 ( .A1(n14721), .A2(n14697), .B1(n15111), .B2(n14723), .ZN(
        n15142) );
  AOI22_X1 U16582 ( .A1(n14885), .A2(n14698), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14699) );
  OAI21_X1 U16583 ( .B1(n15142), .B2(n14700), .A(n14699), .ZN(n14701) );
  AOI21_X1 U16584 ( .B1(n14890), .B2(n14714), .A(n14701), .ZN(n14702) );
  OAI21_X1 U16585 ( .B1(n14703), .B2(n14717), .A(n14702), .ZN(P1_U3240) );
  XNOR2_X1 U16586 ( .A(n14705), .B(n14704), .ZN(n14718) );
  NAND2_X1 U16587 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15481)
         );
  OR2_X1 U16588 ( .A1(n14707), .A2(n14706), .ZN(n14709) );
  NAND2_X1 U16589 ( .A1(n14734), .A2(n15111), .ZN(n14708) );
  NAND2_X1 U16590 ( .A1(n14709), .A2(n14708), .ZN(n15077) );
  NAND2_X1 U16591 ( .A1(n15077), .A2(n14710), .ZN(n14711) );
  OAI211_X1 U16592 ( .C1(n14712), .C2(n15078), .A(n15481), .B(n14711), .ZN(
        n14713) );
  AOI21_X1 U16593 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14716) );
  OAI21_X1 U16594 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(P1_U3241) );
  MUX2_X1 U16595 ( .A(n14719), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14733), .Z(
        P1_U3591) );
  MUX2_X1 U16596 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14841), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16597 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14720), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16598 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14839), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16599 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14721), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16600 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14722), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16601 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14723), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16602 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14724), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16603 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14725), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16604 ( .A(n14726), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14733), .Z(
        P1_U3581) );
  MUX2_X1 U16605 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14727), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16606 ( .A(n14728), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14733), .Z(
        P1_U3579) );
  MUX2_X1 U16607 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14729), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16608 ( .A(n14730), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14733), .Z(
        P1_U3577) );
  MUX2_X1 U16609 ( .A(n14731), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14733), .Z(
        P1_U3576) );
  MUX2_X1 U16610 ( .A(n14732), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14733), .Z(
        P1_U3575) );
  MUX2_X1 U16611 ( .A(n14734), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14733), .Z(
        P1_U3574) );
  MUX2_X1 U16612 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14735), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16613 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14736), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16614 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14737), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16615 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14738), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16616 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14739), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16617 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14740), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16618 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14741), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16619 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14742), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16620 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14743), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16621 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14744), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16622 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14745), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16623 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14746), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16624 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14747), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16625 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15105), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U16626 ( .A(n14748), .ZN(n14763) );
  OAI22_X1 U16627 ( .A1(n15483), .A2(n15316), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14749), .ZN(n14750) );
  AOI21_X1 U16628 ( .B1(n14751), .B2(n15475), .A(n14750), .ZN(n14762) );
  MUX2_X1 U16629 ( .A(n10849), .B(P1_REG2_REG_2__SCAN_IN), .S(n14751), .Z(
        n14754) );
  INV_X1 U16630 ( .A(n14752), .ZN(n14753) );
  NAND2_X1 U16631 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  OAI211_X1 U16632 ( .C1(n14756), .C2(n14755), .A(n15479), .B(n14774), .ZN(
        n14761) );
  OAI211_X1 U16633 ( .C1(n14759), .C2(n14758), .A(n15478), .B(n14757), .ZN(
        n14760) );
  NAND4_X1 U16634 ( .A1(n14763), .A2(n14762), .A3(n14761), .A4(n14760), .ZN(
        P1_U3245) );
  NOR2_X1 U16635 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14764), .ZN(n14767) );
  NOR2_X1 U16636 ( .A1(n14765), .A2(n7034), .ZN(n14766) );
  AOI211_X1 U16637 ( .C1(n14768), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14767), .B(
        n14766), .ZN(n14778) );
  OAI211_X1 U16638 ( .C1(n14771), .C2(n14770), .A(n15478), .B(n14769), .ZN(
        n14777) );
  NAND3_X1 U16639 ( .A1(n14774), .A2(n14773), .A3(n14772), .ZN(n14775) );
  NAND3_X1 U16640 ( .A1(n15479), .A2(n6660), .A3(n14775), .ZN(n14776) );
  NAND3_X1 U16641 ( .A1(n14778), .A2(n14777), .A3(n14776), .ZN(P1_U3246) );
  INV_X1 U16642 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14780) );
  INV_X1 U16643 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15195) );
  XNOR2_X1 U16644 ( .A(n14787), .B(n15195), .ZN(n14782) );
  NAND2_X1 U16645 ( .A1(n14783), .A2(n14782), .ZN(n14796) );
  OAI211_X1 U16646 ( .C1(n14783), .C2(n14782), .A(n14796), .B(n15478), .ZN(
        n14794) );
  INV_X1 U16647 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U16648 ( .B1(n15483), .B2(n14785), .A(n14784), .ZN(n14786) );
  AOI21_X1 U16649 ( .B1(n15475), .B2(n14787), .A(n14786), .ZN(n14793) );
  MUX2_X1 U16650 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n15047), .S(n14787), .Z(
        n14788) );
  OR3_X1 U16651 ( .A1(n14790), .A2(n14789), .A3(n14788), .ZN(n14791) );
  NAND3_X1 U16652 ( .A1(n14795), .A2(n15479), .A3(n14791), .ZN(n14792) );
  NAND3_X1 U16653 ( .A1(n14794), .A2(n14793), .A3(n14792), .ZN(P1_U3260) );
  XNOR2_X1 U16654 ( .A(n14810), .B(n14809), .ZN(n14811) );
  XOR2_X1 U16655 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n14811), .Z(n14806) );
  OAI21_X1 U16656 ( .B1(n14797), .B2(n15195), .A(n14796), .ZN(n14798) );
  OAI211_X1 U16657 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n6553), .A(n6458), .B(
        n15478), .ZN(n14804) );
  INV_X1 U16658 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14801) );
  OAI21_X1 U16659 ( .B1(n15483), .B2(n14801), .A(n14800), .ZN(n14802) );
  AOI21_X1 U16660 ( .B1(n15475), .B2(n14809), .A(n14802), .ZN(n14803) );
  OAI211_X1 U16661 ( .C1(n14806), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        P1_U3261) );
  NAND2_X1 U16662 ( .A1(n14810), .A2(n14809), .ZN(n14814) );
  INV_X1 U16663 ( .A(n14811), .ZN(n14812) );
  NAND2_X1 U16664 ( .A1(n14812), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14813) );
  NAND2_X1 U16665 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  AOI22_X1 U16666 ( .A1(n14818), .A2(n15478), .B1(n15479), .B2(n14816), .ZN(
        n14819) );
  NAND2_X1 U16667 ( .A1(n14821), .A2(n15519), .ZN(n14824) );
  INV_X1 U16668 ( .A(n14822), .ZN(n15124) );
  NOR2_X1 U16669 ( .A1(n15534), .A2(n15124), .ZN(n14829) );
  AOI21_X1 U16670 ( .B1(n15534), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14829), 
        .ZN(n14823) );
  OAI211_X1 U16671 ( .C1(n14825), .C2(n15096), .A(n14824), .B(n14823), .ZN(
        P1_U3263) );
  XNOR2_X1 U16672 ( .A(n14838), .B(n14826), .ZN(n14827) );
  NAND2_X1 U16673 ( .A1(n14827), .A2(n15500), .ZN(n15125) );
  NOR2_X1 U16674 ( .A1(n15249), .A2(n15096), .ZN(n14828) );
  AOI211_X1 U16675 ( .C1(n15534), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14829), 
        .B(n14828), .ZN(n14830) );
  OAI21_X1 U16676 ( .B1(n15125), .B2(n15015), .A(n14830), .ZN(P1_U3264) );
  INV_X1 U16677 ( .A(n14833), .ZN(n14835) );
  NOR2_X1 U16678 ( .A1(n15131), .A2(n15096), .ZN(n14849) );
  NAND2_X1 U16679 ( .A1(n14839), .A2(n15111), .ZN(n15129) );
  NAND2_X1 U16680 ( .A1(n14841), .A2(n14840), .ZN(n15130) );
  NOR2_X1 U16681 ( .A1(n14842), .A2(n15130), .ZN(n14843) );
  AOI21_X1 U16682 ( .B1(n15534), .B2(P1_REG2_REG_29__SCAN_IN), .A(n14843), 
        .ZN(n14847) );
  INV_X1 U16683 ( .A(n14844), .ZN(n14845) );
  NAND3_X1 U16684 ( .A1(n14845), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n15531), 
        .ZN(n14846) );
  OAI211_X1 U16685 ( .C1(n15129), .C2(n15534), .A(n14847), .B(n14846), .ZN(
        n14848) );
  AOI211_X1 U16686 ( .C1(n15128), .C2(n15519), .A(n14849), .B(n14848), .ZN(
        n14855) );
  XNOR2_X1 U16687 ( .A(n14853), .B(n14852), .ZN(n15133) );
  NAND2_X1 U16688 ( .A1(n15133), .A2(n15100), .ZN(n14854) );
  OAI211_X1 U16689 ( .C1(n15134), .C2(n15528), .A(n14855), .B(n14854), .ZN(
        P1_U3356) );
  INV_X1 U16690 ( .A(n14856), .ZN(n14864) );
  NAND2_X1 U16691 ( .A1(n14857), .A2(n15519), .ZN(n14860) );
  AOI22_X1 U16692 ( .A1(n14858), .A2(n15531), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15534), .ZN(n14859) );
  OAI211_X1 U16693 ( .C1(n14861), .C2(n15096), .A(n14860), .B(n14859), .ZN(
        n14862) );
  AOI21_X1 U16694 ( .B1(n6497), .B2(n15100), .A(n14862), .ZN(n14863) );
  OAI21_X1 U16695 ( .B1(n14864), .B2(n15534), .A(n14863), .ZN(P1_U3265) );
  XNOR2_X1 U16696 ( .A(n14865), .B(n14868), .ZN(n15138) );
  INV_X1 U16697 ( .A(n14866), .ZN(n14867) );
  NAND2_X1 U16698 ( .A1(n15513), .A2(n14867), .ZN(n15497) );
  OAI211_X1 U16699 ( .C1(n15138), .C2(n15589), .A(n14873), .B(n14872), .ZN(
        n15140) );
  NAND2_X1 U16700 ( .A1(n15140), .A2(n15513), .ZN(n14882) );
  OAI22_X1 U16701 ( .A1(n14875), .A2(n15511), .B1(n14874), .B2(n15513), .ZN(
        n14879) );
  AOI21_X1 U16702 ( .B1(n14880), .B2(n14887), .A(n15517), .ZN(n14877) );
  NAND2_X1 U16703 ( .A1(n14877), .A2(n14876), .ZN(n15136) );
  NOR2_X1 U16704 ( .A1(n15136), .A2(n15015), .ZN(n14878) );
  AOI211_X1 U16705 ( .C1(n15515), .C2(n14880), .A(n14879), .B(n14878), .ZN(
        n14881) );
  OAI211_X1 U16706 ( .C1(n15138), .C2(n15497), .A(n14882), .B(n14881), .ZN(
        P1_U3266) );
  XNOR2_X1 U16707 ( .A(n14884), .B(n14883), .ZN(n15143) );
  AOI22_X1 U16708 ( .A1(n14885), .A2(n15531), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15534), .ZN(n14886) );
  OAI21_X1 U16709 ( .B1(n15142), .B2(n15534), .A(n14886), .ZN(n14889) );
  OAI211_X1 U16710 ( .C1(n6478), .C2(n15254), .A(n15500), .B(n14887), .ZN(
        n15141) );
  NOR2_X1 U16711 ( .A1(n15141), .A2(n15015), .ZN(n14888) );
  AOI211_X1 U16712 ( .C1(n15515), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        n14894) );
  XNOR2_X1 U16713 ( .A(n14892), .B(n14891), .ZN(n15144) );
  NAND2_X1 U16714 ( .A1(n15144), .A2(n15100), .ZN(n14893) );
  OAI211_X1 U16715 ( .C1(n15143), .C2(n15528), .A(n14894), .B(n14893), .ZN(
        P1_U3267) );
  INV_X1 U16716 ( .A(n15147), .ZN(n14909) );
  INV_X1 U16717 ( .A(n14899), .ZN(n14900) );
  AOI21_X1 U16718 ( .B1(n14902), .B2(n14901), .A(n14900), .ZN(n15149) );
  AOI211_X1 U16719 ( .C1(n14903), .C2(n14919), .A(n15517), .B(n6478), .ZN(
        n15148) );
  NAND2_X1 U16720 ( .A1(n15148), .A2(n15519), .ZN(n14906) );
  AOI22_X1 U16721 ( .A1(n14904), .A2(n15531), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15534), .ZN(n14905) );
  OAI211_X1 U16722 ( .C1(n7641), .C2(n15096), .A(n14906), .B(n14905), .ZN(
        n14907) );
  AOI21_X1 U16723 ( .B1(n15149), .B2(n15100), .A(n14907), .ZN(n14908) );
  OAI21_X1 U16724 ( .B1(n14909), .B2(n15534), .A(n14908), .ZN(P1_U3268) );
  NAND2_X1 U16725 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  NAND2_X1 U16726 ( .A1(n14933), .A2(n14910), .ZN(n14912) );
  OAI21_X1 U16727 ( .B1(n14912), .B2(n14917), .A(n14911), .ZN(n14913) );
  INV_X1 U16728 ( .A(n14913), .ZN(n15157) );
  INV_X1 U16729 ( .A(n14914), .ZN(n14915) );
  AOI211_X1 U16730 ( .C1(n14917), .C2(n14916), .A(n15558), .B(n14915), .ZN(
        n15155) );
  INV_X1 U16731 ( .A(n14918), .ZN(n15152) );
  OAI21_X1 U16732 ( .B1(n15155), .B2(n15152), .A(n15513), .ZN(n14927) );
  AOI21_X1 U16733 ( .B1(n14937), .B2(n14921), .A(n15517), .ZN(n14920) );
  AND2_X1 U16734 ( .A1(n14920), .A2(n14919), .ZN(n15153) );
  INV_X1 U16735 ( .A(n14921), .ZN(n14924) );
  AOI22_X1 U16736 ( .A1(n14922), .A2(n15531), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15534), .ZN(n14923) );
  OAI21_X1 U16737 ( .B1(n14924), .B2(n15096), .A(n14923), .ZN(n14925) );
  AOI21_X1 U16738 ( .B1(n15153), .B2(n15519), .A(n14925), .ZN(n14926) );
  OAI211_X1 U16739 ( .C1(n15157), .C2(n15529), .A(n14927), .B(n14926), .ZN(
        P1_U3269) );
  XNOR2_X1 U16740 ( .A(n14929), .B(n14928), .ZN(n14932) );
  INV_X1 U16741 ( .A(n14930), .ZN(n14931) );
  AOI21_X1 U16742 ( .B1(n14932), .B2(n15604), .A(n14931), .ZN(n15161) );
  OAI21_X1 U16743 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n15160) );
  INV_X1 U16744 ( .A(n14936), .ZN(n14939) );
  INV_X1 U16745 ( .A(n14937), .ZN(n14938) );
  AOI211_X1 U16746 ( .C1(n14940), .C2(n14939), .A(n15517), .B(n14938), .ZN(
        n15159) );
  NAND2_X1 U16747 ( .A1(n15159), .A2(n15519), .ZN(n14943) );
  AOI22_X1 U16748 ( .A1(n14941), .A2(n15531), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15534), .ZN(n14942) );
  OAI211_X1 U16749 ( .C1(n14944), .C2(n15096), .A(n14943), .B(n14942), .ZN(
        n14945) );
  AOI21_X1 U16750 ( .B1(n15160), .B2(n15100), .A(n14945), .ZN(n14946) );
  OAI21_X1 U16751 ( .B1(n15161), .B2(n15534), .A(n14946), .ZN(P1_U3270) );
  INV_X1 U16752 ( .A(n14947), .ZN(n14948) );
  AOI21_X1 U16753 ( .B1(n14954), .B2(n14949), .A(n14948), .ZN(n14952) );
  INV_X1 U16754 ( .A(n14950), .ZN(n14951) );
  OAI21_X1 U16755 ( .B1(n14952), .B2(n15558), .A(n14951), .ZN(n15163) );
  INV_X1 U16756 ( .A(n15163), .ZN(n14964) );
  OAI21_X1 U16757 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(n15165) );
  INV_X1 U16758 ( .A(n14977), .ZN(n14956) );
  AOI211_X1 U16759 ( .C1(n14957), .C2(n14956), .A(n15517), .B(n14936), .ZN(
        n15164) );
  NAND2_X1 U16760 ( .A1(n15164), .A2(n15519), .ZN(n14961) );
  INV_X1 U16761 ( .A(n14958), .ZN(n14959) );
  AOI22_X1 U16762 ( .A1(n14959), .A2(n15531), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15534), .ZN(n14960) );
  OAI211_X1 U16763 ( .C1(n15096), .C2(n15263), .A(n14961), .B(n14960), .ZN(
        n14962) );
  AOI21_X1 U16764 ( .B1(n15165), .B2(n15100), .A(n14962), .ZN(n14963) );
  OAI21_X1 U16765 ( .B1(n14964), .B2(n15534), .A(n14963), .ZN(P1_U3271) );
  XNOR2_X1 U16766 ( .A(n14965), .B(n14967), .ZN(n15170) );
  INV_X1 U16767 ( .A(n15170), .ZN(n14983) );
  NAND3_X1 U16768 ( .A1(n14966), .A2(n10387), .A3(n14968), .ZN(n14969) );
  NAND3_X1 U16769 ( .A1(n14970), .A2(n15604), .A3(n14969), .ZN(n14973) );
  INV_X1 U16770 ( .A(n14971), .ZN(n14972) );
  NAND2_X1 U16771 ( .A1(n14973), .A2(n14972), .ZN(n15168) );
  NAND2_X1 U16772 ( .A1(n6473), .A2(n14974), .ZN(n14975) );
  NAND2_X1 U16773 ( .A1(n14975), .A2(n15500), .ZN(n14976) );
  NOR2_X1 U16774 ( .A1(n14977), .A2(n14976), .ZN(n15169) );
  NAND2_X1 U16775 ( .A1(n15169), .A2(n15519), .ZN(n14980) );
  AOI22_X1 U16776 ( .A1(n14978), .A2(n15531), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15534), .ZN(n14979) );
  OAI211_X1 U16777 ( .C1(n15267), .C2(n15096), .A(n14980), .B(n14979), .ZN(
        n14981) );
  AOI21_X1 U16778 ( .B1(n15168), .B2(n15513), .A(n14981), .ZN(n14982) );
  OAI21_X1 U16779 ( .B1(n14983), .B2(n15529), .A(n14982), .ZN(P1_U3272) );
  NAND2_X1 U16780 ( .A1(n14984), .A2(n10333), .ZN(n14985) );
  NAND2_X1 U16781 ( .A1(n14986), .A2(n14985), .ZN(n15173) );
  NAND2_X1 U16782 ( .A1(n14988), .A2(n14987), .ZN(n14989) );
  NAND3_X1 U16783 ( .A1(n14966), .A2(n15604), .A3(n14989), .ZN(n14991) );
  NAND2_X1 U16784 ( .A1(n14991), .A2(n14990), .ZN(n15176) );
  NOR2_X1 U16785 ( .A1(n14992), .A2(n15511), .ZN(n14993) );
  OAI21_X1 U16786 ( .B1(n15176), .B2(n14993), .A(n15513), .ZN(n14999) );
  AOI21_X1 U16787 ( .B1(n6510), .B2(n14994), .A(n15517), .ZN(n14995) );
  AND2_X1 U16788 ( .A1(n14995), .A2(n6473), .ZN(n15174) );
  INV_X1 U16789 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14996) );
  OAI22_X1 U16790 ( .A1(n15271), .A2(n15096), .B1(n15513), .B2(n14996), .ZN(
        n14997) );
  AOI21_X1 U16791 ( .B1(n15174), .B2(n15519), .A(n14997), .ZN(n14998) );
  OAI211_X1 U16792 ( .C1(n15173), .C2(n15529), .A(n14999), .B(n14998), .ZN(
        P1_U3273) );
  XNOR2_X1 U16793 ( .A(n15000), .B(n15001), .ZN(n15186) );
  AOI21_X1 U16794 ( .B1(n15074), .B2(n15004), .A(n15003), .ZN(n15018) );
  INV_X1 U16795 ( .A(n15005), .ZN(n15007) );
  OAI21_X1 U16796 ( .B1(n15018), .B2(n15007), .A(n15006), .ZN(n15009) );
  NAND2_X1 U16797 ( .A1(n15009), .A2(n15008), .ZN(n15184) );
  OAI211_X1 U16798 ( .C1(n15027), .C2(n15182), .A(n15500), .B(n6510), .ZN(
        n15181) );
  OAI22_X1 U16799 ( .A1(n7036), .A2(n15513), .B1(n15010), .B2(n15511), .ZN(
        n15011) );
  AOI21_X1 U16800 ( .B1(n15179), .B2(n15513), .A(n15011), .ZN(n15014) );
  NAND2_X1 U16801 ( .A1(n15012), .A2(n15515), .ZN(n15013) );
  OAI211_X1 U16802 ( .C1(n15181), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        n15016) );
  AOI21_X1 U16803 ( .B1(n15184), .B2(n15075), .A(n15016), .ZN(n15017) );
  OAI21_X1 U16804 ( .B1(n15529), .B2(n15186), .A(n15017), .ZN(P1_U3274) );
  NOR2_X1 U16805 ( .A1(n15018), .A2(n15558), .ZN(n15026) );
  NOR2_X1 U16806 ( .A1(n15002), .A2(n15019), .ZN(n15023) );
  INV_X1 U16807 ( .A(n15033), .ZN(n15021) );
  OAI211_X1 U16808 ( .C1(n15023), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15025) );
  AOI21_X1 U16809 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15190) );
  INV_X1 U16810 ( .A(n15044), .ZN(n15028) );
  AOI211_X1 U16811 ( .C1(n15188), .C2(n15028), .A(n15517), .B(n15027), .ZN(
        n15187) );
  INV_X1 U16812 ( .A(n15029), .ZN(n15030) );
  AOI22_X1 U16813 ( .A1(n15534), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15030), 
        .B2(n15531), .ZN(n15031) );
  OAI21_X1 U16814 ( .B1(n15032), .B2(n15096), .A(n15031), .ZN(n15035) );
  XNOR2_X1 U16815 ( .A(n6459), .B(n15033), .ZN(n15191) );
  NOR2_X1 U16816 ( .A1(n15191), .A2(n15529), .ZN(n15034) );
  AOI211_X1 U16817 ( .C1(n15187), .C2(n15519), .A(n15035), .B(n15034), .ZN(
        n15036) );
  OAI21_X1 U16818 ( .B1(n15190), .B2(n15534), .A(n15036), .ZN(P1_U3275) );
  XNOR2_X1 U16819 ( .A(n15037), .B(n15041), .ZN(n15194) );
  INV_X1 U16820 ( .A(n15194), .ZN(n15052) );
  NOR2_X1 U16821 ( .A1(n15074), .A2(n15073), .ZN(n15072) );
  INV_X1 U16822 ( .A(n10372), .ZN(n15038) );
  NOR2_X1 U16823 ( .A1(n15072), .A2(n15038), .ZN(n15056) );
  NAND2_X1 U16824 ( .A1(n15056), .A2(n15055), .ZN(n15054) );
  NAND2_X1 U16825 ( .A1(n15054), .A2(n15039), .ZN(n15040) );
  XOR2_X1 U16826 ( .A(n15041), .B(n15040), .Z(n15043) );
  OAI21_X1 U16827 ( .B1(n15043), .B2(n15558), .A(n15042), .ZN(n15192) );
  NAND2_X1 U16828 ( .A1(n15192), .A2(n15513), .ZN(n15051) );
  AOI211_X1 U16829 ( .C1(n15045), .C2(n15058), .A(n15517), .B(n15044), .ZN(
        n15193) );
  NOR2_X1 U16830 ( .A1(n7636), .A2(n15096), .ZN(n15049) );
  OAI22_X1 U16831 ( .A1(n15513), .A2(n15047), .B1(n15046), .B2(n15511), .ZN(
        n15048) );
  AOI211_X1 U16832 ( .C1(n15193), .C2(n15519), .A(n15049), .B(n15048), .ZN(
        n15050) );
  OAI211_X1 U16833 ( .C1(n15052), .C2(n15529), .A(n15051), .B(n15050), .ZN(
        P1_U3276) );
  XNOR2_X1 U16834 ( .A(n15053), .B(n15055), .ZN(n15203) );
  OAI21_X1 U16835 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15197) );
  NAND2_X1 U16836 ( .A1(n15197), .A2(n15075), .ZN(n15067) );
  INV_X1 U16837 ( .A(n15058), .ZN(n15059) );
  AOI211_X1 U16838 ( .C1(n15200), .C2(n15057), .A(n15517), .B(n15059), .ZN(
        n15198) );
  INV_X1 U16839 ( .A(n15060), .ZN(n15199) );
  AOI22_X1 U16840 ( .A1(n15199), .A2(n15513), .B1(n15061), .B2(n15531), .ZN(
        n15063) );
  NAND2_X1 U16841 ( .A1(n15534), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15062) );
  OAI211_X1 U16842 ( .C1(n15064), .C2(n15096), .A(n15063), .B(n15062), .ZN(
        n15065) );
  AOI21_X1 U16843 ( .B1(n15198), .B2(n15519), .A(n15065), .ZN(n15066) );
  OAI211_X1 U16844 ( .C1(n15203), .C2(n15529), .A(n15067), .B(n15066), .ZN(
        P1_U3277) );
  NOR2_X1 U16845 ( .A1(n15068), .A2(n15099), .ZN(n15216) );
  NOR2_X1 U16846 ( .A1(n15216), .A2(n15069), .ZN(n15071) );
  XNOR2_X1 U16847 ( .A(n15071), .B(n15070), .ZN(n15206) );
  AOI21_X1 U16848 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15208) );
  NAND2_X1 U16849 ( .A1(n15208), .A2(n15075), .ZN(n15084) );
  OAI211_X1 U16850 ( .C1(n15076), .C2(n15281), .A(n15500), .B(n15057), .ZN(
        n15204) );
  INV_X1 U16851 ( .A(n15204), .ZN(n15082) );
  INV_X1 U16852 ( .A(n15077), .ZN(n15205) );
  OAI22_X1 U16853 ( .A1(n15205), .A2(n15534), .B1(n15078), .B2(n15511), .ZN(
        n15079) );
  AOI21_X1 U16854 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15534), .A(n15079), 
        .ZN(n15080) );
  OAI21_X1 U16855 ( .B1(n15281), .B2(n15096), .A(n15080), .ZN(n15081) );
  AOI21_X1 U16856 ( .B1(n15082), .B2(n15519), .A(n15081), .ZN(n15083) );
  OAI211_X1 U16857 ( .C1(n15206), .C2(n15529), .A(n15084), .B(n15083), .ZN(
        P1_U3278) );
  INV_X1 U16858 ( .A(n15085), .ZN(n15087) );
  INV_X1 U16859 ( .A(n15099), .ZN(n15086) );
  AOI21_X1 U16860 ( .B1(n15087), .B2(n15086), .A(n15558), .ZN(n15090) );
  AOI21_X1 U16861 ( .B1(n15090), .B2(n15089), .A(n15088), .ZN(n15214) );
  XNOR2_X1 U16862 ( .A(n15091), .B(n15212), .ZN(n15092) );
  NOR2_X1 U16863 ( .A1(n15092), .A2(n15517), .ZN(n15211) );
  INV_X1 U16864 ( .A(n15093), .ZN(n15094) );
  AOI22_X1 U16865 ( .A1(n15534), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15094), 
        .B2(n15531), .ZN(n15095) );
  OAI21_X1 U16866 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15098) );
  AOI21_X1 U16867 ( .B1(n15211), .B2(n15519), .A(n15098), .ZN(n15103) );
  INV_X1 U16868 ( .A(n15216), .ZN(n15101) );
  NAND2_X1 U16869 ( .A1(n15068), .A2(n15099), .ZN(n15210) );
  NAND3_X1 U16870 ( .A1(n15101), .A2(n15100), .A3(n15210), .ZN(n15102) );
  OAI211_X1 U16871 ( .C1(n15214), .C2(n15534), .A(n15103), .B(n15102), .ZN(
        P1_U3279) );
  XNOR2_X1 U16872 ( .A(n15106), .B(n15104), .ZN(n15547) );
  AOI21_X1 U16873 ( .B1(n15106), .B2(n15105), .A(n15558), .ZN(n15112) );
  OAI21_X1 U16874 ( .B1(n15549), .B2(n15525), .A(n15107), .ZN(n15118) );
  XNOR2_X1 U16875 ( .A(n15118), .B(n10301), .ZN(n15109) );
  OAI21_X1 U16876 ( .B1(n15109), .B2(n15558), .A(n15108), .ZN(n15110) );
  OAI21_X1 U16877 ( .B1(n15112), .B2(n15111), .A(n15110), .ZN(n15114) );
  OAI211_X1 U16878 ( .C1(n15547), .C2(n15589), .A(n15114), .B(n15113), .ZN(
        n15550) );
  NAND2_X1 U16879 ( .A1(n15550), .A2(n15513), .ZN(n15123) );
  OAI22_X1 U16880 ( .A1(n15513), .A2(n8213), .B1(n15115), .B2(n15511), .ZN(
        n15116) );
  AOI21_X1 U16881 ( .B1(n15515), .B2(n15117), .A(n15116), .ZN(n15122) );
  OR2_X1 U16882 ( .A1(n15547), .A2(n15497), .ZN(n15121) );
  OR2_X1 U16883 ( .A1(n15118), .A2(n15517), .ZN(n15548) );
  INV_X1 U16884 ( .A(n15548), .ZN(n15119) );
  NAND2_X1 U16885 ( .A1(n15519), .A2(n15119), .ZN(n15120) );
  NAND4_X1 U16886 ( .A1(n15123), .A2(n15122), .A3(n15121), .A4(n15120), .ZN(
        P1_U3292) );
  MUX2_X1 U16887 ( .A(n15126), .B(n15246), .S(n15618), .Z(n15127) );
  OAI21_X1 U16888 ( .B1(n15249), .B2(n15228), .A(n15127), .ZN(P1_U3558) );
  OAI211_X1 U16889 ( .C1(n15131), .C2(n15579), .A(n15130), .B(n15129), .ZN(
        n15132) );
  INV_X1 U16890 ( .A(n15135), .ZN(n15137) );
  OAI211_X1 U16891 ( .C1(n15138), .C2(n15588), .A(n15137), .B(n15136), .ZN(
        n15139) );
  OR2_X2 U16892 ( .A1(n15140), .A2(n15139), .ZN(n15251) );
  MUX2_X1 U16893 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15251), .S(n15618), .Z(
        P1_U3555) );
  MUX2_X1 U16894 ( .A(n15145), .B(n15252), .S(n15618), .Z(n15146) );
  OAI21_X1 U16895 ( .B1(n15254), .B2(n15228), .A(n15146), .ZN(P1_U3554) );
  MUX2_X1 U16896 ( .A(n15150), .B(n15255), .S(n15618), .Z(n15151) );
  OAI21_X1 U16897 ( .B1(n7641), .B2(n15228), .A(n15151), .ZN(P1_U3553) );
  NOR4_X1 U16898 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15156) );
  OAI21_X1 U16899 ( .B1(n15601), .B2(n15157), .A(n15156), .ZN(n15258) );
  MUX2_X1 U16900 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15258), .S(n15618), .Z(
        P1_U3552) );
  AOI211_X1 U16901 ( .C1(n15160), .C2(n15572), .A(n15159), .B(n15158), .ZN(
        n15162) );
  NAND2_X1 U16902 ( .A1(n15162), .A2(n15161), .ZN(n15259) );
  MUX2_X1 U16903 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15259), .S(n15618), .Z(
        P1_U3551) );
  INV_X1 U16904 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15166) );
  AOI211_X1 U16905 ( .C1(n15572), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        n15260) );
  MUX2_X1 U16906 ( .A(n15166), .B(n15260), .S(n15618), .Z(n15167) );
  OAI21_X1 U16907 ( .B1(n15228), .B2(n15263), .A(n15167), .ZN(P1_U3550) );
  AOI211_X1 U16908 ( .C1(n15572), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15264) );
  MUX2_X1 U16909 ( .A(n15171), .B(n15264), .S(n15618), .Z(n15172) );
  OAI21_X1 U16910 ( .B1(n15267), .B2(n15228), .A(n15172), .ZN(P1_U3549) );
  NOR2_X1 U16911 ( .A1(n15173), .A2(n15601), .ZN(n15175) );
  NOR3_X1 U16912 ( .A1(n15176), .A2(n15175), .A3(n15174), .ZN(n15269) );
  MUX2_X1 U16913 ( .A(n15269), .B(n15177), .S(n15615), .Z(n15178) );
  OAI21_X1 U16914 ( .B1(n15271), .B2(n15228), .A(n15178), .ZN(P1_U3548) );
  INV_X1 U16915 ( .A(n15179), .ZN(n15180) );
  OAI211_X1 U16916 ( .C1(n15182), .C2(n15579), .A(n15181), .B(n15180), .ZN(
        n15183) );
  AOI21_X1 U16917 ( .B1(n15184), .B2(n15604), .A(n15183), .ZN(n15185) );
  OAI21_X1 U16918 ( .B1(n15601), .B2(n15186), .A(n15185), .ZN(n15272) );
  MUX2_X1 U16919 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15272), .S(n15618), .Z(
        P1_U3547) );
  AOI21_X1 U16920 ( .B1(n15598), .B2(n15188), .A(n15187), .ZN(n15189) );
  OAI211_X1 U16921 ( .C1(n15601), .C2(n15191), .A(n15190), .B(n15189), .ZN(
        n15273) );
  MUX2_X1 U16922 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15273), .S(n15618), .Z(
        P1_U3546) );
  AOI211_X1 U16923 ( .C1(n15572), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15274) );
  MUX2_X1 U16924 ( .A(n15195), .B(n15274), .S(n15618), .Z(n15196) );
  OAI21_X1 U16925 ( .B1(n7636), .B2(n15228), .A(n15196), .ZN(P1_U3545) );
  NAND2_X1 U16926 ( .A1(n15197), .A2(n15604), .ZN(n15202) );
  AOI211_X1 U16927 ( .C1(n15598), .C2(n15200), .A(n15199), .B(n15198), .ZN(
        n15201) );
  OAI211_X1 U16928 ( .C1(n15601), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15277) );
  MUX2_X1 U16929 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15277), .S(n15618), .Z(
        P1_U3544) );
  OAI211_X1 U16930 ( .C1(n15206), .C2(n15601), .A(n15205), .B(n15204), .ZN(
        n15207) );
  AOI21_X1 U16931 ( .B1(n15208), .B2(n15604), .A(n15207), .ZN(n15278) );
  MUX2_X1 U16932 ( .A(n15473), .B(n15278), .S(n15618), .Z(n15209) );
  OAI21_X1 U16933 ( .B1(n15281), .B2(n15228), .A(n15209), .ZN(P1_U3543) );
  NAND2_X1 U16934 ( .A1(n15210), .A2(n15572), .ZN(n15215) );
  AOI21_X1 U16935 ( .B1(n15598), .B2(n15212), .A(n15211), .ZN(n15213) );
  OAI211_X1 U16936 ( .C1(n15216), .C2(n15215), .A(n15214), .B(n15213), .ZN(
        n15282) );
  MUX2_X1 U16937 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15282), .S(n15618), .Z(
        P1_U3542) );
  AOI211_X1 U16938 ( .C1(n15572), .C2(n15219), .A(n15218), .B(n15217), .ZN(
        n15283) );
  MUX2_X1 U16939 ( .A(n15220), .B(n15283), .S(n15618), .Z(n15221) );
  OAI21_X1 U16940 ( .B1(n15286), .B2(n15228), .A(n15221), .ZN(P1_U3541) );
  NAND2_X1 U16941 ( .A1(n15222), .A2(n15572), .ZN(n15224) );
  OAI211_X1 U16942 ( .C1(n15225), .C2(n15579), .A(n15224), .B(n15223), .ZN(
        n15226) );
  OR2_X1 U16943 ( .A1(n15227), .A2(n15226), .ZN(n15287) );
  MUX2_X1 U16944 ( .A(n15287), .B(P1_REG1_REG_12__SCAN_IN), .S(n15615), .Z(
        P1_U3540) );
  OAI211_X1 U16945 ( .C1(n15601), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        n15289) );
  MUX2_X1 U16946 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15289), .S(n15618), .Z(
        n15232) );
  AOI21_X1 U16947 ( .B1(n10399), .B2(n15291), .A(n15232), .ZN(n15233) );
  INV_X1 U16948 ( .A(n15233), .ZN(P1_U3539) );
  NAND2_X1 U16949 ( .A1(n15234), .A2(n15598), .ZN(n15235) );
  AND4_X1 U16950 ( .A1(n15238), .A2(n15237), .A3(n15236), .A4(n15235), .ZN(
        n15239) );
  OAI21_X1 U16951 ( .B1(n15601), .B2(n15240), .A(n15239), .ZN(n15293) );
  MUX2_X1 U16952 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15293), .S(n15618), .Z(
        P1_U3538) );
  AOI21_X1 U16953 ( .B1(n15598), .B2(n15242), .A(n15241), .ZN(n15243) );
  OAI211_X1 U16954 ( .C1(n15601), .C2(n15245), .A(n15244), .B(n15243), .ZN(
        n15294) );
  MUX2_X1 U16955 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15294), .S(n15618), .Z(
        P1_U3537) );
  INV_X1 U16956 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15247) );
  MUX2_X1 U16957 ( .A(n15247), .B(n15246), .S(n15606), .Z(n15248) );
  OAI21_X1 U16958 ( .B1(n15249), .B2(n15288), .A(n15248), .ZN(P1_U3526) );
  MUX2_X1 U16959 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15250), .S(n15606), .Z(
        P1_U3525) );
  MUX2_X1 U16960 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15251), .S(n15606), .Z(
        P1_U3523) );
  INV_X1 U16961 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15253) );
  INV_X1 U16962 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15256) );
  MUX2_X1 U16963 ( .A(n15256), .B(n15255), .S(n15606), .Z(n15257) );
  OAI21_X1 U16964 ( .B1(n7641), .B2(n15288), .A(n15257), .ZN(P1_U3521) );
  MUX2_X1 U16965 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15258), .S(n15606), .Z(
        P1_U3520) );
  MUX2_X1 U16966 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15259), .S(n15606), .Z(
        P1_U3519) );
  MUX2_X1 U16967 ( .A(n15261), .B(n15260), .S(n15606), .Z(n15262) );
  OAI21_X1 U16968 ( .B1(n15288), .B2(n15263), .A(n15262), .ZN(P1_U3518) );
  INV_X1 U16969 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15265) );
  MUX2_X1 U16970 ( .A(n15265), .B(n15264), .S(n15606), .Z(n15266) );
  OAI21_X1 U16971 ( .B1(n15267), .B2(n15288), .A(n15266), .ZN(P1_U3517) );
  INV_X1 U16972 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15268) );
  MUX2_X1 U16973 ( .A(n15269), .B(n15268), .S(n15605), .Z(n15270) );
  OAI21_X1 U16974 ( .B1(n15271), .B2(n15288), .A(n15270), .ZN(P1_U3516) );
  MUX2_X1 U16975 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15272), .S(n15606), .Z(
        P1_U3515) );
  MUX2_X1 U16976 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15273), .S(n15606), .Z(
        P1_U3513) );
  INV_X1 U16977 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15275) );
  MUX2_X1 U16978 ( .A(n15275), .B(n15274), .S(n15606), .Z(n15276) );
  OAI21_X1 U16979 ( .B1(n7636), .B2(n15288), .A(n15276), .ZN(P1_U3510) );
  MUX2_X1 U16980 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15277), .S(n15606), .Z(
        P1_U3507) );
  MUX2_X1 U16981 ( .A(n15279), .B(n15278), .S(n15606), .Z(n15280) );
  OAI21_X1 U16982 ( .B1(n15281), .B2(n15288), .A(n15280), .ZN(P1_U3504) );
  MUX2_X1 U16983 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15282), .S(n15606), .Z(
        P1_U3501) );
  INV_X1 U16984 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15284) );
  MUX2_X1 U16985 ( .A(n15284), .B(n15283), .S(n15606), .Z(n15285) );
  OAI21_X1 U16986 ( .B1(n15286), .B2(n15288), .A(n15285), .ZN(P1_U3498) );
  MUX2_X1 U16987 ( .A(n15287), .B(P1_REG0_REG_12__SCAN_IN), .S(n15605), .Z(
        P1_U3495) );
  MUX2_X1 U16988 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15289), .S(n15606), .Z(
        n15290) );
  AOI21_X1 U16989 ( .B1(n10118), .B2(n15291), .A(n15290), .ZN(n15292) );
  INV_X1 U16990 ( .A(n15292), .ZN(P1_U3492) );
  MUX2_X1 U16991 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15293), .S(n15606), .Z(
        P1_U3489) );
  MUX2_X1 U16992 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15294), .S(n15606), .Z(
        P1_U3486) );
  INV_X1 U16993 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15296) );
  NOR4_X1 U16994 ( .A1(n15297), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15296), .A4(
        P1_U3086), .ZN(n15298) );
  AOI21_X1 U16995 ( .B1(n15299), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15298), 
        .ZN(n15300) );
  OAI21_X1 U16996 ( .B1(n15301), .B2(n15305), .A(n15300), .ZN(P1_U3324) );
  OAI222_X1 U16997 ( .A1(n15305), .A2(n15303), .B1(n15307), .B2(n15302), .C1(
        P1_U3086), .C2(n10101), .ZN(P1_U3328) );
  OAI222_X1 U16998 ( .A1(P1_U3086), .A2(n15308), .B1(n15307), .B2(n15306), 
        .C1(n15305), .C2(n15304), .ZN(P1_U3329) );
  MUX2_X1 U16999 ( .A(n15309), .B(n12651), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U17000 ( .A(n15310), .ZN(n15311) );
  MUX2_X1 U17001 ( .A(n15311), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U17002 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15484) );
  NOR2_X1 U17003 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15484), .ZN(n15345) );
  INV_X1 U17004 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15343) );
  XOR2_X1 U17005 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n15343), .Z(n15407) );
  INV_X1 U17006 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U17007 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n15339), .ZN(n15312) );
  AOI21_X1 U17008 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15339), .A(n15312), 
        .ZN(n15355) );
  INV_X1 U17009 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15337) );
  INV_X1 U17010 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15333) );
  XOR2_X1 U17011 ( .A(n15333), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n15395) );
  XOR2_X1 U17012 ( .A(n15332), .B(P1_ADDR_REG_8__SCAN_IN), .Z(n15360) );
  NAND2_X1 U17013 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n15313), .ZN(n15327) );
  INV_X1 U17014 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15314) );
  AOI22_X1 U17015 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15314), .B1(
        P3_ADDR_REG_6__SCAN_IN), .B2(n15313), .ZN(n15384) );
  INV_X1 U17016 ( .A(n15369), .ZN(n15315) );
  NAND2_X1 U17017 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15318), .ZN(n15319) );
  NAND2_X1 U17018 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15320), .ZN(n15322) );
  NAND2_X1 U17019 ( .A1(n15363), .A2(n15364), .ZN(n15321) );
  NAND2_X1 U17020 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15323), .ZN(n15325) );
  NAND2_X1 U17021 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15328), .ZN(n15330) );
  INV_X1 U17022 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15389) );
  XOR2_X1 U17023 ( .A(n15337), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n15398) );
  NAND2_X1 U17024 ( .A1(n15399), .A2(n15398), .ZN(n15336) );
  NAND2_X1 U17025 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15402), .ZN(n15340) );
  NAND2_X1 U17026 ( .A1(n15407), .A2(n15406), .ZN(n15342) );
  INV_X1 U17027 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15344) );
  OAI22_X2 U17028 ( .A1(n15345), .A2(n15352), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n15344), .ZN(n15346) );
  NOR2_X1 U17029 ( .A1(n12065), .A2(n15346), .ZN(n15348) );
  XNOR2_X1 U17030 ( .A(n12065), .B(n15346), .ZN(n15409) );
  NOR2_X1 U17031 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15409), .ZN(n15347) );
  NAND2_X1 U17032 ( .A1(n15349), .A2(n14785), .ZN(n15351) );
  XOR2_X1 U17033 ( .A(n14785), .B(n15349), .Z(n15410) );
  NAND2_X1 U17034 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15410), .ZN(n15350) );
  NAND2_X1 U17035 ( .A1(n15351), .A2(n15350), .ZN(n15437) );
  INV_X1 U17036 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15440) );
  XOR2_X1 U17037 ( .A(n15440), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n15438) );
  XOR2_X1 U17038 ( .A(n15484), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n15353) );
  XNOR2_X1 U17039 ( .A(n15353), .B(n15352), .ZN(n15463) );
  XOR2_X1 U17040 ( .A(n15355), .B(n15354), .Z(n15451) );
  INV_X1 U17041 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15359) );
  NOR2_X1 U17042 ( .A1(n15357), .A2(n15356), .ZN(n15358) );
  XNOR2_X1 U17043 ( .A(n15359), .B(n15358), .ZN(n15431) );
  XOR2_X1 U17044 ( .A(n15361), .B(n15360), .Z(n15392) );
  INV_X1 U17045 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15660) );
  NAND2_X1 U17046 ( .A1(n15365), .A2(n15660), .ZN(n15377) );
  INV_X1 U17047 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15632) );
  NOR2_X1 U17048 ( .A1(n15371), .A2(n15632), .ZN(n15372) );
  OAI21_X1 U17049 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n15370), .A(n15369), .ZN(
        n15879) );
  NAND2_X1 U17050 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15879), .ZN(n15888) );
  NAND2_X1 U17051 ( .A1(n15417), .A2(n15416), .ZN(n15373) );
  NOR2_X1 U17052 ( .A1(n15417), .A2(n15416), .ZN(n15415) );
  XOR2_X1 U17053 ( .A(n15375), .B(n15374), .Z(n15883) );
  NAND2_X1 U17054 ( .A1(n15884), .A2(n15883), .ZN(n15882) );
  NAND2_X1 U17055 ( .A1(n15378), .A2(n15380), .ZN(n15381) );
  INV_X1 U17056 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15877) );
  INV_X1 U17057 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15382) );
  NOR2_X1 U17058 ( .A1(n15383), .A2(n15382), .ZN(n15386) );
  XOR2_X1 U17059 ( .A(n15385), .B(n15384), .Z(n15421) );
  INV_X1 U17060 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U17061 ( .A1(n15388), .A2(n15387), .ZN(n15391) );
  XOR2_X1 U17062 ( .A(n15390), .B(n15389), .Z(n15880) );
  INV_X1 U17063 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15424) );
  XOR2_X1 U17064 ( .A(n15396), .B(n15395), .Z(n15426) );
  XNOR2_X1 U17065 ( .A(n15399), .B(n15398), .ZN(n15400) );
  NOR2_X2 U17066 ( .A1(n15401), .A2(n15400), .ZN(n15446) );
  NAND2_X1 U17067 ( .A1(n15451), .A2(n15452), .ZN(n15450) );
  XNOR2_X1 U17068 ( .A(n15402), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n15403) );
  XNOR2_X1 U17069 ( .A(n15404), .B(n15403), .ZN(n15455) );
  INV_X1 U17070 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15405) );
  XNOR2_X1 U17071 ( .A(n15407), .B(n15406), .ZN(n15460) );
  XNOR2_X1 U17072 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15409), .ZN(n15467) );
  XNOR2_X1 U17073 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15410), .ZN(n15411) );
  NOR2_X2 U17074 ( .A1(n15412), .A2(n15411), .ZN(n15434) );
  INV_X1 U17075 ( .A(n15434), .ZN(n15435) );
  INV_X1 U17076 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15714) );
  AOI21_X1 U17077 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15413) );
  OAI21_X1 U17078 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15413), 
        .ZN(U28) );
  AOI21_X1 U17079 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15414) );
  OAI21_X1 U17080 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15414), 
        .ZN(U29) );
  AOI21_X1 U17081 ( .B1(n15417), .B2(n15416), .A(n15415), .ZN(n15418) );
  XOR2_X1 U17082 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n15418), .Z(SUB_1596_U61) );
  AOI21_X1 U17083 ( .B1(n15421), .B2(n15420), .A(n15419), .ZN(SUB_1596_U57) );
  AOI21_X1 U17084 ( .B1(n15424), .B2(n15423), .A(n15422), .ZN(SUB_1596_U55) );
  OAI21_X1 U17085 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15428) );
  XOR2_X1 U17086 ( .A(n15428), .B(n15397), .Z(SUB_1596_U54) );
  OAI21_X1 U17087 ( .B1(n15431), .B2(n15430), .A(n15429), .ZN(n15432) );
  XNOR2_X1 U17088 ( .A(n15432), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI222_X1 U17089 ( .A1(n15714), .A2(n15436), .B1(n15714), .B2(n15435), .C1(
        n15434), .C2(n15433), .ZN(SUB_1596_U63) );
  NAND2_X1 U17090 ( .A1(n15438), .A2(n15437), .ZN(n15439) );
  OAI21_X1 U17091 ( .B1(n15440), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15439), 
        .ZN(n15444) );
  XNOR2_X1 U17092 ( .A(n8040), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15443) );
  OAI222_X1 U17093 ( .A1(n15449), .A2(n15448), .B1(n15449), .B2(n15447), .C1(
        n15446), .C2(n15445), .ZN(SUB_1596_U69) );
  OAI21_X1 U17094 ( .B1(n15452), .B2(n15451), .A(n15450), .ZN(n15453) );
  XOR2_X1 U17095 ( .A(n15453), .B(n7864), .Z(SUB_1596_U68) );
  OAI21_X1 U17096 ( .B1(n15456), .B2(n15455), .A(n15454), .ZN(n15457) );
  XNOR2_X1 U17097 ( .A(n15457), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U17098 ( .B1(n15460), .B2(n15459), .A(n15458), .ZN(n15461) );
  XNOR2_X1 U17099 ( .A(n15461), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U17100 ( .B1(n15463), .B2(n15462), .A(n6531), .ZN(n15464) );
  XOR2_X1 U17101 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15464), .Z(SUB_1596_U65)
         );
  OAI21_X1 U17102 ( .B1(n15467), .B2(n15466), .A(n15465), .ZN(n15468) );
  XNOR2_X1 U17103 ( .A(n15468), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U17104 ( .A(n15469), .ZN(n15472) );
  OAI21_X1 U17105 ( .B1(n15472), .B2(n15471), .A(n15470), .ZN(n15480) );
  XNOR2_X1 U17106 ( .A(n15474), .B(n15473), .ZN(n15477) );
  AOI222_X1 U17107 ( .A1(n15480), .A2(n15479), .B1(n15478), .B2(n15477), .C1(
        n15476), .C2(n15475), .ZN(n15482) );
  OAI211_X1 U17108 ( .C1(n15484), .C2(n15483), .A(n15482), .B(n15481), .ZN(
        P1_U3258) );
  XNOR2_X1 U17109 ( .A(n15485), .B(n15488), .ZN(n15492) );
  NAND2_X1 U17110 ( .A1(n15487), .A2(n15486), .ZN(n15489) );
  XNOR2_X1 U17111 ( .A(n15489), .B(n15488), .ZN(n15496) );
  NOR2_X1 U17112 ( .A1(n15496), .A2(n15589), .ZN(n15490) );
  AOI211_X1 U17113 ( .C1(n15604), .C2(n15492), .A(n15491), .B(n15490), .ZN(
        n15581) );
  INV_X1 U17114 ( .A(n15493), .ZN(n15494) );
  AOI222_X1 U17115 ( .A1(n15495), .A2(n15515), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n15534), .C1(n15494), .C2(n15531), .ZN(n15503) );
  INV_X1 U17116 ( .A(n15496), .ZN(n15584) );
  INV_X1 U17117 ( .A(n15497), .ZN(n15520) );
  OAI211_X1 U17118 ( .C1(n7629), .C2(n15580), .A(n15500), .B(n15499), .ZN(
        n15578) );
  INV_X1 U17119 ( .A(n15578), .ZN(n15501) );
  AOI22_X1 U17120 ( .A1(n15584), .A2(n15520), .B1(n15519), .B2(n15501), .ZN(
        n15502) );
  OAI211_X1 U17121 ( .C1(n15534), .C2(n15581), .A(n15503), .B(n15502), .ZN(
        P1_U3288) );
  OAI21_X1 U17122 ( .B1(n15504), .B2(n15507), .A(n11960), .ZN(n15510) );
  INV_X1 U17123 ( .A(n15505), .ZN(n15509) );
  XNOR2_X1 U17124 ( .A(n15507), .B(n15506), .ZN(n15567) );
  NOR2_X1 U17125 ( .A1(n15567), .A2(n15589), .ZN(n15508) );
  AOI211_X1 U17126 ( .C1(n15604), .C2(n15510), .A(n15509), .B(n15508), .ZN(
        n15566) );
  OAI22_X1 U17127 ( .A1(n15513), .A2(n15512), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15511), .ZN(n15514) );
  AOI21_X1 U17128 ( .B1(n15515), .B2(n15564), .A(n15514), .ZN(n15523) );
  INV_X1 U17129 ( .A(n15567), .ZN(n15521) );
  AOI211_X1 U17130 ( .C1(n15564), .C2(n15518), .A(n15517), .B(n15516), .ZN(
        n15563) );
  AOI22_X1 U17131 ( .A1(n15521), .A2(n15520), .B1(n15563), .B2(n15519), .ZN(
        n15522) );
  OAI211_X1 U17132 ( .C1(n15534), .C2(n15566), .A(n15523), .B(n15522), .ZN(
        P1_U3290) );
  NOR2_X1 U17133 ( .A1(n15525), .A2(n15524), .ZN(n15543) );
  NAND2_X1 U17134 ( .A1(n12652), .A2(n15526), .ZN(n15527) );
  AOI21_X1 U17135 ( .B1(n15543), .B2(n15527), .A(n15544), .ZN(n15533) );
  AOI21_X1 U17136 ( .B1(n15529), .B2(n15528), .A(n15542), .ZN(n15530) );
  AOI21_X1 U17137 ( .B1(n15531), .B2(P1_REG3_REG_0__SCAN_IN), .A(n15530), .ZN(
        n15532) );
  OAI221_X1 U17138 ( .B1(n15534), .B2(n15533), .C1(n15513), .C2(n10879), .A(
        n15532), .ZN(P1_U3293) );
  INV_X1 U17139 ( .A(n15541), .ZN(n15540) );
  NOR2_X1 U17140 ( .A1(n15540), .A2(n15535), .ZN(P1_U3294) );
  NOR2_X1 U17141 ( .A1(n15540), .A2(n15536), .ZN(P1_U3295) );
  AND2_X1 U17142 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15541), .ZN(P1_U3296) );
  AND2_X1 U17143 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15541), .ZN(P1_U3297) );
  AND2_X1 U17144 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15541), .ZN(P1_U3298) );
  AND2_X1 U17145 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15541), .ZN(P1_U3299) );
  AND2_X1 U17146 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15541), .ZN(P1_U3300) );
  AND2_X1 U17147 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15541), .ZN(P1_U3301) );
  AND2_X1 U17148 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15541), .ZN(P1_U3302) );
  AND2_X1 U17149 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15541), .ZN(P1_U3303) );
  NOR2_X1 U17150 ( .A1(n15540), .A2(n15537), .ZN(P1_U3304) );
  AND2_X1 U17151 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15541), .ZN(P1_U3305) );
  AND2_X1 U17152 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15541), .ZN(P1_U3306) );
  AND2_X1 U17153 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15541), .ZN(P1_U3307) );
  AND2_X1 U17154 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15541), .ZN(P1_U3308) );
  AND2_X1 U17155 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15541), .ZN(P1_U3309) );
  AND2_X1 U17156 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15541), .ZN(P1_U3310) );
  AND2_X1 U17157 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15541), .ZN(P1_U3311) );
  NOR2_X1 U17158 ( .A1(n15540), .A2(n15538), .ZN(P1_U3312) );
  AND2_X1 U17159 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15541), .ZN(P1_U3313) );
  AND2_X1 U17160 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15541), .ZN(P1_U3314) );
  NOR2_X1 U17161 ( .A1(n15540), .A2(n15539), .ZN(P1_U3315) );
  AND2_X1 U17162 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15541), .ZN(P1_U3316) );
  AND2_X1 U17163 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15541), .ZN(P1_U3317) );
  AND2_X1 U17164 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15541), .ZN(P1_U3318) );
  AND2_X1 U17165 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15541), .ZN(P1_U3319) );
  AND2_X1 U17166 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15541), .ZN(P1_U3320) );
  AND2_X1 U17167 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15541), .ZN(P1_U3321) );
  AND2_X1 U17168 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15541), .ZN(P1_U3322) );
  AND2_X1 U17169 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15541), .ZN(P1_U3323) );
  AOI21_X1 U17170 ( .B1(n15601), .B2(n15558), .A(n15542), .ZN(n15545) );
  NOR3_X1 U17171 ( .A1(n15545), .A2(n15544), .A3(n15543), .ZN(n15607) );
  INV_X1 U17172 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U17173 ( .A1(n15606), .A2(n15607), .B1(n15546), .B2(n15605), .ZN(
        P1_U3459) );
  INV_X1 U17174 ( .A(n15588), .ZN(n15585) );
  INV_X1 U17175 ( .A(n15547), .ZN(n15552) );
  OAI21_X1 U17176 ( .B1(n15549), .B2(n15579), .A(n15548), .ZN(n15551) );
  AOI211_X1 U17177 ( .C1(n15585), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        n15608) );
  AOI22_X1 U17178 ( .A1(n15606), .A2(n15608), .B1(n6891), .B2(n15605), .ZN(
        P1_U3462) );
  INV_X1 U17179 ( .A(n15589), .ZN(n15561) );
  AOI211_X1 U17180 ( .C1(n15598), .C2(n10303), .A(n15554), .B(n15553), .ZN(
        n15556) );
  NAND2_X1 U17181 ( .A1(n15560), .A2(n15585), .ZN(n15555) );
  OAI211_X1 U17182 ( .C1(n15558), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        n15559) );
  AOI21_X1 U17183 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(n15609) );
  INV_X1 U17184 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U17185 ( .A1(n15606), .A2(n15609), .B1(n15562), .B2(n15605), .ZN(
        P1_U3465) );
  AOI21_X1 U17186 ( .B1(n15598), .B2(n15564), .A(n15563), .ZN(n15565) );
  OAI211_X1 U17187 ( .C1(n15588), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        n15568) );
  INV_X1 U17188 ( .A(n15568), .ZN(n15610) );
  AOI22_X1 U17189 ( .A1(n15606), .A2(n15610), .B1(n8268), .B2(n15605), .ZN(
        P1_U3468) );
  NAND2_X1 U17190 ( .A1(n15569), .A2(n15598), .ZN(n15570) );
  AND2_X1 U17191 ( .A1(n15571), .A2(n15570), .ZN(n15575) );
  NAND2_X1 U17192 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  AND3_X1 U17193 ( .A1(n15576), .A2(n15575), .A3(n15574), .ZN(n15611) );
  INV_X1 U17194 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U17195 ( .A1(n15606), .A2(n15611), .B1(n15577), .B2(n15605), .ZN(
        P1_U3471) );
  OAI21_X1 U17196 ( .B1(n15580), .B2(n15579), .A(n15578), .ZN(n15583) );
  INV_X1 U17197 ( .A(n15581), .ZN(n15582) );
  AOI211_X1 U17198 ( .C1(n15585), .C2(n15584), .A(n15583), .B(n15582), .ZN(
        n15612) );
  INV_X1 U17199 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U17200 ( .A1(n15606), .A2(n15612), .B1(n15586), .B2(n15605), .ZN(
        P1_U3474) );
  OAI21_X1 U17201 ( .B1(n15588), .B2(n15590), .A(n15587), .ZN(n15594) );
  NOR2_X1 U17202 ( .A1(n15590), .A2(n15589), .ZN(n15592) );
  NOR4_X1 U17203 ( .A1(n15594), .A2(n15593), .A3(n15592), .A4(n15591), .ZN(
        n15614) );
  AOI22_X1 U17204 ( .A1(n15606), .A2(n15614), .B1(n8344), .B2(n15605), .ZN(
        P1_U3477) );
  AOI211_X1 U17205 ( .C1(n15598), .C2(n15597), .A(n15596), .B(n15595), .ZN(
        n15599) );
  OAI21_X1 U17206 ( .B1(n15601), .B2(n15600), .A(n15599), .ZN(n15602) );
  AOI21_X1 U17207 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15617) );
  AOI22_X1 U17208 ( .A1(n15606), .A2(n15617), .B1(n8367), .B2(n15605), .ZN(
        P1_U3480) );
  AOI22_X1 U17209 ( .A1(n15618), .A2(n15607), .B1(n8240), .B2(n15615), .ZN(
        P1_U3528) );
  AOI22_X1 U17210 ( .A1(n15618), .A2(n15608), .B1(n10839), .B2(n15615), .ZN(
        P1_U3529) );
  AOI22_X1 U17211 ( .A1(n15618), .A2(n15609), .B1(n10840), .B2(n15615), .ZN(
        P1_U3530) );
  AOI22_X1 U17212 ( .A1(n15618), .A2(n15610), .B1(n10841), .B2(n15615), .ZN(
        P1_U3531) );
  AOI22_X1 U17213 ( .A1(n15618), .A2(n15611), .B1(n10842), .B2(n15615), .ZN(
        P1_U3532) );
  AOI22_X1 U17214 ( .A1(n15618), .A2(n15612), .B1(n10896), .B2(n15615), .ZN(
        P1_U3533) );
  AOI22_X1 U17215 ( .A1(n15618), .A2(n15614), .B1(n15613), .B2(n15615), .ZN(
        P1_U3534) );
  INV_X1 U17216 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U17217 ( .A1(n15618), .A2(n15617), .B1(n15616), .B2(n15615), .ZN(
        P1_U3535) );
  NOR2_X1 U17218 ( .A1(n15634), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17219 ( .A1(n15696), .A2(n15619), .ZN(n15626) );
  INV_X1 U17220 ( .A(n15620), .ZN(n15623) );
  INV_X1 U17221 ( .A(n15621), .ZN(n15622) );
  AOI211_X1 U17222 ( .C1(n15624), .C2(n15623), .A(n15622), .B(n15701), .ZN(
        n15625) );
  AOI211_X1 U17223 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3088), .A(n15626), 
        .B(n15625), .ZN(n15631) );
  OAI211_X1 U17224 ( .C1(n15629), .C2(n15628), .A(n15708), .B(n15627), .ZN(
        n15630) );
  OAI211_X1 U17225 ( .C1(n15715), .C2(n15632), .A(n15631), .B(n15630), .ZN(
        P2_U3215) );
  AOI22_X1 U17226 ( .A1(n15634), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15646) );
  OAI211_X1 U17227 ( .C1(n15637), .C2(n15636), .A(n15690), .B(n15635), .ZN(
        n15638) );
  OAI21_X1 U17228 ( .B1(n15696), .B2(n15639), .A(n15638), .ZN(n15640) );
  INV_X1 U17229 ( .A(n15640), .ZN(n15645) );
  OAI211_X1 U17230 ( .C1(n15643), .C2(n15642), .A(n15708), .B(n15641), .ZN(
        n15644) );
  NAND3_X1 U17231 ( .A1(n15646), .A2(n15645), .A3(n15644), .ZN(P2_U3216) );
  INV_X1 U17232 ( .A(n15647), .ZN(n15653) );
  OAI211_X1 U17233 ( .C1(n15650), .C2(n15649), .A(n15690), .B(n15648), .ZN(
        n15651) );
  INV_X1 U17234 ( .A(n15651), .ZN(n15652) );
  AOI211_X1 U17235 ( .C1(n15707), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        n15659) );
  OAI211_X1 U17236 ( .C1(n15657), .C2(n15656), .A(n15708), .B(n15655), .ZN(
        n15658) );
  OAI211_X1 U17237 ( .C1(n15715), .C2(n15660), .A(n15659), .B(n15658), .ZN(
        P2_U3218) );
  OAI21_X1 U17238 ( .B1(n15663), .B2(n15662), .A(n15661), .ZN(n15664) );
  NAND2_X1 U17239 ( .A1(n15708), .A2(n15664), .ZN(n15674) );
  INV_X1 U17240 ( .A(n15665), .ZN(n15672) );
  INV_X1 U17241 ( .A(n15666), .ZN(n15669) );
  INV_X1 U17242 ( .A(n15667), .ZN(n15668) );
  AOI21_X1 U17243 ( .B1(n15670), .B2(n15669), .A(n15668), .ZN(n15671) );
  OAI21_X1 U17244 ( .B1(n15672), .B2(n15671), .A(n15690), .ZN(n15673) );
  OAI211_X1 U17245 ( .C1(n15696), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n15676) );
  INV_X1 U17246 ( .A(n15676), .ZN(n15678) );
  OAI211_X1 U17247 ( .C1(n15397), .C2(n15715), .A(n15678), .B(n15677), .ZN(
        P2_U3223) );
  INV_X1 U17248 ( .A(n15679), .ZN(n15681) );
  NAND3_X1 U17249 ( .A1(n15682), .A2(n15681), .A3(n15680), .ZN(n15683) );
  NAND2_X1 U17250 ( .A1(n15684), .A2(n15683), .ZN(n15685) );
  NAND2_X1 U17251 ( .A1(n15685), .A2(n15708), .ZN(n15694) );
  INV_X1 U17252 ( .A(n15686), .ZN(n15692) );
  AOI21_X1 U17253 ( .B1(n15689), .B2(n15688), .A(n15687), .ZN(n15691) );
  OAI21_X1 U17254 ( .B1(n15692), .B2(n15691), .A(n15690), .ZN(n15693) );
  OAI211_X1 U17255 ( .C1(n15696), .C2(n15695), .A(n15694), .B(n15693), .ZN(
        n15697) );
  INV_X1 U17256 ( .A(n15697), .ZN(n15699) );
  OAI211_X1 U17257 ( .C1(n7864), .C2(n15715), .A(n15699), .B(n15698), .ZN(
        P2_U3226) );
  AOI211_X1 U17258 ( .C1(n15703), .C2(n15702), .A(n15701), .B(n15700), .ZN(
        n15704) );
  AOI211_X1 U17259 ( .C1(n15707), .C2(n15706), .A(n15705), .B(n15704), .ZN(
        n15713) );
  OAI211_X1 U17260 ( .C1(n15711), .C2(n15710), .A(n15709), .B(n15708), .ZN(
        n15712) );
  OAI211_X1 U17261 ( .C1(n15715), .C2(n15714), .A(n15713), .B(n15712), .ZN(
        P2_U3231) );
  INV_X1 U17262 ( .A(n15722), .ZN(n15724) );
  AND2_X1 U17263 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15719), .ZN(P2_U3266) );
  AND2_X1 U17264 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15719), .ZN(P2_U3267) );
  AND2_X1 U17265 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15719), .ZN(P2_U3268) );
  AND2_X1 U17266 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15719), .ZN(P2_U3269) );
  AND2_X1 U17267 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15719), .ZN(P2_U3270) );
  AND2_X1 U17268 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15719), .ZN(P2_U3271) );
  AND2_X1 U17269 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15719), .ZN(P2_U3272) );
  AND2_X1 U17270 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15719), .ZN(P2_U3273) );
  AND2_X1 U17271 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15719), .ZN(P2_U3274) );
  AND2_X1 U17272 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15719), .ZN(P2_U3275) );
  AND2_X1 U17273 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15719), .ZN(P2_U3276) );
  AND2_X1 U17274 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15719), .ZN(P2_U3277) );
  AND2_X1 U17275 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15719), .ZN(P2_U3278) );
  AND2_X1 U17276 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15719), .ZN(P2_U3279) );
  AND2_X1 U17277 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15719), .ZN(P2_U3280) );
  AND2_X1 U17278 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15719), .ZN(P2_U3281) );
  AND2_X1 U17279 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15719), .ZN(P2_U3282) );
  AND2_X1 U17280 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15719), .ZN(P2_U3283) );
  NOR2_X1 U17281 ( .A1(n15718), .A2(n15717), .ZN(P2_U3284) );
  AND2_X1 U17282 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15719), .ZN(P2_U3285) );
  AND2_X1 U17283 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15719), .ZN(P2_U3286) );
  AND2_X1 U17284 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15719), .ZN(P2_U3287) );
  AND2_X1 U17285 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15719), .ZN(P2_U3288) );
  AND2_X1 U17286 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15719), .ZN(P2_U3289) );
  AND2_X1 U17287 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15719), .ZN(P2_U3290) );
  AND2_X1 U17288 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15719), .ZN(P2_U3291) );
  AND2_X1 U17289 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15719), .ZN(P2_U3292) );
  AND2_X1 U17290 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15719), .ZN(P2_U3293) );
  AND2_X1 U17291 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15719), .ZN(P2_U3294) );
  AND2_X1 U17292 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15719), .ZN(P2_U3295) );
  AOI22_X1 U17293 ( .A1(n15722), .A2(n15721), .B1(n15720), .B2(n15724), .ZN(
        P2_U3416) );
  AOI21_X1 U17294 ( .B1(n15725), .B2(n15724), .A(n15723), .ZN(P2_U3417) );
  NOR3_X1 U17295 ( .A1(n15727), .A2(n15726), .A3(n12534), .ZN(n15730) );
  INV_X1 U17296 ( .A(n15728), .ZN(n15729) );
  AOI211_X1 U17297 ( .C1(n15731), .C2(n6951), .A(n15730), .B(n15729), .ZN(
        n15769) );
  INV_X1 U17298 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U17299 ( .A1(n15767), .A2(n15769), .B1(n15732), .B2(n15765), .ZN(
        P2_U3430) );
  OAI211_X1 U17300 ( .C1(n15736), .C2(n12373), .A(n15735), .B(n15734), .ZN(
        n15737) );
  INV_X1 U17301 ( .A(n15737), .ZN(n15770) );
  AOI22_X1 U17302 ( .A1(n15767), .A2(n15770), .B1(n8892), .B2(n15765), .ZN(
        P2_U3433) );
  AOI22_X1 U17303 ( .A1(n15767), .A2(n15739), .B1(n15738), .B2(n15765), .ZN(
        P2_U3436) );
  AOI211_X1 U17304 ( .C1(n15750), .C2(n15742), .A(n15741), .B(n15740), .ZN(
        n15744) );
  OAI211_X1 U17305 ( .C1(n15748), .C2(n15745), .A(n15744), .B(n15743), .ZN(
        n15746) );
  INV_X1 U17306 ( .A(n15746), .ZN(n15772) );
  INV_X1 U17307 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U17308 ( .A1(n15767), .A2(n15772), .B1(n15747), .B2(n15765), .ZN(
        P2_U3439) );
  NOR2_X1 U17309 ( .A1(n15749), .A2(n15748), .ZN(n15754) );
  INV_X1 U17310 ( .A(n15750), .ZN(n15758) );
  OAI21_X1 U17311 ( .B1(n7888), .B2(n15758), .A(n15751), .ZN(n15752) );
  NOR3_X1 U17312 ( .A1(n15754), .A2(n15753), .A3(n15752), .ZN(n15774) );
  AOI22_X1 U17313 ( .A1(n15767), .A2(n15774), .B1(n15755), .B2(n15765), .ZN(
        P2_U3442) );
  INV_X1 U17314 ( .A(n15756), .ZN(n15763) );
  OAI21_X1 U17315 ( .B1(n15759), .B2(n15758), .A(n15757), .ZN(n15762) );
  INV_X1 U17316 ( .A(n15760), .ZN(n15761) );
  AOI211_X1 U17317 ( .C1(n15764), .C2(n15763), .A(n15762), .B(n15761), .ZN(
        n15777) );
  INV_X1 U17318 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U17319 ( .A1(n15767), .A2(n15777), .B1(n15766), .B2(n15765), .ZN(
        P2_U3445) );
  INV_X1 U17320 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U17321 ( .A1(n15778), .A2(n15769), .B1(n15768), .B2(n15775), .ZN(
        P2_U3499) );
  AOI22_X1 U17322 ( .A1(n15778), .A2(n15770), .B1(n7798), .B2(n15775), .ZN(
        P2_U3500) );
  INV_X1 U17323 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15771) );
  AOI22_X1 U17324 ( .A1(n15778), .A2(n15772), .B1(n15771), .B2(n15775), .ZN(
        P2_U3502) );
  INV_X1 U17325 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15773) );
  AOI22_X1 U17326 ( .A1(n15778), .A2(n15774), .B1(n15773), .B2(n15775), .ZN(
        P2_U3503) );
  INV_X1 U17327 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U17328 ( .A1(n15778), .A2(n15777), .B1(n15776), .B2(n15775), .ZN(
        P2_U3504) );
  NOR2_X1 U17329 ( .A1(P3_U3897), .A2(n15779), .ZN(P3_U3150) );
  XNOR2_X1 U17330 ( .A(n15780), .B(n15781), .ZN(n15788) );
  OAI21_X1 U17331 ( .B1(n15782), .B2(n15781), .A(n11435), .ZN(n15824) );
  OAI22_X1 U17332 ( .A1(n6837), .A2(n15785), .B1(n15784), .B2(n15783), .ZN(
        n15786) );
  AOI21_X1 U17333 ( .B1(n15824), .B2(n15843), .A(n15786), .ZN(n15787) );
  OAI21_X1 U17334 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n15822) );
  INV_X1 U17335 ( .A(n15824), .ZN(n15792) );
  NOR2_X1 U17336 ( .A1(n15790), .A2(n15806), .ZN(n15823) );
  INV_X1 U17337 ( .A(n15823), .ZN(n15791) );
  OAI22_X1 U17338 ( .A1(n15792), .A2(n15810), .B1(n15809), .B2(n15791), .ZN(
        n15793) );
  AOI211_X1 U17339 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15812), .A(n15822), .B(
        n15793), .ZN(n15794) );
  AOI22_X1 U17340 ( .A1(n15816), .A2(n10673), .B1(n15794), .B2(n15813), .ZN(
        P3_U3231) );
  XNOR2_X1 U17341 ( .A(n10442), .B(n15795), .ZN(n15817) );
  AOI22_X1 U17342 ( .A1(n15799), .A2(n15798), .B1(n15797), .B2(n15796), .ZN(
        n15804) );
  XNOR2_X1 U17343 ( .A(n10442), .B(n15800), .ZN(n15802) );
  NAND2_X1 U17344 ( .A1(n15802), .A2(n15801), .ZN(n15803) );
  OAI211_X1 U17345 ( .C1(n15817), .C2(n15805), .A(n15804), .B(n15803), .ZN(
        n15818) );
  NOR2_X1 U17346 ( .A1(n15807), .A2(n15806), .ZN(n15819) );
  INV_X1 U17347 ( .A(n15819), .ZN(n15808) );
  OAI22_X1 U17348 ( .A1(n15817), .A2(n15810), .B1(n15809), .B2(n15808), .ZN(
        n15811) );
  AOI211_X1 U17349 ( .C1(P3_REG3_REG_1__SCAN_IN), .C2(n15812), .A(n15818), .B(
        n15811), .ZN(n15814) );
  AOI22_X1 U17350 ( .A1(n15816), .A2(n15815), .B1(n15814), .B2(n15813), .ZN(
        P3_U3232) );
  INV_X1 U17351 ( .A(n15817), .ZN(n15820) );
  AOI211_X1 U17352 ( .C1(n15856), .C2(n15820), .A(n15819), .B(n15818), .ZN(
        n15862) );
  AOI22_X1 U17353 ( .A1(n15860), .A2(n15862), .B1(n15821), .B2(n15858), .ZN(
        P3_U3393) );
  AOI211_X1 U17354 ( .C1(n15856), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        n15863) );
  INV_X1 U17355 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U17356 ( .A1(n15860), .A2(n15863), .B1(n15825), .B2(n15858), .ZN(
        P3_U3396) );
  INV_X1 U17357 ( .A(n15826), .ZN(n15827) );
  AOI211_X1 U17358 ( .C1(n15829), .C2(n15856), .A(n15828), .B(n15827), .ZN(
        n15865) );
  INV_X1 U17359 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15830) );
  AOI22_X1 U17360 ( .A1(n15860), .A2(n15865), .B1(n15830), .B2(n15858), .ZN(
        P3_U3399) );
  INV_X1 U17361 ( .A(n15831), .ZN(n15834) );
  AOI211_X1 U17362 ( .C1(n15834), .C2(n15856), .A(n15833), .B(n15832), .ZN(
        n15866) );
  INV_X1 U17363 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15835) );
  AOI22_X1 U17364 ( .A1(n15860), .A2(n15866), .B1(n15835), .B2(n15858), .ZN(
        P3_U3402) );
  INV_X1 U17365 ( .A(n15840), .ZN(n15844) );
  NAND2_X1 U17366 ( .A1(n15837), .A2(n15836), .ZN(n15838) );
  OAI211_X1 U17367 ( .C1(n15841), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        n15842) );
  AOI21_X1 U17368 ( .B1(n15844), .B2(n15843), .A(n15842), .ZN(n15868) );
  AOI22_X1 U17369 ( .A1(n15860), .A2(n15868), .B1(n15845), .B2(n15858), .ZN(
        P3_U3408) );
  INV_X1 U17370 ( .A(n15846), .ZN(n15850) );
  INV_X1 U17371 ( .A(n15847), .ZN(n15848) );
  AOI211_X1 U17372 ( .C1(n15851), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15870) );
  INV_X1 U17373 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15852) );
  AOI22_X1 U17374 ( .A1(n15860), .A2(n15870), .B1(n15852), .B2(n15858), .ZN(
        P3_U3411) );
  INV_X1 U17375 ( .A(n15853), .ZN(n15854) );
  AOI211_X1 U17376 ( .C1(n15857), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        n15872) );
  INV_X1 U17377 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15859) );
  AOI22_X1 U17378 ( .A1(n15860), .A2(n15872), .B1(n15859), .B2(n15858), .ZN(
        P3_U3414) );
  AOI22_X1 U17379 ( .A1(n15873), .A2(n15862), .B1(n15861), .B2(n10255), .ZN(
        P3_U3460) );
  AOI22_X1 U17380 ( .A1(n15873), .A2(n15863), .B1(n9487), .B2(n10255), .ZN(
        P3_U3461) );
  AOI22_X1 U17381 ( .A1(n15873), .A2(n15865), .B1(n15864), .B2(n10255), .ZN(
        P3_U3462) );
  AOI22_X1 U17382 ( .A1(n15873), .A2(n15866), .B1(n9505), .B2(n10255), .ZN(
        P3_U3463) );
  AOI22_X1 U17383 ( .A1(n15873), .A2(n15868), .B1(n15867), .B2(n10255), .ZN(
        P3_U3465) );
  AOI22_X1 U17384 ( .A1(n15873), .A2(n15870), .B1(n15869), .B2(n10255), .ZN(
        P3_U3466) );
  AOI22_X1 U17385 ( .A1(n15873), .A2(n15872), .B1(n15871), .B2(n10255), .ZN(
        P3_U3467) );
  OAI21_X1 U17386 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(SUB_1596_U58) );
  XOR2_X1 U17387 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15879), .Z(SUB_1596_U53) );
  OAI21_X1 U17388 ( .B1(n15884), .B2(n15883), .A(n15882), .ZN(n15885) );
  XNOR2_X1 U17389 ( .A(n15885), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17390 ( .B1(n15888), .B2(n15887), .A(n15886), .ZN(SUB_1596_U5) );
  AND2_X1 U12058 ( .A1(n9440), .A2(n9908), .ZN(n9878) );
  AOI21_X1 U9901 ( .B1(n13960), .B2(n7720), .A(n6581), .ZN(n11327) );
  OR2_X1 U7178 ( .A1(n13878), .A2(n6781), .ZN(n6780) );
  CLKBUF_X1 U7434 ( .A(n9014), .Z(n9305) );
endmodule

