

module b22_C_AntiSAT_k_128_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6472, n6473, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n15018;

  AOI21_X1 U7220 ( .B1(n6915), .B2(n12879), .A(n8345), .ZN(n12906) );
  INV_X4 U7221 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7222 ( .A(P3_STATE_REG_SCAN_IN), .ZN(n15018) );
  XNOR2_X1 U7223 ( .A(n13946), .B(n13531), .ZN(n13939) );
  OR2_X1 U7224 ( .A1(n8329), .A2(n6895), .ZN(n6894) );
  OAI21_X1 U7225 ( .B1(n10737), .B2(n8324), .A(n8323), .ZN(n9890) );
  CLKBUF_X2 U7226 ( .A(n11844), .Z(n6828) );
  INV_X4 U7227 ( .A(n11743), .ZN(n11762) );
  INV_X1 U7228 ( .A(n13574), .ZN(n13594) );
  INV_X1 U7229 ( .A(n9795), .ZN(n11209) );
  INV_X1 U7230 ( .A(n9795), .ZN(n13579) );
  INV_X2 U7231 ( .A(n6486), .ZN(n8237) );
  NAND2_X2 U7233 ( .A1(n12971), .A2(n12679), .ZN(n6488) );
  CLKBUF_X2 U7234 ( .A(n7514), .Z(n8190) );
  INV_X2 U7235 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n11301) );
  AND2_X1 U7236 ( .A1(n7515), .A2(n7314), .ZN(n6900) );
  INV_X1 U7237 ( .A(n15018), .ZN(n6472) );
  INV_X1 U7238 ( .A(n6472), .ZN(n6473) );
  INV_X1 U7239 ( .A(n6472), .ZN(P3_U3151) );
  CLKBUF_X3 U7240 ( .A(n6478), .Z(n6486) );
  INV_X1 U7241 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9565) );
  INV_X1 U7242 ( .A(n11613), .ZN(n12310) );
  OAI21_X1 U7244 ( .B1(n12805), .B2(n7217), .A(n7214), .ZN(n12753) );
  OAI21_X1 U7245 ( .B1(n10650), .B2(n7292), .A(n6624), .ZN(n6748) );
  NAND2_X1 U7246 ( .A1(n7606), .A2(n7605), .ZN(n8267) );
  INV_X1 U7247 ( .A(n13311), .ZN(n13064) );
  INV_X1 U7248 ( .A(n13062), .ZN(n13313) );
  INV_X1 U7249 ( .A(n8564), .ZN(n8563) );
  CLKBUF_X3 U7250 ( .A(n10155), .Z(n11454) );
  INV_X1 U7251 ( .A(n12023), .ZN(n12141) );
  NAND2_X1 U7252 ( .A1(n11671), .A2(n6619), .ZN(n12236) );
  NAND2_X2 U7253 ( .A1(n12424), .A2(n9016), .ZN(n11348) );
  INV_X1 U7254 ( .A(n7626), .ZN(n8187) );
  OAI21_X1 U7255 ( .B1(n10678), .B2(n8400), .A(n8399), .ZN(n10650) );
  AND2_X1 U7256 ( .A1(n7868), .A2(n7867), .ZN(n14270) );
  INV_X1 U7258 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U7259 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  AND2_X1 U7260 ( .A1(n6923), .A2(n6922), .ZN(n9912) );
  INV_X1 U7261 ( .A(n9739), .ZN(n11138) );
  INV_X1 U7262 ( .A(n14108), .ZN(n13946) );
  AND2_X1 U7263 ( .A1(n10556), .A2(n13587), .ZN(n13433) );
  INV_X1 U7264 ( .A(n12191), .ZN(n12156) );
  INV_X1 U7265 ( .A(n12178), .ZN(n12206) );
  XNOR2_X1 U7266 ( .A(n11720), .B(n6517), .ZN(n11772) );
  OAI21_X1 U7267 ( .B1(n12907), .B2(n14720), .A(n12905), .ZN(n7047) );
  NAND2_X1 U7268 ( .A1(n6900), .A2(n7553), .ZN(n7556) );
  NAND2_X1 U7269 ( .A1(n11104), .A2(n11103), .ZN(n14116) );
  MUX2_X1 U7270 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14174), .S(n11132), .Z(n14032)
         );
  NAND2_X1 U7271 ( .A1(n7178), .A2(n8757), .ZN(n8579) );
  OAI21_X1 U7272 ( .B1(n10090), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U7273 ( .A1(n7425), .A2(n7556), .ZN(n13003) );
  XNOR2_X1 U7274 ( .A(n6849), .B(n8625), .ZN(n13990) );
  INV_X2 U7275 ( .A(n14228), .ZN(n14908) );
  NAND4_X2 U7276 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n12023) );
  INV_X4 U7277 ( .A(n13063), .ZN(n9725) );
  INV_X1 U7278 ( .A(n7626), .ZN(n6475) );
  NAND2_X2 U7279 ( .A1(n7627), .A2(n7672), .ZN(n7626) );
  NAND2_X2 U7280 ( .A1(n10161), .A2(n11625), .ZN(n10360) );
  OAI222_X1 U7281 ( .A1(P3_U3151), .A2(n8907), .B1(n12423), .B2(n12415), .C1(
        n12414), .C2(n14186), .ZN(P3_U3265) );
  XNOR2_X1 U7282 ( .A(n9095), .B(n9077), .ZN(n12457) );
  INV_X2 U7283 ( .A(n13464), .ZN(n14475) );
  OAI21_X2 U7284 ( .B1(n7328), .B2(n7660), .A(n7326), .ZN(n7697) );
  AOI21_X2 U7286 ( .B1(n10974), .B2(n13624), .A(n6805), .ZN(n10975) );
  OAI21_X2 U7287 ( .B1(n10859), .B2(n13622), .A(n10858), .ZN(n10974) );
  XNOR2_X2 U7288 ( .A(n7984), .B(SI_18_), .ZN(n7983) );
  OR2_X2 U7289 ( .A1(n12457), .A2(n9076), .ZN(n9097) );
  INV_X4 U7290 ( .A(n7528), .ZN(n13022) );
  AOI21_X2 U7291 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n8433), .A(n8432), .ZN(
        n8502) );
  AOI21_X2 U7292 ( .B1(n9975), .B2(n13611), .A(n9974), .ZN(n14393) );
  OAI21_X2 U7293 ( .B1(n12864), .B2(n7232), .A(n7233), .ZN(n12838) );
  OAI222_X1 U7294 ( .A1(n6473), .A2(n12424), .B1(n12423), .B2(n12422), .C1(
        n12421), .C2(n14186), .ZN(P3_U3267) );
  XNOR2_X2 U7295 ( .A(n9011), .B(n9010), .ZN(n12424) );
  NAND2_X1 U7296 ( .A1(n11348), .A2(n6484), .ZN(n10155) );
  XNOR2_X2 U7297 ( .A(n7837), .B(n7836), .ZN(n10573) );
  XNOR2_X2 U7298 ( .A(n8779), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9513) );
  NOR4_X2 U7299 ( .A1(n13634), .A2(n13633), .A3(n13795), .A4(n13632), .ZN(
        n13635) );
  OAI22_X2 U7300 ( .A1(n11922), .A2(n11923), .B1(n11854), .B2(n12024), .ZN(
        n11996) );
  AOI21_X2 U7301 ( .B1(n11873), .B2(n11853), .A(n11852), .ZN(n11922) );
  XNOR2_X2 U7302 ( .A(n8902), .B(n12407), .ZN(n8907) );
  NAND2_X2 U7303 ( .A1(n12406), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8902) );
  AOI21_X2 U7304 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n8449), .A(n8448), .ZN(
        n8451) );
  NAND2_X1 U7305 ( .A1(n12162), .A2(n11599), .ZN(n12161) );
  INV_X1 U7306 ( .A(n12734), .ZN(n12922) );
  NAND2_X1 U7307 ( .A1(n8397), .A2(n8396), .ZN(n10678) );
  OR2_X1 U7308 ( .A1(n10667), .A2(n6594), .ZN(n8397) );
  NAND2_X1 U7309 ( .A1(n10370), .A2(n7419), .ZN(n10942) );
  OR2_X1 U7310 ( .A1(n10140), .A2(n10141), .ZN(n10138) );
  NAND2_X1 U7311 ( .A1(n13447), .A2(n13446), .ZN(n9471) );
  INV_X1 U7312 ( .A(n11892), .ZN(n11844) );
  NAND2_X1 U7313 ( .A1(n9760), .A2(n11501), .ZN(n14866) );
  INV_X1 U7314 ( .A(n10785), .ZN(n14710) );
  NAND2_X2 U7315 ( .A1(n14847), .A2(n11516), .ZN(n9771) );
  INV_X4 U7316 ( .A(n13600), .ZN(n6477) );
  CLKBUF_X2 U7317 ( .A(n8219), .Z(n8235) );
  NAND2_X4 U7318 ( .A1(n13311), .A2(n14076), .ZN(n13062) );
  INV_X1 U7319 ( .A(n8268), .ZN(n8269) );
  INV_X1 U7320 ( .A(n8271), .ZN(n8378) );
  NAND4_X1 U7321 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n12587)
         );
  INV_X2 U7322 ( .A(n8077), .ZN(n8225) );
  BUF_X2 U7323 ( .A(n7647), .Z(n8194) );
  BUF_X2 U7324 ( .A(n9605), .Z(n11466) );
  INV_X2 U7325 ( .A(n7707), .ZN(n6478) );
  OR2_X1 U7326 ( .A1(n8579), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n8549) );
  NAND3_X1 U7327 ( .A1(n8579), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n8577) );
  AND2_X1 U7328 ( .A1(n7385), .A2(n8621), .ZN(n6694) );
  AND2_X1 U7329 ( .A1(n7512), .A2(n7386), .ZN(n7385) );
  AND2_X1 U7330 ( .A1(n14053), .A2(n14052), .ZN(n14054) );
  OR2_X1 U7331 ( .A1(n14067), .A2(n14066), .ZN(n14143) );
  AOI21_X1 U7332 ( .B1(n11217), .B2(n14411), .A(n11216), .ZN(n14060) );
  OAI21_X1 U7333 ( .B1(n7047), .B2(n6741), .A(n14779), .ZN(n6740) );
  AOI211_X1 U7334 ( .C1(n14231), .C2(n12321), .A(n12135), .B(n12134), .ZN(
        n12136) );
  OAI21_X1 U7335 ( .B1(n12122), .B2(n12386), .A(n12118), .ZN(n11806) );
  AND2_X1 U7336 ( .A1(n7422), .A2(n7421), .ZN(n12328) );
  OAI21_X1 U7337 ( .B1(n8062), .B2(n7486), .A(n7487), .ZN(n8140) );
  AOI21_X1 U7338 ( .B1(n12326), .B2(n14878), .A(n11705), .ZN(n7421) );
  NAND2_X1 U7339 ( .A1(n11185), .A2(n13838), .ZN(n13834) );
  AOI21_X1 U7340 ( .B1(n6521), .B2(n7164), .A(n7160), .ZN(n7159) );
  AOI22_X1 U7341 ( .A1(n11996), .A2(n11997), .B1(n12141), .B2(n11856), .ZN(
        n11891) );
  NAND2_X1 U7342 ( .A1(n7423), .A2(n14896), .ZN(n7422) );
  OAI21_X1 U7343 ( .B1(n11698), .B2(n11697), .A(n11704), .ZN(n7423) );
  AOI21_X1 U7344 ( .B1(n11978), .B2(n12206), .A(n11874), .ZN(n11948) );
  OR2_X1 U7345 ( .A1(n11653), .A2(n7027), .ZN(n7026) );
  AND2_X1 U7346 ( .A1(n8410), .A2(n8265), .ZN(n12701) );
  NAND2_X1 U7347 ( .A1(n12137), .A2(n12148), .ZN(n12143) );
  NAND2_X1 U7348 ( .A1(n12161), .A2(n6813), .ZN(n11428) );
  NAND2_X1 U7349 ( .A1(n11199), .A2(n11198), .ZN(n14058) );
  NAND2_X1 U7350 ( .A1(n11786), .A2(n11789), .ZN(n12137) );
  NAND2_X1 U7351 ( .A1(n12793), .A2(n7097), .ZN(n12730) );
  NAND2_X1 U7352 ( .A1(n12153), .A2(n11681), .ZN(n11786) );
  NAND2_X1 U7353 ( .A1(n8189), .A2(n8188), .ZN(n12915) );
  XNOR2_X1 U7354 ( .A(n8167), .B(n8166), .ZN(n11246) );
  OAI21_X1 U7355 ( .B1(n13918), .B2(n13919), .A(n11227), .ZN(n13906) );
  NAND2_X1 U7356 ( .A1(n11188), .A2(n11187), .ZN(n14063) );
  NAND2_X1 U7357 ( .A1(n7315), .A2(n6555), .ZN(n6916) );
  NAND2_X1 U7358 ( .A1(n7336), .A2(n8146), .ZN(n8167) );
  OR2_X1 U7359 ( .A1(n11611), .A2(n7244), .ZN(n7243) );
  OAI21_X1 U7360 ( .B1(n12838), .B2(n6550), .A(n6733), .ZN(n12805) );
  OR2_X1 U7361 ( .A1(n8185), .A2(n8147), .ZN(n7336) );
  NAND2_X1 U7362 ( .A1(n11168), .A2(n11167), .ZN(n14074) );
  NAND2_X1 U7363 ( .A1(n6671), .A2(n11589), .ZN(n12196) );
  INV_X1 U7364 ( .A(n12766), .ZN(n12931) );
  AND2_X1 U7365 ( .A1(n8095), .A2(n8094), .ZN(n12766) );
  AND2_X2 U7366 ( .A1(n11115), .A2(n11114), .ZN(n14108) );
  NAND2_X1 U7367 ( .A1(n8015), .A2(n8014), .ZN(n12951) );
  NOR2_X1 U7368 ( .A1(n11612), .A2(n7144), .ZN(n7143) );
  NAND2_X1 U7369 ( .A1(n11123), .A2(n11122), .ZN(n13923) );
  NAND2_X1 U7370 ( .A1(n13984), .A2(n11089), .ZN(n13963) );
  OAI21_X1 U7371 ( .B1(n13968), .B2(n11223), .A(n11222), .ZN(n13952) );
  INV_X1 U7372 ( .A(n11601), .ZN(n7144) );
  NAND2_X1 U7373 ( .A1(n6727), .A2(n6725), .ZN(n13968) );
  NAND2_X1 U7374 ( .A1(n7295), .A2(n7294), .ZN(n12843) );
  AND2_X1 U7375 ( .A1(n7989), .A2(n7988), .ZN(n12837) );
  NAND2_X1 U7376 ( .A1(n6894), .A2(n6893), .ZN(n7286) );
  NAND2_X1 U7377 ( .A1(n6954), .A2(n6958), .ZN(n8087) );
  NOR2_X1 U7378 ( .A1(n7288), .A2(n12863), .ZN(n7285) );
  AOI21_X1 U7379 ( .B1(n7983), .B2(n6957), .A(n6955), .ZN(n6954) );
  AOI21_X1 U7380 ( .B1(n10806), .B2(n10805), .A(n10804), .ZN(n10859) );
  AND2_X1 U7381 ( .A1(n11718), .A2(n10683), .ZN(n10656) );
  OAI21_X1 U7382 ( .B1(n10586), .B2(n13619), .A(n6749), .ZN(n10806) );
  NAND2_X1 U7383 ( .A1(n10233), .A2(n10454), .ZN(n10457) );
  AOI21_X1 U7384 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n8439), .A(n8438), .ZN(
        n8510) );
  NAND2_X1 U7385 ( .A1(n7051), .A2(n6969), .ZN(n7345) );
  NAND2_X1 U7386 ( .A1(n7803), .A2(n7802), .ZN(n10750) );
  OR2_X1 U7387 ( .A1(n10031), .A2(n11623), .ZN(n10151) );
  NAND2_X1 U7388 ( .A1(n10512), .A2(n10511), .ZN(n13482) );
  AOI21_X1 U7389 ( .B1(n6929), .B2(n9781), .A(n6928), .ZN(n6927) );
  AOI21_X1 U7390 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n13212), .A(n8437), .ZN(
        n8464) );
  NAND2_X1 U7391 ( .A1(n10189), .A2(n10188), .ZN(n13472) );
  OR2_X1 U7392 ( .A1(n9266), .A2(n9261), .ZN(n7402) );
  AND2_X1 U7393 ( .A1(n9306), .A2(n9260), .ZN(n9266) );
  NAND2_X1 U7394 ( .A1(n9384), .A2(n14902), .ZN(n12017) );
  NAND2_X1 U7395 ( .A1(n7752), .A2(n7751), .ZN(n7772) );
  AND2_X2 U7396 ( .A1(n11524), .A2(n11528), .ZN(n11623) );
  NAND2_X1 U7397 ( .A1(n11521), .A2(n11520), .ZN(n14852) );
  INV_X2 U7398 ( .A(n14419), .ZN(n6479) );
  AND2_X1 U7399 ( .A1(n9771), .A2(n9770), .ZN(n7412) );
  AND3_X1 U7400 ( .A1(n7134), .A2(n7133), .A3(n9448), .ZN(n14888) );
  OAI211_X1 U7401 ( .C1(n11132), .C2(n13691), .A(n9787), .B(n9786), .ZN(n14468) );
  INV_X1 U7402 ( .A(n9483), .ZN(n14448) );
  NAND2_X1 U7403 ( .A1(n7650), .A2(n7387), .ZN(n12586) );
  NAND2_X1 U7404 ( .A1(n7634), .A2(n7633), .ZN(n10785) );
  AND2_X2 U7405 ( .A1(n13585), .A2(n13430), .ZN(n13600) );
  NAND4_X2 U7406 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        n12028) );
  AND4_X1 U7407 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n9535)
         );
  AOI222_X2 U7408 ( .A1(n8190), .A2(P2_REG1_REG_31__SCAN_IN), .B1(n8225), .B2(
        P2_REG2_REG_31__SCAN_IN), .C1(n8226), .C2(P2_REG0_REG_31__SCAN_IN), 
        .ZN(n12687) );
  BUF_X2 U7409 ( .A(n6478), .Z(n6481) );
  NAND4_X2 U7410 ( .A1(n9518), .A2(n9520), .A3(n9519), .A4(n9521), .ZN(n14853)
         );
  AND4_X2 U7411 ( .A1(n8912), .A2(n8909), .A3(n8910), .A4(n8911), .ZN(n9769)
         );
  INV_X1 U7412 ( .A(n8267), .ZN(n10309) );
  AND2_X1 U7413 ( .A1(n9377), .A2(n9376), .ZN(n7133) );
  AND3_X1 U7414 ( .A1(n10007), .A2(n10006), .A3(n10005), .ZN(n10146) );
  INV_X2 U7415 ( .A(n9977), .ZN(n13595) );
  AND2_X2 U7416 ( .A1(n9153), .A2(n9152), .ZN(n13311) );
  AND3_X1 U7417 ( .A1(n10021), .A2(n10020), .A3(n10019), .ZN(n10135) );
  OR2_X1 U7418 ( .A1(n9977), .A2(n8760), .ZN(n7509) );
  NAND4_X1 U7419 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .ZN(n8273)
         );
  NAND4_X1 U7420 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), .ZN(n8268)
         );
  AND2_X2 U7421 ( .A1(n11714), .A2(n8563), .ZN(n9739) );
  AND3_X1 U7422 ( .A1(n9516), .A2(n9515), .A3(n9514), .ZN(n9761) );
  NAND2_X1 U7423 ( .A1(n6918), .A2(n7566), .ZN(n14695) );
  NAND2_X1 U7424 ( .A1(n8905), .A2(n8906), .ZN(n9825) );
  OR2_X1 U7425 ( .A1(n11278), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U7426 ( .A1(n6475), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8929), .B2(
        n8939), .ZN(n7605) );
  CLKBUF_X2 U7427 ( .A(n8232), .Z(n6489) );
  XNOR2_X1 U7428 ( .A(n8425), .B(n8424), .ZN(n8486) );
  CLKBUF_X3 U7429 ( .A(n11453), .Z(n11464) );
  INV_X1 U7430 ( .A(n8907), .ZN(n8905) );
  INV_X1 U7431 ( .A(n8906), .ZN(n12419) );
  INV_X1 U7432 ( .A(n8370), .ZN(n10477) );
  XNOR2_X1 U7433 ( .A(n8619), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10556) );
  INV_X1 U7434 ( .A(n6798), .ZN(n8425) );
  INV_X2 U7435 ( .A(n8224), .ZN(n8186) );
  AND2_X2 U7436 ( .A1(n11804), .A2(n9466), .ZN(n11613) );
  NAND2_X1 U7437 ( .A1(n8551), .A2(n8647), .ZN(n9152) );
  BUF_X1 U7438 ( .A(n8632), .Z(n6480) );
  OR2_X1 U7439 ( .A1(n7775), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7777) );
  XNOR2_X1 U7440 ( .A(n8904), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8906) );
  INV_X1 U7441 ( .A(n7627), .ZN(n8929) );
  NOR2_X1 U7442 ( .A1(n10928), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n10953) );
  XNOR2_X1 U7443 ( .A(n7568), .B(n7567), .ZN(n11033) );
  NAND2_X1 U7444 ( .A1(n8692), .A2(n8691), .ZN(n10597) );
  AOI21_X1 U7445 ( .B1(n7597), .B2(n7598), .A(n6994), .ZN(n7621) );
  OR2_X1 U7446 ( .A1(n8290), .A2(n7929), .ZN(n7545) );
  OR2_X1 U7447 ( .A1(n7753), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7775) );
  XNOR2_X1 U7448 ( .A(n8550), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U7450 ( .A1(n8617), .A2(n8537), .ZN(n8623) );
  NAND2_X1 U7451 ( .A1(n8545), .A2(n8549), .ZN(n14170) );
  OR2_X1 U7452 ( .A1(n8903), .A2(n11301), .ZN(n8904) );
  INV_X2 U7453 ( .A(n12092), .ZN(n12069) );
  NAND2_X1 U7454 ( .A1(n7569), .A2(n7319), .ZN(n12996) );
  NOR2_X1 U7455 ( .A1(n8682), .A2(n9012), .ZN(n8800) );
  NAND2_X1 U7456 ( .A1(n8569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U7457 ( .A1(n7569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7568) );
  XNOR2_X1 U7458 ( .A(n8622), .B(n8621), .ZN(n13587) );
  XNOR2_X1 U7459 ( .A(n7670), .B(SI_4_), .ZN(n7669) );
  OR2_X1 U7460 ( .A1(n10823), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U7461 ( .A1(n6746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6745) );
  OR2_X1 U7462 ( .A1(n7729), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7753) );
  XNOR2_X1 U7463 ( .A(n7537), .B(n7539), .ZN(n10555) );
  OAI21_X1 U7464 ( .B1(n6483), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n6839), .ZN(
        n7655) );
  NAND2_X1 U7465 ( .A1(n9009), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9011) );
  NAND2_X1 U7466 ( .A1(n8549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8550) );
  OAI21_X1 U7467 ( .B1(n6483), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n6821), .ZN(
        n7670) );
  NAND2_X1 U7468 ( .A1(n9012), .A2(n9013), .ZN(n9009) );
  BUF_X2 U7469 ( .A(n6483), .Z(n6802) );
  NOR2_X1 U7470 ( .A1(n8579), .A2(n8578), .ZN(n6807) );
  OAI211_X1 U7471 ( .C1(n7036), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n6992), .B(
        n6990), .ZN(n6995) );
  NAND2_X2 U7472 ( .A1(n6484), .A2(P1_U3086), .ZN(n14166) );
  INV_X1 U7473 ( .A(n6717), .ZN(n9012) );
  CLKBUF_X3 U7474 ( .A(n9430), .Z(n6484) );
  NAND3_X1 U7475 ( .A1(n6900), .A2(n7553), .A3(n7554), .ZN(n7095) );
  NAND2_X1 U7476 ( .A1(n7038), .A2(n7036), .ZN(n9430) );
  AND2_X1 U7477 ( .A1(n8695), .A2(n6834), .ZN(n6510) );
  OR2_X1 U7478 ( .A1(n10022), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10070) );
  AND2_X1 U7479 ( .A1(n8558), .A2(n8537), .ZN(n7384) );
  NAND2_X1 U7480 ( .A1(n7037), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U7481 ( .A1(n7039), .A2(n7560), .ZN(n7038) );
  AND2_X1 U7482 ( .A1(n7551), .A2(n7552), .ZN(n7515) );
  AND2_X1 U7483 ( .A1(n8580), .A2(n6921), .ZN(n8582) );
  NAND2_X1 U7484 ( .A1(n8529), .A2(n7507), .ZN(n7506) );
  AND3_X1 U7485 ( .A1(n7662), .A2(n7630), .A3(n7676), .ZN(n7549) );
  AND4_X1 U7486 ( .A1(n8672), .A2(n8671), .A3(n8711), .A4(n8716), .ZN(n8673)
         );
  AND3_X1 U7487 ( .A1(n7534), .A2(n7536), .A3(n7535), .ZN(n7551) );
  AND3_X1 U7488 ( .A1(n8677), .A2(n8675), .A3(n8676), .ZN(n8695) );
  AND4_X1 U7489 ( .A1(n8294), .A2(n7539), .A3(n7864), .A4(n7843), .ZN(n7550)
         );
  AND3_X1 U7490 ( .A1(n7531), .A2(n7529), .A3(n7530), .ZN(n7552) );
  INV_X1 U7491 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8716) );
  INV_X1 U7492 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7179) );
  NOR2_X1 U7493 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8671) );
  INV_X1 U7494 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9564) );
  NOR2_X1 U7495 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7131) );
  INV_X1 U7496 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8711) );
  INV_X1 U7497 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8625) );
  NOR2_X1 U7498 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6803) );
  INV_X1 U7499 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8562) );
  NOR2_X1 U7500 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7132) );
  NOR2_X1 U7501 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7531) );
  INV_X1 U7502 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U7503 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7529) );
  NOR2_X1 U7504 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7530) );
  INV_X4 U7505 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7506 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7630) );
  NOR2_X1 U7507 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8676) );
  NOR2_X1 U7508 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8675) );
  NOR2_X1 U7509 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8677) );
  NOR2_X1 U7510 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7535) );
  NOR2_X1 U7511 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7536) );
  INV_X1 U7512 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7676) );
  NOR2_X1 U7513 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7534) );
  AND3_X2 U7514 ( .A1(n6803), .A2(n7131), .A3(n7132), .ZN(n8710) );
  NAND2_X1 U7515 ( .A1(n12534), .A2(n11738), .ZN(n12532) );
  XNOR2_X1 U7516 ( .A(n11741), .B(n11739), .ZN(n12534) );
  NOR2_X2 U7517 ( .A1(n12904), .A2(n12703), .ZN(n12691) );
  AND2_X2 U7518 ( .A1(n7544), .A2(n7543), .ZN(n8368) );
  AOI21_X2 U7519 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n8445), .A(n8444), .ZN(
        n8512) );
  XNOR2_X1 U7520 ( .A(n8571), .B(n8570), .ZN(n8632) );
  AND2_X2 U7521 ( .A1(n7987), .A2(n10555), .ZN(n8231) );
  INV_X1 U7522 ( .A(n7987), .ZN(n12679) );
  OAI21_X1 U7523 ( .B1(n8469), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6788), .ZN(
        n6798) );
  AND2_X4 U7524 ( .A1(n11714), .A2(n8564), .ZN(n8606) );
  CLKBUF_X2 U7525 ( .A(n6478), .Z(n6482) );
  INV_X2 U7526 ( .A(n9828), .ZN(n11433) );
  XOR2_X2 U7527 ( .A(n10315), .B(n11762), .Z(n6525) );
  OAI21_X2 U7528 ( .B1(n10360), .B2(n6676), .A(n6673), .ZN(n14825) );
  BUF_X4 U7529 ( .A(n9430), .Z(n6483) );
  AOI21_X4 U7530 ( .B1(n10573), .B2(n8186), .A(n6810), .ZN(n10315) );
  NAND2_X1 U7531 ( .A1(n12971), .A2(n12679), .ZN(n6487) );
  INV_X2 U7532 ( .A(n6487), .ZN(n12885) );
  AND2_X1 U7533 ( .A1(n12922), .A2(n12480), .ZN(n7061) );
  OR2_X1 U7534 ( .A1(n7219), .A2(n8407), .ZN(n7217) );
  AOI21_X1 U7535 ( .B1(n7216), .B2(n7222), .A(n7215), .ZN(n7214) );
  NOR2_X1 U7536 ( .A1(n7102), .A2(n12791), .ZN(n7215) );
  INV_X1 U7537 ( .A(n13465), .ZN(n6875) );
  NAND2_X1 U7538 ( .A1(n6870), .A2(n13484), .ZN(n6869) );
  NAND2_X1 U7539 ( .A1(n7278), .A2(n6871), .ZN(n6870) );
  XNOR2_X1 U7540 ( .A(n9014), .B(n9013), .ZN(n9016) );
  NAND2_X1 U7541 ( .A1(n6717), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9014) );
  INV_X1 U7542 ( .A(n6910), .ZN(n6909) );
  NAND2_X1 U7543 ( .A1(n7361), .A2(n6567), .ZN(n7360) );
  NAND2_X1 U7544 ( .A1(n13617), .A2(n6496), .ZN(n7361) );
  NAND2_X1 U7545 ( .A1(n9470), .A2(n8603), .ZN(n8614) );
  XNOR2_X1 U7546 ( .A(n14415), .B(n6747), .ZN(n8628) );
  NAND2_X1 U7547 ( .A1(n7330), .A2(n7329), .ZN(n8221) );
  AOI21_X1 U7548 ( .B1(n7332), .B2(n7335), .A(n6634), .ZN(n7329) );
  NOR2_X1 U7549 ( .A1(n14814), .A2(n7151), .ZN(n7150) );
  INV_X1 U7550 ( .A(n11543), .ZN(n7151) );
  INV_X1 U7551 ( .A(n8194), .ZN(n8023) );
  OAI21_X1 U7552 ( .B1(n12721), .B2(n7207), .A(n6965), .ZN(n12700) );
  INV_X1 U7553 ( .A(n6966), .ZN(n6965) );
  OAI21_X1 U7554 ( .B1(n12720), .B2(n7207), .A(n12701), .ZN(n6966) );
  NAND2_X1 U7555 ( .A1(n7303), .A2(n7302), .ZN(n7063) );
  INV_X1 U7556 ( .A(n7304), .ZN(n7302) );
  INV_X1 U7557 ( .A(n6734), .ZN(n6733) );
  OAI21_X1 U7558 ( .B1(n8405), .B2(n6735), .A(n8406), .ZN(n6734) );
  INV_X1 U7559 ( .A(n13634), .ZN(n7265) );
  AND2_X1 U7560 ( .A1(n7384), .A2(n8570), .ZN(n6502) );
  INV_X1 U7561 ( .A(n7643), .ZN(n6653) );
  OAI22_X1 U7562 ( .A1(n13461), .A2(n7272), .B1(n13462), .B2(n7273), .ZN(
        n13466) );
  INV_X1 U7563 ( .A(n6868), .ZN(n6867) );
  OAI21_X1 U7564 ( .B1(n6869), .B2(n6871), .A(n13483), .ZN(n6868) );
  AND2_X1 U7565 ( .A1(n7877), .A2(n7462), .ZN(n7461) );
  INV_X1 U7566 ( .A(n7878), .ZN(n7462) );
  AND2_X1 U7567 ( .A1(n7253), .A2(n7252), .ZN(n7251) );
  NOR2_X1 U7568 ( .A1(n13500), .A2(n13503), .ZN(n7253) );
  AOI21_X1 U7569 ( .B1(n7494), .B2(n7963), .A(n6583), .ZN(n7491) );
  NOR2_X1 U7570 ( .A1(n7494), .A2(n7493), .ZN(n7492) );
  NAND2_X1 U7571 ( .A1(n6661), .A2(n6660), .ZN(n7490) );
  AOI22_X1 U7572 ( .A1(n12946), .A2(n8235), .B1(n6482), .B2(n12817), .ZN(n8044) );
  NAND2_X1 U7573 ( .A1(n6664), .A2(n8065), .ZN(n8066) );
  INV_X1 U7574 ( .A(n8063), .ZN(n6664) );
  NAND2_X1 U7575 ( .A1(n6858), .A2(n6859), .ZN(n13547) );
  AND2_X1 U7576 ( .A1(n8680), .A2(n8678), .ZN(n7424) );
  INV_X1 U7577 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8680) );
  INV_X1 U7578 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8678) );
  OAI21_X1 U7579 ( .B1(n9758), .B2(n6631), .A(n6778), .ZN(n10844) );
  INV_X1 U7580 ( .A(n6779), .ZN(n6778) );
  NAND2_X1 U7581 ( .A1(n7226), .A2(n6630), .ZN(n7030) );
  NAND2_X1 U7582 ( .A1(n7353), .A2(n10649), .ZN(n6647) );
  XNOR2_X1 U7583 ( .A(n7354), .B(n7987), .ZN(n7353) );
  NAND2_X1 U7584 ( .A1(n12495), .A2(n12862), .ZN(n7296) );
  AND2_X1 U7585 ( .A1(n10754), .A2(n6536), .ZN(n7312) );
  NOR2_X1 U7586 ( .A1(n10651), .A2(n10483), .ZN(n6896) );
  INV_X1 U7587 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7314) );
  INV_X1 U7588 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8294) );
  INV_X1 U7589 ( .A(n9152), .ZN(n9156) );
  NOR2_X1 U7590 ( .A1(n14063), .A2(n7114), .ZN(n7113) );
  INV_X1 U7591 ( .A(n7115), .ZN(n7114) );
  AOI21_X1 U7592 ( .B1(n13891), .B2(n11231), .A(n11230), .ZN(n13872) );
  NOR2_X1 U7593 ( .A1(n13617), .A2(n7190), .ZN(n7189) );
  INV_X1 U7594 ( .A(n10393), .ZN(n7190) );
  INV_X1 U7595 ( .A(n13433), .ZN(n9153) );
  NOR2_X1 U7596 ( .A1(n8564), .A2(n11714), .ZN(n8604) );
  OR2_X1 U7597 ( .A1(n8661), .A2(n10556), .ZN(n9165) );
  OR2_X1 U7598 ( .A1(n8221), .A2(n8220), .ZN(n8223) );
  NAND2_X1 U7599 ( .A1(n8144), .A2(n8143), .ZN(n8185) );
  INV_X1 U7600 ( .A(n6962), .ZN(n6959) );
  NAND2_X1 U7601 ( .A1(n7041), .A2(n8045), .ZN(n6962) );
  INV_X1 U7602 ( .A(n7042), .ZN(n7041) );
  OAI21_X1 U7603 ( .B1(n8012), .B2(n8028), .A(n7043), .ZN(n7042) );
  NAND2_X1 U7604 ( .A1(n7044), .A2(n11361), .ZN(n7043) );
  INV_X1 U7605 ( .A(n8011), .ZN(n7044) );
  NAND2_X1 U7606 ( .A1(n7343), .A2(n7341), .ZN(n7045) );
  NOR2_X1 U7607 ( .A1(n6960), .A2(n8007), .ZN(n7341) );
  NAND2_X1 U7608 ( .A1(n7052), .A2(n7050), .ZN(n7883) );
  AOI21_X1 U7609 ( .B1(n7057), .B2(n7054), .A(n7053), .ZN(n7052) );
  AND2_X1 U7610 ( .A1(n7054), .A2(n7816), .ZN(n7049) );
  NAND2_X1 U7611 ( .A1(n6483), .A2(n8736), .ZN(n6821) );
  OAI21_X1 U7612 ( .B1(n11932), .B2(n11827), .A(n11829), .ZN(n11941) );
  OAI21_X1 U7613 ( .B1(n7078), .B2(n6515), .A(n7074), .ZN(n7073) );
  NAND2_X1 U7614 ( .A1(n6515), .A2(n7075), .ZN(n7074) );
  OR2_X1 U7615 ( .A1(n7078), .A2(n7080), .ZN(n7075) );
  NOR2_X1 U7616 ( .A1(n7093), .A2(n6613), .ZN(n7092) );
  INV_X1 U7617 ( .A(n10998), .ZN(n7093) );
  NAND2_X1 U7618 ( .A1(n6829), .A2(n6613), .ZN(n11810) );
  NAND2_X1 U7619 ( .A1(n10999), .A2(n10998), .ZN(n6829) );
  NOR2_X1 U7620 ( .A1(n11652), .A2(n12309), .ZN(n11653) );
  NOR2_X1 U7621 ( .A1(n7033), .A2(n11647), .ZN(n11648) );
  NAND2_X1 U7622 ( .A1(n8907), .A2(n12419), .ZN(n9605) );
  NOR2_X1 U7623 ( .A1(n10851), .A2(n10597), .ZN(n8693) );
  NAND2_X1 U7624 ( .A1(n9238), .A2(n9239), .ZN(n9287) );
  XNOR2_X1 U7625 ( .A(n9667), .B(n10018), .ZN(n9288) );
  NAND2_X1 U7626 ( .A1(n9963), .A2(n9964), .ZN(n10099) );
  AND2_X1 U7627 ( .A1(n6712), .A2(n6711), .ZN(n6710) );
  OR2_X1 U7628 ( .A1(n6713), .A2(n9952), .ZN(n6712) );
  INV_X1 U7629 ( .A(n10093), .ZN(n6711) );
  XNOR2_X1 U7630 ( .A(n10211), .B(n10922), .ZN(n10101) );
  OR2_X1 U7631 ( .A1(n9953), .A2(n6708), .ZN(n6707) );
  INV_X1 U7632 ( .A(n6709), .ZN(n6708) );
  AOI21_X1 U7633 ( .B1(n6706), .B2(n6709), .A(n6705), .ZN(n6704) );
  INV_X1 U7634 ( .A(n10206), .ZN(n6705) );
  INV_X1 U7635 ( .A(n6710), .ZN(n6706) );
  NAND2_X1 U7636 ( .A1(n11790), .A2(n11786), .ZN(n6777) );
  OR2_X1 U7637 ( .A1(n11612), .A2(n11603), .ZN(n11683) );
  AOI21_X1 U7638 ( .B1(n11624), .B2(n6675), .A(n6674), .ZN(n6673) );
  INV_X1 U7639 ( .A(n11539), .ZN(n6674) );
  INV_X1 U7640 ( .A(n11533), .ZN(n6675) );
  AND3_X1 U7641 ( .A1(n10065), .A2(n10064), .A3(n10063), .ZN(n14841) );
  NAND2_X1 U7642 ( .A1(n6476), .A2(n8799), .ZN(n9364) );
  INV_X1 U7643 ( .A(n9016), .ZN(n12092) );
  NAND2_X1 U7644 ( .A1(n6752), .A2(n6755), .ZN(n11261) );
  INV_X1 U7645 ( .A(n6756), .ZN(n6755) );
  NAND2_X1 U7646 ( .A1(n10894), .A2(n6753), .ZN(n6752) );
  OAI21_X1 U7647 ( .B1(n11248), .B2(n6636), .A(n7240), .ZN(n6756) );
  NAND2_X1 U7648 ( .A1(n10894), .A2(n10893), .ZN(n6757) );
  NOR2_X1 U7649 ( .A1(n11008), .A2(n8696), .ZN(n9344) );
  XNOR2_X1 U7650 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n10600) );
  XNOR2_X1 U7651 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8718) );
  NAND2_X1 U7652 ( .A1(n9901), .A2(n7400), .ZN(n7399) );
  NAND2_X1 U7653 ( .A1(n11730), .A2(n6987), .ZN(n6986) );
  INV_X1 U7654 ( .A(n11733), .ZN(n6987) );
  INV_X1 U7655 ( .A(n6643), .ZN(n6649) );
  INV_X1 U7656 ( .A(n7646), .ZN(n8077) );
  AND2_X1 U7657 ( .A1(n7578), .A2(n7570), .ZN(n7647) );
  AND2_X1 U7658 ( .A1(n7578), .A2(n12996), .ZN(n7646) );
  AND2_X1 U7659 ( .A1(n7570), .A2(n11033), .ZN(n7514) );
  AOI21_X1 U7660 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n12721) );
  NAND2_X1 U7661 ( .A1(n12922), .A2(n12747), .ZN(n7209) );
  NOR2_X1 U7662 ( .A1(n12747), .A2(n12922), .ZN(n7208) );
  AND2_X1 U7663 ( .A1(n12951), .A2(n12465), .ZN(n7316) );
  NAND2_X1 U7664 ( .A1(n8335), .A2(n12802), .ZN(n7317) );
  INV_X1 U7665 ( .A(n12815), .ZN(n7318) );
  AOI21_X1 U7666 ( .B1(n7234), .B2(n7237), .A(n6558), .ZN(n7233) );
  INV_X1 U7667 ( .A(n7234), .ZN(n7232) );
  NOR2_X1 U7668 ( .A1(n9648), .A2(n7309), .ZN(n7308) );
  INV_X1 U7669 ( .A(n8319), .ZN(n7309) );
  NAND2_X1 U7670 ( .A1(n10258), .A2(n10262), .ZN(n7212) );
  AOI21_X1 U7671 ( .B1(n6907), .B2(n6903), .A(n6577), .ZN(n6902) );
  INV_X1 U7672 ( .A(n6912), .ZN(n6903) );
  AND2_X1 U7673 ( .A1(n8553), .A2(n8930), .ZN(n9083) );
  AND2_X1 U7674 ( .A1(n8348), .A2(n13004), .ZN(n14681) );
  OR2_X1 U7675 ( .A1(n8297), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U7676 ( .A1(n10351), .A2(n10350), .ZN(n6946) );
  AOI22_X1 U7677 ( .A1(n13571), .A2(n13570), .B1(n13569), .B2(n13568), .ZN(
        n13591) );
  INV_X1 U7678 ( .A(n13590), .ZN(n7266) );
  AND2_X1 U7679 ( .A1(n8643), .A2(n9152), .ZN(n8644) );
  AND2_X1 U7680 ( .A1(n13793), .A2(n11205), .ZN(n13631) );
  AND4_X1 U7681 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n14001) );
  OAI21_X1 U7682 ( .B1(n13666), .B2(n14426), .A(n7382), .ZN(n9975) );
  NAND2_X1 U7683 ( .A1(n9812), .A2(n9811), .ZN(n14410) );
  NAND2_X1 U7684 ( .A1(n8631), .A2(n8630), .ZN(n14411) );
  NAND2_X1 U7685 ( .A1(n10391), .A2(n10390), .ZN(n14498) );
  INV_X1 U7686 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8555) );
  XNOR2_X1 U7687 ( .A(n8087), .B(n11383), .ZN(n11130) );
  INV_X1 U7688 ( .A(n8700), .ZN(n6696) );
  NOR2_X1 U7689 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8531) );
  AND2_X1 U7690 ( .A1(n8533), .A2(n8534), .ZN(n6695) );
  NAND2_X1 U7691 ( .A1(n6850), .A2(n8536), .ZN(n10090) );
  INV_X1 U7692 ( .A(n9821), .ZN(n6850) );
  NOR2_X1 U7693 ( .A1(n7506), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n6841) );
  INV_X1 U7694 ( .A(n6784), .ZN(n8489) );
  OAI21_X1 U7695 ( .B1(n14971), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6564), .ZN(
        n6784) );
  NAND2_X1 U7696 ( .A1(n6678), .A2(n6537), .ZN(n11480) );
  INV_X1 U7697 ( .A(n6637), .ZN(n6713) );
  NOR2_X1 U7698 ( .A1(n12072), .A2(n12073), .ZN(n12093) );
  NAND2_X1 U7699 ( .A1(n6650), .A2(n7503), .ZN(n7694) );
  NAND2_X1 U7700 ( .A1(n7668), .A2(n7504), .ZN(n7503) );
  INV_X1 U7701 ( .A(n7667), .ZN(n7504) );
  NAND2_X1 U7702 ( .A1(n7723), .A2(n7722), .ZN(n6666) );
  NOR2_X1 U7703 ( .A1(n13468), .A2(n13471), .ZN(n7271) );
  NAND2_X1 U7704 ( .A1(n13468), .A2(n13471), .ZN(n7270) );
  NAND2_X1 U7705 ( .A1(n7833), .A2(n7832), .ZN(n6655) );
  NOR2_X1 U7706 ( .A1(n6867), .A2(n6865), .ZN(n6864) );
  NOR2_X1 U7707 ( .A1(n6866), .A2(n13484), .ZN(n6865) );
  INV_X1 U7708 ( .A(n6871), .ZN(n6866) );
  AOI21_X1 U7709 ( .B1(n6867), .B2(n6869), .A(n6506), .ZN(n6863) );
  NAND2_X1 U7710 ( .A1(n7461), .A2(n7459), .ZN(n7458) );
  OAI21_X1 U7711 ( .B1(n7454), .B2(n7457), .A(n7456), .ZN(n7451) );
  INV_X1 U7712 ( .A(n7895), .ZN(n7454) );
  NAND2_X1 U7713 ( .A1(n7455), .A2(n7461), .ZN(n7453) );
  NOR2_X1 U7714 ( .A1(n7496), .A2(n7979), .ZN(n7495) );
  INV_X1 U7715 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U7716 ( .B1(n6495), .B2(n7252), .A(n7254), .ZN(n7250) );
  INV_X1 U7717 ( .A(n13511), .ZN(n7254) );
  INV_X1 U7718 ( .A(n13510), .ZN(n7248) );
  NAND2_X1 U7719 ( .A1(n13543), .A2(n6860), .ZN(n6859) );
  AOI21_X1 U7720 ( .B1(n6575), .B2(n7501), .A(n7499), .ZN(n7498) );
  AND2_X1 U7721 ( .A1(n8043), .A2(n8044), .ZN(n7499) );
  INV_X1 U7722 ( .A(n8081), .ZN(n7489) );
  INV_X1 U7723 ( .A(n8082), .ZN(n7488) );
  NOR2_X1 U7724 ( .A1(n13546), .A2(n13549), .ZN(n7260) );
  NAND2_X1 U7725 ( .A1(n13549), .A2(n13546), .ZN(n7259) );
  OAI22_X1 U7726 ( .A1(n13540), .A2(n7277), .B1(n7276), .B2(n13541), .ZN(
        n13544) );
  INV_X1 U7727 ( .A(n13539), .ZN(n7276) );
  NOR2_X1 U7728 ( .A1(n13542), .A2(n13539), .ZN(n7277) );
  AND2_X1 U7729 ( .A1(n13545), .A2(n6862), .ZN(n6861) );
  INV_X1 U7730 ( .A(n13543), .ZN(n6862) );
  NOR2_X1 U7731 ( .A1(n7260), .A2(n6857), .ZN(n6856) );
  INV_X1 U7732 ( .A(n6859), .ZN(n6857) );
  AOI211_X1 U7733 ( .C1(n8248), .C2(n8246), .A(n8247), .B(n8245), .ZN(n8215)
         );
  NAND2_X1 U7734 ( .A1(n7243), .A2(n11614), .ZN(n7242) );
  NOR2_X1 U7735 ( .A1(n6491), .A2(n7032), .ZN(n7031) );
  INV_X1 U7736 ( .A(n6763), .ZN(n6762) );
  OAI21_X1 U7737 ( .B1(n11329), .B2(n6764), .A(n9637), .ZN(n6763) );
  INV_X1 U7738 ( .A(n7191), .ZN(n6764) );
  INV_X1 U7739 ( .A(n10487), .ZN(n7394) );
  NAND2_X1 U7740 ( .A1(n13560), .A2(n6845), .ZN(n6844) );
  INV_X1 U7741 ( .A(n7275), .ZN(n6845) );
  NAND2_X1 U7742 ( .A1(n7275), .A2(n7274), .ZN(n6847) );
  NOR2_X1 U7743 ( .A1(n6490), .A2(n6848), .ZN(n6843) );
  NOR2_X1 U7744 ( .A1(n13560), .A2(n6846), .ZN(n6848) );
  AOI21_X1 U7745 ( .B1(n7055), .B2(n7347), .A(n6581), .ZN(n7054) );
  AND2_X1 U7746 ( .A1(n7350), .A2(n7879), .ZN(n7055) );
  AND2_X1 U7747 ( .A1(n7352), .A2(n7520), .ZN(n7351) );
  INV_X1 U7748 ( .A(n7324), .ZN(n7323) );
  OAI21_X1 U7749 ( .B1(n7771), .B2(n7325), .A(n7798), .ZN(n7324) );
  INV_X1 U7750 ( .A(n7774), .ZN(n7325) );
  OAI21_X1 U7751 ( .B1(n8482), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6524), .ZN(
        n6789) );
  INV_X1 U7752 ( .A(n11484), .ZN(n7148) );
  NAND2_X1 U7753 ( .A1(n14781), .A2(n6881), .ZN(n9703) );
  NAND2_X1 U7754 ( .A1(n14796), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U7755 ( .A1(n9847), .A2(n6880), .ZN(n9960) );
  OR2_X1 U7756 ( .A1(n9849), .A2(n9848), .ZN(n6880) );
  NAND2_X1 U7757 ( .A1(n10095), .A2(n10096), .ZN(n10216) );
  INV_X1 U7758 ( .A(n7416), .ZN(n7415) );
  OR2_X1 U7759 ( .A1(n12346), .A2(n12206), .ZN(n11486) );
  NOR2_X1 U7760 ( .A1(n12204), .A2(n7417), .ZN(n7416) );
  INV_X1 U7761 ( .A(n11675), .ZN(n7417) );
  OR2_X1 U7762 ( .A1(n12351), .A2(n11961), .ZN(n11589) );
  OR2_X1 U7763 ( .A1(n11359), .A2(n7155), .ZN(n7154) );
  INV_X1 U7764 ( .A(n11492), .ZN(n7155) );
  AND2_X1 U7765 ( .A1(n12242), .A2(n11496), .ZN(n7156) );
  INV_X1 U7766 ( .A(n7407), .ZN(n7406) );
  OAI21_X1 U7767 ( .B1(n12290), .B2(n7408), .A(n11665), .ZN(n7407) );
  INV_X1 U7768 ( .A(n11664), .ZN(n7408) );
  OR2_X1 U7769 ( .A1(n14235), .A2(n11812), .ZN(n11556) );
  INV_X1 U7770 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9013) );
  INV_X1 U7771 ( .A(n9111), .ZN(n6768) );
  INV_X1 U7772 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U7773 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n9001), .ZN(n9108) );
  AOI21_X1 U7774 ( .B1(n7014), .B2(n7016), .A(n6582), .ZN(n7011) );
  NAND2_X1 U7775 ( .A1(n8731), .A2(n7014), .ZN(n7012) );
  INV_X1 U7776 ( .A(n12996), .ZN(n7570) );
  NOR2_X1 U7777 ( .A1(n12730), .A2(n12915), .ZN(n6823) );
  NOR2_X1 U7778 ( .A1(n12931), .A2(n7102), .ZN(n7101) );
  NAND2_X1 U7779 ( .A1(n6964), .A2(n12757), .ZN(n12755) );
  NAND2_X1 U7780 ( .A1(n6500), .A2(n7223), .ZN(n7222) );
  NAND2_X1 U7781 ( .A1(n9890), .A2(n9889), .ZN(n7313) );
  INV_X1 U7782 ( .A(n7300), .ZN(n7299) );
  OAI21_X1 U7783 ( .B1(n10259), .B2(n7301), .A(n8311), .ZN(n7300) );
  INV_X1 U7784 ( .A(n8310), .ZN(n7301) );
  NOR2_X1 U7785 ( .A1(n7061), .A2(n6913), .ZN(n6912) );
  NAND2_X1 U7786 ( .A1(n6823), .A2(n6822), .ZN(n12703) );
  INV_X1 U7787 ( .A(n12909), .ZN(n6822) );
  AND2_X1 U7788 ( .A1(n6898), .A2(n6531), .ZN(n7290) );
  OR2_X1 U7789 ( .A1(n8329), .A2(n6899), .ZN(n6898) );
  INV_X1 U7790 ( .A(n6748), .ZN(n12892) );
  NOR2_X1 U7791 ( .A1(n13839), .A2(n14074), .ZN(n7115) );
  NAND2_X1 U7792 ( .A1(n13939), .A2(n11120), .ZN(n7184) );
  NOR2_X1 U7793 ( .A1(n13520), .A2(n6729), .ZN(n6728) );
  INV_X1 U7794 ( .A(n6731), .ZN(n6729) );
  NOR2_X1 U7795 ( .A1(n14291), .A2(n13499), .ZN(n7120) );
  OR2_X1 U7796 ( .A1(n13620), .A2(n7169), .ZN(n7168) );
  INV_X1 U7797 ( .A(n10795), .ZN(n7169) );
  INV_X1 U7798 ( .A(n7363), .ZN(n7358) );
  NAND2_X1 U7799 ( .A1(n10355), .A2(n10192), .ZN(n7370) );
  AND2_X1 U7800 ( .A1(n7370), .A2(n9976), .ZN(n7363) );
  AND2_X1 U7801 ( .A1(n7366), .A2(n7365), .ZN(n7364) );
  INV_X1 U7802 ( .A(n13614), .ZN(n7365) );
  NAND2_X1 U7803 ( .A1(n7045), .A2(n8011), .ZN(n7040) );
  NAND2_X1 U7804 ( .A1(n7983), .A2(n7982), .ZN(n7343) );
  AND2_X1 U7805 ( .A1(n7942), .A2(n7927), .ZN(n7940) );
  NAND2_X1 U7806 ( .A1(n7345), .A2(n7344), .ZN(n7905) );
  INV_X1 U7807 ( .A(n7897), .ZN(n7346) );
  AOI21_X1 U7808 ( .B1(n7351), .B2(n7349), .A(n7348), .ZN(n7347) );
  INV_X1 U7809 ( .A(n7838), .ZN(n7349) );
  INV_X1 U7810 ( .A(n7862), .ZN(n7348) );
  INV_X1 U7811 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7507) );
  NOR2_X1 U7812 ( .A1(n6995), .A2(n9431), .ZN(n6994) );
  INV_X1 U7813 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8419) );
  OAI22_X1 U7814 ( .A1(n8490), .A2(n8428), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14805), .ZN(n8429) );
  INV_X1 U7815 ( .A(n11817), .ZN(n7067) );
  AOI21_X1 U7816 ( .B1(n7083), .B2(n7082), .A(n6616), .ZN(n7081) );
  INV_X1 U7817 ( .A(n11958), .ZN(n7082) );
  NAND2_X1 U7818 ( .A1(n10128), .A2(n10127), .ZN(n7091) );
  INV_X1 U7819 ( .A(n11988), .ZN(n12013) );
  AND4_X1 U7820 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11929) );
  NAND2_X1 U7821 ( .A1(n9287), .A2(n6540), .ZN(n9667) );
  OAI21_X1 U7822 ( .B1(n9677), .B2(n14958), .A(n14784), .ZN(n9698) );
  XNOR2_X1 U7823 ( .A(n9703), .B(n10156), .ZN(n9671) );
  NAND2_X1 U7824 ( .A1(n9707), .A2(n9708), .ZN(n9847) );
  XNOR2_X1 U7825 ( .A(n9960), .B(n10602), .ZN(n9850) );
  NAND2_X1 U7826 ( .A1(n9957), .A2(n9958), .ZN(n10095) );
  NAND2_X1 U7827 ( .A1(n10099), .A2(n10100), .ZN(n10211) );
  NAND2_X1 U7828 ( .A1(n10723), .A2(n10724), .ZN(n10726) );
  NAND2_X1 U7829 ( .A1(n10726), .A2(n10725), .ZN(n11017) );
  XNOR2_X1 U7830 ( .A(n12032), .B(n6882), .ZN(n11019) );
  NAND2_X1 U7831 ( .A1(n11017), .A2(n11018), .ZN(n12032) );
  OR2_X1 U7832 ( .A1(n12321), .A2(n11795), .ZN(n11484) );
  NAND2_X1 U7833 ( .A1(n11791), .A2(n6554), .ZN(n6776) );
  AND2_X1 U7834 ( .A1(n11396), .A2(n11395), .ZN(n11845) );
  NAND2_X1 U7835 ( .A1(n11393), .A2(n11464), .ZN(n11396) );
  NAND2_X1 U7836 ( .A1(n7418), .A2(n7416), .ZN(n12201) );
  NAND2_X1 U7837 ( .A1(n12212), .A2(n11674), .ZN(n7418) );
  AND2_X1 U7838 ( .A1(n11589), .A2(n11588), .ZN(n12204) );
  NAND2_X1 U7839 ( .A1(n12219), .A2(n12218), .ZN(n12217) );
  OR2_X1 U7840 ( .A1(n12362), .A2(n12224), .ZN(n11492) );
  NAND2_X1 U7841 ( .A1(n12236), .A2(n6505), .ZN(n12227) );
  NAND2_X1 U7842 ( .A1(n12249), .A2(n7156), .ZN(n12241) );
  AND2_X1 U7843 ( .A1(n11570), .A2(n11575), .ZN(n12276) );
  NAND2_X1 U7844 ( .A1(n12281), .A2(n12290), .ZN(n12280) );
  NAND2_X1 U7845 ( .A1(n14188), .A2(n11464), .ZN(n11271) );
  NAND2_X1 U7846 ( .A1(n10942), .A2(n6546), .ZN(n14821) );
  AND4_X1 U7847 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n14818) );
  AOI21_X1 U7848 ( .B1(n7412), .B2(n7410), .A(n6571), .ZN(n7409) );
  NAND2_X1 U7849 ( .A1(n9391), .A2(n11613), .ZN(n14867) );
  INV_X1 U7850 ( .A(n14890), .ZN(n14869) );
  AND3_X1 U7851 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n14887) );
  NAND2_X1 U7852 ( .A1(n11453), .A2(n9429), .ZN(n9435) );
  AND2_X1 U7853 ( .A1(n11656), .A2(n11499), .ZN(n14916) );
  AND2_X1 U7854 ( .A1(n9368), .A2(n9015), .ZN(n9619) );
  INV_X1 U7855 ( .A(n14916), .ZN(n14886) );
  AOI21_X1 U7856 ( .B1(n11261), .B2(n11249), .A(n7239), .ZN(n11444) );
  AND2_X1 U7857 ( .A1(n14162), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7239) );
  MUX2_X1 U7858 ( .A(n11301), .B(n8679), .S(P3_IR_REG_26__SCAN_IN), .Z(n8682)
         );
  NAND2_X1 U7859 ( .A1(n10846), .A2(n10847), .ZN(n10894) );
  NOR2_X1 U7860 ( .A1(n10121), .A2(n7229), .ZN(n7228) );
  INV_X1 U7861 ( .A(n7230), .ZN(n7229) );
  NAND2_X1 U7862 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n7231), .ZN(n7230) );
  NAND2_X1 U7863 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  NAND2_X1 U7864 ( .A1(n9758), .A2(n9757), .ZN(n9859) );
  INV_X1 U7865 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8697) );
  XNOR2_X1 U7866 ( .A(n9756), .B(n10553), .ZN(n9755) );
  NAND2_X1 U7867 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7192), .ZN(n7191) );
  NAND2_X1 U7868 ( .A1(n9217), .A2(n9216), .ZN(n11331) );
  NAND2_X1 U7869 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n9824), .ZN(n9216) );
  NAND2_X1 U7870 ( .A1(n9115), .A2(n9114), .ZN(n11300) );
  INV_X1 U7871 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U7872 ( .A1(n8789), .A2(n6530), .ZN(n11008) );
  AND2_X1 U7873 ( .A1(n8673), .A2(n8710), .ZN(n8789) );
  INV_X1 U7874 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8674) );
  XNOR2_X1 U7875 ( .A(n9109), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n11267) );
  XNOR2_X1 U7876 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8765) );
  NAND2_X1 U7877 ( .A1(n7012), .A2(n7011), .ZN(n8766) );
  XNOR2_X1 U7878 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8729) );
  NOR2_X1 U7879 ( .A1(n6609), .A2(n7204), .ZN(n7203) );
  INV_X1 U7880 ( .A(n8709), .ZN(n7204) );
  NAND2_X1 U7881 ( .A1(n8777), .A2(n8776), .ZN(n7205) );
  NAND2_X1 U7882 ( .A1(n6771), .A2(n8708), .ZN(n8777) );
  NAND2_X1 U7883 ( .A1(n8753), .A2(n8752), .ZN(n6771) );
  INV_X1 U7884 ( .A(n8750), .ZN(n7413) );
  INV_X1 U7885 ( .A(n12915), .ZN(n12432) );
  AND2_X1 U7886 ( .A1(n12450), .A2(n11731), .ZN(n11732) );
  NOR2_X1 U7887 ( .A1(n12426), .A2(n7391), .ZN(n7390) );
  INV_X1 U7888 ( .A(n11757), .ZN(n7391) );
  INV_X1 U7889 ( .A(n7399), .ZN(n7398) );
  NAND2_X1 U7890 ( .A1(n9640), .A2(n9641), .ZN(n9902) );
  OR2_X1 U7891 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  NAND2_X1 U7892 ( .A1(n6641), .A2(n6640), .ZN(n6643) );
  INV_X1 U7893 ( .A(n8262), .ZN(n6640) );
  NAND2_X1 U7894 ( .A1(n8264), .A2(n8263), .ZN(n6641) );
  NAND2_X1 U7895 ( .A1(n6647), .A2(n6638), .ZN(n6644) );
  INV_X1 U7896 ( .A(n6647), .ZN(n6646) );
  AND2_X1 U7897 ( .A1(n7999), .A2(n7998), .ZN(n12525) );
  NOR2_X1 U7898 ( .A1(n12432), .A2(n12576), .ZN(n6905) );
  NAND2_X1 U7899 ( .A1(n6911), .A2(n6907), .ZN(n6906) );
  OR2_X1 U7900 ( .A1(n7061), .A2(n8338), .ZN(n6910) );
  NAND2_X1 U7901 ( .A1(n12745), .A2(n6912), .ZN(n6911) );
  XNOR2_X1 U7902 ( .A(n12783), .B(n12791), .ZN(n12784) );
  NAND2_X1 U7903 ( .A1(n7224), .A2(n12536), .ZN(n7223) );
  NOR2_X1 U7904 ( .A1(n12805), .A2(n8407), .ZN(n7225) );
  NAND2_X1 U7905 ( .A1(n12801), .A2(n6542), .ZN(n7315) );
  INV_X1 U7906 ( .A(n12863), .ZN(n7237) );
  NOR2_X1 U7907 ( .A1(n12845), .A2(n7235), .ZN(n7234) );
  INV_X1 U7908 ( .A(n8402), .ZN(n7235) );
  INV_X1 U7909 ( .A(n7296), .ZN(n7289) );
  AOI21_X1 U7910 ( .B1(n6896), .B2(n14264), .A(n6587), .ZN(n6893) );
  NAND2_X1 U7911 ( .A1(n8329), .A2(n10687), .ZN(n6897) );
  INV_X1 U7912 ( .A(n12883), .ZN(n11719) );
  NAND2_X1 U7913 ( .A1(n6892), .A2(n7310), .ZN(n10662) );
  OR2_X1 U7914 ( .A1(n7312), .A2(n6498), .ZN(n7310) );
  NOR2_X1 U7915 ( .A1(n6498), .A2(n8325), .ZN(n7311) );
  OR2_X1 U7916 ( .A1(n7825), .A2(n7824), .ZN(n7849) );
  NAND2_X1 U7917 ( .A1(n10766), .A2(n14276), .ZN(n10765) );
  NOR2_X1 U7918 ( .A1(n10694), .A2(n7194), .ZN(n7193) );
  INV_X1 U7919 ( .A(n8387), .ZN(n7194) );
  INV_X1 U7920 ( .A(n12773), .ZN(n12882) );
  NAND2_X1 U7921 ( .A1(n9494), .A2(n9493), .ZN(n9492) );
  AND2_X1 U7922 ( .A1(n10337), .A2(n10284), .ZN(n10281) );
  NOR2_X2 U7923 ( .A1(n10334), .A2(n14727), .ZN(n10337) );
  XNOR2_X1 U7924 ( .A(n12586), .B(n6738), .ZN(n10262) );
  NAND2_X1 U7925 ( .A1(n8309), .A2(n10259), .ZN(n10264) );
  NAND2_X1 U7926 ( .A1(n10774), .A2(n8383), .ZN(n6739) );
  INV_X1 U7927 ( .A(n12586), .ZN(n10779) );
  NAND2_X1 U7928 ( .A1(n6724), .A2(n8379), .ZN(n10300) );
  NAND2_X1 U7929 ( .A1(n7197), .A2(n9075), .ZN(n6724) );
  INV_X1 U7930 ( .A(n9080), .ZN(n9487) );
  INV_X1 U7931 ( .A(n12879), .ZN(n12774) );
  INV_X1 U7932 ( .A(n10315), .ZN(n9894) );
  INV_X1 U7933 ( .A(n10324), .ZN(n9655) );
  OR2_X1 U7934 ( .A1(n9731), .A2(n8224), .ZN(n7665) );
  OR2_X1 U7935 ( .A1(n8601), .A2(n8224), .ZN(n7606) );
  NAND2_X1 U7936 ( .A1(n7556), .A2(n6534), .ZN(n6901) );
  XNOR2_X1 U7937 ( .A(n8301), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U7938 ( .A1(n8294), .A2(n8295), .ZN(n8297) );
  XNOR2_X1 U7939 ( .A(n8294), .B(n8292), .ZN(n8930) );
  OR2_X1 U7940 ( .A1(n7673), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7675) );
  AND2_X1 U7941 ( .A1(n6518), .A2(n13099), .ZN(n7476) );
  NAND2_X1 U7942 ( .A1(n7475), .A2(n6518), .ZN(n7474) );
  INV_X1 U7943 ( .A(n13406), .ZN(n7475) );
  AOI22_X1 U7944 ( .A1(n9721), .A2(n9720), .B1(n9719), .B2(n9718), .ZN(n14369)
         );
  AOI21_X1 U7945 ( .B1(n6950), .B2(n6952), .A(n6507), .ZN(n6949) );
  NOR2_X1 U7946 ( .A1(n6557), .A2(n13026), .ZN(n7430) );
  OR2_X1 U7947 ( .A1(n13029), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U7948 ( .A1(n7433), .A2(n13026), .ZN(n7429) );
  AND2_X1 U7949 ( .A1(n13029), .A2(n13417), .ZN(n7433) );
  AND2_X1 U7950 ( .A1(n13118), .A2(n7481), .ZN(n7480) );
  OR2_X1 U7951 ( .A1(n13385), .A2(n7482), .ZN(n7481) );
  INV_X1 U7952 ( .A(n13079), .ZN(n7482) );
  INV_X1 U7953 ( .A(n6945), .ZN(n6943) );
  NAND2_X1 U7954 ( .A1(n13394), .A2(n6522), .ZN(n13298) );
  NOR2_X1 U7955 ( .A1(n14170), .A2(n10994), .ZN(n8551) );
  NOR2_X1 U7956 ( .A1(n11055), .A2(n6983), .ZN(n8853) );
  NOR2_X1 U7957 ( .A1(n11059), .A2(n8850), .ZN(n6983) );
  OR2_X1 U7958 ( .A1(n8853), .A2(n8852), .ZN(n6982) );
  NOR2_X1 U7959 ( .A1(n13735), .A2(n6976), .ZN(n13739) );
  AND2_X1 U7960 ( .A1(n13736), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6976) );
  OR2_X1 U7961 ( .A1(n13739), .A2(n13738), .ZN(n6975) );
  NAND2_X1 U7962 ( .A1(n6852), .A2(n6851), .ZN(n9821) );
  INV_X1 U7963 ( .A(n9661), .ZN(n6852) );
  XNOR2_X1 U7964 ( .A(n6973), .B(n13767), .ZN(n13753) );
  NAND2_X1 U7965 ( .A1(n6975), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U7966 ( .A1(n13752), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U7967 ( .A1(n13818), .A2(n7383), .ZN(n13800) );
  AND2_X1 U7968 ( .A1(n11237), .A2(n11236), .ZN(n7383) );
  NAND2_X1 U7969 ( .A1(n13834), .A2(n11186), .ZN(n13821) );
  NAND2_X1 U7970 ( .A1(n13821), .A2(n13822), .ZN(n13820) );
  AOI21_X1 U7971 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n7371) );
  INV_X1 U7972 ( .A(n11233), .ZN(n7372) );
  AND2_X1 U7973 ( .A1(n11186), .A2(n11184), .ZN(n13838) );
  NAND2_X1 U7974 ( .A1(n13872), .A2(n13871), .ZN(n13870) );
  NAND2_X1 U7975 ( .A1(n13873), .A2(n6543), .ZN(n13849) );
  NAND2_X1 U7976 ( .A1(n13897), .A2(n6697), .ZN(n13873) );
  NOR2_X1 U7977 ( .A1(n13871), .A2(n6698), .ZN(n6697) );
  INV_X1 U7978 ( .A(n11154), .ZN(n6698) );
  OAI21_X1 U7979 ( .B1(n13951), .B2(n11112), .A(n11111), .ZN(n13938) );
  OR2_X1 U7980 ( .A1(n13938), .A2(n13939), .ZN(n13936) );
  OR2_X1 U7981 ( .A1(n14116), .A2(n13965), .ZN(n11224) );
  NAND2_X1 U7982 ( .A1(n13952), .A2(n11112), .ZN(n11225) );
  NAND2_X1 U7983 ( .A1(n13996), .A2(n7185), .ZN(n13984) );
  NOR2_X1 U7984 ( .A1(n13980), .A2(n7186), .ZN(n7185) );
  INV_X1 U7985 ( .A(n11077), .ZN(n7186) );
  NAND2_X1 U7986 ( .A1(n14008), .A2(n14014), .ZN(n6731) );
  NAND2_X1 U7987 ( .A1(n11069), .A2(n6699), .ZN(n13996) );
  AND2_X1 U7988 ( .A1(n13626), .A2(n13509), .ZN(n6699) );
  OR2_X1 U7989 ( .A1(n14307), .A2(n14001), .ZN(n13509) );
  NAND2_X1 U7990 ( .A1(n7377), .A2(n6528), .ZN(n7376) );
  INV_X1 U7991 ( .A(n7380), .ZN(n7377) );
  NOR2_X1 U7992 ( .A1(n14024), .A2(n7381), .ZN(n7380) );
  INV_X1 U7993 ( .A(n7513), .ZN(n7381) );
  AND4_X1 U7994 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n14016) );
  AND2_X1 U7995 ( .A1(n13509), .A2(n13508), .ZN(n14024) );
  NOR2_X1 U7996 ( .A1(n13499), .A2(n13658), .ZN(n6805) );
  NAND2_X1 U7997 ( .A1(n10975), .A2(n13504), .ZN(n11218) );
  NAND2_X1 U7998 ( .A1(n10793), .A2(n10792), .ZN(n13490) );
  AOI21_X1 U7999 ( .B1(n6692), .B2(n7187), .A(n6568), .ZN(n6691) );
  INV_X1 U8000 ( .A(n7187), .ZN(n6693) );
  OR2_X1 U8001 ( .A1(n13482), .A2(n13661), .ZN(n6749) );
  NOR2_X1 U8002 ( .A1(n10513), .A2(n7188), .ZN(n7187) );
  INV_X1 U8003 ( .A(n10507), .ZN(n7188) );
  NAND2_X1 U8004 ( .A1(n10394), .A2(n7189), .ZN(n10508) );
  NOR2_X1 U8005 ( .A1(n6538), .A2(n7175), .ZN(n7174) );
  OAI211_X1 U8006 ( .C1(n13574), .C2(n9919), .A(n9918), .B(n9917), .ZN(n13464)
         );
  XNOR2_X1 U8007 ( .A(n13665), .B(n14475), .ZN(n14396) );
  NAND2_X1 U8008 ( .A1(n9985), .A2(n6688), .ZN(n6687) );
  NOR2_X1 U8009 ( .A1(n14410), .A2(n6690), .ZN(n6685) );
  INV_X1 U8010 ( .A(n14396), .ZN(n14394) );
  XNOR2_X1 U8011 ( .A(n14414), .B(n9973), .ZN(n13611) );
  AND2_X1 U8012 ( .A1(n8626), .A2(n13022), .ZN(n9805) );
  OAI211_X1 U8013 ( .C1(n9474), .C2(n7173), .A(n7172), .B(n13616), .ZN(n9812)
         );
  INV_X1 U8014 ( .A(n13446), .ZN(n7173) );
  INV_X1 U8015 ( .A(n8628), .ZN(n13616) );
  AND4_X2 U8016 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n13431)
         );
  INV_X1 U8017 ( .A(n14291), .ZN(n14315) );
  AND3_X1 U8018 ( .A1(n9736), .A2(n9735), .A3(n9734), .ZN(n14461) );
  AND2_X1 U8019 ( .A1(n8223), .A2(n8222), .ZN(n13572) );
  AND2_X1 U8020 ( .A1(n8539), .A2(n6533), .ZN(n7177) );
  NAND2_X1 U8021 ( .A1(n6960), .A2(n6959), .ZN(n6958) );
  NOR2_X1 U8022 ( .A1(n6962), .A2(n7981), .ZN(n6957) );
  NAND2_X1 U8023 ( .A1(n7345), .A2(n7883), .ZN(n7898) );
  NAND2_X1 U8024 ( .A1(n7322), .A2(n7774), .ZN(n7799) );
  AOI21_X1 U8025 ( .B1(n7327), .B2(n7669), .A(n6580), .ZN(n7326) );
  INV_X1 U8026 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6921) );
  INV_X1 U8027 ( .A(n6827), .ZN(n8473) );
  NAND2_X1 U8028 ( .A1(n8484), .A2(n8485), .ZN(n8488) );
  NAND2_X1 U8029 ( .A1(n7125), .A2(n8492), .ZN(n8495) );
  NOR2_X1 U8030 ( .A1(n8500), .A2(n8501), .ZN(n8504) );
  NAND2_X1 U8031 ( .A1(n14209), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6796) );
  INV_X1 U8032 ( .A(n14353), .ZN(n7123) );
  AOI21_X1 U8033 ( .B1(n14632), .B2(n8514), .A(n14356), .ZN(n8515) );
  OAI21_X1 U8034 ( .B1(n10128), .B2(n7089), .A(n7086), .ZN(n10233) );
  AOI21_X1 U8035 ( .B1(n7088), .B2(n7087), .A(n6541), .ZN(n7086) );
  INV_X1 U8036 ( .A(n10127), .ZN(n7087) );
  NAND2_X1 U8037 ( .A1(n11453), .A2(n10154), .ZN(n10159) );
  AND4_X1 U8038 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10919) );
  AOI21_X1 U8039 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9604) );
  NOR2_X1 U8040 ( .A1(n6516), .A2(n12019), .ZN(n7070) );
  INV_X1 U8041 ( .A(n7080), .ZN(n7076) );
  NAND2_X1 U8042 ( .A1(n7073), .A2(n7077), .ZN(n7072) );
  NAND2_X1 U8043 ( .A1(n6515), .A2(n7079), .ZN(n7077) );
  AND3_X1 U8044 ( .A1(n10605), .A2(n10604), .A3(n10603), .ZN(n10943) );
  XNOR2_X1 U8045 ( .A(n11873), .B(n11871), .ZN(n11978) );
  AND3_X1 U8046 ( .A1(n10925), .A2(n10924), .A3(n10923), .ZN(n11005) );
  NAND2_X1 U8047 ( .A1(n10921), .A2(n11464), .ZN(n10925) );
  NOR2_X1 U8048 ( .A1(n11653), .A2(n7141), .ZN(n7022) );
  NAND2_X1 U8049 ( .A1(n7025), .A2(n11660), .ZN(n7023) );
  INV_X1 U8050 ( .A(n11655), .ZN(n7027) );
  INV_X1 U8051 ( .A(n12224), .ZN(n12247) );
  INV_X1 U8052 ( .A(n11929), .ZN(n12270) );
  AOI22_X1 U8053 ( .A1(n9060), .A2(n9059), .B1(n9058), .B2(n9057), .ZN(n9136)
         );
  NAND2_X1 U8054 ( .A1(n14782), .A2(n14783), .ZN(n14781) );
  NAND2_X1 U8055 ( .A1(n9696), .A2(n9695), .ZN(n9836) );
  AOI21_X1 U8056 ( .B1(n6710), .B2(n6713), .A(n6716), .ZN(n6709) );
  NAND2_X1 U8057 ( .A1(n9953), .A2(n6710), .ZN(n6703) );
  NAND2_X1 U8058 ( .A1(n10214), .A2(n10215), .ZN(n10540) );
  NOR2_X1 U8059 ( .A1(n10538), .A2(n10539), .ZN(n10709) );
  AOI21_X1 U8060 ( .B1(n12111), .B2(n14788), .A(n12110), .ZN(n6883) );
  NAND2_X1 U8061 ( .A1(n6885), .A2(n14801), .ZN(n6884) );
  XNOR2_X1 U8062 ( .A(n6887), .B(n6886), .ZN(n6885) );
  INV_X1 U8063 ( .A(n12108), .ZN(n6886) );
  OAI22_X1 U8064 ( .A1(n12107), .A2(n12106), .B1(n12105), .B2(n13209), .ZN(
        n6887) );
  NOR2_X1 U8065 ( .A1(n12093), .A2(n6831), .ZN(n6721) );
  NAND2_X1 U8066 ( .A1(n12411), .A2(n11464), .ZN(n11456) );
  NAND2_X1 U8067 ( .A1(n11263), .A2(n11262), .ZN(n12325) );
  OR2_X1 U8068 ( .A1(n11454), .A2(n11712), .ZN(n11262) );
  NAND2_X1 U8069 ( .A1(n11711), .A2(n11464), .ZN(n11263) );
  NAND2_X1 U8070 ( .A1(n11428), .A2(n11601), .ZN(n11684) );
  NAND2_X1 U8071 ( .A1(n11432), .A2(n11431), .ZN(n12329) );
  OR2_X1 U8072 ( .A1(n11454), .A2(n11430), .ZN(n11431) );
  NAND2_X1 U8073 ( .A1(n11409), .A2(n11408), .ZN(n12337) );
  NAND2_X1 U8074 ( .A1(n11406), .A2(n11464), .ZN(n11409) );
  NAND2_X1 U8075 ( .A1(n11385), .A2(n11384), .ZN(n12346) );
  OR2_X1 U8076 ( .A1(n11454), .A2(n11383), .ZN(n11384) );
  NAND2_X1 U8077 ( .A1(n11382), .A2(n11464), .ZN(n11385) );
  NAND2_X1 U8078 ( .A1(n14194), .A2(n11464), .ZN(n11276) );
  INV_X1 U8079 ( .A(n14884), .ZN(n14902) );
  INV_X1 U8080 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9218) );
  OAI21_X1 U8081 ( .B1(n11332), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U8082 ( .A1(n12427), .A2(n12426), .ZN(n6809) );
  NOR2_X1 U8083 ( .A1(n12432), .A2(n12516), .ZN(n6837) );
  AND4_X1 U8084 ( .A1(n7789), .A2(n7788), .A3(n7787), .A4(n7786), .ZN(n10738)
         );
  AND2_X1 U8085 ( .A1(n7978), .A2(n7977), .ZN(n12443) );
  NAND2_X1 U8086 ( .A1(n7953), .A2(n7952), .ZN(n12966) );
  NAND2_X1 U8087 ( .A1(n8051), .A2(n8050), .ZN(n12940) );
  OAI21_X1 U8088 ( .B1(n12821), .B2(n8023), .A(n8022), .ZN(n12802) );
  NAND2_X1 U8089 ( .A1(n12700), .A2(n8410), .ZN(n8411) );
  INV_X1 U8090 ( .A(n11718), .ZN(n11779) );
  NAND2_X1 U8091 ( .A1(n8365), .A2(n8364), .ZN(n14684) );
  NOR2_X1 U8092 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7401) );
  OAI22_X1 U8093 ( .A1(n10112), .A2(n10111), .B1(n10109), .B2(n10110), .ZN(
        n10351) );
  NAND2_X1 U8094 ( .A1(n11145), .A2(n11144), .ZN(n14087) );
  NAND2_X1 U8095 ( .A1(n11080), .A2(n11079), .ZN(n14126) );
  NAND2_X1 U8096 ( .A1(n11158), .A2(n11157), .ZN(n14083) );
  NAND2_X1 U8097 ( .A1(n10576), .A2(n10575), .ZN(n14301) );
  NAND2_X1 U8098 ( .A1(n6874), .A2(n7261), .ZN(n13644) );
  NAND2_X1 U8099 ( .A1(n7264), .A2(n6508), .ZN(n7261) );
  NAND2_X1 U8100 ( .A1(n13591), .A2(n7262), .ZN(n6874) );
  NOR2_X1 U8101 ( .A1(n13637), .A2(n13606), .ZN(n6873) );
  OR2_X1 U8102 ( .A1(n9172), .A2(P1_U3086), .ZN(n14136) );
  NOR2_X1 U8103 ( .A1(n11056), .A2(n11057), .ZN(n11055) );
  NAND2_X1 U8104 ( .A1(n8602), .A2(n7170), .ZN(n9483) );
  INV_X1 U8105 ( .A(n7171), .ZN(n7170) );
  OAI22_X1 U8106 ( .A1(n13574), .A2(n7600), .B1(n11059), .B2(n11132), .ZN(
        n7171) );
  INV_X1 U8107 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8108 ( .A1(n8623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8624) );
  AOI21_X1 U8109 ( .B1(n8481), .B2(n8480), .A(n14178), .ZN(n14978) );
  AND2_X1 U8110 ( .A1(n6790), .A2(n6818), .ZN(n14342) );
  AND2_X1 U8111 ( .A1(n6819), .A2(n8509), .ZN(n6790) );
  AND2_X1 U8112 ( .A1(n6818), .A2(n6819), .ZN(n6792) );
  NAND2_X1 U8113 ( .A1(n7124), .A2(n7123), .ZN(n7122) );
  OAI21_X1 U8114 ( .B1(n6786), .B2(n6785), .A(n6787), .ZN(n7124) );
  OR2_X1 U8115 ( .A1(n14350), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6787) );
  INV_X1 U8116 ( .A(n14345), .ZN(n6786) );
  NAND2_X1 U8117 ( .A1(n6800), .A2(n6551), .ZN(n6785) );
  NOR2_X1 U8118 ( .A1(n8515), .A2(n8516), .ZN(n14361) );
  NAND2_X1 U8119 ( .A1(n8515), .A2(n8516), .ZN(n6799) );
  INV_X1 U8120 ( .A(n7128), .ZN(n8518) );
  NAND2_X1 U8121 ( .A1(n6657), .A2(n7615), .ZN(n7613) );
  INV_X1 U8122 ( .A(n7616), .ZN(n6657) );
  NAND2_X1 U8123 ( .A1(n6659), .A2(n6658), .ZN(n7616) );
  NAND2_X1 U8124 ( .A1(n6481), .A2(n8268), .ZN(n6658) );
  NAND2_X1 U8125 ( .A1(n8219), .A2(n8267), .ZN(n6659) );
  NAND2_X1 U8126 ( .A1(n6652), .A2(n7667), .ZN(n6651) );
  INV_X1 U8127 ( .A(n7668), .ZN(n6652) );
  AOI21_X1 U8128 ( .B1(n7694), .B2(n7693), .A(n7691), .ZN(n7692) );
  NAND2_X1 U8129 ( .A1(n13434), .A2(n13433), .ZN(n13437) );
  OAI22_X1 U8130 ( .A1(n7505), .A2(n7746), .B1(n7768), .B2(n7766), .ZN(n7791)
         );
  NOR2_X1 U8131 ( .A1(n13460), .A2(n13463), .ZN(n7272) );
  INV_X1 U8132 ( .A(n13460), .ZN(n7273) );
  NAND2_X1 U8133 ( .A1(n6656), .A2(n7442), .ZN(n7833) );
  NAND2_X1 U8134 ( .A1(n7810), .A2(n7443), .ZN(n7442) );
  OAI21_X1 U8135 ( .B1(n13469), .B2(n7271), .A(n7270), .ZN(n13475) );
  AOI21_X1 U8136 ( .B1(n7271), .B2(n7270), .A(n7268), .ZN(n7267) );
  NOR2_X1 U8137 ( .A1(n6872), .A2(n13480), .ZN(n7278) );
  NAND2_X1 U8138 ( .A1(n13480), .A2(n6872), .ZN(n6871) );
  OAI22_X1 U8139 ( .A1(n13487), .A2(n7280), .B1(n7279), .B2(n13488), .ZN(
        n13493) );
  INV_X1 U8140 ( .A(n13486), .ZN(n7279) );
  NOR2_X1 U8141 ( .A1(n13489), .A2(n13486), .ZN(n7280) );
  NAND2_X1 U8142 ( .A1(n6588), .A2(n7895), .ZN(n7452) );
  NAND2_X1 U8143 ( .A1(n13500), .A2(n13503), .ZN(n7252) );
  NAND2_X1 U8144 ( .A1(n7938), .A2(n6663), .ZN(n6660) );
  NOR2_X1 U8145 ( .A1(n7495), .A2(n7497), .ZN(n7493) );
  NOR2_X1 U8146 ( .A1(n7495), .A2(n7964), .ZN(n7494) );
  AOI21_X1 U8147 ( .B1(n7249), .B2(n6495), .A(n7248), .ZN(n7247) );
  NOR2_X1 U8148 ( .A1(n8002), .A2(n8000), .ZN(n8006) );
  INV_X1 U8149 ( .A(n7501), .ZN(n7500) );
  OR2_X1 U8150 ( .A1(n8044), .A2(n8043), .ZN(n7501) );
  NAND2_X1 U8151 ( .A1(n13538), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U8152 ( .A1(n7489), .A2(n7488), .ZN(n7487) );
  NOR2_X1 U8153 ( .A1(n13558), .A2(n13556), .ZN(n7275) );
  AND2_X1 U8154 ( .A1(n7257), .A2(n13552), .ZN(n7256) );
  NAND2_X1 U8155 ( .A1(n7260), .A2(n7259), .ZN(n7257) );
  AOI21_X1 U8156 ( .B1(n6856), .B2(n6861), .A(n6854), .ZN(n6853) );
  INV_X1 U8157 ( .A(n7259), .ZN(n6854) );
  NAND2_X1 U8158 ( .A1(n12133), .A2(n7245), .ZN(n7244) );
  NAND2_X1 U8159 ( .A1(n11612), .A2(n11613), .ZN(n7245) );
  NAND2_X1 U8160 ( .A1(n11701), .A2(n6783), .ZN(n11700) );
  INV_X1 U8161 ( .A(n11699), .ZN(n6783) );
  INV_X1 U8162 ( .A(n10594), .ZN(n7227) );
  INV_X1 U8163 ( .A(n8724), .ZN(n7016) );
  INV_X1 U8164 ( .A(n7015), .ZN(n7014) );
  OAI21_X1 U8165 ( .B1(n8729), .B2(n7016), .A(n10600), .ZN(n7015) );
  AND2_X1 U8166 ( .A1(n7017), .A2(n6773), .ZN(n6772) );
  NAND2_X1 U8167 ( .A1(n6774), .A2(n8708), .ZN(n6773) );
  NOR2_X1 U8168 ( .A1(n6492), .A2(n7018), .ZN(n7017) );
  NAND4_X1 U8169 ( .A1(n8285), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(n8252)
         );
  AND2_X1 U8170 ( .A1(n8215), .A2(n8209), .ZN(n8210) );
  AND2_X1 U8171 ( .A1(n8284), .A2(n8412), .ZN(n7355) );
  INV_X1 U8172 ( .A(n12784), .ZN(n8337) );
  NAND2_X1 U8173 ( .A1(n6573), .A2(n8408), .ZN(n7219) );
  INV_X1 U8174 ( .A(n7219), .ZN(n7216) );
  AOI21_X1 U8175 ( .B1(n7337), .B2(n7334), .A(n7333), .ZN(n7332) );
  INV_X1 U8176 ( .A(n8174), .ZN(n7333) );
  INV_X1 U8177 ( .A(n7339), .ZN(n7334) );
  NAND2_X1 U8178 ( .A1(n8093), .A2(n8092), .ZN(n8108) );
  INV_X1 U8179 ( .A(n11842), .ZN(n7085) );
  NAND2_X1 U8180 ( .A1(n14245), .A2(n11477), .ZN(n11645) );
  NAND2_X1 U8181 ( .A1(n9285), .A2(n6539), .ZN(n9663) );
  OAI21_X1 U8182 ( .B1(n9849), .B2(n14961), .A(n9845), .ZN(n9954) );
  NAND2_X1 U8183 ( .A1(n10540), .A2(n10541), .ZN(n10722) );
  XNOR2_X1 U8184 ( .A(n12037), .B(n6882), .ZN(n11022) );
  NAND2_X1 U8185 ( .A1(n11020), .A2(n11021), .ZN(n12037) );
  NAND2_X1 U8186 ( .A1(n12056), .A2(n12057), .ZN(n12076) );
  NAND2_X1 U8187 ( .A1(n11700), .A2(n6782), .ZN(n11787) );
  NAND2_X1 U8188 ( .A1(n11701), .A2(n11702), .ZN(n6782) );
  INV_X1 U8189 ( .A(n11524), .ZN(n7139) );
  OAI21_X1 U8190 ( .B1(n7139), .B2(n11623), .A(n11630), .ZN(n6824) );
  NAND2_X1 U8191 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n7241), .ZN(n7240) );
  NOR2_X1 U8192 ( .A1(n11248), .A2(n6754), .ZN(n6753) );
  INV_X1 U8193 ( .A(n10893), .ZN(n6754) );
  AND2_X1 U8194 ( .A1(n6530), .A2(n8689), .ZN(n7157) );
  AND2_X1 U8195 ( .A1(n6669), .A2(n6668), .ZN(n6834) );
  NOR2_X1 U8196 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n6669) );
  NOR2_X1 U8197 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n6668) );
  NAND2_X1 U8198 ( .A1(n6760), .A2(n6759), .ZN(n9756) );
  AOI21_X1 U8199 ( .B1(n6762), .B2(n6764), .A(n6635), .ZN(n6759) );
  NAND2_X1 U8200 ( .A1(n11331), .A2(n6762), .ZN(n6760) );
  INV_X1 U8201 ( .A(n8768), .ZN(n7202) );
  NAND2_X1 U8202 ( .A1(n8753), .A2(n6772), .ZN(n6770) );
  INV_X1 U8203 ( .A(n7021), .ZN(n7020) );
  OAI21_X1 U8204 ( .B1(n7203), .B2(n6492), .A(n8718), .ZN(n7021) );
  NAND2_X1 U8205 ( .A1(n6772), .A2(n6775), .ZN(n6769) );
  INV_X1 U8206 ( .A(n8708), .ZN(n6775) );
  OR2_X1 U8207 ( .A1(n8715), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U8208 ( .A1(n6523), .A2(n7394), .ZN(n7393) );
  NAND2_X1 U8209 ( .A1(n10251), .A2(n6523), .ZN(n7392) );
  AND2_X1 U8210 ( .A1(n8153), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8154) );
  INV_X1 U8211 ( .A(n8154), .ZN(n8193) );
  AOI21_X1 U8212 ( .B1(n6559), .B2(n12752), .A(n12743), .ZN(n7303) );
  NOR2_X1 U8213 ( .A1(n7305), .A2(n12757), .ZN(n7304) );
  INV_X1 U8214 ( .A(n7307), .ZN(n7305) );
  NAND2_X1 U8215 ( .A1(n12783), .A2(n12791), .ZN(n7307) );
  OR2_X1 U8216 ( .A1(n12771), .A2(n12784), .ZN(n7306) );
  AND2_X1 U8217 ( .A1(n8052), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U8218 ( .A1(n6526), .A2(n6500), .ZN(n6917) );
  NAND2_X1 U8219 ( .A1(n6736), .A2(n8404), .ZN(n6735) );
  INV_X1 U8220 ( .A(n8403), .ZN(n6736) );
  INV_X1 U8221 ( .A(n8404), .ZN(n6737) );
  OR2_X1 U8222 ( .A1(n7993), .A2(n7992), .ZN(n8016) );
  NOR2_X1 U8223 ( .A1(n7293), .A2(n6896), .ZN(n6895) );
  NAND2_X1 U8224 ( .A1(n9073), .A2(n8271), .ZN(n8272) );
  AND2_X1 U8225 ( .A1(n7526), .A2(n8385), .ZN(n7211) );
  NOR2_X1 U8226 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7548) );
  INV_X1 U8227 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7946) );
  INV_X1 U8228 ( .A(n13068), .ZN(n7485) );
  INV_X1 U8229 ( .A(n13417), .ZN(n7435) );
  NAND2_X1 U8230 ( .A1(n6532), .A2(n10353), .ZN(n6945) );
  NAND2_X1 U8231 ( .A1(n13561), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U8232 ( .A1(n6490), .A2(n6844), .ZN(n6842) );
  OR2_X1 U8233 ( .A1(n13429), .A2(n13587), .ZN(n13430) );
  NOR2_X1 U8234 ( .A1(n13923), .A2(n13940), .ZN(n7108) );
  AND2_X1 U8235 ( .A1(n6528), .A2(n13504), .ZN(n7379) );
  INV_X1 U8236 ( .A(n7189), .ZN(n6692) );
  INV_X1 U8237 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U8238 ( .A1(n10195), .A2(n13472), .ZN(n7110) );
  INV_X1 U8239 ( .A(n9990), .ZN(n7175) );
  AND2_X1 U8240 ( .A1(n14405), .A2(n14475), .ZN(n9982) );
  INV_X1 U8241 ( .A(n9814), .ZN(n6690) );
  NAND2_X1 U8242 ( .A1(n6689), .A2(n9814), .ZN(n6688) );
  INV_X1 U8243 ( .A(n9813), .ZN(n6689) );
  NOR2_X1 U8244 ( .A1(n14058), .A2(n7112), .ZN(n7111) );
  INV_X1 U8245 ( .A(n7113), .ZN(n7112) );
  INV_X1 U8246 ( .A(n7108), .ZN(n13924) );
  AND2_X1 U8247 ( .A1(n10867), .A2(n7116), .ZN(n14003) );
  NOR2_X1 U8248 ( .A1(n14132), .A2(n7118), .ZN(n7116) );
  NAND2_X1 U8249 ( .A1(n10867), .A2(n14325), .ZN(n10987) );
  NOR2_X1 U8250 ( .A1(n8166), .A2(n7340), .ZN(n7339) );
  INV_X1 U8251 ( .A(n8146), .ZN(n7340) );
  AOI21_X1 U8252 ( .B1(n7339), .B2(n8147), .A(n7338), .ZN(n7337) );
  INV_X1 U8253 ( .A(n8165), .ZN(n7338) );
  INV_X1 U8254 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U8255 ( .A(n8108), .B(SI_24_), .ZN(n8105) );
  NAND2_X1 U8256 ( .A1(n6956), .A2(n8048), .ZN(n6955) );
  NAND2_X1 U8257 ( .A1(n6959), .A2(n6499), .ZN(n6956) );
  INV_X1 U8258 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8537) );
  INV_X1 U8259 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8534) );
  INV_X1 U8260 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8533) );
  INV_X1 U8261 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8530) );
  AND2_X1 U8262 ( .A1(n7967), .A2(n7945), .ZN(n7965) );
  AND2_X1 U8263 ( .A1(n7054), .A2(n7053), .ZN(n6969) );
  NAND2_X1 U8264 ( .A1(n7837), .A2(n7056), .ZN(n7051) );
  NAND2_X1 U8265 ( .A1(n7818), .A2(n8769), .ZN(n7838) );
  NAND2_X1 U8266 ( .A1(n6967), .A2(n7321), .ZN(n7814) );
  AOI21_X1 U8267 ( .B1(n7323), .B2(n7325), .A(n6576), .ZN(n7321) );
  NAND2_X1 U8268 ( .A1(n6953), .A2(n7728), .ZN(n7749) );
  OAI21_X1 U8269 ( .B1(n6484), .B2(P2_DATAO_REG_5__SCAN_IN), .A(n6817), .ZN(
        n7698) );
  NAND2_X1 U8270 ( .A1(n6484), .A2(n8759), .ZN(n6817) );
  INV_X1 U8271 ( .A(n7657), .ZN(n7654) );
  OAI21_X1 U8272 ( .B1(n6483), .B2(n7600), .A(n7599), .ZN(n7657) );
  NAND2_X1 U8273 ( .A1(n6483), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7599) );
  INV_X1 U8274 ( .A(n7038), .ZN(n6993) );
  NOR2_X1 U8275 ( .A1(n8421), .A2(n8420), .ZN(n8423) );
  AND2_X1 U8276 ( .A1(n8419), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n8420) );
  INV_X1 U8277 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8422) );
  XNOR2_X1 U8278 ( .A(n6789), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n8469) );
  NOR2_X1 U8279 ( .A1(n8431), .A2(n8430), .ZN(n8468) );
  INV_X1 U8280 ( .A(n10066), .ZN(n7090) );
  NAND2_X1 U8281 ( .A1(n11846), .A2(n12156), .ZN(n7080) );
  NAND2_X1 U8282 ( .A1(n7068), .A2(n11813), .ZN(n11909) );
  INV_X1 U8283 ( .A(n11911), .ZN(n7068) );
  NAND2_X1 U8284 ( .A1(n9453), .A2(n9450), .ZN(n9511) );
  NAND2_X1 U8285 ( .A1(n11620), .A2(n7147), .ZN(n7146) );
  NOR2_X1 U8286 ( .A1(n11481), .A2(n7148), .ZN(n7147) );
  INV_X1 U8287 ( .A(n11645), .ZN(n11617) );
  AND4_X1 U8288 ( .A1(n11259), .A2(n11258), .A3(n11257), .A4(n11256), .ZN(
        n11795) );
  AND4_X1 U8289 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11961) );
  NAND2_X1 U8290 ( .A1(n6804), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9377) );
  OAI21_X1 U8291 ( .B1(n12069), .B2(n9633), .A(n6720), .ZN(n6719) );
  NAND2_X1 U8292 ( .A1(n12069), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U8293 ( .A1(n9236), .A2(n9237), .ZN(n9238) );
  XNOR2_X1 U8294 ( .A(n9663), .B(n10018), .ZN(n9286) );
  AOI21_X1 U8295 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(n14794) );
  NAND2_X1 U8296 ( .A1(n9705), .A2(n9706), .ZN(n9707) );
  NAND2_X1 U8297 ( .A1(n9699), .A2(n9700), .ZN(n9701) );
  NAND2_X1 U8298 ( .A1(n9961), .A2(n9962), .ZN(n9963) );
  NAND2_X1 U8299 ( .A1(n10218), .A2(n10219), .ZN(n10222) );
  XNOR2_X1 U8300 ( .A(n10722), .B(n11268), .ZN(n10542) );
  NAND2_X1 U8301 ( .A1(n11012), .A2(n11011), .ZN(n12047) );
  NAND2_X1 U8302 ( .A1(n12054), .A2(n6889), .ZN(n12083) );
  NAND2_X1 U8303 ( .A1(n14202), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U8304 ( .A(n12076), .B(n6888), .ZN(n12075) );
  OR2_X1 U8305 ( .A1(n12333), .A2(n12155), .ZN(n11601) );
  NOR2_X1 U8306 ( .A1(n6815), .A2(n6814), .ZN(n6813) );
  INV_X1 U8307 ( .A(n11600), .ZN(n6815) );
  INV_X1 U8308 ( .A(n12147), .ZN(n6814) );
  INV_X1 U8309 ( .A(n12138), .ZN(n12148) );
  AND2_X1 U8310 ( .A1(n11601), .A2(n11600), .ZN(n12138) );
  INV_X1 U8311 ( .A(n12177), .ZN(n12140) );
  NAND2_X1 U8312 ( .A1(n6670), .A2(n11486), .ZN(n12175) );
  OR2_X1 U8313 ( .A1(n6503), .A2(n6599), .ZN(n7414) );
  INV_X1 U8314 ( .A(n11678), .ZN(n12174) );
  INV_X1 U8315 ( .A(SI_22_), .ZN(n11383) );
  AND2_X1 U8316 ( .A1(n6825), .A2(n12250), .ZN(n6677) );
  INV_X1 U8317 ( .A(n7154), .ZN(n6825) );
  INV_X1 U8318 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13126) );
  INV_X1 U8319 ( .A(n11669), .ZN(n12250) );
  INV_X1 U8320 ( .A(SI_16_), .ZN(n11307) );
  AOI21_X1 U8321 ( .B1(n7406), .B2(n7408), .A(n6614), .ZN(n7405) );
  INV_X1 U8322 ( .A(SI_15_), .ZN(n11287) );
  NOR2_X1 U8323 ( .A1(n14234), .A2(n10948), .ZN(n10949) );
  NAND2_X1 U8324 ( .A1(n11464), .A2(n10937), .ZN(n10938) );
  INV_X1 U8325 ( .A(n11632), .ZN(n10926) );
  INV_X1 U8326 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10372) );
  INV_X1 U8327 ( .A(n11538), .ZN(n14826) );
  NOR2_X1 U8328 ( .A1(n11624), .A2(n7420), .ZN(n7419) );
  INV_X1 U8329 ( .A(n10369), .ZN(n7420) );
  NAND2_X1 U8330 ( .A1(n10360), .A2(n11533), .ZN(n10918) );
  NAND2_X1 U8331 ( .A1(n7137), .A2(n11524), .ZN(n14831) );
  NAND2_X1 U8332 ( .A1(n10160), .A2(n11623), .ZN(n7137) );
  NAND2_X1 U8333 ( .A1(n11453), .A2(n9599), .ZN(n9602) );
  AND2_X1 U8334 ( .A1(n14875), .A2(n9770), .ZN(n9772) );
  NOR2_X1 U8335 ( .A1(n14886), .A2(n6672), .ZN(n14933) );
  INV_X1 U8336 ( .A(n9364), .ZN(n11031) );
  NOR2_X1 U8337 ( .A1(n13573), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7029) );
  NOR2_X2 U8338 ( .A1(n9009), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U8339 ( .A1(n8694), .A2(n6510), .ZN(n8688) );
  INV_X1 U8340 ( .A(n11008), .ZN(n8694) );
  INV_X1 U8341 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10596) );
  XNOR2_X1 U8342 ( .A(n8699), .B(n8698), .ZN(n9020) );
  INV_X1 U8343 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8698) );
  OAI21_X1 U8344 ( .B1(n9017), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8699) );
  OR2_X1 U8345 ( .A1(n9347), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U8346 ( .A(n9019), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9466) );
  OR2_X1 U8347 ( .A1(n11305), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U8348 ( .A1(n6758), .A2(n6811), .ZN(n9215) );
  NAND2_X1 U8349 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n6812), .ZN(n6811) );
  INV_X1 U8350 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U8351 ( .A1(n9113), .A2(n9112), .ZN(n11286) );
  AOI21_X1 U8352 ( .B1(n9111), .B2(n6767), .A(n6629), .ZN(n6765) );
  INV_X1 U8353 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n10711) );
  OAI21_X1 U8354 ( .B1(n7012), .B2(n7201), .A(n6780), .ZN(n9105) );
  INV_X1 U8355 ( .A(n6781), .ZN(n6780) );
  OAI21_X1 U8356 ( .B1(n7011), .B2(n7201), .A(n7198), .ZN(n6781) );
  AOI21_X1 U8357 ( .B1(n7200), .B2(n7202), .A(n6579), .ZN(n7198) );
  NOR2_X1 U8358 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7130) );
  INV_X1 U8359 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8670) );
  XNOR2_X1 U8360 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8785) );
  NAND2_X1 U8361 ( .A1(n8742), .A2(n8703), .ZN(n8782) );
  AND2_X1 U8362 ( .A1(n8833), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8743) );
  XNOR2_X1 U8363 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8744) );
  NAND2_X1 U8364 ( .A1(n8744), .A2(n8743), .ZN(n8742) );
  INV_X1 U8365 ( .A(n9333), .ZN(n7009) );
  NOR2_X1 U8366 ( .A1(n8034), .A2(n12464), .ZN(n8052) );
  OR2_X1 U8367 ( .A1(n8016), .A2(n12524), .ZN(n8034) );
  AND2_X1 U8368 ( .A1(n10084), .A2(n9581), .ZN(n6997) );
  CLKBUF_X1 U8369 ( .A(n12486), .Z(n12499) );
  NOR2_X1 U8370 ( .A1(n7785), .A2(n7784), .ZN(n7804) );
  OR2_X1 U8371 ( .A1(n12519), .A2(n11734), .ZN(n12518) );
  NAND2_X1 U8372 ( .A1(n12462), .A2(n6988), .ZN(n11741) );
  NAND2_X1 U8373 ( .A1(n11736), .A2(n6989), .ZN(n6988) );
  INV_X1 U8374 ( .A(n11737), .ZN(n6989) );
  NAND2_X1 U8375 ( .A1(n6493), .A2(n7397), .ZN(n7395) );
  NAND2_X1 U8376 ( .A1(n12507), .A2(n6560), .ZN(n12440) );
  NAND2_X1 U8377 ( .A1(n9320), .A2(n9319), .ZN(n9334) );
  OR2_X1 U8378 ( .A1(n7891), .A2(n7890), .ZN(n7913) );
  INV_X1 U8379 ( .A(n8231), .ZN(n7484) );
  OR2_X1 U8380 ( .A1(n14592), .A2(n14591), .ZN(n14593) );
  AND2_X1 U8381 ( .A1(n8154), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8371) );
  AND2_X1 U8382 ( .A1(n8169), .A2(n8168), .ZN(n8373) );
  INV_X1 U8383 ( .A(n6823), .ZN(n12714) );
  AND4_X1 U8384 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), .ZN(n12728)
         );
  NOR2_X1 U8385 ( .A1(n12922), .A2(n7099), .ZN(n7097) );
  NAND2_X1 U8386 ( .A1(n12793), .A2(n7101), .ZN(n12762) );
  NAND2_X1 U8387 ( .A1(n7306), .A2(n7307), .ZN(n12756) );
  AND2_X1 U8388 ( .A1(n12755), .A2(n12754), .ZN(n12767) );
  NAND2_X1 U8389 ( .A1(n12793), .A2(n12783), .ZN(n12779) );
  NAND2_X1 U8390 ( .A1(n6916), .A2(n6917), .ZN(n12771) );
  OR2_X1 U8391 ( .A1(n12833), .A2(n12951), .ZN(n12823) );
  NAND2_X1 U8392 ( .A1(n12850), .A2(n12837), .ZN(n12833) );
  NOR2_X1 U8393 ( .A1(n7913), .A2(n11775), .ZN(n7933) );
  NOR2_X1 U8394 ( .A1(n7849), .A2(n7848), .ZN(n7869) );
  AND2_X1 U8395 ( .A1(n7313), .A2(n7312), .ZN(n10756) );
  AND2_X1 U8396 ( .A1(n7313), .A2(n6536), .ZN(n10755) );
  OR2_X1 U8397 ( .A1(n10750), .A2(n12580), .ZN(n7213) );
  AND4_X1 U8398 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n10758)
         );
  NAND2_X1 U8399 ( .A1(n7195), .A2(n6556), .ZN(n9647) );
  OR2_X1 U8400 ( .A1(n7758), .A2(n7757), .ZN(n7785) );
  OR2_X1 U8401 ( .A1(n7735), .A2(n9338), .ZN(n7758) );
  NAND2_X1 U8402 ( .A1(n7299), .A2(n7301), .ZN(n7297) );
  INV_X1 U8403 ( .A(n10782), .ZN(n7096) );
  NOR2_X2 U8404 ( .A1(n8267), .A2(n10475), .ZN(n10783) );
  NAND2_X1 U8405 ( .A1(n10467), .A2(n8307), .ZN(n10304) );
  INV_X1 U8406 ( .A(n9075), .ZN(n12456) );
  NAND2_X1 U8407 ( .A1(n9073), .A2(n8370), .ZN(n10475) );
  INV_X1 U8408 ( .A(n12971), .ZN(n12865) );
  NAND2_X1 U8409 ( .A1(n9066), .A2(n8302), .ZN(n12773) );
  INV_X1 U8410 ( .A(n8373), .ZN(n12904) );
  INV_X1 U8411 ( .A(n8408), .ZN(n7218) );
  NAND2_X1 U8412 ( .A1(n7290), .A2(n7291), .ZN(n12877) );
  NAND2_X1 U8413 ( .A1(n6897), .A2(n6896), .ZN(n7291) );
  AND2_X1 U8414 ( .A1(n7912), .A2(n7911), .ZN(n11718) );
  OR2_X1 U8415 ( .A1(n9068), .A2(n9067), .ZN(n14756) );
  AND2_X1 U8416 ( .A1(n6485), .A2(n14740), .ZN(n14720) );
  INV_X1 U8417 ( .A(n14756), .ZN(n14738) );
  INV_X1 U8418 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7284) );
  NOR2_X2 U8419 ( .A1(n7542), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8290) );
  INV_X1 U8420 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7969) );
  OR2_X1 U8421 ( .A1(n7949), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n7968) );
  INV_X1 U8422 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7885) );
  INV_X1 U8423 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7864) );
  INV_X1 U8424 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6890) );
  INV_X1 U8425 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U8426 ( .A1(n10179), .A2(n10178), .ZN(n10400) );
  OR2_X1 U8427 ( .A1(n8761), .A2(n9977), .ZN(n6702) );
  NAND2_X1 U8428 ( .A1(n7474), .A2(n7471), .ZN(n7470) );
  INV_X1 U8429 ( .A(n7476), .ZN(n7471) );
  OR2_X1 U8430 ( .A1(n13308), .A2(n13307), .ZN(n7477) );
  NOR2_X1 U8431 ( .A1(n7472), .A2(n7466), .ZN(n7465) );
  INV_X1 U8432 ( .A(n13337), .ZN(n7466) );
  NAND2_X1 U8433 ( .A1(n7473), .A2(n7474), .ZN(n7472) );
  INV_X1 U8434 ( .A(n13309), .ZN(n7473) );
  NOR2_X1 U8435 ( .A1(n6925), .A2(n9781), .ZN(n6924) );
  OR2_X1 U8436 ( .A1(n9534), .A2(n13063), .ZN(n9155) );
  NAND2_X1 U8437 ( .A1(n9157), .A2(n6936), .ZN(n9398) );
  NAND2_X1 U8438 ( .A1(n6938), .A2(n6937), .ZN(n6936) );
  INV_X1 U8439 ( .A(n13062), .ZN(n6937) );
  OR2_X1 U8440 ( .A1(n11107), .A2(n13130), .ZN(n11116) );
  OR2_X1 U8441 ( .A1(n11116), .A2(n13379), .ZN(n11125) );
  INV_X1 U8442 ( .A(n6951), .ZN(n6950) );
  OAI21_X1 U8443 ( .B1(n6522), .B2(n6952), .A(n13377), .ZN(n6951) );
  INV_X1 U8444 ( .A(n13061), .ZN(n6952) );
  NAND2_X1 U8445 ( .A1(n13384), .A2(n13385), .ZN(n13383) );
  NOR2_X1 U8446 ( .A1(n7445), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U8447 ( .A1(n7448), .A2(n7447), .ZN(n7445) );
  NAND2_X1 U8448 ( .A1(n6944), .A2(n6941), .ZN(n6940) );
  INV_X1 U8449 ( .A(n10350), .ZN(n6941) );
  XNOR2_X1 U8450 ( .A(n9159), .B(n13022), .ZN(n9222) );
  OAI22_X1 U8451 ( .A1(n13431), .A2(n13063), .B1(n9158), .B2(n13064), .ZN(
        n9159) );
  OAI21_X1 U8452 ( .B1(n9730), .B2(n6935), .A(n6931), .ZN(n6928) );
  NAND2_X1 U8453 ( .A1(n14288), .A2(n13027), .ZN(n7439) );
  NAND2_X1 U8454 ( .A1(n7263), .A2(n13593), .ZN(n7262) );
  AND2_X1 U8455 ( .A1(n6982), .A2(n6981), .ZN(n9413) );
  NAND2_X1 U8456 ( .A1(n8869), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6981) );
  NOR2_X1 U8457 ( .A1(n9194), .A2(n6971), .ZN(n13702) );
  NOR2_X1 U8458 ( .A1(n6972), .A2(n8970), .ZN(n6971) );
  INV_X1 U8459 ( .A(n9979), .ZN(n6972) );
  NAND2_X1 U8460 ( .A1(n13702), .A2(n13701), .ZN(n13700) );
  NAND2_X1 U8461 ( .A1(n13700), .A2(n6970), .ZN(n13715) );
  OR2_X1 U8462 ( .A1(n13709), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8463 ( .A1(n13715), .A2(n13716), .ZN(n13714) );
  NOR2_X1 U8464 ( .A1(n9419), .A2(n6978), .ZN(n9422) );
  AND2_X1 U8465 ( .A1(n10510), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8466 ( .A1(n9422), .A2(n9421), .ZN(n9553) );
  NAND2_X1 U8467 ( .A1(n9553), .A2(n6977), .ZN(n9554) );
  OR2_X1 U8468 ( .A1(n10574), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8469 ( .A1(n9554), .A2(n9555), .ZN(n9866) );
  NOR2_X1 U8470 ( .A1(n9943), .A2(n6985), .ZN(n9944) );
  AND2_X1 U8471 ( .A1(n10855), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U8472 ( .A1(n9944), .A2(n9945), .ZN(n10627) );
  NAND2_X1 U8473 ( .A1(n10627), .A2(n6984), .ZN(n10629) );
  OR2_X1 U8474 ( .A1(n10970), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U8475 ( .A1(n8539), .A2(n8757), .ZN(n9661) );
  NAND2_X1 U8476 ( .A1(n7163), .A2(n11197), .ZN(n7162) );
  INV_X1 U8477 ( .A(n13793), .ZN(n7160) );
  INV_X1 U8478 ( .A(n13795), .ZN(n13801) );
  NAND2_X1 U8479 ( .A1(n13820), .A2(n6801), .ZN(n11206) );
  NOR2_X1 U8480 ( .A1(n13631), .A2(n7164), .ZN(n6801) );
  NAND2_X1 U8481 ( .A1(n13880), .A2(n7115), .ZN(n13840) );
  OAI21_X1 U8482 ( .B1(n14065), .B2(n13824), .A(n13823), .ZN(n6682) );
  NAND2_X1 U8483 ( .A1(n11177), .A2(n11176), .ZN(n13839) );
  NAND2_X1 U8484 ( .A1(n13849), .A2(n13831), .ZN(n11185) );
  NAND2_X1 U8485 ( .A1(n13880), .A2(n13855), .ZN(n13857) );
  OR2_X1 U8486 ( .A1(n13909), .A2(n14087), .ZN(n13881) );
  AND2_X1 U8487 ( .A1(n13897), .A2(n11154), .ZN(n13874) );
  NAND2_X1 U8488 ( .A1(n7108), .A2(n13915), .ZN(n13909) );
  NOR2_X1 U8489 ( .A1(n14094), .A2(n13651), .ZN(n11229) );
  INV_X1 U8490 ( .A(n13876), .ZN(n13388) );
  AOI21_X1 U8491 ( .B1(n7182), .B2(n7181), .A(n6569), .ZN(n7180) );
  INV_X1 U8492 ( .A(n11120), .ZN(n7181) );
  NAND2_X1 U8493 ( .A1(n13953), .A2(n14108), .ZN(n13940) );
  NAND2_X1 U8494 ( .A1(n11092), .A2(n11091), .ZN(n13972) );
  NOR2_X1 U8495 ( .A1(n11083), .A2(n11082), .ZN(n11093) );
  AOI21_X1 U8496 ( .B1(n6728), .B2(n13626), .A(n6726), .ZN(n6725) );
  NAND2_X1 U8497 ( .A1(n13995), .A2(n6728), .ZN(n6727) );
  INV_X1 U8498 ( .A(n11220), .ZN(n6726) );
  OR2_X1 U8499 ( .A1(n10977), .A2(n10976), .ZN(n11083) );
  NAND2_X1 U8500 ( .A1(n10867), .A2(n7120), .ZN(n14012) );
  AOI21_X1 U8501 ( .B1(n6494), .B2(n7169), .A(n6570), .ZN(n7166) );
  NAND2_X1 U8502 ( .A1(n10794), .A2(n6494), .ZN(n7165) );
  OR2_X1 U8503 ( .A1(n13490), .A2(n13659), .ZN(n10858) );
  NOR2_X1 U8504 ( .A1(n10578), .A2(n10577), .ZN(n10796) );
  OR2_X1 U8505 ( .A1(n10518), .A2(n10517), .ZN(n10578) );
  AND2_X1 U8506 ( .A1(n10807), .A2(n14216), .ZN(n10867) );
  NOR2_X1 U8507 ( .A1(n10524), .A2(n13482), .ZN(n10588) );
  AND2_X1 U8508 ( .A1(n10588), .A2(n14331), .ZN(n10807) );
  INV_X1 U8509 ( .A(n13620), .ZN(n10805) );
  NAND2_X1 U8510 ( .A1(n7357), .A2(n14393), .ZN(n6750) );
  NAND2_X1 U8511 ( .A1(n7110), .A2(n7109), .ZN(n10524) );
  INV_X1 U8512 ( .A(n7110), .ZN(n10399) );
  OR2_X1 U8513 ( .A1(n9923), .A2(n9922), .ZN(n9992) );
  OR2_X1 U8514 ( .A1(n9992), .A2(n9991), .ZN(n10179) );
  INV_X1 U8515 ( .A(n14484), .ZN(n10192) );
  OR2_X1 U8516 ( .A1(n14427), .A2(n13608), .ZN(n14428) );
  NAND2_X1 U8517 ( .A1(n9479), .A2(n6747), .ZN(n14427) );
  NAND2_X1 U8518 ( .A1(n9473), .A2(n13446), .ZN(n8629) );
  INV_X1 U8519 ( .A(n9471), .ZN(n13610) );
  NAND2_X1 U8520 ( .A1(n13610), .A2(n9474), .ZN(n9473) );
  NAND2_X1 U8521 ( .A1(n8663), .A2(n9163), .ZN(n14421) );
  INV_X1 U8522 ( .A(n14076), .ZN(n14429) );
  INV_X1 U8523 ( .A(n7359), .ZN(n10516) );
  AOI21_X1 U8524 ( .B1(n7367), .B2(n7364), .A(n6496), .ZN(n7359) );
  NOR2_X2 U8525 ( .A1(n9166), .A2(n9165), .ZN(n14499) );
  INV_X1 U8526 ( .A(n14499), .ZN(n14512) );
  OR2_X1 U8527 ( .A1(n8818), .A2(P1_U3086), .ZN(n8808) );
  XNOR2_X1 U8528 ( .A(n8182), .B(n8181), .ZN(n12992) );
  XNOR2_X1 U8529 ( .A(n8185), .B(n8184), .ZN(n13001) );
  INV_X1 U8530 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8573) );
  XNOR2_X1 U8531 ( .A(n8538), .B(P1_IR_REG_23__SCAN_IN), .ZN(n8818) );
  OAI21_X1 U8532 ( .B1(n8623), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U8533 ( .A1(n6961), .A2(n7041), .ZN(n8049) );
  NAND2_X1 U8534 ( .A1(n6578), .A2(n7343), .ZN(n6961) );
  INV_X1 U8535 ( .A(n7506), .ZN(n7386) );
  INV_X1 U8536 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U8537 ( .A1(n7045), .A2(n8012), .ZN(n8030) );
  NAND2_X1 U8538 ( .A1(n7040), .A2(n11361), .ZN(n8031) );
  OAI21_X1 U8539 ( .B1(n7837), .B2(n7350), .A(n7347), .ZN(n7882) );
  OR2_X1 U8540 ( .A1(n8814), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8822) );
  XNOR2_X1 U8541 ( .A(n7772), .B(n7770), .ZN(n10187) );
  NAND2_X1 U8542 ( .A1(n6484), .A2(n8733), .ZN(n6839) );
  AND2_X1 U8543 ( .A1(n6793), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8475) );
  INV_X1 U8544 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n8476) );
  AOI21_X1 U8545 ( .B1(n6827), .B2(n8475), .A(n7121), .ZN(n8472) );
  AND2_X1 U8546 ( .A1(n8418), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U8547 ( .A(n8419), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U8548 ( .A(n8469), .B(n7129), .ZN(n8470) );
  XNOR2_X1 U8549 ( .A(n8486), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n8487) );
  NOR2_X1 U8550 ( .A1(n8427), .A2(n8426), .ZN(n8490) );
  NAND2_X1 U8551 ( .A1(n8496), .A2(n8497), .ZN(n8498) );
  OAI21_X1 U8552 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n8435), .A(n8434), .ZN(
        n8466) );
  OAI21_X1 U8553 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n8441), .A(n8440), .ZN(
        n8461) );
  AOI21_X1 U8554 ( .B1(n14223), .B2(n14222), .A(n6565), .ZN(n7128) );
  AOI21_X1 U8555 ( .B1(n7066), .B2(n11912), .A(n6623), .ZN(n7065) );
  AND2_X1 U8556 ( .A1(n10821), .A2(n10814), .ZN(n7094) );
  AND2_X1 U8557 ( .A1(n10815), .A2(n10814), .ZN(n10822) );
  AND3_X1 U8558 ( .A1(n10820), .A2(n10819), .A3(n10818), .ZN(n10945) );
  NAND2_X1 U8559 ( .A1(n11453), .A2(n10816), .ZN(n10820) );
  NAND2_X1 U8560 ( .A1(n11453), .A2(n10361), .ZN(n10364) );
  OR2_X1 U8561 ( .A1(n9605), .A2(n8908), .ZN(n8909) );
  NAND2_X1 U8562 ( .A1(n11957), .A2(n11842), .ZN(n11902) );
  NAND2_X1 U8563 ( .A1(n11826), .A2(n11825), .ZN(n11932) );
  NAND2_X1 U8564 ( .A1(n11453), .A2(n10003), .ZN(n10007) );
  AND4_X1 U8565 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n14819) );
  NAND2_X1 U8566 ( .A1(n11881), .A2(n11839), .ZN(n11959) );
  NAND2_X1 U8567 ( .A1(n11959), .A2(n11958), .ZN(n11957) );
  NAND2_X1 U8568 ( .A1(n11909), .A2(n11817), .ZN(n11970) );
  INV_X1 U8569 ( .A(n14807), .ZN(n11913) );
  OR2_X1 U8570 ( .A1(n9458), .A2(n11659), .ZN(n12009) );
  OR2_X1 U8571 ( .A1(n9458), .A2(n9392), .ZN(n11988) );
  NAND2_X1 U8572 ( .A1(n7091), .A2(n10060), .ZN(n10067) );
  NAND2_X1 U8573 ( .A1(n7091), .A2(n7088), .ZN(n10232) );
  CLKBUF_X1 U8574 ( .A(n12003), .Z(n12015) );
  INV_X1 U8575 ( .A(n12124), .ZN(n11998) );
  INV_X1 U8576 ( .A(n14818), .ZN(n14237) );
  INV_X1 U8577 ( .A(n10919), .ZN(n14809) );
  OR2_X1 U8578 ( .A1(n11466), .A2(n14931), .ZN(n10026) );
  INV_X1 U8579 ( .A(n14833), .ZN(n14854) );
  INV_X1 U8580 ( .A(n10131), .ZN(n12029) );
  OR2_X1 U8581 ( .A1(n11468), .A2(n9776), .ZN(n9518) );
  NAND4_X2 U8582 ( .A1(n9390), .A2(n9387), .A3(n9388), .A4(n9389), .ZN(n12030)
         );
  OR2_X1 U8583 ( .A1(n9605), .A2(n9386), .ZN(n9387) );
  OR2_X1 U8584 ( .A1(n11468), .A2(n9385), .ZN(n9390) );
  OR2_X1 U8585 ( .A1(n9368), .A2(n12404), .ZN(n12031) );
  NAND2_X1 U8586 ( .A1(n14792), .A2(n6719), .ZN(n9189) );
  AOI22_X1 U8587 ( .A1(n9234), .A2(n9233), .B1(n9600), .B2(n9232), .ZN(n9280)
         );
  INV_X1 U8588 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U8589 ( .A1(n9669), .A2(n9670), .ZN(n14782) );
  OAI21_X1 U8590 ( .B1(n14794), .B2(n9687), .A(n9686), .ZN(n9694) );
  NAND2_X1 U8591 ( .A1(n9694), .A2(n9693), .ZN(n9696) );
  AND2_X1 U8592 ( .A1(n6715), .A2(n6714), .ZN(n10209) );
  NAND2_X1 U8593 ( .A1(n10205), .A2(n10922), .ZN(n6714) );
  NAND2_X1 U8594 ( .A1(n6707), .A2(n6704), .ZN(n6715) );
  NAND2_X1 U8595 ( .A1(n10212), .A2(n10213), .ZN(n10214) );
  NAND2_X1 U8596 ( .A1(n10209), .A2(n10208), .ZN(n10535) );
  NOR2_X1 U8597 ( .A1(n10709), .A2(n6723), .ZN(n10716) );
  AND2_X1 U8598 ( .A1(n10710), .A2(n11268), .ZN(n6723) );
  NAND2_X1 U8599 ( .A1(n10716), .A2(n10715), .ZN(n11012) );
  NAND2_X1 U8600 ( .A1(n12033), .A2(n12034), .ZN(n12035) );
  NAND2_X1 U8601 ( .A1(n12035), .A2(n12036), .ZN(n12054) );
  XNOR2_X1 U8602 ( .A(n12083), .B(n6888), .ZN(n12085) );
  AOI21_X1 U8603 ( .B1(n12062), .B2(n14202), .A(n12061), .ZN(n12064) );
  XNOR2_X1 U8604 ( .A(n6722), .B(n14208), .ZN(n12072) );
  INV_X1 U8605 ( .A(n12094), .ZN(n6722) );
  AND2_X1 U8606 ( .A1(n12116), .A2(n11255), .ZN(n12129) );
  NAND2_X1 U8607 ( .A1(n11252), .A2(n11251), .ZN(n12321) );
  NAND2_X1 U8608 ( .A1(n6777), .A2(n6776), .ZN(n12123) );
  INV_X1 U8609 ( .A(n11688), .ZN(n12332) );
  AOI21_X1 U8610 ( .B1(n12330), .B2(n14878), .A(n11685), .ZN(n11686) );
  NAND2_X1 U8611 ( .A1(n11420), .A2(n11419), .ZN(n12333) );
  OR2_X1 U8612 ( .A1(n11454), .A2(n11418), .ZN(n11419) );
  NAND2_X1 U8613 ( .A1(n11417), .A2(n11464), .ZN(n11420) );
  INV_X1 U8614 ( .A(n11845), .ZN(n12341) );
  NAND2_X1 U8615 ( .A1(n7418), .A2(n11675), .ZN(n12203) );
  NAND2_X1 U8616 ( .A1(n11374), .A2(n11373), .ZN(n12351) );
  NAND2_X1 U8617 ( .A1(n11371), .A2(n11464), .ZN(n11374) );
  NAND2_X1 U8618 ( .A1(n11363), .A2(n11362), .ZN(n12354) );
  OR2_X1 U8619 ( .A1(n11454), .A2(n11361), .ZN(n11362) );
  NAND2_X1 U8620 ( .A1(n12241), .A2(n11492), .ZN(n12231) );
  NAND2_X1 U8621 ( .A1(n12236), .A2(n11672), .ZN(n12223) );
  NAND2_X1 U8622 ( .A1(n11338), .A2(n11337), .ZN(n12362) );
  NAND2_X1 U8623 ( .A1(n12280), .A2(n11664), .ZN(n12269) );
  AND2_X1 U8624 ( .A1(n14904), .A2(n10917), .ZN(n12305) );
  NAND2_X1 U8625 ( .A1(n7152), .A2(n11543), .ZN(n14813) );
  INV_X1 U8626 ( .A(n12252), .ZN(n14231) );
  AND2_X1 U8627 ( .A1(n9619), .A2(n9383), .ZN(n14884) );
  AND2_X2 U8628 ( .A1(n12317), .A2(n12316), .ZN(n14968) );
  NAND2_X1 U8629 ( .A1(n12328), .A2(n12327), .ZN(n12389) );
  INV_X2 U8630 ( .A(n14949), .ZN(n14948) );
  AND2_X1 U8631 ( .A1(n9020), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9015) );
  OAI21_X1 U8632 ( .B1(n9364), .B2(P3_D_REG_0__SCAN_IN), .A(n9351), .ZN(n9352)
         );
  INV_X1 U8633 ( .A(n9015), .ZN(n12404) );
  XNOR2_X1 U8634 ( .A(n7028), .B(n11452), .ZN(n12411) );
  AOI21_X1 U8635 ( .B1(n11462), .B2(n11461), .A(n7029), .ZN(n7028) );
  INV_X1 U8636 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12407) );
  INV_X1 U8637 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9010) );
  XNOR2_X1 U8638 ( .A(n11261), .B(n11260), .ZN(n11711) );
  AND2_X1 U8639 ( .A1(n6757), .A2(n6636), .ZN(n11247) );
  NAND2_X1 U8640 ( .A1(n8687), .A2(n8686), .ZN(n10851) );
  INV_X1 U8641 ( .A(n8685), .ZN(n8687) );
  AOI21_X1 U8642 ( .B1(n9860), .B2(n7228), .A(n6491), .ZN(n10595) );
  XNOR2_X1 U8643 ( .A(n9018), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U8644 ( .A1(n9017), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U8645 ( .A1(n9860), .A2(n7230), .ZN(n10122) );
  INV_X1 U8646 ( .A(n9466), .ZN(n11499) );
  NAND2_X1 U8647 ( .A1(n9348), .A2(n9347), .ZN(n9639) );
  NAND2_X1 U8648 ( .A1(n6761), .A2(n7191), .ZN(n9636) );
  NAND2_X1 U8649 ( .A1(n11331), .A2(n11329), .ZN(n6761) );
  NAND2_X1 U8650 ( .A1(n6766), .A2(n9111), .ZN(n11273) );
  NAND2_X1 U8651 ( .A1(n11267), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8652 ( .A1(n8789), .A2(n8674), .ZN(n10531) );
  INV_X1 U8653 ( .A(SI_11_), .ZN(n8769) );
  NAND2_X1 U8654 ( .A1(n7199), .A2(n8768), .ZN(n8792) );
  NAND2_X1 U8655 ( .A1(n8766), .A2(n8765), .ZN(n7199) );
  NAND2_X1 U8656 ( .A1(n7013), .A2(n8724), .ZN(n10601) );
  NAND2_X1 U8657 ( .A1(n8731), .A2(n8729), .ZN(n7013) );
  INV_X1 U8658 ( .A(n7019), .ZN(n8719) );
  AOI21_X1 U8659 ( .B1(n7205), .B2(n7203), .A(n6492), .ZN(n7019) );
  NAND2_X1 U8660 ( .A1(n7205), .A2(n8709), .ZN(n8748) );
  NAND2_X1 U8661 ( .A1(n8741), .A2(n8740), .ZN(n9432) );
  NOR2_X1 U8662 ( .A1(n8553), .A2(n8552), .ZN(n8932) );
  NAND2_X1 U8663 ( .A1(n7008), .A2(n9335), .ZN(n9575) );
  NAND2_X1 U8664 ( .A1(n9334), .A2(n9333), .ZN(n7008) );
  NAND2_X1 U8665 ( .A1(n12791), .A2(n6487), .ZN(n6820) );
  NAND2_X1 U8666 ( .A1(n9902), .A2(n7399), .ZN(n9904) );
  OR2_X1 U8667 ( .A1(n12571), .A2(n12885), .ZN(n12476) );
  INV_X1 U8668 ( .A(n7390), .ZN(n7005) );
  INV_X1 U8669 ( .A(n11760), .ZN(n7003) );
  NAND2_X1 U8670 ( .A1(n12518), .A2(n12520), .ZN(n12517) );
  NAND2_X1 U8671 ( .A1(n12517), .A2(n12463), .ZN(n12462) );
  NOR2_X1 U8672 ( .A1(n7875), .A2(n7874), .ZN(n10759) );
  NAND2_X2 U8673 ( .A1(n7847), .A2(n7846), .ZN(n10768) );
  AND4_X1 U8674 ( .A1(n8103), .A2(n8102), .A3(n8101), .A4(n8100), .ZN(n12776)
         );
  AND2_X1 U8675 ( .A1(n7932), .A2(n7931), .ZN(n12495) );
  NOR2_X1 U8676 ( .A1(n10486), .A2(n10487), .ZN(n10485) );
  INV_X1 U8677 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U8678 ( .A1(n7000), .A2(n7395), .ZN(n10086) );
  NAND2_X1 U8679 ( .A1(n9640), .A2(n6529), .ZN(n7000) );
  NAND2_X1 U8680 ( .A1(n12507), .A2(n11727), .ZN(n12550) );
  NAND2_X1 U8681 ( .A1(n9129), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12538) );
  INV_X1 U8682 ( .A(n12476), .ZN(n12563) );
  NAND2_X1 U8683 ( .A1(n9088), .A2(n12886), .ZN(n12569) );
  NAND2_X1 U8684 ( .A1(n6646), .A2(n7484), .ZN(n6645) );
  NAND2_X1 U8685 ( .A1(n6644), .A2(n6643), .ZN(n6642) );
  INV_X1 U8686 ( .A(n12728), .ZN(n12758) );
  INV_X1 U8687 ( .A(n12776), .ZN(n12746) );
  INV_X1 U8688 ( .A(n10758), .ZN(n12579) );
  INV_X1 U8689 ( .A(n7388), .ZN(n7387) );
  OAI211_X1 U8690 ( .C1(n8077), .C2(n7389), .A(n7651), .B(n7649), .ZN(n7388)
         );
  NAND2_X1 U8691 ( .A1(n7646), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7582) );
  INV_X1 U8692 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12684) );
  AND2_X1 U8693 ( .A1(n8956), .A2(n8955), .ZN(n14657) );
  CLKBUF_X1 U8694 ( .A(n8216), .Z(n8217) );
  INV_X1 U8695 ( .A(n8236), .ZN(n12902) );
  NAND2_X1 U8696 ( .A1(n12913), .A2(n7206), .ZN(n12702) );
  NAND2_X1 U8697 ( .A1(n6906), .A2(n6904), .ZN(n12695) );
  INV_X1 U8698 ( .A(n6905), .ZN(n6904) );
  NAND2_X1 U8699 ( .A1(n6911), .A2(n6910), .ZN(n12710) );
  INV_X1 U8700 ( .A(n12767), .ZN(n12934) );
  INV_X1 U8701 ( .A(n7221), .ZN(n12797) );
  INV_X1 U8702 ( .A(n7223), .ZN(n7220) );
  INV_X1 U8703 ( .A(n12940), .ZN(n12796) );
  NAND2_X1 U8704 ( .A1(n7315), .A2(n8336), .ZN(n12789) );
  NAND2_X1 U8705 ( .A1(n6732), .A2(n8404), .ZN(n12819) );
  NAND2_X1 U8706 ( .A1(n12838), .A2(n8403), .ZN(n6732) );
  NAND2_X1 U8707 ( .A1(n7236), .A2(n8402), .ZN(n12844) );
  OR2_X1 U8708 ( .A1(n7238), .A2(n7237), .ZN(n7236) );
  NAND2_X1 U8709 ( .A1(n7286), .A2(n7287), .ZN(n12859) );
  INV_X1 U8710 ( .A(n12495), .ZN(n12970) );
  AND2_X1 U8711 ( .A1(n6897), .A2(n12577), .ZN(n8330) );
  INV_X1 U8712 ( .A(n7823), .ZN(n6810) );
  AND2_X1 U8713 ( .A1(n7783), .A2(n7782), .ZN(n10324) );
  NAND2_X1 U8714 ( .A1(n8320), .A2(n8319), .ZN(n9649) );
  NAND2_X1 U8715 ( .A1(n9492), .A2(n8387), .ZN(n10692) );
  NAND2_X1 U8716 ( .A1(n10264), .A2(n8310), .ZN(n10331) );
  NAND2_X1 U8717 ( .A1(n7212), .A2(n8385), .ZN(n10343) );
  INV_X1 U8718 ( .A(n14667), .ZN(n12811) );
  NAND2_X1 U8719 ( .A1(n12889), .A2(n9086), .ZN(n14673) );
  INV_X1 U8720 ( .A(n14673), .ZN(n12896) );
  NAND2_X1 U8721 ( .A1(n14685), .A2(n9487), .ZN(n12886) );
  NOR2_X2 U8722 ( .A1(n12858), .A2(n7987), .ZN(n14667) );
  AND2_X1 U8723 ( .A1(n9083), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14685) );
  NOR2_X1 U8724 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7320) );
  XNOR2_X1 U8725 ( .A(n8296), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13004) );
  AND2_X1 U8726 ( .A1(n8299), .A2(n8300), .ZN(n10905) );
  INV_X1 U8727 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10553) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9562) );
  INV_X1 U8729 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8844) );
  INV_X1 U8730 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8771) );
  INV_X1 U8731 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8759) );
  INV_X1 U8732 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8736) );
  INV_X1 U8733 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U8734 ( .A1(n7467), .A2(n7474), .ZN(n13310) );
  NAND2_X1 U8735 ( .A1(n7478), .A2(n7476), .ZN(n7467) );
  NAND2_X1 U8736 ( .A1(n13383), .A2(n13079), .ZN(n13117) );
  NAND2_X1 U8737 ( .A1(n10558), .A2(n7448), .ZN(n10876) );
  NAND2_X1 U8738 ( .A1(n13394), .A2(n13052), .ZN(n13300) );
  NAND2_X1 U8739 ( .A1(n7464), .A2(n7468), .ZN(n13317) );
  INV_X1 U8740 ( .A(n7469), .ZN(n7468) );
  NAND2_X1 U8741 ( .A1(n13336), .A2(n7465), .ZN(n7464) );
  OAI21_X1 U8742 ( .B1(n13309), .B2(n7470), .A(n7477), .ZN(n7469) );
  AND2_X1 U8743 ( .A1(n6946), .A2(n6532), .ZN(n10352) );
  NAND2_X1 U8744 ( .A1(n13376), .A2(n13068), .ZN(n13328) );
  INV_X1 U8745 ( .A(n7433), .ZN(n7431) );
  AND2_X1 U8746 ( .A1(n13348), .A2(n7429), .ZN(n7428) );
  AND2_X1 U8747 ( .A1(n7437), .A2(n7438), .ZN(n13347) );
  NAND2_X1 U8748 ( .A1(n7432), .A2(n13029), .ZN(n7438) );
  NAND2_X1 U8749 ( .A1(n13418), .A2(n13417), .ZN(n7437) );
  INV_X1 U8750 ( .A(n7439), .ZN(n7432) );
  AOI21_X1 U8751 ( .B1(n7480), .B2(n7482), .A(n6561), .ZN(n7479) );
  INV_X1 U8752 ( .A(n6926), .ZN(n6934) );
  NAND2_X1 U8753 ( .A1(n10499), .A2(n10498), .ZN(n10558) );
  OAI21_X1 U8754 ( .B1(n13394), .B2(n6952), .A(n6950), .ZN(n13376) );
  NAND2_X1 U8755 ( .A1(n13298), .A2(n13061), .ZN(n13378) );
  OAI21_X1 U8756 ( .B1(n10351), .B2(n6942), .A(n6939), .ZN(n14298) );
  INV_X1 U8757 ( .A(n6944), .ZN(n6942) );
  AND2_X1 U8758 ( .A1(n6947), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U8759 ( .A1(n7446), .A2(n7447), .ZN(n6947) );
  NAND2_X1 U8760 ( .A1(n14298), .A2(n14299), .ZN(n14297) );
  INV_X1 U8761 ( .A(n13425), .ZN(n14366) );
  NAND2_X1 U8762 ( .A1(n9738), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14376) );
  XNOR2_X1 U8763 ( .A(n7439), .B(n13029), .ZN(n13418) );
  AND2_X1 U8764 ( .A1(n14364), .A2(n14499), .ZN(n14300) );
  NAND2_X1 U8765 ( .A1(n9739), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8610) );
  OR2_X2 U8766 ( .A1(n8808), .A2(n9152), .ZN(n13668) );
  INV_X1 U8767 ( .A(n6982), .ZN(n8868) );
  XNOR2_X1 U8768 ( .A(n10629), .B(n14384), .ZN(n14382) );
  INV_X1 U8769 ( .A(n6975), .ZN(n13751) );
  AND2_X1 U8770 ( .A1(n9823), .A2(n10090), .ZN(n13752) );
  XNOR2_X1 U8771 ( .A(n13764), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13771) );
  INV_X1 U8772 ( .A(n6973), .ZN(n13761) );
  OAI21_X1 U8773 ( .B1(n13771), .B2(n13737), .A(n6979), .ZN(n13775) );
  INV_X1 U8774 ( .A(n6980), .ZN(n6979) );
  OAI21_X1 U8775 ( .B1(n13774), .B2(n13773), .A(n13772), .ZN(n6980) );
  AOI22_X1 U8776 ( .A1(n12992), .A2(n13595), .B1(n13594), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U8777 ( .A1(n7106), .A2(n14429), .ZN(n14040) );
  XNOR2_X1 U8778 ( .A(n13785), .B(n7107), .ZN(n7106) );
  INV_X1 U8779 ( .A(n14041), .ZN(n7107) );
  NAND2_X1 U8780 ( .A1(n13576), .A2(n13575), .ZN(n13791) );
  NAND2_X1 U8781 ( .A1(n13565), .A2(n13564), .ZN(n14049) );
  NAND2_X1 U8782 ( .A1(n13818), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U8783 ( .A1(n6683), .A2(n6681), .ZN(n14067) );
  NAND2_X1 U8784 ( .A1(n6684), .A2(n14411), .ZN(n6683) );
  INV_X1 U8785 ( .A(n6682), .ZN(n6681) );
  OAI21_X1 U8786 ( .B1(n13822), .B2(n13821), .A(n13820), .ZN(n6684) );
  NAND2_X1 U8787 ( .A1(n13870), .A2(n11232), .ZN(n13853) );
  NAND2_X1 U8788 ( .A1(n13873), .A2(n11166), .ZN(n13851) );
  INV_X1 U8789 ( .A(n14087), .ZN(n13896) );
  NAND2_X1 U8790 ( .A1(n13936), .A2(n11120), .ZN(n13920) );
  NAND2_X1 U8791 ( .A1(n13996), .A2(n11077), .ZN(n13981) );
  NAND2_X1 U8792 ( .A1(n6730), .A2(n6731), .ZN(n13978) );
  OR2_X1 U8793 ( .A1(n13995), .A2(n13626), .ZN(n6730) );
  NAND2_X1 U8794 ( .A1(n11069), .A2(n13509), .ZN(n13998) );
  NAND2_X1 U8795 ( .A1(n11218), .A2(n7513), .ZN(n14023) );
  NAND2_X1 U8796 ( .A1(n10972), .A2(n10971), .ZN(n14291) );
  NAND2_X1 U8797 ( .A1(n7167), .A2(n10795), .ZN(n10852) );
  NAND2_X1 U8798 ( .A1(n10794), .A2(n13620), .ZN(n7167) );
  NAND2_X1 U8799 ( .A1(n10508), .A2(n7187), .ZN(n10572) );
  NAND2_X1 U8800 ( .A1(n10508), .A2(n10507), .ZN(n10514) );
  NAND2_X1 U8801 ( .A1(n10394), .A2(n10393), .ZN(n10396) );
  NAND2_X1 U8802 ( .A1(n7366), .A2(n7367), .ZN(n10397) );
  NAND2_X1 U8803 ( .A1(n7176), .A2(n9990), .ZN(n10184) );
  NAND2_X1 U8804 ( .A1(n7368), .A2(n9976), .ZN(n10194) );
  OR2_X1 U8805 ( .A1(n14393), .A2(n14394), .ZN(n7368) );
  OR2_X1 U8806 ( .A1(n6479), .A2(n8665), .ZN(n14422) );
  NAND2_X1 U8807 ( .A1(n6686), .A2(n9814), .ZN(n9986) );
  NAND2_X1 U8808 ( .A1(n14410), .A2(n9813), .ZN(n6686) );
  OR2_X1 U8809 ( .A1(n6479), .A2(n9806), .ZN(n14025) );
  INV_X1 U8810 ( .A(n14422), .ZN(n14033) );
  OR2_X1 U8811 ( .A1(n13807), .A2(n13928), .ZN(n14022) );
  INV_X1 U8812 ( .A(n14421), .ZN(n14400) );
  INV_X1 U8813 ( .A(n14534), .ZN(n14532) );
  NAND2_X1 U8814 ( .A1(n14040), .A2(n7104), .ZN(n14139) );
  INV_X1 U8815 ( .A(n7105), .ZN(n7104) );
  OAI21_X1 U8816 ( .B1(n14041), .B2(n14512), .A(n14042), .ZN(n7105) );
  INV_X1 U8817 ( .A(n13572), .ZN(n11715) );
  NAND2_X1 U8818 ( .A1(n8616), .A2(n6502), .ZN(n8559) );
  INV_X1 U8819 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14162) );
  INV_X1 U8820 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14172) );
  NAND2_X1 U8821 ( .A1(n8548), .A2(n8579), .ZN(n10994) );
  NAND2_X1 U8822 ( .A1(n7177), .A2(n8757), .ZN(n8546) );
  XNOR2_X1 U8823 ( .A(n8070), .B(n8069), .ZN(n11142) );
  INV_X1 U8824 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9571) );
  INV_X1 U8825 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9276) );
  INV_X1 U8826 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8842) );
  AND2_X1 U8827 ( .A1(n8825), .A2(n8829), .ZN(n13725) );
  INV_X1 U8828 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U8829 ( .A1(n7660), .A2(n7058), .ZN(n7001) );
  OR2_X1 U8830 ( .A1(n8582), .A2(n14155), .ZN(n8600) );
  INV_X1 U8831 ( .A(n8582), .ZN(n8583) );
  NAND2_X1 U8832 ( .A1(n8478), .A2(n8479), .ZN(n14180) );
  OAI21_X1 U8833 ( .B1(n8483), .B2(n14980), .A(n14977), .ZN(n14969) );
  XNOR2_X1 U8834 ( .A(n8470), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n14970) );
  XNOR2_X1 U8835 ( .A(n8487), .B(n8488), .ZN(n14971) );
  INV_X1 U8836 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7126) );
  XNOR2_X1 U8837 ( .A(n8495), .B(n12634), .ZN(n14975) );
  INV_X1 U8838 ( .A(n8505), .ZN(n7127) );
  AND2_X1 U8839 ( .A1(n6796), .A2(n6794), .ZN(n14210) );
  AND2_X1 U8840 ( .A1(n8506), .A2(n6795), .ZN(n6794) );
  INV_X1 U8841 ( .A(n14212), .ZN(n6795) );
  NOR2_X1 U8842 ( .A1(n6791), .A2(n14343), .ZN(n14346) );
  OAI21_X1 U8843 ( .B1(n14346), .B2(n14347), .A(P2_ADDR_REG_12__SCAN_IN), .ZN(
        n6800) );
  NAND2_X1 U8844 ( .A1(n14346), .A2(n14347), .ZN(n14345) );
  AND2_X1 U8845 ( .A1(n6797), .A2(n7122), .ZN(n14358) );
  OAI21_X1 U8846 ( .B1(n7124), .B2(n7123), .A(n14619), .ZN(n6797) );
  NOR2_X1 U8847 ( .A1(n14358), .A2(n14357), .ZN(n14356) );
  AOI21_X1 U8848 ( .B1(n6799), .B2(n14647), .A(n14361), .ZN(n14222) );
  INV_X1 U8849 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U8850 ( .A1(n7072), .A2(n11984), .ZN(n7071) );
  INV_X1 U8851 ( .A(n6679), .ZN(P3_U3296) );
  OAI21_X1 U8852 ( .B1(n7140), .B2(n6680), .A(n7023), .ZN(n6679) );
  NAND2_X1 U8853 ( .A1(n7022), .A2(n7024), .ZN(n6680) );
  AOI21_X1 U8854 ( .B1(n9953), .B2(n9952), .A(n6713), .ZN(n10094) );
  NAND2_X1 U8855 ( .A1(n6703), .A2(n6709), .ZN(n10207) );
  XNOR2_X1 U8856 ( .A(n6721), .B(n6830), .ZN(n12114) );
  AND2_X1 U8857 ( .A1(n6884), .A2(n6883), .ZN(n12112) );
  INV_X1 U8858 ( .A(n12095), .ZN(n6830) );
  NOR2_X1 U8859 ( .A1(n6837), .A2(n6836), .ZN(n6835) );
  INV_X1 U8860 ( .A(n12431), .ZN(n6836) );
  NAND2_X1 U8861 ( .A1(n6740), .A2(n6914), .ZN(P2_U3528) );
  NAND2_X1 U8862 ( .A1(n14777), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6914) );
  INV_X1 U8863 ( .A(n12906), .ZN(n6741) );
  NAND2_X1 U8864 ( .A1(n14762), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U8865 ( .A1(n7047), .A2(n14764), .ZN(n7046) );
  AND2_X1 U8866 ( .A1(n13644), .A2(n6873), .ZN(n13649) );
  INV_X1 U8867 ( .A(n7124), .ZN(n14354) );
  INV_X1 U8868 ( .A(n7122), .ZN(n14352) );
  INV_X1 U8869 ( .A(n6799), .ZN(n14360) );
  XNOR2_X1 U8870 ( .A(n7519), .B(n12104), .ZN(n8525) );
  AND2_X1 U8871 ( .A1(n6509), .A2(n13559), .ZN(n6490) );
  AND2_X1 U8872 ( .A1(n11785), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6491) );
  CLKBUF_X3 U8873 ( .A(n9825), .Z(n11400) );
  INV_X1 U8874 ( .A(n13871), .ZN(n7373) );
  AND2_X1 U8875 ( .A1(n9919), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6492) );
  AND2_X1 U8876 ( .A1(n10050), .A2(n10043), .ZN(n6493) );
  AND2_X1 U8877 ( .A1(n13622), .A2(n7168), .ZN(n6494) );
  OR2_X1 U8878 ( .A1(n7251), .A2(n13504), .ZN(n6495) );
  INV_X1 U8879 ( .A(n6483), .ZN(n7672) );
  NOR2_X1 U8880 ( .A1(n13472), .A2(n13663), .ZN(n6496) );
  OR2_X1 U8881 ( .A1(n12874), .A2(n12966), .ZN(n6497) );
  AND2_X1 U8882 ( .A1(n14276), .A2(n12578), .ZN(n6498) );
  NAND2_X1 U8883 ( .A1(n7342), .A2(n6615), .ZN(n6499) );
  INV_X1 U8884 ( .A(n7986), .ZN(n6960) );
  XOR2_X1 U8885 ( .A(n12940), .B(n6968), .Z(n6500) );
  AND2_X1 U8886 ( .A1(n9810), .A2(n6747), .ZN(n6501) );
  NAND2_X1 U8887 ( .A1(n8033), .A2(n8032), .ZN(n12946) );
  INV_X1 U8888 ( .A(n12946), .ZN(n7224) );
  INV_X1 U8889 ( .A(n10651), .ZN(n7292) );
  NOR2_X1 U8890 ( .A1(n12174), .A2(n12171), .ZN(n6503) );
  NAND2_X1 U8891 ( .A1(n7413), .A2(n8670), .ZN(n8772) );
  INV_X1 U8892 ( .A(n13499), .ZN(n14325) );
  NAND2_X1 U8893 ( .A1(n10857), .A2(n10856), .ZN(n13499) );
  OR2_X1 U8894 ( .A1(n13560), .A2(n6847), .ZN(n6504) );
  AND2_X1 U8895 ( .A1(n8128), .A2(n8127), .ZN(n12734) );
  AND2_X1 U8896 ( .A1(n11640), .A2(n11672), .ZN(n6505) );
  AND3_X1 U8897 ( .A1(n13485), .A2(n6871), .A3(n7278), .ZN(n6506) );
  NAND2_X1 U8898 ( .A1(n7878), .A2(n7460), .ZN(n7459) );
  INV_X1 U8899 ( .A(n7459), .ZN(n7457) );
  NAND2_X1 U8900 ( .A1(n10873), .A2(n10874), .ZN(n7447) );
  OR2_X1 U8901 ( .A1(n13329), .A2(n7485), .ZN(n6507) );
  NAND2_X1 U8902 ( .A1(n7265), .A2(n13593), .ZN(n6508) );
  INV_X1 U8903 ( .A(n7118), .ZN(n7117) );
  NAND2_X1 U8904 ( .A1(n7120), .A2(n7119), .ZN(n7118) );
  NAND2_X1 U8905 ( .A1(n13560), .A2(n6846), .ZN(n6509) );
  NOR2_X1 U8906 ( .A1(n6602), .A2(n7500), .ZN(n6511) );
  AND2_X1 U8907 ( .A1(n11671), .A2(n11670), .ZN(n6512) );
  AND2_X1 U8908 ( .A1(n6612), .A2(n6504), .ZN(n6513) );
  INV_X1 U8909 ( .A(n14832), .ZN(n12027) );
  AND4_X1 U8910 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n14832) );
  AND2_X1 U8911 ( .A1(n7149), .A2(n7146), .ZN(n6514) );
  XOR2_X1 U8912 ( .A(n11951), .B(n12140), .Z(n6515) );
  AND2_X1 U8913 ( .A1(n7073), .A2(n6618), .ZN(n6516) );
  INV_X1 U8914 ( .A(n9858), .ZN(n7032) );
  AND2_X1 U8915 ( .A1(n11539), .A2(n11540), .ZN(n11624) );
  INV_X1 U8916 ( .A(n11624), .ZN(n6676) );
  AND2_X1 U8917 ( .A1(n8080), .A2(n8079), .ZN(n12539) );
  INV_X1 U8918 ( .A(n12539), .ZN(n12791) );
  OAI21_X1 U8919 ( .B1(n7228), .B2(n6491), .A(n7227), .ZN(n7226) );
  NOR2_X1 U8920 ( .A1(n7225), .A2(n7222), .ZN(n7221) );
  XOR2_X1 U8921 ( .A(n11718), .B(n11762), .Z(n6517) );
  NAND4_X1 U8922 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n14415)
         );
  OR2_X1 U8923 ( .A1(n13105), .A2(n13104), .ZN(n6518) );
  NOR2_X1 U8924 ( .A1(n11322), .A2(n11313), .ZN(n6519) );
  NAND2_X1 U8925 ( .A1(n12251), .A2(n12250), .ZN(n12249) );
  NAND2_X1 U8926 ( .A1(n6746), .A2(n8561), .ZN(n8564) );
  OR2_X1 U8927 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9024), .ZN(n6520) );
  AND2_X1 U8928 ( .A1(n13631), .A2(n7162), .ZN(n6521) );
  AND2_X1 U8929 ( .A1(n11033), .A2(n12996), .ZN(n7635) );
  AND2_X1 U8930 ( .A1(n13057), .A2(n13052), .ZN(n6522) );
  NOR2_X1 U8931 ( .A1(n10559), .A2(n10560), .ZN(n7449) );
  INV_X1 U8932 ( .A(n7201), .ZN(n7200) );
  OAI21_X1 U8933 ( .B1(n8765), .B2(n7202), .A(n8791), .ZN(n7201) );
  INV_X1 U8934 ( .A(n7207), .ZN(n7206) );
  NOR2_X1 U8935 ( .A1(n12432), .A2(n12729), .ZN(n7207) );
  NAND2_X1 U8936 ( .A1(n11717), .A2(n11716), .ZN(n6523) );
  BUF_X1 U8937 ( .A(n8586), .Z(n13432) );
  INV_X1 U8938 ( .A(n7810), .ZN(n7444) );
  OR2_X1 U8939 ( .A1(n8423), .A2(n8422), .ZN(n6524) );
  NAND2_X1 U8940 ( .A1(n12796), .A2(n6968), .ZN(n6526) );
  AND2_X1 U8941 ( .A1(n13880), .A2(n7113), .ZN(n6527) );
  NAND2_X1 U8942 ( .A1(n6919), .A2(n13092), .ZN(n13336) );
  NOR2_X1 U8943 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8739) );
  NAND2_X1 U8944 ( .A1(n7119), .A2(n14001), .ZN(n6528) );
  AND2_X1 U8945 ( .A1(n6493), .A2(n9641), .ZN(n6529) );
  AND2_X1 U8946 ( .A1(n8674), .A2(n7158), .ZN(n6530) );
  INV_X1 U8947 ( .A(n7896), .ZN(n7463) );
  NAND2_X1 U8948 ( .A1(n13934), .A2(n7527), .ZN(n13918) );
  OR2_X1 U8949 ( .A1(n11779), .A2(n11719), .ZN(n6531) );
  INV_X1 U8950 ( .A(n14498), .ZN(n7109) );
  OR2_X1 U8951 ( .A1(n10349), .A2(n10348), .ZN(n6532) );
  INV_X1 U8952 ( .A(n13504), .ZN(n7255) );
  NAND2_X1 U8953 ( .A1(n6702), .A2(n6700), .ZN(n14363) );
  INV_X1 U8954 ( .A(n14363), .ZN(n6747) );
  AND4_X1 U8955 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n6533)
         );
  INV_X1 U8956 ( .A(n11197), .ZN(n7164) );
  INV_X1 U8957 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6767) );
  INV_X1 U8958 ( .A(n7197), .ZN(n8380) );
  AND2_X1 U8959 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6534) );
  AND2_X1 U8960 ( .A1(n8072), .A2(n8071), .ZN(n12783) );
  INV_X1 U8961 ( .A(n12783), .ZN(n7102) );
  NAND2_X1 U8962 ( .A1(n11068), .A2(n11067), .ZN(n14307) );
  INV_X1 U8963 ( .A(n14307), .ZN(n7119) );
  AND3_X2 U8964 ( .A1(n6890), .A2(n8964), .A3(n6891), .ZN(n7603) );
  NAND2_X1 U8965 ( .A1(n8115), .A2(n8114), .ZN(n12926) );
  INV_X1 U8966 ( .A(n12926), .ZN(n7100) );
  NOR2_X1 U8967 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7601) );
  NOR2_X1 U8968 ( .A1(n8700), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8755) );
  AND3_X1 U8969 ( .A1(n6510), .A2(n8789), .A3(n7157), .ZN(n8683) );
  OR3_X1 U8970 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6535) );
  INV_X1 U8971 ( .A(n13562), .ZN(n7283) );
  INV_X1 U8972 ( .A(n13481), .ZN(n6872) );
  OR2_X1 U8973 ( .A1(n10315), .A2(n12579), .ZN(n6536) );
  INV_X1 U8974 ( .A(n8325), .ZN(n9889) );
  XNOR2_X1 U8975 ( .A(n14498), .B(n10565), .ZN(n13617) );
  AND2_X1 U8976 ( .A1(n14173), .A2(n11132), .ZN(n14094) );
  NOR2_X1 U8977 ( .A1(n11617), .A2(n11479), .ZN(n6537) );
  NOR2_X1 U8978 ( .A1(n13664), .A2(n10192), .ZN(n6538) );
  INV_X1 U8979 ( .A(n9448), .ZN(n9635) );
  OR2_X1 U8980 ( .A1(n10004), .A2(n14955), .ZN(n6539) );
  OR2_X1 U8981 ( .A1(n10004), .A2(n14863), .ZN(n6540) );
  AND2_X1 U8982 ( .A1(n8528), .A2(n6841), .ZN(n8757) );
  AND2_X1 U8983 ( .A1(n10231), .A2(n12028), .ZN(n6541) );
  OR2_X1 U8984 ( .A1(n7224), .A2(n12817), .ZN(n6542) );
  AND2_X1 U8985 ( .A1(n13854), .A2(n11166), .ZN(n6543) );
  AND4_X1 U8986 ( .A1(n7548), .A2(n7547), .A3(n7546), .A4(n7284), .ZN(n6544)
         );
  NOR2_X1 U8987 ( .A1(n7225), .A2(n7220), .ZN(n6545) );
  AND2_X1 U8988 ( .A1(n11538), .A2(n10941), .ZN(n6546) );
  NAND2_X1 U8989 ( .A1(n12793), .A2(n7098), .ZN(n7103) );
  AND2_X1 U8990 ( .A1(n7973), .A2(n7972), .ZN(n12853) );
  INV_X1 U8991 ( .A(n12853), .ZN(n12961) );
  NAND2_X1 U8992 ( .A1(n8528), .A2(n8527), .ZN(n8700) );
  OR2_X1 U8993 ( .A1(n7767), .A2(n7769), .ZN(n6547) );
  AND2_X1 U8994 ( .A1(n13479), .A2(n13478), .ZN(n6548) );
  NAND2_X1 U8995 ( .A1(n9727), .A2(n9729), .ZN(n9730) );
  INV_X1 U8996 ( .A(n9730), .ZN(n6925) );
  OR2_X1 U8997 ( .A1(n7694), .A2(n7693), .ZN(n6549) );
  OR2_X1 U8998 ( .A1(n8405), .A2(n6737), .ZN(n6550) );
  OR2_X1 U8999 ( .A1(n6808), .A2(n14605), .ZN(n6551) );
  AND2_X1 U9000 ( .A1(n11720), .A2(n6517), .ZN(n6552) );
  AND2_X1 U9001 ( .A1(n7236), .A2(n7234), .ZN(n6553) );
  INV_X1 U9002 ( .A(n13454), .ZN(n13666) );
  AND4_X1 U9003 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n13454)
         );
  NAND2_X1 U9004 ( .A1(n11793), .A2(n11792), .ZN(n6554) );
  AND2_X1 U9005 ( .A1(n6526), .A2(n8336), .ZN(n6555) );
  NAND2_X1 U9006 ( .A1(n10705), .A2(n12582), .ZN(n6556) );
  AND2_X1 U9007 ( .A1(n7436), .A2(n7434), .ZN(n6557) );
  AND2_X1 U9008 ( .A1(n12853), .A2(n12443), .ZN(n6558) );
  AND2_X1 U9009 ( .A1(n7307), .A2(n12784), .ZN(n6559) );
  AND2_X1 U9010 ( .A1(n11729), .A2(n11727), .ZN(n6560) );
  INV_X1 U9011 ( .A(n7288), .ZN(n7287) );
  NOR2_X1 U9012 ( .A1(n8331), .A2(n7289), .ZN(n7288) );
  AND2_X1 U9013 ( .A1(n13085), .A2(n13084), .ZN(n6561) );
  AND2_X1 U9014 ( .A1(n11957), .A2(n7083), .ZN(n6562) );
  AND2_X1 U9015 ( .A1(n13870), .A2(n7374), .ZN(n6563) );
  OR2_X1 U9016 ( .A1(n8488), .A2(n8487), .ZN(n6564) );
  AND2_X1 U9017 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n8456), .ZN(n6565) );
  XNOR2_X1 U9018 ( .A(n8624), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8661) );
  AND2_X1 U9019 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6566) );
  OR2_X1 U9020 ( .A1(n14498), .A2(n13662), .ZN(n6567) );
  NOR2_X1 U9021 ( .A1(n13482), .A2(n10584), .ZN(n6568) );
  NOR2_X1 U9022 ( .A1(n13387), .A2(n13923), .ZN(n6569) );
  NOR2_X1 U9023 ( .A1(n13490), .A2(n10853), .ZN(n6570) );
  INV_X1 U9024 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14155) );
  INV_X1 U9025 ( .A(n7811), .ZN(n7443) );
  AND2_X1 U9026 ( .A1(n14853), .A2(n14917), .ZN(n6571) );
  AND2_X1 U9027 ( .A1(n13555), .A2(n13554), .ZN(n6572) );
  AND4_X1 U9028 ( .A1(n8590), .A2(n8589), .A3(n8588), .A4(n8587), .ZN(n9534)
         );
  INV_X1 U9029 ( .A(n9534), .ZN(n6938) );
  OR2_X1 U9030 ( .A1(n12783), .A2(n12539), .ZN(n6573) );
  AND2_X1 U9031 ( .A1(n6855), .A2(n6853), .ZN(n6574) );
  AND2_X1 U9032 ( .A1(n7502), .A2(n8024), .ZN(n6575) );
  INV_X1 U9033 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8964) );
  INV_X1 U9034 ( .A(n7099), .ZN(n7098) );
  NAND2_X1 U9035 ( .A1(n7100), .A2(n7101), .ZN(n7099) );
  AND2_X1 U9036 ( .A1(n7800), .A2(SI_9_), .ZN(n6576) );
  OR2_X1 U9037 ( .A1(n12701), .A2(n6905), .ZN(n6577) );
  INV_X1 U9038 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U9039 ( .A1(n8739), .A2(n7130), .ZN(n8750) );
  NOR2_X1 U9040 ( .A1(n6960), .A2(n6499), .ZN(n6578) );
  INV_X1 U9041 ( .A(n7089), .ZN(n7088) );
  NAND2_X1 U9042 ( .A1(n7090), .A2(n10060), .ZN(n7089) );
  NAND2_X1 U9043 ( .A1(n11608), .A2(n12131), .ZN(n11701) );
  AND2_X1 U9044 ( .A1(n8842), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6579) );
  AND2_X1 U9045 ( .A1(n7671), .A2(SI_4_), .ZN(n6580) );
  AND2_X1 U9046 ( .A1(n7881), .A2(SI_13_), .ZN(n6581) );
  AND2_X1 U9047 ( .A1(n8725), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6582) );
  AND2_X1 U9048 ( .A1(n7979), .A2(n7496), .ZN(n6583) );
  OR2_X1 U9049 ( .A1(n6501), .A2(n13454), .ZN(n6584) );
  AND4_X1 U9050 ( .A1(n8530), .A2(n9564), .A3(n9565), .A4(n9566), .ZN(n6585)
         );
  INV_X1 U9051 ( .A(n7456), .ZN(n7455) );
  OR2_X1 U9052 ( .A1(n7463), .A2(n7457), .ZN(n7456) );
  AND2_X1 U9053 ( .A1(n11622), .A2(n11621), .ZN(n12232) );
  INV_X1 U9054 ( .A(n7057), .ZN(n7056) );
  NAND2_X1 U9055 ( .A1(n7347), .A2(n7879), .ZN(n7057) );
  AND2_X1 U9056 ( .A1(n11233), .A2(n11175), .ZN(n13852) );
  AND2_X1 U9057 ( .A1(n7306), .A2(n7304), .ZN(n6586) );
  OAI21_X1 U9058 ( .B1(n10498), .B2(n7449), .A(n10875), .ZN(n7446) );
  OAI21_X1 U9059 ( .B1(n7156), .B2(n7154), .A(n11622), .ZN(n7153) );
  NAND2_X1 U9060 ( .A1(n6531), .A2(n7296), .ZN(n6587) );
  NAND2_X1 U9061 ( .A1(n7463), .A2(n7458), .ZN(n6588) );
  INV_X1 U9062 ( .A(n7449), .ZN(n7448) );
  AND2_X1 U9063 ( .A1(n11072), .A2(n11071), .ZN(n14008) );
  INV_X1 U9064 ( .A(n14008), .ZN(n14132) );
  INV_X1 U9065 ( .A(n7264), .ZN(n7263) );
  NAND2_X1 U9066 ( .A1(n7265), .A2(n7266), .ZN(n7264) );
  INV_X1 U9067 ( .A(n7877), .ZN(n7460) );
  AND2_X1 U9068 ( .A1(n9574), .A2(n9573), .ZN(n6589) );
  OR2_X1 U9069 ( .A1(n7645), .A2(n7644), .ZN(n6590) );
  OR2_X1 U9070 ( .A1(n6525), .A2(n10082), .ZN(n6591) );
  OR2_X1 U9071 ( .A1(n7221), .A2(n7218), .ZN(n6592) );
  AND2_X1 U9072 ( .A1(n7303), .A2(n6917), .ZN(n6593) );
  NOR2_X1 U9073 ( .A1(n14270), .A2(n10759), .ZN(n6594) );
  NAND2_X1 U9074 ( .A1(n13558), .A2(n13556), .ZN(n7274) );
  INV_X1 U9075 ( .A(n7274), .ZN(n6846) );
  AND3_X1 U9076 ( .A1(n8673), .A2(n7424), .A3(n8710), .ZN(n6595) );
  AND2_X1 U9077 ( .A1(n11484), .A2(n11483), .ZN(n12133) );
  NOR2_X1 U9078 ( .A1(n11646), .A2(n11794), .ZN(n6596) );
  AND2_X1 U9079 ( .A1(n11679), .A2(n11674), .ZN(n6597) );
  AND2_X1 U9080 ( .A1(n8576), .A2(n8575), .ZN(n6598) );
  AND2_X1 U9081 ( .A1(n11679), .A2(n7415), .ZN(n6599) );
  OR2_X1 U9082 ( .A1(n12766), .A2(n12776), .ZN(n6600) );
  AND2_X1 U9083 ( .A1(n7672), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6601) );
  AND2_X1 U9084 ( .A1(n11197), .A2(n11196), .ZN(n13822) );
  INV_X1 U9085 ( .A(n13822), .ZN(n7163) );
  NOR2_X1 U9086 ( .A1(n7502), .A2(n8024), .ZN(n6602) );
  INV_X1 U9087 ( .A(n13545), .ZN(n6860) );
  AND2_X1 U9088 ( .A1(n6502), .A2(n6744), .ZN(n6603) );
  NAND2_X1 U9089 ( .A1(n9911), .A2(n9910), .ZN(n6604) );
  AND2_X1 U9090 ( .A1(n7453), .A2(n7452), .ZN(n6605) );
  NAND2_X1 U9091 ( .A1(n14727), .A2(n10266), .ZN(n6606) );
  INV_X1 U9092 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U9093 ( .A1(n7811), .A2(n7444), .ZN(n6607) );
  AND2_X1 U9094 ( .A1(n13467), .A2(n6875), .ZN(n6608) );
  AND2_X1 U9095 ( .A1(n8771), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U9096 ( .A1(n8081), .A2(n8082), .ZN(n6610) );
  INV_X1 U9097 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7843) );
  INV_X1 U9098 ( .A(n7375), .ZN(n7374) );
  NAND2_X1 U9099 ( .A1(n13852), .A2(n11232), .ZN(n7375) );
  AND2_X1 U9100 ( .A1(n14727), .A2(n12585), .ZN(n6611) );
  INV_X1 U9101 ( .A(n6908), .ZN(n6907) );
  OR2_X1 U9102 ( .A1(n12720), .A2(n6909), .ZN(n6908) );
  INV_X1 U9103 ( .A(n7183), .ZN(n7182) );
  NAND2_X1 U9104 ( .A1(n7184), .A2(n13919), .ZN(n7183) );
  INV_X1 U9105 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7539) );
  INV_X1 U9106 ( .A(n8528), .ZN(n8612) );
  OR2_X1 U9107 ( .A1(n7283), .A2(n13561), .ZN(n6612) );
  INV_X1 U9108 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6851) );
  INV_X1 U9109 ( .A(n8606), .ZN(n13584) );
  INV_X1 U9110 ( .A(n8607), .ZN(n9795) );
  INV_X1 U9111 ( .A(n7937), .ZN(n6663) );
  NAND4_X1 U9112 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n12191) );
  INV_X1 U9113 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U9114 ( .A1(n6946), .A2(n6943), .ZN(n10499) );
  INV_X1 U9115 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7231) );
  OAI21_X1 U9116 ( .B1(n10394), .B2(n6693), .A(n6691), .ZN(n10794) );
  AND2_X1 U9117 ( .A1(n11492), .A2(n11491), .ZN(n12242) );
  INV_X1 U9118 ( .A(n12242), .ZN(n12237) );
  OAI21_X1 U9119 ( .B1(n12293), .B2(n11272), .A(n11561), .ZN(n12289) );
  XOR2_X1 U9120 ( .A(n11005), .B(n6828), .Z(n6613) );
  XNOR2_X1 U9121 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8752) );
  INV_X1 U9122 ( .A(n8752), .ZN(n6774) );
  XNOR2_X1 U9123 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8776) );
  INV_X1 U9124 ( .A(n8776), .ZN(n7018) );
  INV_X1 U9125 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7192) );
  AND2_X1 U9126 ( .A1(n8059), .A2(n8058), .ZN(n12772) );
  INV_X1 U9127 ( .A(n12772), .ZN(n6968) );
  NAND2_X1 U9128 ( .A1(n8041), .A2(n8040), .ZN(n12817) );
  AND2_X1 U9129 ( .A1(n12374), .A2(n12283), .ZN(n6614) );
  INV_X1 U9130 ( .A(n13476), .ZN(n7268) );
  INV_X1 U9131 ( .A(n14014), .ZN(n13655) );
  OR2_X1 U9132 ( .A1(n8029), .A2(n11361), .ZN(n6615) );
  INV_X1 U9133 ( .A(n8007), .ZN(n7342) );
  AND4_X1 U9134 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8134), .ZN(n12480)
         );
  INV_X1 U9135 ( .A(n12480), .ZN(n12747) );
  AND2_X1 U9136 ( .A1(n11843), .A2(n11961), .ZN(n6616) );
  AND2_X1 U9137 ( .A1(n10867), .A2(n7117), .ZN(n6617) );
  OR2_X1 U9138 ( .A1(n6515), .A2(n7076), .ZN(n6618) );
  AND2_X1 U9139 ( .A1(n12237), .A2(n11670), .ZN(n6619) );
  OR2_X1 U9140 ( .A1(n11719), .A2(n12885), .ZN(n6620) );
  NAND2_X1 U9141 ( .A1(n10942), .A2(n10941), .ZN(n6621) );
  INV_X1 U9142 ( .A(n7079), .ZN(n7078) );
  NAND2_X1 U9143 ( .A1(n11949), .A2(n12191), .ZN(n7079) );
  AND2_X1 U9144 ( .A1(n11218), .A2(n7380), .ZN(n6622) );
  INV_X1 U9145 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8536) );
  NOR2_X1 U9146 ( .A1(n11968), .A2(n11967), .ZN(n6623) );
  INV_X1 U9147 ( .A(n7084), .ZN(n7083) );
  OR2_X1 U9148 ( .A1(n11903), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U9149 ( .A1(n11718), .A2(n11719), .ZN(n6624) );
  INV_X1 U9150 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6812) );
  INV_X1 U9151 ( .A(n14350), .ZN(n6808) );
  NOR2_X1 U9152 ( .A1(n14349), .A2(n14350), .ZN(n6625) );
  INV_X1 U9153 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7389) );
  AND2_X1 U9154 ( .A1(n12249), .A2(n11496), .ZN(n6626) );
  NOR2_X1 U9155 ( .A1(n11818), .A2(n7067), .ZN(n7066) );
  INV_X1 U9156 ( .A(SI_14_), .ZN(n7053) );
  NAND2_X1 U9157 ( .A1(n11620), .A2(n11484), .ZN(n6627) );
  NAND2_X1 U9158 ( .A1(n14393), .A2(n7363), .ZN(n7367) );
  AND2_X1 U9159 ( .A1(n9580), .A2(n9581), .ZN(n9640) );
  AND2_X1 U9160 ( .A1(n9902), .A2(n7396), .ZN(n6628) );
  XOR2_X1 U9161 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .Z(n6629) );
  NAND2_X1 U9162 ( .A1(n10904), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U9163 ( .A1(n7031), .A2(n6630), .ZN(n6631) );
  INV_X1 U9164 ( .A(n13029), .ZN(n7436) );
  INV_X1 U9165 ( .A(n9605), .ZN(n6804) );
  AND2_X1 U9166 ( .A1(n10370), .A2(n10369), .ZN(n6632) );
  INV_X1 U9167 ( .A(n7635), .ZN(n7708) );
  NOR2_X1 U9168 ( .A1(n10485), .A2(n10251), .ZN(n6633) );
  AND2_X1 U9169 ( .A1(n8177), .A2(n12417), .ZN(n6634) );
  INV_X1 U9170 ( .A(n11660), .ZN(n7141) );
  NAND2_X1 U9171 ( .A1(n9492), .A2(n7193), .ZN(n7195) );
  AND2_X1 U9172 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10203), .ZN(n6635) );
  INV_X1 U9173 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10126) );
  INV_X1 U9174 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9752) );
  INV_X1 U9175 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10646) );
  INV_X1 U9176 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7241) );
  INV_X1 U9177 ( .A(n12019), .ZN(n11984) );
  NAND2_X1 U9178 ( .A1(n12308), .A2(n11655), .ZN(n14896) );
  INV_X1 U9179 ( .A(n12084), .ZN(n6888) );
  AND2_X2 U9180 ( .A1(n9506), .A2(n14684), .ZN(n14764) );
  AND3_X1 U9181 ( .A1(n10159), .A2(n10158), .A3(n10157), .ZN(n10368) );
  NAND2_X1 U9182 ( .A1(n14172), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U9183 ( .A1(n9381), .A2(n9619), .ZN(n12019) );
  INV_X1 U9184 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13006) );
  INV_X1 U9185 ( .A(n14199), .ZN(n6882) );
  INV_X1 U9186 ( .A(n6718), .ZN(n9059) );
  OR2_X1 U9187 ( .A1(n6719), .A2(n9033), .ZN(n6718) );
  XNOR2_X1 U9188 ( .A(n9219), .B(n9218), .ZN(n12091) );
  OR2_X1 U9189 ( .A1(n9843), .A2(n14185), .ZN(n6637) );
  INV_X1 U9190 ( .A(n8368), .ZN(n10649) );
  NAND2_X1 U9191 ( .A1(n8289), .A2(n7987), .ZN(n6638) );
  INV_X1 U9192 ( .A(n10123), .ZN(n11657) );
  INV_X1 U9193 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6793) );
  INV_X1 U9194 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U9195 ( .A1(n8217), .A2(n12687), .ZN(n8218) );
  XNOR2_X2 U9196 ( .A(n6639), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7987) );
  OAI21_X2 U9197 ( .B1(n7928), .B2(n7533), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6639) );
  NAND2_X1 U9198 ( .A1(n7907), .A2(n7908), .ZN(n7928) );
  NAND3_X1 U9199 ( .A1(n6648), .A2(n6645), .A3(n6642), .ZN(n7483) );
  NAND2_X1 U9200 ( .A1(n6649), .A2(n8288), .ZN(n6648) );
  NAND3_X1 U9201 ( .A1(n6653), .A2(n6590), .A3(n6651), .ZN(n6650) );
  AOI22_X1 U9202 ( .A1(n7835), .A2(n7834), .B1(n6655), .B2(n6654), .ZN(n7857)
         );
  INV_X1 U9203 ( .A(n7831), .ZN(n6654) );
  NAND3_X1 U9204 ( .A1(n7441), .A2(n6607), .A3(n7440), .ZN(n6656) );
  NAND2_X1 U9205 ( .A1(n6662), .A2(n7939), .ZN(n6661) );
  OR2_X1 U9206 ( .A1(n7938), .A2(n6663), .ZN(n6662) );
  NAND3_X1 U9207 ( .A1(n7552), .A2(n7549), .A3(n7603), .ZN(n7842) );
  NAND4_X1 U9208 ( .A1(n7552), .A2(n7549), .A3(n7603), .A4(n7843), .ZN(n7863)
         );
  NAND2_X1 U9209 ( .A1(n6665), .A2(n7498), .ZN(n8063) );
  NAND2_X1 U9210 ( .A1(n8026), .A2(n6511), .ZN(n6665) );
  OAI21_X1 U9211 ( .B1(n7745), .B2(n7744), .A(n6547), .ZN(n7505) );
  NAND2_X1 U9212 ( .A1(n6667), .A2(n6666), .ZN(n7745) );
  NAND2_X1 U9213 ( .A1(n7719), .A2(n7718), .ZN(n6667) );
  NAND2_X1 U9214 ( .A1(n12196), .A2(n11485), .ZN(n6670) );
  NAND2_X1 U9215 ( .A1(n12200), .A2(n11588), .ZN(n6671) );
  INV_X1 U9216 ( .A(n10368), .ZN(n6672) );
  NAND2_X1 U9217 ( .A1(n6672), .A2(n12027), .ZN(n11534) );
  AOI21_X2 U9218 ( .B1(n12251), .B2(n6677), .A(n7153), .ZN(n12219) );
  OAI21_X1 U9219 ( .B1(n12132), .B2(n6627), .A(n6514), .ZN(n6678) );
  NAND2_X2 U9220 ( .A1(n11693), .A2(n11696), .ZN(n12132) );
  NAND3_X1 U9221 ( .A1(n6595), .A2(n7157), .A3(n6510), .ZN(n6717) );
  OAI21_X1 U9222 ( .B1(n6687), .B2(n6685), .A(n9988), .ZN(n14395) );
  NAND3_X1 U9223 ( .A1(n6696), .A2(n8539), .A3(n7385), .ZN(n8620) );
  AND3_X2 U9224 ( .A1(n6696), .A2(n8539), .A3(n6694), .ZN(n8616) );
  AND4_X2 U9225 ( .A1(n6585), .A2(n8531), .A3(n6695), .A4(n8532), .ZN(n8539)
         );
  INV_X1 U9226 ( .A(n6701), .ZN(n6700) );
  OAI22_X1 U9227 ( .A1(n13574), .A2(n8762), .B1(n11132), .B2(n8873), .ZN(n6701) );
  NAND2_X4 U9228 ( .A1(n11132), .A2(n6483), .ZN(n13574) );
  XNOR2_X1 U9229 ( .A(n7625), .B(n7624), .ZN(n8761) );
  NOR2_X1 U9230 ( .A1(n10092), .A2(n10098), .ZN(n6716) );
  NAND2_X1 U9231 ( .A1(n9647), .A2(n9648), .ZN(n8389) );
  NAND2_X1 U9232 ( .A1(n8272), .A2(n8307), .ZN(n7197) );
  NAND2_X1 U9233 ( .A1(n8378), .A2(n14695), .ZN(n8307) );
  AND2_X2 U9234 ( .A1(n13817), .A2(n13818), .ZN(n14065) );
  OR2_X2 U9235 ( .A1(n13816), .A2(n13822), .ZN(n13818) );
  AOI21_X1 U9236 ( .B1(n7212), .B2(n7211), .A(n6611), .ZN(n10276) );
  NAND2_X1 U9237 ( .A1(n6739), .A2(n8384), .ZN(n10258) );
  INV_X1 U9238 ( .A(n10262), .ZN(n10259) );
  INV_X1 U9239 ( .A(n14717), .ZN(n6738) );
  INV_X1 U9240 ( .A(n6742), .ZN(n6918) );
  OAI21_X1 U9241 ( .B1(n8224), .B2(n8760), .A(n6743), .ZN(n6742) );
  NAND2_X2 U9242 ( .A1(n7627), .A2(n6483), .ZN(n8224) );
  NAND2_X4 U9243 ( .A1(n13003), .A2(n8933), .ZN(n7627) );
  NAND2_X1 U9244 ( .A1(n7627), .A2(n6601), .ZN(n6743) );
  NAND2_X1 U9245 ( .A1(n8616), .A2(n6603), .ZN(n6746) );
  XNOR2_X2 U9246 ( .A(n6745), .B(n8562), .ZN(n11714) );
  NOR2_X1 U9247 ( .A1(n9804), .A2(n6501), .ZN(n14426) );
  AND2_X1 U9248 ( .A1(n8614), .A2(n8628), .ZN(n9804) );
  NAND2_X1 U9249 ( .A1(n9472), .A2(n9471), .ZN(n9470) );
  NAND2_X1 U9250 ( .A1(n6751), .A2(n6750), .ZN(n10586) );
  OR2_X1 U9251 ( .A1(n7362), .A2(n7360), .ZN(n6751) );
  AOI21_X2 U9252 ( .B1(n13906), .B2(n13907), .A(n11229), .ZN(n13891) );
  NAND2_X1 U9253 ( .A1(n9215), .A2(n9214), .ZN(n9217) );
  NAND2_X1 U9254 ( .A1(n11300), .A2(n11298), .ZN(n6758) );
  OAI21_X1 U9255 ( .B1(n6768), .B2(n11267), .A(n6765), .ZN(n9113) );
  NAND3_X1 U9256 ( .A1(n6770), .A2(n7020), .A3(n6769), .ZN(n8722) );
  NAND3_X1 U9257 ( .A1(n6777), .A2(n6776), .A3(n11794), .ZN(n12127) );
  OAI21_X1 U9258 ( .B1(n9757), .B2(n6631), .A(n7030), .ZN(n6779) );
  XNOR2_X1 U9259 ( .A(n10844), .B(n10596), .ZN(n10845) );
  NAND2_X1 U9260 ( .A1(n9105), .A2(n9106), .ZN(n7010) );
  NAND2_X1 U9261 ( .A1(n6800), .A2(n14345), .ZN(n14349) );
  NAND2_X1 U9262 ( .A1(n6789), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U9263 ( .A1(n6792), .A2(n8509), .ZN(n14343) );
  NOR2_X1 U9264 ( .A1(n14342), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6791) );
  XNOR2_X1 U9265 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n6827) );
  XNOR2_X1 U9266 ( .A(n8504), .B(n7127), .ZN(n14209) );
  NAND2_X1 U9267 ( .A1(n6796), .A2(n8506), .ZN(n14211) );
  XNOR2_X1 U9268 ( .A(n7128), .B(n8517), .ZN(n14175) );
  NAND2_X1 U9269 ( .A1(n8507), .A2(n8508), .ZN(n6818) );
  NAND2_X1 U9270 ( .A1(n14395), .A2(n14394), .ZN(n7176) );
  NAND2_X1 U9271 ( .A1(n11065), .A2(n13505), .ZN(n14011) );
  NAND2_X1 U9272 ( .A1(n10186), .A2(n10185), .ZN(n10392) );
  NAND2_X1 U9273 ( .A1(n7905), .A2(n7904), .ZN(n7924) );
  NAND2_X1 U9274 ( .A1(n6999), .A2(n10084), .ZN(n6998) );
  NAND2_X1 U9275 ( .A1(n12440), .A2(n11732), .ZN(n12446) );
  INV_X1 U9276 ( .A(n7351), .ZN(n7350) );
  NAND2_X1 U9277 ( .A1(n8110), .A2(n8109), .ZN(n8125) );
  NAND2_X1 U9278 ( .A1(n12488), .A2(n12487), .ZN(n12486) );
  XOR2_X2 U9279 ( .A(n12576), .B(n12915), .Z(n12720) );
  OAI21_X1 U9280 ( .B1(n12745), .B2(n6908), .A(n6902), .ZN(n12697) );
  NAND2_X1 U9281 ( .A1(n12029), .A2(n14858), .ZN(n11521) );
  NAND2_X1 U9282 ( .A1(n14825), .A2(n11544), .ZN(n7152) );
  NAND2_X1 U9283 ( .A1(n12265), .A2(n12266), .ZN(n12264) );
  NAND2_X2 U9284 ( .A1(n12175), .A2(n12174), .ZN(n12162) );
  NAND2_X1 U9285 ( .A1(n10008), .A2(n11518), .ZN(n14850) );
  OAI21_X2 U9286 ( .B1(n12289), .B2(n12290), .A(n11566), .ZN(n12277) );
  NAND2_X1 U9287 ( .A1(n14240), .A2(n11552), .ZN(n11265) );
  NAND2_X1 U9288 ( .A1(n14865), .A2(n11508), .ZN(n9763) );
  INV_X1 U9289 ( .A(n6824), .ZN(n7138) );
  NAND2_X1 U9290 ( .A1(n9763), .A2(n11629), .ZN(n14848) );
  NAND2_X1 U9291 ( .A1(n12264), .A2(n11576), .ZN(n12251) );
  AND2_X1 U9292 ( .A1(n9374), .A2(n9373), .ZN(n7134) );
  NAND2_X1 U9293 ( .A1(n14850), .A2(n11520), .ZN(n10160) );
  XNOR2_X1 U9294 ( .A(n6826), .B(n11803), .ZN(n12122) );
  NAND2_X1 U9295 ( .A1(n7142), .A2(n11602), .ZN(n11693) );
  NAND2_X1 U9296 ( .A1(n7152), .A2(n7150), .ZN(n14811) );
  NAND2_X1 U9297 ( .A1(n7138), .A2(n7139), .ZN(n7136) );
  NAND2_X1 U9298 ( .A1(n7196), .A2(n8382), .ZN(n10774) );
  OAI21_X1 U9299 ( .B1(n9888), .B2(n8391), .A(n8392), .ZN(n10753) );
  NAND2_X1 U9300 ( .A1(n7060), .A2(n7059), .ZN(n7327) );
  OAI21_X1 U9301 ( .B1(n7654), .B2(n8783), .A(n8788), .ZN(n7659) );
  OAI21_X1 U9302 ( .B1(n13908), .B2(n13907), .A(n11141), .ZN(n13899) );
  NOR2_X1 U9303 ( .A1(n6807), .A2(n6598), .ZN(n6806) );
  NAND2_X1 U9304 ( .A1(n9535), .A2(n9483), .ZN(n13446) );
  NAND2_X2 U9305 ( .A1(n8577), .A2(n6806), .ZN(n14163) );
  OR2_X1 U9306 ( .A1(n9534), .A2(n11038), .ZN(n9533) );
  NAND2_X1 U9307 ( .A1(n7772), .A2(n7771), .ZN(n7322) );
  OAI21_X1 U9308 ( .B1(n13872), .B2(n7375), .A(n7371), .ZN(n13837) );
  NOR2_X1 U9309 ( .A1(n7360), .A2(n7358), .ZN(n7357) );
  NAND2_X1 U9310 ( .A1(n7369), .A2(n7370), .ZN(n7366) );
  NAND2_X2 U9311 ( .A1(n10242), .A2(n6840), .ZN(n10486) );
  AND2_X2 U9312 ( .A1(n6996), .A2(n6998), .ZN(n10242) );
  NAND3_X1 U9313 ( .A1(n6809), .A2(n12428), .A3(n12533), .ZN(n6838) );
  XNOR2_X1 U9314 ( .A(n11745), .B(n11744), .ZN(n12433) );
  NAND2_X1 U9315 ( .A1(n12446), .A2(n6986), .ZN(n12519) );
  XNOR2_X1 U9316 ( .A(n6525), .B(n10081), .ZN(n10050) );
  NAND2_X2 U9317 ( .A1(n11751), .A2(n11750), .ZN(n12554) );
  NAND2_X1 U9318 ( .A1(n14241), .A2(n10926), .ZN(n14240) );
  INV_X1 U9319 ( .A(n14210), .ZN(n6819) );
  NAND2_X1 U9320 ( .A1(n7010), .A2(n9108), .ZN(n9109) );
  INV_X1 U9321 ( .A(n7556), .ZN(n7555) );
  XNOR2_X1 U9322 ( .A(n8411), .B(n8339), .ZN(n12907) );
  NAND2_X1 U9323 ( .A1(n10300), .A2(n8381), .ZN(n7196) );
  NAND2_X1 U9324 ( .A1(n12755), .A2(n6600), .ZN(n12738) );
  NAND2_X1 U9325 ( .A1(n7515), .A2(n7553), .ZN(n7557) );
  NAND2_X1 U9326 ( .A1(n7145), .A2(n11484), .ZN(n6826) );
  NAND2_X1 U9327 ( .A1(n11507), .A2(n14888), .ZN(n9760) );
  XNOR2_X1 U9328 ( .A(n6816), .B(n11794), .ZN(n12324) );
  NAND2_X1 U9329 ( .A1(n12132), .A2(n12131), .ZN(n6816) );
  NAND2_X1 U9330 ( .A1(n6963), .A2(n7518), .ZN(n12724) );
  INV_X1 U9331 ( .A(n12753), .ZN(n6964) );
  NAND2_X1 U9332 ( .A1(n14394), .A2(n9976), .ZN(n7356) );
  INV_X1 U9333 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7558) );
  XNOR2_X1 U9334 ( .A(n8498), .B(n8499), .ZN(n14203) );
  NAND2_X1 U9335 ( .A1(n7814), .A2(n7813), .ZN(n7817) );
  OR2_X2 U9336 ( .A1(n12433), .A2(n6820), .ZN(n12471) );
  INV_X1 U9337 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9338 ( .A1(n7772), .A2(n7323), .ZN(n6967) );
  NAND2_X1 U9339 ( .A1(n7395), .A2(n6591), .ZN(n6999) );
  NOR2_X2 U9340 ( .A1(n10745), .A2(n10750), .ZN(n9893) );
  NOR2_X2 U9341 ( .A1(n6497), .A2(n12961), .ZN(n12850) );
  NAND2_X2 U9342 ( .A1(n11532), .A2(n11530), .ZN(n14836) );
  NAND3_X1 U9343 ( .A1(n7135), .A2(n7136), .A3(n11532), .ZN(n10161) );
  NAND2_X1 U9344 ( .A1(n11266), .A2(n11556), .ZN(n12293) );
  NOR2_X1 U9345 ( .A1(n11806), .A2(n12115), .ZN(n12318) );
  XNOR2_X1 U9346 ( .A(n8489), .B(n7126), .ZN(n14193) );
  NAND2_X1 U9347 ( .A1(n14193), .A2(n14192), .ZN(n7125) );
  NAND2_X1 U9348 ( .A1(n14975), .A2(n14976), .ZN(n8496) );
  XNOR2_X1 U9349 ( .A(n8423), .B(n8422), .ZN(n8482) );
  INV_X1 U9350 ( .A(n11941), .ZN(n11831) );
  OR2_X1 U9351 ( .A1(n11468), .A2(n9043), .ZN(n8912) );
  AND2_X1 U9352 ( .A1(n12094), .A2(n12105), .ZN(n6831) );
  NAND2_X1 U9353 ( .A1(n12738), .A2(n8409), .ZN(n6963) );
  INV_X1 U9354 ( .A(n12724), .ZN(n7210) );
  NAND3_X1 U9355 ( .A1(n7562), .A2(n7561), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7037) );
  NAND2_X1 U9356 ( .A1(n7701), .A2(n7700), .ZN(n7725) );
  OAI21_X1 U9357 ( .B1(n10735), .B2(n8390), .A(n7213), .ZN(n9888) );
  NAND2_X1 U9358 ( .A1(n7378), .A2(n7376), .ZN(n13995) );
  NAND3_X1 U9359 ( .A1(n14060), .A2(n14061), .A3(n14059), .ZN(n14142) );
  NAND2_X1 U9360 ( .A1(n7034), .A2(n7967), .ZN(n7984) );
  NAND2_X1 U9361 ( .A1(n7035), .A2(n7942), .ZN(n7966) );
  NAND2_X1 U9362 ( .A1(n13794), .A2(n11206), .ZN(n11217) );
  NAND2_X1 U9363 ( .A1(n6833), .A2(n8519), .ZN(n8526) );
  NAND2_X1 U9364 ( .A1(n14175), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U9365 ( .A1(n8472), .A2(n8471), .ZN(n8421) );
  MUX2_X1 U9366 ( .A(n11807), .B(n12318), .S(n14948), .Z(n11808) );
  MUX2_X1 U9367 ( .A(n12319), .B(n12318), .S(n14968), .Z(n12320) );
  NAND2_X1 U9368 ( .A1(n6838), .A2(n6835), .ZN(P2_U3186) );
  NAND2_X1 U9369 ( .A1(n12555), .A2(n11757), .ZN(n12427) );
  NAND2_X1 U9370 ( .A1(n7653), .A2(n7652), .ZN(n7660) );
  NOR2_X2 U9371 ( .A1(n11782), .A2(n6552), .ZN(n12488) );
  NOR2_X2 U9372 ( .A1(n11772), .A2(n6620), .ZN(n11782) );
  OR2_X1 U9373 ( .A1(n10243), .A2(n10244), .ZN(n6840) );
  AND2_X2 U9374 ( .A1(n8582), .A2(n8599), .ZN(n8528) );
  OAI211_X1 U9375 ( .C1(n6572), .C2(n6843), .A(n6842), .B(n6513), .ZN(n7281)
         );
  OR2_X1 U9376 ( .A1(n13544), .A2(n6861), .ZN(n6858) );
  NAND2_X1 U9377 ( .A1(n13544), .A2(n6856), .ZN(n6855) );
  OAI21_X1 U9378 ( .B1(n6548), .B2(n6864), .A(n6863), .ZN(n13487) );
  OAI22_X1 U9379 ( .A1(n13466), .A2(n6608), .B1(n13467), .B2(n6875), .ZN(
        n13469) );
  INV_X1 U9380 ( .A(n13536), .ZN(n6877) );
  NAND2_X1 U9381 ( .A1(n13535), .A2(n6878), .ZN(n6876) );
  OAI22_X1 U9382 ( .A1(n6877), .A2(n6876), .B1(n13538), .B2(n6879), .ZN(n13540) );
  INV_X1 U9383 ( .A(n13537), .ZN(n6879) );
  NAND2_X1 U9384 ( .A1(n9890), .A2(n7311), .ZN(n6892) );
  NAND2_X1 U9385 ( .A1(n9652), .A2(n8321), .ZN(n10737) );
  NAND3_X1 U9386 ( .A1(n8307), .A2(n8272), .A3(n10468), .ZN(n10467) );
  INV_X1 U9387 ( .A(n8329), .ZN(n10676) );
  INV_X1 U9388 ( .A(n7293), .ZN(n6899) );
  OAI211_X2 U9389 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(P2_IR_REG_28__SCAN_IN), 
        .A(n7095), .B(n6901), .ZN(n8933) );
  NAND2_X1 U9390 ( .A1(n12745), .A2(n7517), .ZN(n12726) );
  INV_X1 U9391 ( .A(n7517), .ZN(n6913) );
  XNOR2_X1 U9392 ( .A(n8340), .B(n8339), .ZN(n6915) );
  NAND2_X1 U9393 ( .A1(n6916), .A2(n6593), .ZN(n7062) );
  INV_X2 U9394 ( .A(n14695), .ZN(n9073) );
  NAND2_X1 U9395 ( .A1(n13368), .A2(n13369), .ZN(n6919) );
  NAND2_X1 U9396 ( .A1(n6920), .A2(n7479), .ZN(n13368) );
  NAND2_X1 U9397 ( .A1(n13384), .A2(n7480), .ZN(n6920) );
  NAND2_X1 U9398 ( .A1(n6923), .A2(n6930), .ZN(n9909) );
  AND2_X1 U9399 ( .A1(n6930), .A2(n6604), .ZN(n6922) );
  NAND2_X1 U9400 ( .A1(n6927), .A2(n6932), .ZN(n6923) );
  NAND2_X1 U9401 ( .A1(n14367), .A2(n6924), .ZN(n6930) );
  AOI21_X1 U9402 ( .B1(n14367), .B2(n9730), .A(n6935), .ZN(n6926) );
  NAND2_X1 U9403 ( .A1(n14367), .A2(n6933), .ZN(n6932) );
  INV_X1 U9404 ( .A(n14367), .ZN(n6929) );
  NAND2_X1 U9405 ( .A1(n6934), .A2(n6932), .ZN(n9783) );
  INV_X1 U9406 ( .A(n9782), .ZN(n6931) );
  NOR2_X1 U9407 ( .A1(n6925), .A2(n9781), .ZN(n6933) );
  INV_X1 U9408 ( .A(n9781), .ZN(n6935) );
  OR2_X2 U9409 ( .A1(n13596), .A2(n10556), .ZN(n14076) );
  NAND2_X1 U9410 ( .A1(n13394), .A2(n6950), .ZN(n6948) );
  NAND2_X1 U9411 ( .A1(n6948), .A2(n6949), .ZN(n13326) );
  NAND2_X1 U9412 ( .A1(n7749), .A2(n7748), .ZN(n7752) );
  NAND2_X1 U9413 ( .A1(n7725), .A2(n7724), .ZN(n6953) );
  NAND2_X1 U9414 ( .A1(n12721), .A2(n12720), .ZN(n12913) );
  NAND2_X2 U9415 ( .A1(n7817), .A2(n7816), .ZN(n7837) );
  NAND2_X2 U9416 ( .A1(n11723), .A2(n12501), .ZN(n12507) );
  NAND3_X1 U9417 ( .A1(n7036), .A2(n7038), .A3(n6991), .ZN(n6990) );
  NAND2_X1 U9418 ( .A1(n6993), .A2(n8735), .ZN(n6992) );
  XNOR2_X1 U9419 ( .A(n6995), .B(SI_1_), .ZN(n7597) );
  NAND3_X1 U9420 ( .A1(n6529), .A2(n9580), .A3(n6997), .ZN(n6996) );
  XNOR2_X1 U9421 ( .A(n7001), .B(n7669), .ZN(n9731) );
  OAI21_X1 U9422 ( .B1(n12554), .B2(n7005), .A(n7002), .ZN(n11765) );
  AOI21_X1 U9423 ( .B1(n7390), .B2(n7004), .A(n7003), .ZN(n7002) );
  INV_X1 U9424 ( .A(n11754), .ZN(n7004) );
  NAND2_X1 U9425 ( .A1(n12555), .A2(n7390), .ZN(n12428) );
  NAND2_X2 U9426 ( .A1(n12554), .A2(n11754), .ZN(n12555) );
  NAND3_X1 U9427 ( .A1(n9320), .A2(n9319), .A3(n9335), .ZN(n7007) );
  NAND2_X1 U9428 ( .A1(n7007), .A2(n7006), .ZN(n9583) );
  AOI21_X1 U9429 ( .B1(n7009), .B2(n9335), .A(n6589), .ZN(n7006) );
  INV_X1 U9430 ( .A(n11654), .ZN(n7024) );
  OAI21_X1 U9431 ( .B1(n11654), .B2(n7026), .A(n11657), .ZN(n7025) );
  NAND4_X1 U9432 ( .A1(n11645), .A2(n11644), .A3(n11803), .A4(n6596), .ZN(
        n7033) );
  NAND2_X1 U9433 ( .A1(n7966), .A2(n7965), .ZN(n7034) );
  NAND2_X1 U9434 ( .A1(n7941), .A2(n7940), .ZN(n7035) );
  NAND3_X1 U9435 ( .A1(n7559), .A2(n7558), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7039) );
  OAI211_X1 U9436 ( .C1(n12906), .C2(n14762), .A(n7046), .B(n7048), .ZN(
        P2_U3496) );
  NAND2_X1 U9437 ( .A1(n7817), .A2(n7049), .ZN(n7050) );
  INV_X1 U9438 ( .A(n7327), .ZN(n7058) );
  NAND2_X1 U9439 ( .A1(n6832), .A2(n7656), .ZN(n7059) );
  NAND2_X1 U9440 ( .A1(n7659), .A2(n7658), .ZN(n7060) );
  NAND3_X1 U9441 ( .A1(n7063), .A2(n7062), .A3(n12742), .ZN(n12745) );
  NAND2_X1 U9442 ( .A1(n11911), .A2(n7066), .ZN(n7064) );
  NAND2_X1 U9443 ( .A1(n7064), .A2(n7065), .ZN(n11864) );
  NAND2_X1 U9444 ( .A1(n11948), .A2(n7070), .ZN(n7069) );
  OAI211_X1 U9445 ( .C1(n11948), .C2(n7071), .A(n11956), .B(n7069), .ZN(
        P3_U3169) );
  XNOR2_X1 U9446 ( .A(n11948), .B(n11949), .ZN(n11950) );
  OAI21_X2 U9447 ( .B1(n11959), .B2(n7084), .A(n7081), .ZN(n11873) );
  NAND2_X2 U9448 ( .A1(n10815), .A2(n7094), .ZN(n10999) );
  NAND2_X1 U9449 ( .A1(n10999), .A2(n7092), .ZN(n11809) );
  AOI21_X1 U9450 ( .B1(n7095), .B2(n6566), .A(n7320), .ZN(n7319) );
  NOR2_X2 U9451 ( .A1(n10680), .A2(n10687), .ZN(n10683) );
  OR2_X2 U9452 ( .A1(n10765), .A2(n10671), .ZN(n10680) );
  AND2_X2 U9453 ( .A1(n9893), .A2(n10315), .ZN(n10766) );
  NOR2_X2 U9454 ( .A1(n12823), .A2(n12946), .ZN(n12807) );
  AND2_X2 U9455 ( .A1(n10281), .A2(n14674), .ZN(n10702) );
  NAND2_X1 U9456 ( .A1(n7096), .A2(n6738), .ZN(n10334) );
  INV_X1 U9457 ( .A(n7103), .ZN(n12739) );
  NOR2_X2 U9458 ( .A1(n14428), .A2(n14468), .ZN(n14405) );
  NOR2_X2 U9459 ( .A1(n13810), .A2(n13791), .ZN(n13785) );
  NOR2_X2 U9460 ( .A1(n13969), .A2(n14116), .ZN(n13953) );
  NAND2_X1 U9461 ( .A1(n13880), .A2(n7111), .ZN(n13808) );
  NAND2_X1 U9462 ( .A1(n7134), .A2(n7133), .ZN(n14889) );
  NAND2_X1 U9463 ( .A1(n10160), .A2(n7138), .ZN(n7135) );
  XNOR2_X1 U9464 ( .A(n11480), .B(n12100), .ZN(n7140) );
  NAND2_X1 U9465 ( .A1(n11428), .A2(n7143), .ZN(n7142) );
  NAND2_X1 U9466 ( .A1(n12132), .A2(n11481), .ZN(n7145) );
  NOR2_X1 U9467 ( .A1(n11647), .A2(n11476), .ZN(n7149) );
  OAI21_X1 U9468 ( .B1(n13821), .B2(n7164), .A(n6521), .ZN(n13794) );
  NAND2_X1 U9469 ( .A1(n7161), .A2(n7159), .ZN(n13796) );
  NAND2_X1 U9470 ( .A1(n13821), .A2(n6521), .ZN(n7161) );
  NAND2_X1 U9471 ( .A1(n7165), .A2(n7166), .ZN(n10966) );
  NAND2_X4 U9472 ( .A1(n14163), .A2(n8632), .ZN(n11132) );
  NAND2_X1 U9473 ( .A1(n9471), .A2(n13446), .ZN(n7172) );
  NAND2_X1 U9474 ( .A1(n7176), .A2(n7174), .ZN(n10186) );
  AND3_X2 U9475 ( .A1(n8539), .A2(n6533), .A3(n7179), .ZN(n7178) );
  OAI21_X1 U9476 ( .B1(n13938), .B2(n7183), .A(n7180), .ZN(n13908) );
  AND4_X2 U9477 ( .A1(n6544), .A2(n7550), .A3(n7549), .A4(n7603), .ZN(n7553)
         );
  INV_X1 U9478 ( .A(n12864), .ZN(n7238) );
  OAI21_X1 U9479 ( .B1(n7243), .B2(n11613), .A(n7242), .ZN(n11616) );
  NAND2_X1 U9480 ( .A1(n7246), .A2(n7247), .ZN(n13513) );
  NAND2_X1 U9481 ( .A1(n13501), .A2(n7249), .ZN(n7246) );
  NAND2_X1 U9482 ( .A1(n7258), .A2(n7256), .ZN(n13551) );
  NAND2_X1 U9483 ( .A1(n13547), .A2(n7259), .ZN(n7258) );
  NAND2_X1 U9484 ( .A1(n7269), .A2(n7267), .ZN(n13474) );
  NAND2_X1 U9485 ( .A1(n13469), .A2(n7270), .ZN(n7269) );
  NAND2_X1 U9486 ( .A1(n13493), .A2(n13494), .ZN(n13492) );
  NAND2_X1 U9487 ( .A1(n7281), .A2(n7282), .ZN(n13566) );
  AND2_X1 U9488 ( .A1(n8290), .A2(n7284), .ZN(n8295) );
  XNOR2_X1 U9489 ( .A(n7545), .B(n7284), .ZN(n8232) );
  NAND2_X1 U9490 ( .A1(n7286), .A2(n7285), .ZN(n7295) );
  AOI21_X1 U9491 ( .B1(n10676), .B2(n14264), .A(n8330), .ZN(n10652) );
  NOR2_X1 U9492 ( .A1(n10651), .A2(n10687), .ZN(n7293) );
  OR2_X1 U9493 ( .A1(n12966), .A2(n12547), .ZN(n7294) );
  NAND3_X1 U9494 ( .A1(n7298), .A2(n7297), .A3(n6606), .ZN(n10278) );
  NAND2_X1 U9495 ( .A1(n8309), .A2(n7299), .ZN(n7298) );
  NAND2_X1 U9496 ( .A1(n8320), .A2(n7308), .ZN(n9652) );
  AOI21_X2 U9497 ( .B1(n7318), .B2(n7317), .A(n7316), .ZN(n12801) );
  INV_X1 U9498 ( .A(n7669), .ZN(n7328) );
  NAND2_X1 U9499 ( .A1(n7697), .A2(n7696), .ZN(n7701) );
  NAND2_X1 U9500 ( .A1(n8185), .A2(n7332), .ZN(n7330) );
  NAND2_X1 U9501 ( .A1(n7331), .A2(n7337), .ZN(n8175) );
  NAND2_X1 U9502 ( .A1(n8185), .A2(n7339), .ZN(n7331) );
  INV_X1 U9503 ( .A(n7337), .ZN(n7335) );
  NAND2_X1 U9504 ( .A1(n7343), .A2(n7986), .ZN(n8008) );
  NAND2_X1 U9505 ( .A1(n7883), .A2(n7346), .ZN(n7344) );
  OAI21_X1 U9506 ( .B1(n7837), .B2(n7836), .A(n7838), .ZN(n7861) );
  NAND2_X1 U9507 ( .A1(n7836), .A2(n7838), .ZN(n7352) );
  NAND3_X1 U9508 ( .A1(n8285), .A2(n8283), .A3(n7355), .ZN(n7354) );
  NAND2_X1 U9509 ( .A1(n7356), .A2(n10193), .ZN(n7369) );
  AND2_X1 U9510 ( .A1(n7364), .A2(n13617), .ZN(n7362) );
  NAND2_X1 U9511 ( .A1(n10975), .A2(n7379), .ZN(n7378) );
  OAI21_X1 U9512 ( .B1(n9804), .B2(n6584), .A(n14461), .ZN(n7382) );
  NAND2_X1 U9513 ( .A1(n8616), .A2(n7384), .ZN(n8569) );
  OAI21_X2 U9514 ( .B1(n10486), .B2(n7393), .A(n7392), .ZN(n11720) );
  OR2_X1 U9515 ( .A1(n9905), .A2(n7398), .ZN(n7397) );
  INV_X1 U9516 ( .A(n9903), .ZN(n7400) );
  NAND2_X1 U9517 ( .A1(n7555), .A2(n7401), .ZN(n7569) );
  NAND3_X1 U9518 ( .A1(n7403), .A2(n9264), .A3(n7402), .ZN(n9318) );
  NAND3_X1 U9519 ( .A1(n9256), .A2(n9258), .A3(n9257), .ZN(n7403) );
  NAND2_X2 U9520 ( .A1(n9079), .A2(n9096), .ZN(n9257) );
  AND2_X1 U9521 ( .A1(n9125), .A2(n9124), .ZN(n9256) );
  NAND2_X1 U9522 ( .A1(n12281), .A2(n7406), .ZN(n7404) );
  NAND2_X1 U9523 ( .A1(n7404), .A2(n7405), .ZN(n12259) );
  OAI21_X1 U9524 ( .B1(n9768), .B2(n7411), .A(n7409), .ZN(n14851) );
  INV_X1 U9525 ( .A(n11627), .ZN(n7410) );
  INV_X1 U9526 ( .A(n7412), .ZN(n7411) );
  NAND2_X1 U9527 ( .A1(n14875), .A2(n7412), .ZN(n10028) );
  NAND2_X1 U9528 ( .A1(n9768), .A2(n11627), .ZN(n14875) );
  AOI21_X1 U9529 ( .B1(n12212), .B2(n6597), .A(n7414), .ZN(n12181) );
  AND2_X1 U9530 ( .A1(n8683), .A2(n8678), .ZN(n8681) );
  MUX2_X1 U9531 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7426), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n7425) );
  NAND2_X1 U9532 ( .A1(n7557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9533 ( .A1(n14288), .A2(n7430), .ZN(n7427) );
  OAI211_X1 U9534 ( .C1(n14288), .C2(n7431), .A(n7427), .B(n7428), .ZN(n13346)
         );
  NAND2_X1 U9535 ( .A1(n7796), .A2(n7795), .ZN(n7440) );
  NAND2_X1 U9536 ( .A1(n7794), .A2(n7793), .ZN(n7441) );
  NAND2_X1 U9537 ( .A1(n7876), .A2(n7451), .ZN(n7450) );
  NAND2_X1 U9538 ( .A1(n7450), .A2(n6605), .ZN(n7917) );
  NAND2_X1 U9539 ( .A1(n13336), .A2(n13337), .ZN(n7478) );
  NAND2_X1 U9540 ( .A1(n7478), .A2(n13099), .ZN(n13407) );
  NAND2_X1 U9541 ( .A1(n7483), .A2(n8293), .ZN(n8306) );
  NAND2_X1 U9542 ( .A1(n8066), .A2(n6610), .ZN(n7486) );
  OAI21_X1 U9543 ( .B1(n7490), .B2(n7492), .A(n7491), .ZN(n8002) );
  INV_X1 U9544 ( .A(n7980), .ZN(n7496) );
  INV_X1 U9545 ( .A(n7963), .ZN(n7497) );
  INV_X1 U9546 ( .A(n8027), .ZN(n7502) );
  OAI211_X1 U9547 ( .C1(n13574), .C2(n6991), .A(n7509), .B(n7508), .ZN(n8586)
         );
  OR2_X1 U9548 ( .A1(n11132), .A2(n8855), .ZN(n7508) );
  NAND2_X2 U9549 ( .A1(n11132), .A2(n8585), .ZN(n9977) );
  OAI21_X1 U9550 ( .B1(n11687), .B2(n14873), .A(n11686), .ZN(n11688) );
  NAND2_X1 U9551 ( .A1(n9445), .A2(n9444), .ZN(n9510) );
  OR2_X1 U9552 ( .A1(n9364), .A2(n9363), .ZN(n9618) );
  INV_X1 U9553 ( .A(n12405), .ZN(n12313) );
  NAND2_X2 U9554 ( .A1(n10138), .A2(n10057), .ZN(n10128) );
  NAND2_X1 U9555 ( .A1(n14871), .A2(n11892), .ZN(n9445) );
  NOR2_X2 U9556 ( .A1(n13881), .A2(n14083), .ZN(n13880) );
  NAND2_X1 U9557 ( .A1(n7647), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7572) );
  OR2_X1 U9558 ( .A1(n8661), .A2(n13990), .ZN(n13427) );
  OR2_X1 U9559 ( .A1(n14076), .A2(n13990), .ZN(n11048) );
  INV_X1 U9560 ( .A(n13990), .ZN(n13928) );
  NOR2_X1 U9561 ( .A1(n12906), .A2(n12858), .ZN(n8377) );
  AND2_X1 U9562 ( .A1(n8413), .A2(n8368), .ZN(n9066) );
  INV_X1 U9563 ( .A(n8232), .ZN(n8413) );
  AND2_X1 U9564 ( .A1(n13800), .A2(n11239), .ZN(n14056) );
  NAND2_X1 U9565 ( .A1(n7647), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9566 ( .A1(n9066), .A2(n8933), .ZN(n12777) );
  AND2_X1 U9567 ( .A1(n7884), .A2(n7885), .ZN(n7907) );
  NAND2_X1 U9568 ( .A1(n8906), .A2(n8907), .ZN(n9828) );
  INV_X1 U9569 ( .A(n7608), .ZN(n7611) );
  XNOR2_X1 U9570 ( .A(n13431), .B(n8586), .ZN(n9528) );
  INV_X1 U9571 ( .A(n13432), .ZN(n9158) );
  NAND2_X1 U9572 ( .A1(n12532), .A2(n11742), .ZN(n11745) );
  AND2_X2 U9573 ( .A1(n10151), .A2(n10150), .ZN(n14837) );
  NAND2_X1 U9574 ( .A1(n11501), .A2(n11844), .ZN(n9444) );
  NAND2_X1 U9575 ( .A1(n14870), .A2(n14887), .ZN(n14871) );
  AND3_X1 U9576 ( .A1(n11348), .A2(n9437), .A3(n11613), .ZN(n14890) );
  INV_X1 U9577 ( .A(n14301), .ZN(n14331) );
  INV_X1 U9578 ( .A(n14094), .ZN(n13915) );
  INV_X1 U9579 ( .A(n6478), .ZN(n8219) );
  INV_X1 U9580 ( .A(n14680), .ZN(n12889) );
  AND2_X2 U9581 ( .A1(n8369), .A2(n12886), .ZN(n14680) );
  OR3_X1 U9582 ( .A1(n9089), .A2(n13003), .A3(n12773), .ZN(n7510) );
  AND2_X1 U9583 ( .A1(n11913), .A2(n14242), .ZN(n7511) );
  AND4_X1 U9584 ( .A1(n8536), .A2(n6851), .A3(n8535), .A4(n8625), .ZN(n7512)
         );
  OR2_X1 U9585 ( .A1(n14315), .A2(n14016), .ZN(n7513) );
  INV_X1 U9586 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9107) );
  OR2_X1 U9587 ( .A1(n12907), .A2(n12893), .ZN(n7516) );
  OR2_X1 U9588 ( .A1(n7100), .A2(n12758), .ZN(n7517) );
  OR2_X1 U9589 ( .A1(n7100), .A2(n12728), .ZN(n7518) );
  XOR2_X1 U9590 ( .A(n8524), .B(n8523), .Z(n7519) );
  AND2_X1 U9591 ( .A1(n7862), .A2(n7841), .ZN(n7520) );
  INV_X1 U9592 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9001) );
  INV_X1 U9593 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10201) );
  INV_X1 U9594 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9835) );
  INV_X1 U9595 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9824) );
  INV_X1 U9596 ( .A(n14270), .ZN(n10671) );
  INV_X1 U9597 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10481) );
  INV_X1 U9598 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7600) );
  OAI21_X1 U9599 ( .B1(n13911), .B2(n11153), .A(n11140), .ZN(n13651) );
  INV_X1 U9600 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8494) );
  AND2_X1 U9601 ( .A1(n7785), .A2(n7784), .ZN(n7521) );
  NAND2_X2 U9602 ( .A1(n9631), .A2(n14902), .ZN(n14228) );
  AND3_X1 U9603 ( .A1(n13525), .A2(n13950), .A3(n13524), .ZN(n7522) );
  INV_X1 U9604 ( .A(n12091), .ZN(n12100) );
  AND3_X1 U9605 ( .A1(n8215), .A2(n8214), .A3(n8213), .ZN(n7523) );
  AND2_X1 U9606 ( .A1(n10179), .A2(n10178), .ZN(n7524) );
  NOR2_X1 U9607 ( .A1(n10860), .A2(n10797), .ZN(n7525) );
  OR2_X1 U9608 ( .A1(n14727), .A2(n12585), .ZN(n7526) );
  OR2_X1 U9609 ( .A1(n14108), .A2(n13531), .ZN(n7527) );
  AND2_X1 U9610 ( .A1(n13428), .A2(n9153), .ZN(n7528) );
  INV_X1 U9611 ( .A(n14814), .ZN(n10920) );
  AND2_X1 U9612 ( .A1(n13438), .A2(n13600), .ZN(n13435) );
  AOI21_X1 U9613 ( .B1(n6477), .B2(n13431), .A(n9158), .ZN(n13444) );
  INV_X1 U9614 ( .A(n7609), .ZN(n7610) );
  AOI22_X1 U9615 ( .A1(n10785), .A2(n6486), .B1(n7707), .B2(n12587), .ZN(n7642) );
  NAND2_X1 U9616 ( .A1(n13498), .A2(n13497), .ZN(n13501) );
  INV_X1 U9617 ( .A(n7792), .ZN(n7793) );
  OAI21_X1 U9618 ( .B1(n7857), .B2(n7856), .A(n7855), .ZN(n7858) );
  INV_X1 U9619 ( .A(n7962), .ZN(n7964) );
  INV_X1 U9620 ( .A(n8060), .ZN(n8061) );
  OAI21_X1 U9621 ( .B1(n8217), .B2(n8219), .A(n8218), .ZN(n8244) );
  INV_X1 U9622 ( .A(n10759), .ZN(n8326) );
  INV_X1 U9623 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8554) );
  AND2_X1 U9624 ( .A1(n14245), .A2(n11646), .ZN(n11479) );
  NAND2_X1 U9625 ( .A1(n11792), .A2(n11788), .ZN(n11791) );
  INV_X1 U9626 ( .A(n14872), .ZN(n11627) );
  NOR2_X1 U9627 ( .A1(n7523), .A2(n8254), .ZN(n8255) );
  AND4_X1 U9628 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n8558)
         );
  INV_X1 U9629 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11933) );
  INV_X1 U9630 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n11952) );
  INV_X1 U9631 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n11340) );
  INV_X1 U9632 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n10952) );
  INV_X1 U9633 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8901) );
  INV_X1 U9634 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7848) );
  INV_X1 U9635 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7554) );
  INV_X1 U9636 ( .A(n9728), .ZN(n9729) );
  INV_X1 U9637 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10577) );
  NOR2_X1 U9638 ( .A1(n14301), .A2(n13660), .ZN(n10804) );
  INV_X1 U9639 ( .A(n8183), .ZN(n8145) );
  INV_X1 U9640 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8529) );
  INV_X1 U9641 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10163) );
  INV_X1 U9642 ( .A(n11912), .ZN(n11813) );
  INV_X1 U9643 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10010) );
  INV_X1 U9644 ( .A(n9639), .ZN(n9622) );
  NOR2_X1 U9645 ( .A1(n10949), .A2(n7511), .ZN(n10950) );
  OR2_X1 U9646 ( .A1(n9623), .A2(n12100), .ZN(n9766) );
  INV_X1 U9647 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7784) );
  INV_X1 U9648 ( .A(n9323), .ZN(n9319) );
  NAND2_X1 U9649 ( .A1(n7954), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7993) );
  NOR2_X1 U9650 ( .A1(n12996), .A2(n7576), .ZN(n7577) );
  OR2_X1 U9651 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  OR2_X1 U9652 ( .A1(n12946), .A2(n12536), .ZN(n8336) );
  NOR2_X1 U9653 ( .A1(n12853), .A2(n12861), .ZN(n8332) );
  NOR2_X1 U9654 ( .A1(n11125), .A2(n11124), .ZN(n11133) );
  INV_X1 U9655 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9991) );
  INV_X1 U9656 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8570) );
  OR2_X1 U9657 ( .A1(n9568), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9000) );
  INV_X1 U9658 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7560) );
  INV_X1 U9659 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n8435) );
  AND2_X1 U9660 ( .A1(n10164), .A2(n10163), .ZN(n10373) );
  INV_X1 U9661 ( .A(n11940), .ZN(n11830) );
  OR2_X1 U9662 ( .A1(n9461), .A2(n9382), .ZN(n9384) );
  INV_X1 U9663 ( .A(n10217), .ZN(n10922) );
  INV_X1 U9664 ( .A(n14191), .ZN(n11268) );
  AND2_X1 U9665 ( .A1(n9029), .A2(n9028), .ZN(n9037) );
  AND4_X1 U9666 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n12124)
         );
  INV_X1 U9667 ( .A(n11666), .ZN(n12266) );
  OR2_X1 U9668 ( .A1(n10613), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10823) );
  NOR2_X1 U9669 ( .A1(n14886), .A2(n14901), .ZN(n9383) );
  INV_X1 U9670 ( .A(n11804), .ZN(n11656) );
  AND2_X1 U9671 ( .A1(n10939), .A2(n10938), .ZN(n11812) );
  INV_X1 U9672 ( .A(n14896), .ZN(n14873) );
  AND2_X1 U9673 ( .A1(n9767), .A2(n9766), .ZN(n14900) );
  INV_X1 U9674 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9338) );
  OR2_X1 U9675 ( .A1(n10250), .A2(n10249), .ZN(n10251) );
  AND2_X1 U9676 ( .A1(n12477), .A2(n11749), .ZN(n12473) );
  INV_X1 U9677 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12524) );
  INV_X1 U9678 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11775) );
  AND2_X1 U9679 ( .A1(n8157), .A2(n8156), .ZN(n11766) );
  AND2_X1 U9680 ( .A1(n7933), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7954) );
  OAI21_X1 U9681 ( .B1(n8300), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8296) );
  AND2_X1 U9682 ( .A1(n10796), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10860) );
  INV_X1 U9683 ( .A(n13835), .ZN(n13321) );
  INV_X1 U9684 ( .A(n13858), .ZN(n13340) );
  INV_X1 U9685 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10517) );
  AND2_X1 U9686 ( .A1(n11191), .A2(n11207), .ZN(n13825) );
  AND2_X1 U9687 ( .A1(n11133), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11146) );
  INV_X1 U9688 ( .A(n14136), .ZN(n9170) );
  NAND2_X1 U9689 ( .A1(n13835), .A2(n14416), .ZN(n11214) );
  INV_X1 U9690 ( .A(n13658), .ZN(n10973) );
  INV_X1 U9691 ( .A(n13662), .ZN(n10565) );
  NAND2_X1 U9692 ( .A1(n7924), .A2(n7923), .ZN(n7941) );
  OR2_X1 U9693 ( .A1(n9619), .A2(n11657), .ZN(n9029) );
  NOR2_X1 U9694 ( .A1(n10070), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U9695 ( .A1(n11811), .A2(n11810), .ZN(n11911) );
  INV_X1 U9696 ( .A(n12009), .ZN(n11999) );
  OR2_X1 U9697 ( .A1(n9825), .A2(n12116), .ZN(n11472) );
  AND4_X1 U9698 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n12155) );
  AND4_X1 U9699 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n12224) );
  AND4_X1 U9700 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n12010) );
  INV_X1 U9701 ( .A(n12113), .ZN(n14792) );
  AND2_X1 U9702 ( .A1(n9037), .A2(n9036), .ZN(n14801) );
  AND2_X1 U9703 ( .A1(n9037), .A2(n12069), .ZN(n14788) );
  AND2_X1 U9704 ( .A1(n11620), .A2(n11619), .ZN(n11803) );
  INV_X1 U9705 ( .A(n14900), .ZN(n14878) );
  NAND2_X1 U9706 ( .A1(n11290), .A2(n11289), .ZN(n12374) );
  INV_X1 U9707 ( .A(n14867), .ZN(n14891) );
  INV_X1 U9708 ( .A(n12117), .ZN(n14861) );
  NAND2_X1 U9709 ( .A1(n12100), .A2(n9639), .ZN(n14901) );
  AND2_X1 U9710 ( .A1(n9621), .A2(n9620), .ZN(n12317) );
  AND2_X1 U9711 ( .A1(n14225), .A2(n14224), .ZN(n14247) );
  OR2_X1 U9712 ( .A1(n14901), .A2(n11804), .ZN(n12344) );
  AND2_X1 U9713 ( .A1(n14900), .A2(n12344), .ZN(n12386) );
  INV_X1 U9714 ( .A(n12386), .ZN(n14946) );
  INV_X1 U9715 ( .A(n12344), .ZN(n14937) );
  NAND2_X1 U9716 ( .A1(n9344), .A2(n8697), .ZN(n9347) );
  AND2_X1 U9717 ( .A1(n8193), .A2(n8192), .ZN(n12716) );
  INV_X1 U9718 ( .A(n12837), .ZN(n12956) );
  INV_X1 U9719 ( .A(n12538), .ZN(n12558) );
  INV_X1 U9720 ( .A(n12444), .ZN(n12429) );
  INV_X1 U9721 ( .A(n12571), .ZN(n12533) );
  AND4_X1 U9722 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n12729)
         );
  INV_X1 U9723 ( .A(n14633), .ZN(n14652) );
  NAND2_X1 U9724 ( .A1(n8935), .A2(n8934), .ZN(n14661) );
  INV_X1 U9725 ( .A(n14657), .ZN(n14637) );
  INV_X1 U9726 ( .A(n12777), .ZN(n12880) );
  INV_X1 U9727 ( .A(n12893), .ZN(n14677) );
  NAND2_X1 U9728 ( .A1(n8342), .A2(n8341), .ZN(n12879) );
  INV_X1 U9729 ( .A(n14684), .ZN(n9491) );
  NAND2_X1 U9730 ( .A1(n8231), .A2(n6489), .ZN(n14740) );
  INV_X1 U9731 ( .A(n6485), .ZN(n14745) );
  AND2_X1 U9732 ( .A1(n9490), .A2(n14686), .ZN(n9506) );
  INV_X1 U9733 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7908) );
  INV_X1 U9734 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7662) );
  INV_X1 U9735 ( .A(n14461), .ZN(n13608) );
  INV_X1 U9736 ( .A(n13332), .ZN(n14373) );
  NAND2_X1 U9737 ( .A1(n8642), .A2(n8848), .ZN(n14015) );
  INV_X1 U9738 ( .A(n11208), .ZN(n11153) );
  AND4_X1 U9739 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n11073), .ZN(
        n14014) );
  INV_X1 U9740 ( .A(n14386), .ZN(n13737) );
  INV_X1 U9741 ( .A(n13772), .ZN(n14383) );
  AND2_X1 U9742 ( .A1(n8899), .A2(n14163), .ZN(n14386) );
  INV_X1 U9743 ( .A(n14013), .ZN(n14413) );
  INV_X1 U9744 ( .A(n14015), .ZN(n14416) );
  INV_X1 U9745 ( .A(n14022), .ZN(n14432) );
  NAND2_X1 U9746 ( .A1(n13807), .A2(n14421), .ZN(n14419) );
  INV_X1 U9747 ( .A(n14025), .ZN(n14433) );
  NOR2_X1 U9748 ( .A1(n14136), .A2(n11041), .ZN(n11049) );
  INV_X1 U9749 ( .A(n14411), .ZN(n14501) );
  INV_X1 U9750 ( .A(n14515), .ZN(n14316) );
  NAND2_X1 U9751 ( .A1(n13824), .A2(n14503), .ZN(n14515) );
  AND2_X1 U9752 ( .A1(n11048), .A2(n11047), .ZN(n14137) );
  OAI211_X1 U9753 ( .C1(P1_B_REG_SCAN_IN), .C2(n10994), .A(n8646), .B(n8647), 
        .ZN(n8807) );
  INV_X1 U9754 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8621) );
  AND2_X1 U9755 ( .A1(n9274), .A2(n9006), .ZN(n10855) );
  INV_X1 U9756 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8599) );
  AND2_X1 U9757 ( .A1(n9030), .A2(n9029), .ZN(n14780) );
  NOR2_X1 U9758 ( .A1(n9593), .A2(n11657), .ZN(n12003) );
  INV_X1 U9759 ( .A(n12017), .ZN(n11994) );
  INV_X1 U9760 ( .A(n12155), .ZN(n12024) );
  INV_X1 U9761 ( .A(n11961), .ZN(n12213) );
  INV_X1 U9762 ( .A(n12010), .ZN(n12297) );
  INV_X1 U9763 ( .A(n14780), .ZN(n14804) );
  INV_X1 U9764 ( .A(n14801), .ZN(n12109) );
  OR2_X1 U9765 ( .A1(n12031), .A2(n9022), .ZN(n12113) );
  AND2_X1 U9766 ( .A1(n12285), .A2(n12284), .ZN(n12381) );
  INV_X1 U9767 ( .A(n14968), .ZN(n14965) );
  AND2_X1 U9768 ( .A1(n9465), .A2(n9464), .ZN(n14949) );
  OR2_X1 U9769 ( .A1(n11031), .A2(n12404), .ZN(n11032) );
  INV_X1 U9770 ( .A(n9352), .ZN(n12405) );
  INV_X1 U9771 ( .A(SI_26_), .ZN(n11430) );
  INV_X1 U9772 ( .A(SI_20_), .ZN(n11361) );
  INV_X1 U9773 ( .A(SI_12_), .ZN(n10935) );
  NAND2_X1 U9774 ( .A1(n9091), .A2(n9070), .ZN(n12571) );
  INV_X1 U9775 ( .A(n12729), .ZN(n12576) );
  INV_X1 U9776 ( .A(n12525), .ZN(n12846) );
  INV_X1 U9777 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14562) );
  OR2_X1 U9778 ( .A1(n8954), .A2(n8955), .ZN(n14633) );
  OR2_X1 U9779 ( .A1(n8935), .A2(P2_U3088), .ZN(n14665) );
  INV_X1 U9780 ( .A(n12889), .ZN(n12858) );
  NAND2_X1 U9781 ( .A1(n12889), .A2(n8416), .ZN(n12893) );
  INV_X1 U9782 ( .A(n14779), .ZN(n14777) );
  AND2_X2 U9783 ( .A1(n9506), .A2(n9491), .ZN(n14779) );
  AND2_X1 U9784 ( .A1(n14280), .A2(n14279), .ZN(n14287) );
  AND3_X1 U9785 ( .A1(n14724), .A2(n14723), .A3(n14722), .ZN(n14770) );
  INV_X1 U9786 ( .A(n14764), .ZN(n14762) );
  OR2_X1 U9787 ( .A1(n14687), .A2(n14681), .ZN(n14682) );
  INV_X1 U9788 ( .A(n13490), .ZN(n14216) );
  NAND2_X1 U9789 ( .A1(n9168), .A2(n9167), .ZN(n13425) );
  OAI21_X1 U9790 ( .B1(n13893), .B2(n11153), .A(n11152), .ZN(n13876) );
  OR2_X1 U9791 ( .A1(n11110), .A2(n11109), .ZN(n13965) );
  OR2_X1 U9792 ( .A1(n8849), .A2(n8848), .ZN(n13772) );
  INV_X1 U9793 ( .A(n14387), .ZN(n13773) );
  NAND2_X1 U9794 ( .A1(n8847), .A2(n8845), .ZN(n14391) );
  AND2_X2 U9795 ( .A1(n11049), .A2(n14137), .ZN(n14534) );
  INV_X1 U9796 ( .A(n14519), .ZN(n14517) );
  AND2_X2 U9797 ( .A1(n14138), .A2(n14137), .ZN(n14519) );
  INV_X1 U9798 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n11042) );
  INV_X1 U9799 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11156) );
  INV_X1 U9800 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10203) );
  INV_X1 U9801 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9110) );
  INV_X1 U9802 ( .A(n12031), .ZN(P3_U3897) );
  AND2_X1 U9803 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8932), .ZN(P2_U3947) );
  INV_X1 U9804 ( .A(n13668), .ZN(P1_U4016) );
  OR4_X1 U9805 ( .A1(n8669), .A2(n8668), .A3(n8667), .A4(n8666), .ZN(P1_U3290)
         );
  XNOR2_X1 U9806 ( .A(n8526), .B(n8525), .ZN(SUB_1596_U4) );
  NOR2_X2 U9807 ( .A1(n7863), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7884) );
  INV_X1 U9808 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7532) );
  NAND3_X1 U9809 ( .A1(n7946), .A2(n7532), .A3(n7969), .ZN(n7533) );
  NAND2_X1 U9810 ( .A1(n7884), .A2(n7551), .ZN(n7538) );
  NAND2_X1 U9811 ( .A1(n7538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7537) );
  INV_X1 U9812 ( .A(n7538), .ZN(n7540) );
  NAND2_X1 U9813 ( .A1(n7540), .A2(n7539), .ZN(n7542) );
  NAND2_X1 U9814 ( .A1(n7542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7541) );
  MUX2_X1 U9815 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7541), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7544) );
  INV_X1 U9816 ( .A(n8290), .ZN(n7543) );
  AND3_X2 U9817 ( .A1(n8231), .A2(n8368), .A3(n6489), .ZN(n7707) );
  INV_X1 U9818 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7547) );
  INV_X1 U9819 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7546) );
  INV_X1 U9820 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7559) );
  INV_X1 U9821 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7561) );
  INV_X1 U9822 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8735) );
  INV_X1 U9823 ( .A(n6483), .ZN(n8585) );
  AND2_X1 U9824 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U9825 ( .A1(n8585), .A2(n7563), .ZN(n8593) );
  AND2_X1 U9826 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9827 ( .A1(n6483), .A2(n7564), .ZN(n7584) );
  NAND2_X1 U9828 ( .A1(n8593), .A2(n7584), .ZN(n7598) );
  XNOR2_X1 U9829 ( .A(n7597), .B(n7598), .ZN(n8760) );
  NAND2_X1 U9830 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7565) );
  XNOR2_X1 U9831 ( .A(n7565), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U9832 ( .A1(n8929), .A2(n8937), .ZN(n7566) );
  INV_X1 U9833 ( .A(n11033), .ZN(n7578) );
  NAND2_X1 U9834 ( .A1(n7646), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U9835 ( .A1(n7635), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U9836 ( .A1(n7514), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7571) );
  NAND4_X2 U9837 ( .A1(n7574), .A2(n7573), .A3(n7572), .A4(n7571), .ZN(n8271)
         );
  NAND2_X1 U9838 ( .A1(n6481), .A2(n8271), .ZN(n7575) );
  OAI21_X1 U9839 ( .B1(n6482), .B2(n9073), .A(n7575), .ZN(n7609) );
  NAND2_X1 U9840 ( .A1(n7514), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9841 ( .A1(n7635), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7580) );
  INV_X1 U9842 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9843 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  NAND2_X1 U9844 ( .A1(n6484), .A2(SI_0_), .ZN(n7583) );
  NAND2_X1 U9845 ( .A1(n7583), .A2(n8833), .ZN(n7585) );
  NAND2_X1 U9846 ( .A1(n7585), .A2(n7584), .ZN(n13014) );
  MUX2_X1 U9847 ( .A(n8964), .B(n13014), .S(n7627), .Z(n8370) );
  NAND2_X1 U9848 ( .A1(n8273), .A2(n8370), .ZN(n7586) );
  NAND2_X1 U9849 ( .A1(n7586), .A2(n7707), .ZN(n7590) );
  NAND2_X1 U9850 ( .A1(n8368), .A2(n10555), .ZN(n9071) );
  AND2_X1 U9851 ( .A1(n8370), .A2(n9071), .ZN(n7588) );
  INV_X1 U9852 ( .A(n9071), .ZN(n8415) );
  NAND2_X1 U9853 ( .A1(n8415), .A2(n10477), .ZN(n7587) );
  OAI211_X1 U9854 ( .C1(n8273), .C2(n7588), .A(n6478), .B(n7587), .ZN(n7589)
         );
  NAND2_X1 U9855 ( .A1(n7590), .A2(n7589), .ZN(n7608) );
  NAND2_X1 U9856 ( .A1(n7609), .A2(n7608), .ZN(n7592) );
  OAI22_X1 U9857 ( .A1(n6482), .A2(n8378), .B1(n8219), .B2(n9073), .ZN(n7591)
         );
  NAND2_X1 U9858 ( .A1(n7592), .A2(n7591), .ZN(n7614) );
  NAND2_X1 U9859 ( .A1(n7514), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9860 ( .A1(n7635), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9861 ( .A1(n7646), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7593) );
  INV_X1 U9862 ( .A(SI_1_), .ZN(n9431) );
  XNOR2_X1 U9863 ( .A(n7621), .B(n6832), .ZN(n7620) );
  XNOR2_X1 U9864 ( .A(n7620), .B(SI_2_), .ZN(n8601) );
  NOR2_X1 U9865 ( .A1(n7601), .A2(n7929), .ZN(n7602) );
  MUX2_X1 U9866 ( .A(n7929), .B(n7602), .S(P2_IR_REG_2__SCAN_IN), .Z(n7604) );
  NOR2_X1 U9867 ( .A1(n7604), .A2(n7603), .ZN(n8939) );
  NAND2_X1 U9868 ( .A1(n8267), .A2(n6482), .ZN(n7607) );
  OAI21_X1 U9869 ( .B1(n6481), .B2(n8269), .A(n7607), .ZN(n7615) );
  NAND2_X1 U9870 ( .A1(n7611), .A2(n7610), .ZN(n7612) );
  NAND3_X1 U9871 ( .A1(n7614), .A2(n7613), .A3(n7612), .ZN(n7619) );
  INV_X1 U9872 ( .A(n7615), .ZN(n7617) );
  NAND2_X1 U9873 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  NAND2_X1 U9874 ( .A1(n7619), .A2(n7618), .ZN(n7645) );
  NAND2_X1 U9875 ( .A1(n7620), .A2(SI_2_), .ZN(n7623) );
  INV_X1 U9876 ( .A(n7621), .ZN(n7653) );
  NAND2_X1 U9877 ( .A1(n7653), .A2(n6832), .ZN(n7622) );
  NAND2_X1 U9878 ( .A1(n7623), .A2(n7622), .ZN(n7625) );
  INV_X1 U9879 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8762) );
  XNOR2_X1 U9880 ( .A(n7655), .B(SI_3_), .ZN(n7624) );
  OR2_X1 U9881 ( .A1(n8761), .A2(n8224), .ZN(n7634) );
  NOR2_X1 U9882 ( .A1(n7603), .A2(n7929), .ZN(n7628) );
  MUX2_X1 U9883 ( .A(n7929), .B(n7628), .S(P2_IR_REG_3__SCAN_IN), .Z(n7629) );
  INV_X1 U9884 ( .A(n7629), .ZN(n7631) );
  NAND2_X1 U9885 ( .A1(n7603), .A2(n7630), .ZN(n7673) );
  NAND2_X1 U9886 ( .A1(n7631), .A2(n7673), .ZN(n14545) );
  OAI22_X1 U9887 ( .A1(n7626), .A2(n8733), .B1(n7627), .B2(n14545), .ZN(n7632)
         );
  INV_X1 U9888 ( .A(n7632), .ZN(n7633) );
  NAND2_X1 U9889 ( .A1(n10785), .A2(n7707), .ZN(n7641) );
  INV_X1 U9890 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U9891 ( .A1(n8194), .A2(n10784), .ZN(n7639) );
  NAND2_X1 U9892 ( .A1(n7635), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9893 ( .A1(n7646), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U9894 ( .A1(n7514), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9895 ( .A1(n6486), .A2(n12587), .ZN(n7640) );
  NAND2_X1 U9896 ( .A1(n7641), .A2(n7640), .ZN(n7644) );
  AOI21_X1 U9897 ( .B1(n7645), .B2(n7644), .A(n7642), .ZN(n7643) );
  NAND2_X1 U9898 ( .A1(n7635), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9899 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7683) );
  OAI21_X1 U9900 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7683), .ZN(n7648) );
  INV_X1 U9901 ( .A(n7648), .ZN(n10269) );
  NAND2_X1 U9902 ( .A1(n8194), .A2(n10269), .ZN(n7650) );
  NAND2_X1 U9903 ( .A1(n7514), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7649) );
  INV_X1 U9904 ( .A(SI_2_), .ZN(n8783) );
  INV_X1 U9905 ( .A(SI_3_), .ZN(n8788) );
  AOI22_X1 U9906 ( .A1(n8783), .A2(n7654), .B1(n7655), .B2(n8788), .ZN(n7652)
         );
  INV_X1 U9907 ( .A(n7655), .ZN(n7658) );
  AND2_X1 U9908 ( .A1(SI_2_), .A2(SI_3_), .ZN(n7656) );
  INV_X1 U9909 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U9910 ( .A1(n7673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7661) );
  XNOR2_X1 U9911 ( .A(n7662), .B(n7661), .ZN(n14556) );
  OAI22_X1 U9912 ( .A1(n7626), .A2(n8736), .B1(n7627), .B2(n14556), .ZN(n7663)
         );
  INV_X1 U9913 ( .A(n7663), .ZN(n7664) );
  NAND2_X1 U9914 ( .A1(n7665), .A2(n7664), .ZN(n14717) );
  NAND2_X1 U9915 ( .A1(n14717), .A2(n6481), .ZN(n7666) );
  OAI21_X1 U9916 ( .B1(n6486), .B2(n10779), .A(n7666), .ZN(n7667) );
  OAI22_X1 U9917 ( .A1(n6486), .A2(n6738), .B1(n7707), .B2(n10779), .ZN(n7668)
         );
  INV_X1 U9918 ( .A(n7670), .ZN(n7671) );
  INV_X1 U9919 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9785) );
  XNOR2_X1 U9920 ( .A(n7698), .B(SI_5_), .ZN(n7696) );
  XNOR2_X1 U9921 ( .A(n7697), .B(n7696), .ZN(n9784) );
  OR2_X1 U9922 ( .A1(n9784), .A2(n8224), .ZN(n7681) );
  NAND2_X1 U9923 ( .A1(n7675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7674) );
  MUX2_X1 U9924 ( .A(n7674), .B(P2_IR_REG_31__SCAN_IN), .S(n7676), .Z(n7678)
         );
  INV_X1 U9925 ( .A(n7675), .ZN(n7677) );
  NAND2_X1 U9926 ( .A1(n7677), .A2(n7676), .ZN(n7729) );
  NAND2_X1 U9927 ( .A1(n7678), .A2(n7729), .ZN(n14570) );
  OAI22_X1 U9928 ( .A1(n7626), .A2(n8759), .B1(n7627), .B2(n14570), .ZN(n7679)
         );
  INV_X1 U9929 ( .A(n7679), .ZN(n7680) );
  NAND2_X1 U9930 ( .A1(n7681), .A2(n7680), .ZN(n14727) );
  NAND2_X1 U9931 ( .A1(n14727), .A2(n8235), .ZN(n7690) );
  INV_X2 U9932 ( .A(n7708), .ZN(n8226) );
  NAND2_X1 U9933 ( .A1(n8226), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9934 ( .A1(n8190), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7687) );
  INV_X1 U9935 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7682) );
  NOR2_X1 U9936 ( .A1(n7683), .A2(n7682), .ZN(n7709) );
  AND2_X1 U9937 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NOR2_X1 U9938 ( .A1(n7709), .A2(n7684), .ZN(n10338) );
  NAND2_X1 U9939 ( .A1(n8194), .A2(n10338), .ZN(n7686) );
  NAND2_X1 U9940 ( .A1(n8225), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7685) );
  NAND4_X1 U9941 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n12585)
         );
  NAND2_X1 U9942 ( .A1(n6486), .A2(n12585), .ZN(n7689) );
  NAND2_X1 U9943 ( .A1(n7690), .A2(n7689), .ZN(n7693) );
  AOI22_X1 U9944 ( .A1(n6486), .A2(n14727), .B1(n8235), .B2(n12585), .ZN(n7691) );
  INV_X1 U9945 ( .A(n7692), .ZN(n7695) );
  NAND2_X1 U9946 ( .A1(n7695), .A2(n6549), .ZN(n7720) );
  INV_X1 U9947 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9948 ( .A1(n7699), .A2(SI_5_), .ZN(n7700) );
  MUX2_X1 U9949 ( .A(n9919), .B(n8771), .S(n6484), .Z(n7726) );
  XNOR2_X1 U9950 ( .A(n7726), .B(SI_6_), .ZN(n7724) );
  XNOR2_X1 U9951 ( .A(n7725), .B(n7724), .ZN(n9915) );
  OR2_X1 U9952 ( .A1(n9915), .A2(n8224), .ZN(n7706) );
  NAND2_X1 U9953 ( .A1(n7729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7703) );
  INV_X1 U9954 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U9955 ( .A(n7703), .B(n7702), .ZN(n12614) );
  OAI22_X1 U9956 ( .A1(n7626), .A2(n8771), .B1(n7627), .B2(n12614), .ZN(n7704)
         );
  INV_X1 U9957 ( .A(n7704), .ZN(n7705) );
  NAND2_X1 U9958 ( .A1(n7706), .A2(n7705), .ZN(n14737) );
  NAND2_X1 U9959 ( .A1(n14737), .A2(n6486), .ZN(n7716) );
  NAND2_X1 U9960 ( .A1(n8190), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U9961 ( .A1(n8226), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9962 ( .A1(n7709), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7735) );
  OR2_X1 U9963 ( .A1(n7709), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7710) );
  AND2_X1 U9964 ( .A1(n7735), .A2(n7710), .ZN(n9324) );
  NAND2_X1 U9965 ( .A1(n8194), .A2(n9324), .ZN(n7712) );
  NAND2_X1 U9966 ( .A1(n8225), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7711) );
  NAND4_X1 U9967 ( .A1(n7714), .A2(n7713), .A3(n7712), .A4(n7711), .ZN(n12584)
         );
  NAND2_X1 U9968 ( .A1(n8237), .A2(n12584), .ZN(n7715) );
  NAND2_X1 U9969 ( .A1(n7716), .A2(n7715), .ZN(n7721) );
  NAND2_X1 U9970 ( .A1(n7720), .A2(n7721), .ZN(n7719) );
  INV_X1 U9971 ( .A(n12584), .ZN(n9332) );
  NAND2_X1 U9972 ( .A1(n14737), .A2(n8235), .ZN(n7717) );
  OAI21_X1 U9973 ( .B1(n8235), .B2(n9332), .A(n7717), .ZN(n7718) );
  INV_X1 U9974 ( .A(n7720), .ZN(n7723) );
  INV_X1 U9975 ( .A(n7721), .ZN(n7722) );
  INV_X1 U9976 ( .A(n7726), .ZN(n7727) );
  NAND2_X1 U9977 ( .A1(n7727), .A2(SI_6_), .ZN(n7728) );
  MUX2_X1 U9978 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6484), .Z(n7750) );
  XNOR2_X1 U9979 ( .A(n7750), .B(SI_7_), .ZN(n7747) );
  XNOR2_X1 U9980 ( .A(n7749), .B(n7747), .ZN(n9978) );
  NAND2_X1 U9981 ( .A1(n9978), .A2(n8186), .ZN(n7734) );
  INV_X1 U9982 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U9983 ( .A1(n7753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7731) );
  INV_X1 U9984 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7730) );
  XNOR2_X1 U9985 ( .A(n7731), .B(n7730), .ZN(n12631) );
  OAI22_X1 U9986 ( .A1(n7626), .A2(n8805), .B1(n7627), .B2(n12631), .ZN(n7732)
         );
  INV_X1 U9987 ( .A(n7732), .ZN(n7733) );
  NAND2_X1 U9988 ( .A1(n7734), .A2(n7733), .ZN(n9501) );
  NAND2_X1 U9989 ( .A1(n9501), .A2(n8235), .ZN(n7742) );
  NAND2_X1 U9990 ( .A1(n8190), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U9991 ( .A1(n8226), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U9992 ( .A1(n7735), .A2(n9338), .ZN(n7736) );
  AND2_X1 U9993 ( .A1(n7758), .A2(n7736), .ZN(n14670) );
  NAND2_X1 U9994 ( .A1(n8194), .A2(n14670), .ZN(n7738) );
  NAND2_X1 U9995 ( .A1(n8225), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7737) );
  NAND4_X1 U9996 ( .A1(n7740), .A2(n7739), .A3(n7738), .A4(n7737), .ZN(n12583)
         );
  NAND2_X1 U9997 ( .A1(n6486), .A2(n12583), .ZN(n7741) );
  NAND2_X1 U9998 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  AOI22_X1 U9999 ( .A1(n9501), .A2(n6486), .B1(n8235), .B2(n12583), .ZN(n7743)
         );
  AOI21_X1 U10000 ( .B1(n7745), .B2(n7744), .A(n7743), .ZN(n7746) );
  INV_X1 U10001 ( .A(n7747), .ZN(n7748) );
  NAND2_X1 U10002 ( .A1(n7750), .A2(SI_7_), .ZN(n7751) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6484), .Z(n7773) );
  XNOR2_X1 U10004 ( .A(n7773), .B(SI_8_), .ZN(n7770) );
  NAND2_X1 U10005 ( .A1(n10187), .A2(n8186), .ZN(n7756) );
  NAND2_X1 U10006 ( .A1(n7775), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U10007 ( .A(n7754), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8950) );
  AOI22_X1 U10008 ( .A1(n8187), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8950), .B2(
        n8929), .ZN(n7755) );
  NAND2_X1 U10009 ( .A1(n7756), .A2(n7755), .ZN(n10705) );
  NAND2_X1 U10010 ( .A1(n10705), .A2(n6486), .ZN(n7765) );
  NAND2_X1 U10011 ( .A1(n8190), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U10012 ( .A1(n8226), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7762) );
  INV_X1 U10013 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10014 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U10015 ( .A1(n7785), .A2(n7759), .ZN(n10699) );
  INV_X1 U10016 ( .A(n10699), .ZN(n9586) );
  NAND2_X1 U10017 ( .A1(n8194), .A2(n9586), .ZN(n7761) );
  NAND2_X1 U10018 ( .A1(n8225), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7760) );
  NAND4_X1 U10019 ( .A1(n7763), .A2(n7762), .A3(n7761), .A4(n7760), .ZN(n12582) );
  NAND2_X1 U10020 ( .A1(n8237), .A2(n12582), .ZN(n7764) );
  NAND2_X1 U10021 ( .A1(n7765), .A2(n7764), .ZN(n7768) );
  AOI22_X1 U10022 ( .A1(n10705), .A2(n8235), .B1(n6482), .B2(n12582), .ZN(
        n7766) );
  INV_X1 U10023 ( .A(n7766), .ZN(n7767) );
  INV_X1 U10024 ( .A(n7768), .ZN(n7769) );
  INV_X1 U10025 ( .A(n7791), .ZN(n7796) );
  INV_X1 U10026 ( .A(n7770), .ZN(n7771) );
  NAND2_X1 U10027 ( .A1(n7773), .A2(SI_8_), .ZN(n7774) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6483), .Z(n7800) );
  XNOR2_X1 U10029 ( .A(n7800), .B(SI_9_), .ZN(n7797) );
  XNOR2_X1 U10030 ( .A(n7799), .B(n7797), .ZN(n10389) );
  NAND2_X1 U10031 ( .A1(n10389), .A2(n8186), .ZN(n7783) );
  NAND2_X1 U10032 ( .A1(n7777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U10033 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7776), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7780) );
  INV_X1 U10034 ( .A(n7777), .ZN(n7779) );
  INV_X1 U10035 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U10036 ( .A1(n7779), .A2(n7778), .ZN(n7821) );
  NAND2_X1 U10037 ( .A1(n7780), .A2(n7821), .ZN(n8989) );
  INV_X1 U10038 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8828) );
  OAI22_X1 U10039 ( .A1(n8989), .A2(n7627), .B1(n7626), .B2(n8828), .ZN(n7781)
         );
  INV_X1 U10040 ( .A(n7781), .ZN(n7782) );
  NAND2_X1 U10041 ( .A1(n8226), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10042 ( .A1(n8190), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7788) );
  NOR2_X1 U10043 ( .A1(n7804), .A2(n7521), .ZN(n10322) );
  NAND2_X1 U10044 ( .A1(n8194), .A2(n10322), .ZN(n7787) );
  NAND2_X1 U10045 ( .A1(n8225), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7786) );
  OAI22_X1 U10046 ( .A1(n10324), .A2(n6486), .B1(n8235), .B2(n10738), .ZN(
        n7790) );
  INV_X1 U10047 ( .A(n7790), .ZN(n7795) );
  NAND2_X1 U10048 ( .A1(n7791), .A2(n7790), .ZN(n7794) );
  INV_X1 U10049 ( .A(n10738), .ZN(n12581) );
  AOI22_X1 U10050 ( .A1(n9655), .A2(n6486), .B1(n8237), .B2(n12581), .ZN(n7792) );
  INV_X1 U10051 ( .A(n7797), .ZN(n7798) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6802), .Z(n7815) );
  XNOR2_X1 U10053 ( .A(n7815), .B(SI_10_), .ZN(n7812) );
  XNOR2_X1 U10054 ( .A(n7814), .B(n7812), .ZN(n10509) );
  NAND2_X1 U10055 ( .A1(n10509), .A2(n8186), .ZN(n7803) );
  NAND2_X1 U10056 ( .A1(n7821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7801) );
  XNOR2_X1 U10057 ( .A(n7801), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U10058 ( .A1(n10432), .A2(n8929), .B1(n8187), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10059 ( .A1(n8190), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10060 ( .A1(n8226), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7808) );
  OR2_X1 U10061 ( .A1(n7804), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10062 ( .A1(n7804), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7825) );
  AND2_X1 U10063 ( .A1(n7805), .A2(n7825), .ZN(n10742) );
  NAND2_X1 U10064 ( .A1(n8194), .A2(n10742), .ZN(n7807) );
  NAND2_X1 U10065 ( .A1(n8225), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7806) );
  NAND4_X1 U10066 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n12580) );
  AOI22_X1 U10067 ( .A1(n10750), .A2(n6486), .B1(n8237), .B2(n12580), .ZN(
        n7810) );
  AOI22_X1 U10068 ( .A1(n10750), .A2(n8237), .B1(n6482), .B2(n12580), .ZN(
        n7811) );
  INV_X1 U10069 ( .A(n7833), .ZN(n7835) );
  INV_X1 U10070 ( .A(n7812), .ZN(n7813) );
  NAND2_X1 U10071 ( .A1(n7815), .A2(SI_10_), .ZN(n7816) );
  MUX2_X1 U10072 ( .A(n8842), .B(n8844), .S(n6484), .Z(n7818) );
  INV_X1 U10073 ( .A(n7818), .ZN(n7819) );
  NAND2_X1 U10074 ( .A1(n7819), .A2(SI_11_), .ZN(n7820) );
  NAND2_X1 U10075 ( .A1(n7838), .A2(n7820), .ZN(n7836) );
  OAI21_X1 U10076 ( .B1(n7821), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7822) );
  XNOR2_X1 U10077 ( .A(n7822), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U10078 ( .A1(n10435), .A2(n8929), .B1(n8187), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10079 ( .A1(n8190), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10080 ( .A1(n8226), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7829) );
  INV_X1 U10081 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10082 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  AND2_X1 U10083 ( .A1(n7849), .A2(n7826), .ZN(n10313) );
  NAND2_X1 U10084 ( .A1(n8194), .A2(n10313), .ZN(n7828) );
  NAND2_X1 U10085 ( .A1(n8225), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7827) );
  OAI22_X1 U10086 ( .A1(n10315), .A2(n6486), .B1(n8235), .B2(n10758), .ZN(
        n7832) );
  INV_X1 U10087 ( .A(n7832), .ZN(n7834) );
  AOI22_X1 U10088 ( .A1(n9894), .A2(n6486), .B1(n8235), .B2(n12579), .ZN(n7831) );
  INV_X1 U10089 ( .A(n7857), .ZN(n7860) );
  MUX2_X1 U10090 ( .A(n9001), .B(n9107), .S(n6484), .Z(n7839) );
  NAND2_X1 U10091 ( .A1(n7839), .A2(n10935), .ZN(n7862) );
  INV_X1 U10092 ( .A(n7839), .ZN(n7840) );
  NAND2_X1 U10093 ( .A1(n7840), .A2(SI_12_), .ZN(n7841) );
  XNOR2_X1 U10094 ( .A(n7861), .B(n7520), .ZN(n10790) );
  NAND2_X1 U10095 ( .A1(n10790), .A2(n8186), .ZN(n7847) );
  NAND2_X1 U10096 ( .A1(n7842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7844) );
  XNOR2_X1 U10097 ( .A(n7844), .B(n7843), .ZN(n14586) );
  OAI22_X1 U10098 ( .A1(n7626), .A2(n9107), .B1(n7627), .B2(n14586), .ZN(n7845) );
  INV_X1 U10099 ( .A(n7845), .ZN(n7846) );
  AND2_X1 U10100 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  NOR2_X1 U10101 ( .A1(n7869), .A2(n7850), .ZN(n10767) );
  NAND2_X1 U10102 ( .A1(n10767), .A2(n8194), .ZN(n7854) );
  NAND2_X1 U10103 ( .A1(n8190), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10104 ( .A1(n8226), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10105 ( .A1(n8225), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7851) );
  NAND4_X1 U10106 ( .A1(n7854), .A2(n7853), .A3(n7852), .A4(n7851), .ZN(n12578) );
  AOI22_X1 U10107 ( .A1(n10768), .A2(n6486), .B1(n8235), .B2(n12578), .ZN(
        n7856) );
  INV_X1 U10108 ( .A(n7856), .ZN(n7859) );
  INV_X1 U10109 ( .A(n10768), .ZN(n14276) );
  INV_X1 U10110 ( .A(n12578), .ZN(n10482) );
  OAI22_X1 U10111 ( .A1(n14276), .A2(n6486), .B1(n8235), .B2(n10482), .ZN(
        n7855) );
  OAI21_X1 U10112 ( .B1(n7860), .B2(n7859), .A(n7858), .ZN(n7876) );
  MUX2_X1 U10113 ( .A(n9110), .B(n6767), .S(n6484), .Z(n7880) );
  XNOR2_X1 U10114 ( .A(n7880), .B(SI_13_), .ZN(n7879) );
  XNOR2_X1 U10115 ( .A(n7882), .B(n7879), .ZN(n10854) );
  NAND2_X1 U10116 ( .A1(n10854), .A2(n8186), .ZN(n7868) );
  NAND2_X1 U10117 ( .A1(n7863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7865) );
  XNOR2_X1 U10118 ( .A(n7865), .B(n7864), .ZN(n14601) );
  OAI22_X1 U10119 ( .A1(n7626), .A2(n6767), .B1(n7627), .B2(n14601), .ZN(n7866) );
  INV_X1 U10120 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U10121 ( .A1(n7869), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7891) );
  OR2_X1 U10122 ( .A1(n7869), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10123 ( .A1(n7891), .A2(n7870), .ZN(n10669) );
  NAND2_X1 U10124 ( .A1(n8226), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7871) );
  OAI21_X1 U10125 ( .B1(n10669), .B2(n8023), .A(n7871), .ZN(n7875) );
  NAND2_X1 U10126 ( .A1(n8225), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U10127 ( .A1(n8190), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10128 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  OAI22_X1 U10129 ( .A1(n14270), .A2(n6486), .B1(n8235), .B2(n10759), .ZN(
        n7877) );
  OAI22_X1 U10130 ( .A1(n14270), .A2(n8237), .B1(n10759), .B2(n6486), .ZN(
        n7878) );
  INV_X1 U10131 ( .A(n7880), .ZN(n7881) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6802), .Z(n7897) );
  XNOR2_X1 U10133 ( .A(n7898), .B(n7897), .ZN(n10969) );
  NAND2_X1 U10134 ( .A1(n10969), .A2(n8186), .ZN(n7889) );
  INV_X1 U10135 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9343) );
  OR2_X1 U10136 ( .A1(n7884), .A2(n7929), .ZN(n7886) );
  XNOR2_X1 U10137 ( .A(n7886), .B(n7885), .ZN(n14611) );
  OAI22_X1 U10138 ( .A1(n7626), .A2(n9343), .B1(n7627), .B2(n14611), .ZN(n7887) );
  INV_X1 U10139 ( .A(n7887), .ZN(n7888) );
  NAND2_X2 U10140 ( .A1(n7889), .A2(n7888), .ZN(n10687) );
  INV_X1 U10141 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10142 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NAND2_X1 U10143 ( .A1(n7913), .A2(n7892), .ZN(n10685) );
  AOI22_X1 U10144 ( .A1(n8190), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n8226), .B2(
        P2_REG0_REG_14__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10145 ( .A1(n8225), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7893) );
  OAI211_X1 U10146 ( .C1(n10685), .C2(n8023), .A(n7894), .B(n7893), .ZN(n12577) );
  AOI22_X1 U10147 ( .A1(n10687), .A2(n6486), .B1(n8235), .B2(n12577), .ZN(
        n7896) );
  INV_X1 U10148 ( .A(n10687), .ZN(n14264) );
  INV_X1 U10149 ( .A(n12577), .ZN(n10483) );
  OAI22_X1 U10150 ( .A1(n14264), .A2(n6486), .B1(n8235), .B2(n10483), .ZN(
        n7895) );
  INV_X1 U10151 ( .A(n7905), .ZN(n7902) );
  MUX2_X1 U10152 ( .A(n9571), .B(n9562), .S(n6802), .Z(n7899) );
  NAND2_X1 U10153 ( .A1(n7899), .A2(n11287), .ZN(n7923) );
  INV_X1 U10154 ( .A(n7899), .ZN(n7900) );
  NAND2_X1 U10155 ( .A1(n7900), .A2(SI_15_), .ZN(n7901) );
  NAND2_X1 U10156 ( .A1(n7923), .A2(n7901), .ZN(n7903) );
  NAND2_X1 U10157 ( .A1(n7902), .A2(n7903), .ZN(n7906) );
  INV_X1 U10158 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U10159 ( .A1(n7906), .A2(n7924), .ZN(n11066) );
  NAND2_X1 U10160 ( .A1(n11066), .A2(n8186), .ZN(n7912) );
  OR2_X1 U10161 ( .A1(n7907), .A2(n7929), .ZN(n7909) );
  XNOR2_X1 U10162 ( .A(n7909), .B(n7908), .ZN(n10445) );
  OAI22_X1 U10163 ( .A1(n7627), .A2(n10445), .B1(n7626), .B2(n9562), .ZN(n7910) );
  INV_X1 U10164 ( .A(n7910), .ZN(n7911) );
  AND2_X1 U10165 ( .A1(n7913), .A2(n11775), .ZN(n7914) );
  OR2_X1 U10166 ( .A1(n7914), .A2(n7933), .ZN(n11774) );
  AOI22_X1 U10167 ( .A1(n8225), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8226), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10168 ( .A1(n8190), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7915) );
  OAI211_X1 U10169 ( .C1(n11774), .C2(n8023), .A(n7916), .B(n7915), .ZN(n12883) );
  OAI22_X1 U10170 ( .A1(n11718), .A2(n6486), .B1(n8237), .B2(n11719), .ZN(
        n7918) );
  NAND2_X1 U10171 ( .A1(n7917), .A2(n7918), .ZN(n7922) );
  OAI22_X1 U10172 ( .A1(n11718), .A2(n8237), .B1(n11719), .B2(n6482), .ZN(
        n7921) );
  INV_X1 U10173 ( .A(n7917), .ZN(n7920) );
  INV_X1 U10174 ( .A(n7918), .ZN(n7919) );
  AOI22_X1 U10175 ( .A1(n7922), .A2(n7921), .B1(n7920), .B2(n7919), .ZN(n7938)
         );
  MUX2_X1 U10176 ( .A(n6812), .B(n9752), .S(n6802), .Z(n7925) );
  NAND2_X1 U10177 ( .A1(n7925), .A2(n11307), .ZN(n7942) );
  INV_X1 U10178 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U10179 ( .A1(n7926), .A2(SI_16_), .ZN(n7927) );
  XNOR2_X1 U10180 ( .A(n7941), .B(n7940), .ZN(n11070) );
  NAND2_X1 U10181 ( .A1(n11070), .A2(n8186), .ZN(n7932) );
  INV_X1 U10182 ( .A(n7928), .ZN(n7947) );
  OR2_X1 U10183 ( .A1(n7947), .A2(n7929), .ZN(n7930) );
  XNOR2_X1 U10184 ( .A(n7930), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14643) );
  AOI22_X1 U10185 ( .A1(n14643), .A2(n8929), .B1(n8187), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7931) );
  NOR2_X1 U10186 ( .A1(n7933), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7934) );
  OR2_X1 U10187 ( .A1(n7954), .A2(n7934), .ZN(n12887) );
  AOI22_X1 U10188 ( .A1(n8190), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8226), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10189 ( .A1(n8225), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7935) );
  OAI211_X1 U10190 ( .C1(n12887), .C2(n8023), .A(n7936), .B(n7935), .ZN(n12862) );
  INV_X1 U10191 ( .A(n12862), .ZN(n12498) );
  OAI22_X1 U10192 ( .A1(n12495), .A2(n8237), .B1(n12498), .B2(n6486), .ZN(
        n7937) );
  OAI22_X1 U10193 ( .A1(n12495), .A2(n6486), .B1(n8235), .B2(n12498), .ZN(
        n7939) );
  MUX2_X1 U10194 ( .A(n9824), .B(n9835), .S(n6802), .Z(n7943) );
  INV_X1 U10195 ( .A(SI_17_), .ZN(n11318) );
  NAND2_X1 U10196 ( .A1(n7943), .A2(n11318), .ZN(n7967) );
  INV_X1 U10197 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U10198 ( .A1(n7944), .A2(SI_17_), .ZN(n7945) );
  XNOR2_X1 U10199 ( .A(n7966), .B(n7965), .ZN(n11078) );
  NAND2_X1 U10200 ( .A1(n11078), .A2(n8186), .ZN(n7953) );
  NAND2_X1 U10201 ( .A1(n7947), .A2(n7946), .ZN(n7949) );
  NAND2_X1 U10202 ( .A1(n7949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7948) );
  MUX2_X1 U10203 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7948), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7950) );
  AND2_X1 U10204 ( .A1(n7950), .A2(n7968), .ZN(n12670) );
  NOR2_X1 U10205 ( .A1(n7626), .A2(n9835), .ZN(n7951) );
  AOI21_X1 U10206 ( .B1(n12670), .B2(n8929), .A(n7951), .ZN(n7952) );
  OR2_X1 U10207 ( .A1(n7954), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7955) );
  AND2_X1 U10208 ( .A1(n7993), .A2(n7955), .ZN(n12867) );
  NAND2_X1 U10209 ( .A1(n12867), .A2(n8194), .ZN(n7961) );
  INV_X1 U10210 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10211 ( .A1(n8190), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10212 ( .A1(n8226), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7956) );
  OAI211_X1 U10213 ( .C1(n7958), .C2(n8077), .A(n7957), .B(n7956), .ZN(n7959)
         );
  INV_X1 U10214 ( .A(n7959), .ZN(n7960) );
  NAND2_X1 U10215 ( .A1(n7961), .A2(n7960), .ZN(n12881) );
  AOI22_X1 U10216 ( .A1(n12966), .A2(n8235), .B1(n6482), .B2(n12881), .ZN(
        n7963) );
  INV_X1 U10217 ( .A(n12966), .ZN(n12870) );
  INV_X1 U10218 ( .A(n12881), .ZN(n12547) );
  OAI22_X1 U10219 ( .A1(n12870), .A2(n8237), .B1(n12547), .B2(n6486), .ZN(
        n7962) );
  MUX2_X1 U10220 ( .A(n7192), .B(n10126), .S(n6802), .Z(n7981) );
  XNOR2_X1 U10221 ( .A(n7983), .B(n7981), .ZN(n11090) );
  NAND2_X1 U10222 ( .A1(n11090), .A2(n8186), .ZN(n7973) );
  NAND2_X1 U10223 ( .A1(n7968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7970) );
  XNOR2_X1 U10224 ( .A(n7970), .B(n7969), .ZN(n14660) );
  OAI22_X1 U10225 ( .A1(n14660), .A2(n7627), .B1(n7626), .B2(n10126), .ZN(
        n7971) );
  INV_X1 U10226 ( .A(n7971), .ZN(n7972) );
  XNOR2_X1 U10227 ( .A(n7993), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U10228 ( .A1(n12851), .A2(n8194), .ZN(n7978) );
  INV_X1 U10229 ( .A(n8190), .ZN(n8230) );
  INV_X1 U10230 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U10231 ( .A1(n8225), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10232 ( .A1(n8226), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7974) );
  OAI211_X1 U10233 ( .C1(n8230), .C2(n14649), .A(n7975), .B(n7974), .ZN(n7976)
         );
  INV_X1 U10234 ( .A(n7976), .ZN(n7977) );
  OAI22_X1 U10235 ( .A1(n12853), .A2(n8237), .B1(n12443), .B2(n6486), .ZN(
        n7979) );
  OAI22_X1 U10236 ( .A1(n12853), .A2(n6481), .B1(n8237), .B2(n12443), .ZN(
        n7980) );
  INV_X1 U10237 ( .A(n7981), .ZN(n7982) );
  INV_X1 U10238 ( .A(n7984), .ZN(n7985) );
  NAND2_X1 U10239 ( .A1(n7985), .A2(SI_18_), .ZN(n7986) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6802), .Z(n8009) );
  XNOR2_X1 U10241 ( .A(n8009), .B(SI_19_), .ZN(n8007) );
  XNOR2_X1 U10242 ( .A(n8008), .B(n8007), .ZN(n11101) );
  NAND2_X1 U10243 ( .A1(n11101), .A2(n8186), .ZN(n7989) );
  AOI22_X1 U10244 ( .A1(n7987), .A2(n8929), .B1(n8187), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n7988) );
  INV_X1 U10245 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7991) );
  INV_X1 U10246 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7990) );
  OAI21_X1 U10247 ( .B1(n7993), .B2(n7991), .A(n7990), .ZN(n7994) );
  NAND2_X1 U10248 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n7992) );
  NAND2_X1 U10249 ( .A1(n7994), .A2(n8016), .ZN(n12834) );
  OR2_X1 U10250 ( .A1(n12834), .A2(n8023), .ZN(n7999) );
  INV_X1 U10251 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U10252 ( .A1(n8226), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10253 ( .A1(n8225), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7995) );
  OAI211_X1 U10254 ( .C1(n8230), .C2(n12673), .A(n7996), .B(n7995), .ZN(n7997)
         );
  INV_X1 U10255 ( .A(n7997), .ZN(n7998) );
  OAI22_X1 U10256 ( .A1(n12837), .A2(n6486), .B1(n8237), .B2(n12525), .ZN(
        n8003) );
  INV_X1 U10257 ( .A(n8003), .ZN(n8000) );
  OAI22_X1 U10258 ( .A1(n12837), .A2(n8237), .B1(n12525), .B2(n6486), .ZN(
        n8001) );
  INV_X1 U10259 ( .A(n8001), .ZN(n8005) );
  INV_X1 U10260 ( .A(n8002), .ZN(n8004) );
  OAI22_X1 U10261 ( .A1(n8006), .A2(n8005), .B1(n8004), .B2(n8003), .ZN(n8026)
         );
  INV_X1 U10262 ( .A(n8009), .ZN(n8010) );
  INV_X1 U10263 ( .A(SI_19_), .ZN(n9220) );
  NAND2_X1 U10264 ( .A1(n8010), .A2(n9220), .ZN(n8011) );
  AND2_X1 U10265 ( .A1(n8011), .A2(SI_20_), .ZN(n8012) );
  NAND2_X1 U10266 ( .A1(n8031), .A2(n8030), .ZN(n8013) );
  MUX2_X1 U10267 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6802), .Z(n8028) );
  XNOR2_X1 U10268 ( .A(n8013), .B(n8028), .ZN(n11113) );
  NAND2_X1 U10269 ( .A1(n11113), .A2(n8186), .ZN(n8015) );
  NAND2_X1 U10270 ( .A1(n8187), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10271 ( .A1(n8016), .A2(n12524), .ZN(n8017) );
  NAND2_X1 U10272 ( .A1(n8034), .A2(n8017), .ZN(n12821) );
  INV_X1 U10273 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10274 ( .A1(n8226), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10275 ( .A1(n8190), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8018) );
  OAI211_X1 U10276 ( .C1(n8077), .C2(n8020), .A(n8019), .B(n8018), .ZN(n8021)
         );
  INV_X1 U10277 ( .A(n8021), .ZN(n8022) );
  AOI22_X1 U10278 ( .A1(n12951), .A2(n6481), .B1(n8235), .B2(n12802), .ZN(
        n8025) );
  INV_X1 U10279 ( .A(n8025), .ZN(n8024) );
  INV_X1 U10280 ( .A(n12951), .ZN(n8335) );
  INV_X1 U10281 ( .A(n12802), .ZN(n12465) );
  OAI22_X1 U10282 ( .A1(n8335), .A2(n6486), .B1(n8237), .B2(n12465), .ZN(n8027) );
  INV_X1 U10283 ( .A(n8028), .ZN(n8029) );
  MUX2_X1 U10284 ( .A(n7231), .B(n10646), .S(n6802), .Z(n8046) );
  XNOR2_X1 U10285 ( .A(n8046), .B(SI_21_), .ZN(n8045) );
  XNOR2_X1 U10286 ( .A(n8049), .B(n8045), .ZN(n11121) );
  NAND2_X1 U10287 ( .A1(n11121), .A2(n8186), .ZN(n8033) );
  NAND2_X1 U10288 ( .A1(n8187), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8032) );
  INV_X1 U10289 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12464) );
  AND2_X1 U10290 ( .A1(n8034), .A2(n12464), .ZN(n8035) );
  NOR2_X1 U10291 ( .A1(n8052), .A2(n8035), .ZN(n12808) );
  NAND2_X1 U10292 ( .A1(n12808), .A2(n8194), .ZN(n8041) );
  INV_X1 U10293 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10294 ( .A1(n8225), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10295 ( .A1(n8226), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8036) );
  OAI211_X1 U10296 ( .C1(n8230), .C2(n8038), .A(n8037), .B(n8036), .ZN(n8039)
         );
  INV_X1 U10297 ( .A(n8039), .ZN(n8040) );
  AOI22_X1 U10298 ( .A1(n12946), .A2(n6486), .B1(n8235), .B2(n12817), .ZN(
        n8042) );
  INV_X1 U10299 ( .A(n8042), .ZN(n8043) );
  INV_X1 U10300 ( .A(n8046), .ZN(n8047) );
  NAND2_X1 U10301 ( .A1(n8047), .A2(SI_21_), .ZN(n8048) );
  MUX2_X1 U10302 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6802), .Z(n8084) );
  INV_X1 U10303 ( .A(n8084), .ZN(n8088) );
  XNOR2_X1 U10304 ( .A(n11130), .B(n8088), .ZN(n11783) );
  NAND2_X1 U10305 ( .A1(n11783), .A2(n8186), .ZN(n8051) );
  NAND2_X1 U10306 ( .A1(n8187), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8050) );
  NOR2_X1 U10307 ( .A1(n8052), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8053) );
  OR2_X1 U10308 ( .A1(n8073), .A2(n8053), .ZN(n12537) );
  INV_X1 U10309 ( .A(n12537), .ZN(n12794) );
  NAND2_X1 U10310 ( .A1(n12794), .A2(n8194), .ZN(n8059) );
  INV_X1 U10311 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U10312 ( .A1(n8190), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10313 ( .A1(n8225), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8054) );
  OAI211_X1 U10314 ( .C1(n7708), .C2(n8056), .A(n8055), .B(n8054), .ZN(n8057)
         );
  INV_X1 U10315 ( .A(n8057), .ZN(n8058) );
  OAI22_X1 U10316 ( .A1(n12796), .A2(n8237), .B1(n12772), .B2(n6482), .ZN(
        n8064) );
  OAI22_X1 U10317 ( .A1(n12796), .A2(n6482), .B1(n8237), .B2(n12772), .ZN(
        n8060) );
  AOI21_X1 U10318 ( .B1(n8063), .B2(n8064), .A(n8061), .ZN(n8062) );
  INV_X1 U10319 ( .A(n8064), .ZN(n8065) );
  NAND2_X1 U10320 ( .A1(n11130), .A2(n8084), .ZN(n8068) );
  NAND2_X1 U10321 ( .A1(n8087), .A2(SI_22_), .ZN(n8067) );
  NAND2_X1 U10322 ( .A1(n8068), .A2(n8067), .ZN(n8070) );
  MUX2_X1 U10323 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6802), .Z(n8089) );
  XNOR2_X1 U10324 ( .A(n8089), .B(SI_23_), .ZN(n8069) );
  NAND2_X1 U10325 ( .A1(n11142), .A2(n8186), .ZN(n8072) );
  NAND2_X1 U10326 ( .A1(n8187), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8071) );
  OR2_X1 U10327 ( .A1(n8073), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10328 ( .A1(n8073), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10329 ( .A1(n8074), .A2(n8097), .ZN(n12435) );
  INV_X1 U10330 ( .A(n12435), .ZN(n12778) );
  NAND2_X1 U10331 ( .A1(n12778), .A2(n8194), .ZN(n8080) );
  INV_X1 U10332 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U10333 ( .A1(n8226), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10334 ( .A1(n8190), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8075) );
  OAI211_X1 U10335 ( .C1(n8077), .C2(n12782), .A(n8076), .B(n8075), .ZN(n8078)
         );
  INV_X1 U10336 ( .A(n8078), .ZN(n8079) );
  OAI22_X1 U10337 ( .A1(n12783), .A2(n6486), .B1(n8237), .B2(n12539), .ZN(
        n8082) );
  AOI22_X1 U10338 ( .A1(n7102), .A2(n6486), .B1(n8235), .B2(n12791), .ZN(n8081) );
  INV_X1 U10339 ( .A(n8089), .ZN(n8083) );
  INV_X1 U10340 ( .A(SI_23_), .ZN(n11394) );
  NAND2_X1 U10341 ( .A1(n8083), .A2(n11394), .ZN(n8090) );
  OAI21_X1 U10342 ( .B1(SI_22_), .B2(n8084), .A(n8090), .ZN(n8085) );
  INV_X1 U10343 ( .A(n8085), .ZN(n8086) );
  NAND2_X1 U10344 ( .A1(n8087), .A2(n8086), .ZN(n8093) );
  NOR2_X1 U10345 ( .A1(n8088), .A2(n11383), .ZN(n8091) );
  AOI22_X1 U10346 ( .A1(n8091), .A2(n8090), .B1(n8089), .B2(SI_23_), .ZN(n8092) );
  MUX2_X1 U10347 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6802), .Z(n8106) );
  XNOR2_X1 U10348 ( .A(n8105), .B(n8106), .ZN(n11155) );
  NAND2_X1 U10349 ( .A1(n11155), .A2(n8186), .ZN(n8095) );
  NAND2_X1 U10350 ( .A1(n8187), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10351 ( .A1(n8226), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10352 ( .A1(n8225), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8102) );
  INV_X1 U10353 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10354 ( .A1(n8096), .A2(n8097), .ZN(n8099) );
  INV_X1 U10355 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U10356 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8098), .ZN(n8132) );
  AND2_X1 U10357 ( .A1(n8099), .A2(n8132), .ZN(n12764) );
  NAND2_X1 U10358 ( .A1(n8194), .A2(n12764), .ZN(n8101) );
  NAND2_X1 U10359 ( .A1(n8190), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8100) );
  OAI22_X1 U10360 ( .A1(n12766), .A2(n8237), .B1(n12776), .B2(n6481), .ZN(
        n8139) );
  AOI22_X1 U10361 ( .A1(n12931), .A2(n8235), .B1(n6481), .B2(n12746), .ZN(
        n8104) );
  AOI21_X1 U10362 ( .B1(n8140), .B2(n8139), .A(n8104), .ZN(n8212) );
  INV_X1 U10363 ( .A(n8105), .ZN(n8107) );
  NAND2_X1 U10364 ( .A1(n8107), .A2(n8106), .ZN(n8110) );
  NAND2_X1 U10365 ( .A1(n8108), .A2(SI_24_), .ZN(n8109) );
  INV_X1 U10366 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13011) );
  MUX2_X1 U10367 ( .A(n14172), .B(n13011), .S(n6802), .Z(n8111) );
  INV_X1 U10368 ( .A(SI_25_), .ZN(n11418) );
  NAND2_X1 U10369 ( .A1(n8111), .A2(n11418), .ZN(n8123) );
  INV_X1 U10370 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U10371 ( .A1(n8112), .A2(SI_25_), .ZN(n8113) );
  NAND2_X1 U10372 ( .A1(n8123), .A2(n8113), .ZN(n8124) );
  XNOR2_X1 U10373 ( .A(n8125), .B(n8124), .ZN(n13009) );
  NAND2_X1 U10374 ( .A1(n13009), .A2(n8186), .ZN(n8115) );
  NAND2_X1 U10375 ( .A1(n8187), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10376 ( .A1(n8190), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10377 ( .A1(n8226), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8118) );
  XNOR2_X1 U10378 ( .A(n8132), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U10379 ( .A1(n8194), .A2(n12740), .ZN(n8117) );
  NAND2_X1 U10380 ( .A1(n8225), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8116) );
  NOR2_X1 U10381 ( .A1(n6482), .A2(n12728), .ZN(n8120) );
  AOI21_X1 U10382 ( .B1(n12926), .B2(n6486), .A(n8120), .ZN(n8203) );
  NAND2_X1 U10383 ( .A1(n12926), .A2(n8237), .ZN(n8122) );
  NAND2_X1 U10384 ( .A1(n6481), .A2(n12758), .ZN(n8121) );
  NAND2_X1 U10385 ( .A1(n8122), .A2(n8121), .ZN(n8202) );
  OAI21_X2 U10386 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8142) );
  MUX2_X1 U10387 ( .A(n7241), .B(n13006), .S(n6802), .Z(n8141) );
  XNOR2_X1 U10388 ( .A(n8141), .B(SI_26_), .ZN(n8126) );
  XNOR2_X1 U10389 ( .A(n8142), .B(n8126), .ZN(n13005) );
  NAND2_X1 U10390 ( .A1(n13005), .A2(n8186), .ZN(n8128) );
  NAND2_X1 U10391 ( .A1(n8187), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10392 ( .A1(n8190), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10393 ( .A1(n8226), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8136) );
  INV_X1 U10394 ( .A(n8132), .ZN(n8130) );
  AND2_X1 U10395 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8129) );
  NAND2_X1 U10396 ( .A1(n8130), .A2(n8129), .ZN(n8191) );
  INV_X1 U10397 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12481) );
  INV_X1 U10398 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8131) );
  OAI21_X1 U10399 ( .B1(n8132), .B2(n12481), .A(n8131), .ZN(n8133) );
  AND2_X1 U10400 ( .A1(n8191), .A2(n8133), .ZN(n12732) );
  NAND2_X1 U10401 ( .A1(n8194), .A2(n12732), .ZN(n8135) );
  NAND2_X1 U10402 ( .A1(n8225), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8134) );
  OAI22_X1 U10403 ( .A1(n12734), .A2(n8237), .B1(n12480), .B2(n6481), .ZN(
        n8207) );
  AOI22_X1 U10404 ( .A1(n12922), .A2(n8235), .B1(n6482), .B2(n12747), .ZN(
        n8208) );
  NOR2_X1 U10405 ( .A1(n8207), .A2(n8208), .ZN(n8204) );
  AOI21_X1 U10406 ( .B1(n8203), .B2(n8202), .A(n8204), .ZN(n8138) );
  OAI21_X1 U10407 ( .B1(n8140), .B2(n8139), .A(n8138), .ZN(n8211) );
  OAI21_X1 U10408 ( .B1(n8142), .B2(n11430), .A(n8141), .ZN(n8144) );
  NAND2_X1 U10409 ( .A1(n8142), .A2(n11430), .ZN(n8143) );
  INV_X1 U10410 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13002) );
  MUX2_X1 U10411 ( .A(n14162), .B(n13002), .S(n6802), .Z(n8183) );
  NOR2_X1 U10412 ( .A1(n8145), .A2(SI_27_), .ZN(n8147) );
  NAND2_X1 U10413 ( .A1(n8145), .A2(SI_27_), .ZN(n8146) );
  INV_X1 U10414 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11442) );
  INV_X1 U10415 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11443) );
  MUX2_X1 U10416 ( .A(n11442), .B(n11443), .S(n6802), .Z(n8148) );
  INV_X1 U10417 ( .A(SI_28_), .ZN(n12421) );
  NAND2_X1 U10418 ( .A1(n8148), .A2(n12421), .ZN(n8165) );
  INV_X1 U10419 ( .A(n8148), .ZN(n8149) );
  NAND2_X1 U10420 ( .A1(n8149), .A2(SI_28_), .ZN(n8150) );
  NAND2_X1 U10421 ( .A1(n8165), .A2(n8150), .ZN(n8166) );
  NAND2_X1 U10422 ( .A1(n11246), .A2(n8186), .ZN(n8152) );
  NAND2_X1 U10423 ( .A1(n8187), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8151) );
  NAND2_X2 U10424 ( .A1(n8152), .A2(n8151), .ZN(n12909) );
  NAND2_X1 U10425 ( .A1(n8190), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10426 ( .A1(n8226), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8160) );
  INV_X1 U10427 ( .A(n8191), .ZN(n8153) );
  INV_X1 U10428 ( .A(n8371), .ZN(n8157) );
  INV_X1 U10429 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10430 ( .A1(n8193), .A2(n8155), .ZN(n8156) );
  NAND2_X1 U10431 ( .A1(n8194), .A2(n11766), .ZN(n8159) );
  NAND2_X1 U10432 ( .A1(n8225), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8158) );
  NAND4_X1 U10433 ( .A1(n8161), .A2(n8160), .A3(n8159), .A4(n8158), .ZN(n12575) );
  AND2_X1 U10434 ( .A1(n6482), .A2(n12575), .ZN(n8162) );
  AOI21_X1 U10435 ( .B1(n12909), .B2(n8237), .A(n8162), .ZN(n8248) );
  NAND2_X1 U10436 ( .A1(n12909), .A2(n6486), .ZN(n8164) );
  NAND2_X1 U10437 ( .A1(n8237), .A2(n12575), .ZN(n8163) );
  NAND2_X1 U10438 ( .A1(n8164), .A2(n8163), .ZN(n8246) );
  MUX2_X1 U10439 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6802), .Z(n8176) );
  INV_X1 U10440 ( .A(SI_29_), .ZN(n12417) );
  XNOR2_X1 U10441 ( .A(n8176), .B(n12417), .ZN(n8174) );
  XNOR2_X1 U10442 ( .A(n8175), .B(n8174), .ZN(n13563) );
  NAND2_X1 U10443 ( .A1(n13563), .A2(n8186), .ZN(n8169) );
  NAND2_X1 U10444 ( .A1(n8187), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10445 ( .A1(n8190), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U10446 ( .A1(n8226), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10447 ( .A1(n8194), .A2(n8371), .ZN(n8171) );
  NAND2_X1 U10448 ( .A1(n8225), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8170) );
  AND4_X1 U10449 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n8170), .ZN(n11767)
         );
  OAI22_X1 U10450 ( .A1(n8373), .A2(n6481), .B1(n8237), .B2(n11767), .ZN(n8238) );
  INV_X1 U10451 ( .A(n11767), .ZN(n12574) );
  AOI22_X1 U10452 ( .A1(n12904), .A2(n6486), .B1(n8235), .B2(n12574), .ZN(
        n8239) );
  NOR2_X1 U10453 ( .A1(n8238), .A2(n8239), .ZN(n8247) );
  INV_X1 U10454 ( .A(n8176), .ZN(n8177) );
  MUX2_X1 U10455 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6802), .Z(n8178) );
  NAND2_X1 U10456 ( .A1(n8178), .A2(SI_30_), .ZN(n8179) );
  OAI21_X1 U10457 ( .B1(n8178), .B2(SI_30_), .A(n8179), .ZN(n8220) );
  NAND2_X1 U10458 ( .A1(n8223), .A2(n8179), .ZN(n8182) );
  MUX2_X1 U10459 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6802), .Z(n8180) );
  XNOR2_X1 U10460 ( .A(n8180), .B(SI_31_), .ZN(n8181) );
  AOI22_X1 U10461 ( .A1(n12992), .A2(n8186), .B1(n8187), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8216) );
  XOR2_X1 U10462 ( .A(n12687), .B(n8216), .Z(n8245) );
  XNOR2_X1 U10463 ( .A(n8183), .B(SI_27_), .ZN(n8184) );
  NAND2_X1 U10464 ( .A1(n13001), .A2(n8186), .ZN(n8189) );
  NAND2_X1 U10465 ( .A1(n8187), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10466 ( .A1(n8190), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10467 ( .A1(n8226), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8197) );
  INV_X1 U10468 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U10469 ( .A1(n8191), .A2(n13214), .ZN(n8192) );
  NAND2_X1 U10470 ( .A1(n8194), .A2(n12716), .ZN(n8196) );
  NAND2_X1 U10471 ( .A1(n8225), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8195) );
  NOR2_X1 U10472 ( .A1(n6486), .A2(n12729), .ZN(n8199) );
  AOI21_X1 U10473 ( .B1(n12915), .B2(n6482), .A(n8199), .ZN(n8214) );
  NAND2_X1 U10474 ( .A1(n12915), .A2(n8237), .ZN(n8201) );
  NAND2_X1 U10475 ( .A1(n6481), .A2(n12576), .ZN(n8200) );
  NAND2_X1 U10476 ( .A1(n8201), .A2(n8200), .ZN(n8213) );
  NOR2_X1 U10477 ( .A1(n8214), .A2(n8213), .ZN(n8206) );
  NOR3_X1 U10478 ( .A1(n8204), .A2(n8203), .A3(n8202), .ZN(n8205) );
  AOI211_X1 U10479 ( .C1(n8208), .C2(n8207), .A(n8206), .B(n8205), .ZN(n8209)
         );
  OAI21_X1 U10480 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8256) );
  NOR2_X1 U10481 ( .A1(n12687), .A2(n6482), .ZN(n8243) );
  NAND2_X1 U10482 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  INV_X1 U10483 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11447) );
  OAI22_X1 U10484 ( .A1(n11715), .A2(n8224), .B1(n7626), .B2(n11447), .ZN(
        n8236) );
  INV_X1 U10485 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10486 ( .A1(n8225), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10487 ( .A1(n8226), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8227) );
  OAI211_X1 U10488 ( .C1(n8230), .C2(n8229), .A(n8228), .B(n8227), .ZN(n12573)
         );
  INV_X1 U10489 ( .A(n12687), .ZN(n8834) );
  NAND2_X1 U10490 ( .A1(n8834), .A2(n6486), .ZN(n8259) );
  NAND2_X1 U10491 ( .A1(n12679), .A2(n10555), .ZN(n8359) );
  NAND2_X1 U10492 ( .A1(n8231), .A2(n8413), .ZN(n8233) );
  NAND4_X1 U10493 ( .A1(n8259), .A2(n8368), .A3(n8359), .A4(n8233), .ZN(n8234)
         );
  AOI22_X1 U10494 ( .A1(n8236), .A2(n8235), .B1(n12573), .B2(n8234), .ZN(n8258) );
  INV_X1 U10495 ( .A(n12573), .ZN(n8344) );
  OAI22_X1 U10496 ( .A1(n12902), .A2(n8237), .B1(n8344), .B2(n6486), .ZN(n8257) );
  INV_X1 U10497 ( .A(n8238), .ZN(n8241) );
  INV_X1 U10498 ( .A(n8239), .ZN(n8240) );
  OAI22_X1 U10499 ( .A1(n8258), .A2(n8257), .B1(n8241), .B2(n8240), .ZN(n8242)
         );
  OAI21_X1 U10500 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8253) );
  INV_X1 U10501 ( .A(n8245), .ZN(n8285) );
  INV_X1 U10502 ( .A(n8246), .ZN(n8251) );
  INV_X1 U10503 ( .A(n8247), .ZN(n8250) );
  INV_X1 U10504 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U10505 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  NAND2_X1 U10506 ( .A1(n8256), .A2(n8255), .ZN(n8264) );
  NAND2_X1 U10507 ( .A1(n8258), .A2(n8257), .ZN(n8263) );
  INV_X1 U10508 ( .A(n8259), .ZN(n8261) );
  NOR2_X1 U10509 ( .A1(n8217), .A2(n6486), .ZN(n8260) );
  AOI211_X1 U10510 ( .C1(n12687), .C2(n8217), .A(n8261), .B(n8260), .ZN(n8262)
         );
  NAND2_X1 U10511 ( .A1(n12909), .A2(n12575), .ZN(n8410) );
  OR2_X1 U10512 ( .A1(n12909), .A2(n12575), .ZN(n8265) );
  XNOR2_X1 U10513 ( .A(n12922), .B(n12480), .ZN(n12725) );
  XNOR2_X1 U10514 ( .A(n12926), .B(n12758), .ZN(n12742) );
  INV_X1 U10515 ( .A(n12817), .ZN(n12536) );
  XNOR2_X1 U10516 ( .A(n12946), .B(n12536), .ZN(n12804) );
  XNOR2_X1 U10517 ( .A(n12951), .B(n12802), .ZN(n12818) );
  XNOR2_X1 U10518 ( .A(n12966), .B(n12547), .ZN(n12863) );
  XNOR2_X1 U10519 ( .A(n12970), .B(n12498), .ZN(n12891) );
  XNOR2_X1 U10520 ( .A(n11779), .B(n11719), .ZN(n10651) );
  OR2_X1 U10521 ( .A1(n10687), .A2(n12577), .ZN(n8398) );
  NAND2_X1 U10522 ( .A1(n10687), .A2(n12577), .ZN(n8399) );
  NAND2_X1 U10523 ( .A1(n8398), .A2(n8399), .ZN(n10679) );
  XNOR2_X1 U10524 ( .A(n9894), .B(n10758), .ZN(n8325) );
  XNOR2_X1 U10525 ( .A(n9655), .B(n10738), .ZN(n9648) );
  INV_X1 U10526 ( .A(n12580), .ZN(n10040) );
  OR2_X1 U10527 ( .A1(n10750), .A2(n10040), .ZN(n8322) );
  NAND2_X1 U10528 ( .A1(n10750), .A2(n10040), .ZN(n8323) );
  NAND2_X1 U10529 ( .A1(n8322), .A2(n8323), .ZN(n10736) );
  NAND2_X1 U10530 ( .A1(n14710), .A2(n12587), .ZN(n8266) );
  INV_X1 U10531 ( .A(n12587), .ZN(n10265) );
  NAND2_X1 U10532 ( .A1(n10785), .A2(n10265), .ZN(n10261) );
  NAND2_X1 U10533 ( .A1(n8266), .A2(n10261), .ZN(n8383) );
  INV_X1 U10534 ( .A(n12585), .ZN(n10266) );
  XNOR2_X1 U10535 ( .A(n14727), .B(n10266), .ZN(n10341) );
  NAND2_X1 U10536 ( .A1(n10309), .A2(n8268), .ZN(n8270) );
  NAND2_X1 U10537 ( .A1(n8267), .A2(n8269), .ZN(n8308) );
  NAND2_X1 U10538 ( .A1(n8270), .A2(n8308), .ZN(n8381) );
  INV_X1 U10539 ( .A(n10555), .ZN(n10288) );
  XNOR2_X1 U10540 ( .A(n8273), .B(n10477), .ZN(n14691) );
  NAND4_X1 U10541 ( .A1(n10259), .A2(n10288), .A3(n8380), .A4(n14691), .ZN(
        n8274) );
  NOR4_X1 U10542 ( .A1(n8383), .A2(n10341), .A3(n8381), .A4(n8274), .ZN(n8275)
         );
  XNOR2_X1 U10543 ( .A(n10705), .B(n12582), .ZN(n10694) );
  XNOR2_X1 U10544 ( .A(n14737), .B(n12584), .ZN(n10277) );
  XNOR2_X1 U10545 ( .A(n9501), .B(n12583), .ZN(n9495) );
  NAND4_X1 U10546 ( .A1(n8275), .A2(n10694), .A3(n10277), .A4(n9495), .ZN(
        n8276) );
  NOR4_X1 U10547 ( .A1(n8325), .A2(n9648), .A3(n10736), .A4(n8276), .ZN(n8277)
         );
  XNOR2_X1 U10548 ( .A(n10671), .B(n8326), .ZN(n10666) );
  XNOR2_X1 U10549 ( .A(n10768), .B(n12578), .ZN(n10754) );
  NAND4_X1 U10550 ( .A1(n10679), .A2(n8277), .A3(n10666), .A4(n10754), .ZN(
        n8278) );
  NOR4_X1 U10551 ( .A1(n12863), .A2(n12891), .A3(n10651), .A4(n8278), .ZN(
        n8279) );
  XNOR2_X1 U10552 ( .A(n12956), .B(n12846), .ZN(n12839) );
  INV_X1 U10553 ( .A(n12443), .ZN(n12861) );
  XNOR2_X1 U10554 ( .A(n12961), .B(n12861), .ZN(n12845) );
  NAND4_X1 U10555 ( .A1(n12818), .A2(n8279), .A3(n12839), .A4(n12845), .ZN(
        n8280) );
  NOR3_X1 U10556 ( .A1(n6500), .A2(n12804), .A3(n8280), .ZN(n8281) );
  XNOR2_X1 U10557 ( .A(n12931), .B(n12746), .ZN(n12752) );
  NAND4_X1 U10558 ( .A1(n12742), .A2(n8281), .A3(n12752), .A4(n8337), .ZN(
        n8282) );
  NOR4_X1 U10559 ( .A1(n12720), .A2(n12701), .A3(n12725), .A4(n8282), .ZN(
        n8284) );
  XNOR2_X1 U10560 ( .A(n12904), .B(n12574), .ZN(n8412) );
  XOR2_X1 U10561 ( .A(n12573), .B(n12902), .Z(n8283) );
  OAI21_X1 U10562 ( .B1(n7987), .B2(n10649), .A(n8359), .ZN(n8286) );
  AOI21_X1 U10563 ( .B1(n8415), .B2(n6489), .A(n8286), .ZN(n8287) );
  INV_X1 U10564 ( .A(n8287), .ZN(n8288) );
  MUX2_X1 U10565 ( .A(n8413), .B(n8368), .S(n10288), .Z(n8289) );
  INV_X1 U10566 ( .A(n8295), .ZN(n8291) );
  NAND2_X1 U10567 ( .A1(n8291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8292) );
  OR2_X1 U10568 ( .A1(n8930), .A2(P2_U3088), .ZN(n10902) );
  INV_X1 U10569 ( .A(n10902), .ZN(n8293) );
  NAND2_X1 U10570 ( .A1(n8297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8298) );
  MUX2_X1 U10571 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8298), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8299) );
  NAND2_X1 U10572 ( .A1(n8300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8301) );
  NAND3_X1 U10573 ( .A1(n13004), .A2(n10905), .A3(n8361), .ZN(n8553) );
  INV_X1 U10574 ( .A(n8359), .ZN(n9067) );
  NAND2_X1 U10575 ( .A1(n14685), .A2(n9067), .ZN(n9089) );
  INV_X1 U10576 ( .A(n8933), .ZN(n8302) );
  OAI21_X1 U10577 ( .B1(n10902), .B2(n8413), .A(P2_B_REG_SCAN_IN), .ZN(n8303)
         );
  INV_X1 U10578 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U10579 ( .A1(n7510), .A2(n8304), .ZN(n8305) );
  NAND2_X1 U10580 ( .A1(n8306), .A2(n8305), .ZN(P2_U3328) );
  INV_X1 U10581 ( .A(n12575), .ZN(n8343) );
  NOR2_X1 U10582 ( .A1(n8273), .A2(n8370), .ZN(n10468) );
  INV_X1 U10583 ( .A(n8381), .ZN(n10305) );
  NAND2_X1 U10584 ( .A1(n10304), .A2(n10305), .ZN(n10303) );
  NAND2_X1 U10585 ( .A1(n10303), .A2(n8308), .ZN(n10776) );
  INV_X1 U10586 ( .A(n8383), .ZN(n10775) );
  NAND2_X1 U10587 ( .A1(n10776), .A2(n10775), .ZN(n10778) );
  NAND2_X1 U10588 ( .A1(n10778), .A2(n10261), .ZN(n8309) );
  NAND2_X1 U10589 ( .A1(n10779), .A2(n14717), .ZN(n8310) );
  INV_X1 U10590 ( .A(n14727), .ZN(n10340) );
  NAND2_X1 U10591 ( .A1(n10340), .A2(n12585), .ZN(n8311) );
  NAND2_X1 U10592 ( .A1(n10278), .A2(n10277), .ZN(n8313) );
  NAND2_X1 U10593 ( .A1(n14737), .A2(n9332), .ZN(n8312) );
  NAND2_X1 U10594 ( .A1(n8313), .A2(n8312), .ZN(n9496) );
  INV_X1 U10595 ( .A(n12583), .ZN(n9588) );
  OR2_X1 U10596 ( .A1(n9501), .A2(n9588), .ZN(n8314) );
  NAND2_X1 U10597 ( .A1(n9496), .A2(n8314), .ZN(n8316) );
  NAND2_X1 U10598 ( .A1(n9501), .A2(n9588), .ZN(n8315) );
  NAND2_X1 U10599 ( .A1(n8316), .A2(n8315), .ZN(n10695) );
  INV_X1 U10600 ( .A(n12582), .ZN(n8318) );
  OR2_X1 U10601 ( .A1(n10705), .A2(n8318), .ZN(n8317) );
  NAND2_X1 U10602 ( .A1(n10695), .A2(n8317), .ZN(n8320) );
  NAND2_X1 U10603 ( .A1(n10705), .A2(n8318), .ZN(n8319) );
  NAND2_X1 U10604 ( .A1(n10324), .A2(n12581), .ZN(n8321) );
  INV_X1 U10605 ( .A(n8322), .ZN(n8324) );
  NAND2_X1 U10606 ( .A1(n14270), .A2(n8326), .ZN(n8327) );
  NAND2_X1 U10607 ( .A1(n10662), .A2(n8327), .ZN(n8328) );
  OAI21_X1 U10608 ( .B1(n14270), .B2(n8326), .A(n8328), .ZN(n8329) );
  INV_X1 U10609 ( .A(n12891), .ZN(n8331) );
  INV_X1 U10610 ( .A(n12843), .ZN(n8333) );
  OAI22_X2 U10611 ( .A1(n8333), .A2(n8332), .B1(n12443), .B2(n12961), .ZN(
        n12829) );
  OAI21_X1 U10612 ( .B1(n12837), .B2(n12846), .A(n12829), .ZN(n8334) );
  OAI21_X1 U10613 ( .B1(n12525), .B2(n12956), .A(n8334), .ZN(n12815) );
  INV_X1 U10614 ( .A(n12752), .ZN(n12757) );
  NOR2_X1 U10615 ( .A1(n12766), .A2(n12746), .ZN(n12743) );
  NAND2_X1 U10616 ( .A1(n12734), .A2(n12747), .ZN(n8338) );
  OAI21_X1 U10617 ( .B1(n8343), .B2(n12909), .A(n12697), .ZN(n8340) );
  INV_X1 U10618 ( .A(n8412), .ZN(n8339) );
  OR2_X1 U10619 ( .A1(n6489), .A2(n12679), .ZN(n8342) );
  NAND2_X1 U10620 ( .A1(n8368), .A2(n10288), .ZN(n8341) );
  INV_X1 U10621 ( .A(P2_B_REG_SCAN_IN), .ZN(n8346) );
  OAI21_X1 U10622 ( .B1(n13003), .B2(n8346), .A(n12880), .ZN(n12686) );
  OAI22_X1 U10623 ( .A1(n12686), .A2(n8344), .B1(n8343), .B2(n12773), .ZN(
        n8345) );
  XNOR2_X1 U10624 ( .A(n10905), .B(n8346), .ZN(n8347) );
  INV_X1 U10625 ( .A(n8361), .ZN(n13013) );
  NAND2_X1 U10626 ( .A1(n8347), .A2(n13013), .ZN(n8348) );
  NOR4_X1 U10627 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8357) );
  OR4_X1 U10628 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8354) );
  NOR4_X1 U10629 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8352) );
  NOR4_X1 U10630 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8351) );
  NOR4_X1 U10631 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8350) );
  NOR4_X1 U10632 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8349) );
  NAND4_X1 U10633 ( .A1(n8352), .A2(n8351), .A3(n8350), .A4(n8349), .ZN(n8353)
         );
  NOR4_X1 U10634 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8354), .A4(n8353), .ZN(n8356) );
  NOR4_X1 U10635 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8355) );
  NAND3_X1 U10636 ( .A1(n8357), .A2(n8356), .A3(n8355), .ZN(n8358) );
  AND2_X1 U10637 ( .A1(n14681), .A2(n8358), .ZN(n9064) );
  NAND2_X1 U10638 ( .A1(n9066), .A2(n8359), .ZN(n9082) );
  INV_X1 U10639 ( .A(n9082), .ZN(n8360) );
  OR2_X1 U10640 ( .A1(n9064), .A2(n8360), .ZN(n9488) );
  INV_X1 U10641 ( .A(n9488), .ZN(n8367) );
  INV_X1 U10642 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14688) );
  NAND2_X1 U10643 ( .A1(n14681), .A2(n14688), .ZN(n8363) );
  OR2_X1 U10644 ( .A1(n13004), .A2(n8361), .ZN(n8362) );
  NAND2_X1 U10645 ( .A1(n8363), .A2(n8362), .ZN(n9489) );
  INV_X1 U10646 ( .A(n9489), .ZN(n8366) );
  INV_X1 U10647 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14683) );
  NAND2_X1 U10648 ( .A1(n14681), .A2(n14683), .ZN(n8365) );
  OR2_X1 U10649 ( .A1(n13004), .A2(n10905), .ZN(n8364) );
  NAND4_X1 U10650 ( .A1(n8367), .A2(n14685), .A3(n8366), .A4(n14684), .ZN(
        n8369) );
  OR2_X1 U10651 ( .A1(n14740), .A2(n8368), .ZN(n9080) );
  NAND2_X1 U10652 ( .A1(n14710), .A2(n10783), .ZN(n10782) );
  INV_X1 U10653 ( .A(n14737), .ZN(n10284) );
  INV_X1 U10654 ( .A(n9501), .ZN(n14674) );
  INV_X1 U10655 ( .A(n10705), .ZN(n14749) );
  NAND2_X1 U10656 ( .A1(n10702), .A2(n14749), .ZN(n10701) );
  OR2_X1 U10657 ( .A1(n10701), .A2(n9655), .ZN(n10745) );
  NAND2_X1 U10658 ( .A1(n12495), .A2(n10656), .ZN(n12874) );
  AND2_X2 U10659 ( .A1(n12796), .A2(n12807), .ZN(n12793) );
  AND2_X2 U10660 ( .A1(n6489), .A2(n10649), .ZN(n10289) );
  AND2_X4 U10661 ( .A1(n10289), .A2(n10555), .ZN(n12971) );
  AOI211_X1 U10662 ( .C1(n12904), .C2(n12703), .A(n12865), .B(n12691), .ZN(
        n12903) );
  AND2_X1 U10663 ( .A1(n10289), .A2(n10288), .ZN(n9086) );
  INV_X1 U10664 ( .A(n12886), .ZN(n14669) );
  AOI22_X1 U10665 ( .A1(n14680), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8371), 
        .B2(n14669), .ZN(n8372) );
  OAI21_X1 U10666 ( .B1(n8373), .B2(n14673), .A(n8372), .ZN(n8374) );
  AOI21_X1 U10667 ( .B1(n12903), .B2(n14667), .A(n8374), .ZN(n8375) );
  INV_X1 U10668 ( .A(n8375), .ZN(n8376) );
  NOR2_X1 U10669 ( .A1(n8377), .A2(n8376), .ZN(n8417) );
  NAND2_X1 U10670 ( .A1(n8273), .A2(n10477), .ZN(n9075) );
  NAND2_X1 U10671 ( .A1(n8378), .A2(n9073), .ZN(n8379) );
  NAND2_X1 U10672 ( .A1(n10309), .A2(n8269), .ZN(n8382) );
  NAND2_X1 U10673 ( .A1(n14710), .A2(n10265), .ZN(n8384) );
  NAND2_X1 U10674 ( .A1(n6738), .A2(n10779), .ZN(n8385) );
  INV_X1 U10675 ( .A(n10277), .ZN(n10275) );
  NAND2_X1 U10676 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  OR2_X1 U10677 ( .A1(n14737), .A2(n12584), .ZN(n8386) );
  NAND2_X1 U10678 ( .A1(n10274), .A2(n8386), .ZN(n9494) );
  INV_X1 U10679 ( .A(n9495), .ZN(n9493) );
  OR2_X1 U10680 ( .A1(n9501), .A2(n12583), .ZN(n8387) );
  OR2_X1 U10681 ( .A1(n10324), .A2(n10738), .ZN(n8388) );
  NAND2_X1 U10682 ( .A1(n8389), .A2(n8388), .ZN(n10735) );
  AND2_X1 U10683 ( .A1(n10750), .A2(n12580), .ZN(n8390) );
  AND2_X1 U10684 ( .A1(n10315), .A2(n10758), .ZN(n8391) );
  OR2_X1 U10685 ( .A1(n10315), .A2(n10758), .ZN(n8392) );
  INV_X1 U10686 ( .A(n10754), .ZN(n8393) );
  NAND2_X1 U10687 ( .A1(n10753), .A2(n8393), .ZN(n8395) );
  NAND2_X1 U10688 ( .A1(n10768), .A2(n12578), .ZN(n8394) );
  NAND2_X1 U10689 ( .A1(n8395), .A2(n8394), .ZN(n10667) );
  NAND2_X1 U10690 ( .A1(n14270), .A2(n10759), .ZN(n8396) );
  INV_X1 U10691 ( .A(n8398), .ZN(n8400) );
  NAND2_X1 U10692 ( .A1(n12892), .A2(n12891), .ZN(n12890) );
  OR2_X1 U10693 ( .A1(n12495), .A2(n12498), .ZN(n8401) );
  NAND2_X1 U10694 ( .A1(n12890), .A2(n8401), .ZN(n12864) );
  NAND2_X1 U10695 ( .A1(n12966), .A2(n12881), .ZN(n8402) );
  OR2_X1 U10696 ( .A1(n12837), .A2(n12525), .ZN(n8403) );
  NAND2_X1 U10697 ( .A1(n12837), .A2(n12525), .ZN(n8404) );
  NOR2_X1 U10698 ( .A1(n12951), .A2(n12802), .ZN(n8405) );
  NAND2_X1 U10699 ( .A1(n12951), .A2(n12802), .ZN(n8406) );
  INV_X1 U10700 ( .A(n12804), .ZN(n8407) );
  OR2_X1 U10701 ( .A1(n12796), .A2(n12772), .ZN(n8408) );
  OR2_X1 U10702 ( .A1(n12926), .A2(n12758), .ZN(n8409) );
  XNOR2_X1 U10703 ( .A(n8413), .B(n9071), .ZN(n8414) );
  NAND2_X1 U10704 ( .A1(n8414), .A2(n12679), .ZN(n9072) );
  NAND2_X1 U10705 ( .A1(n8415), .A2(n7987), .ZN(n10294) );
  NAND2_X1 U10706 ( .A1(n6485), .A2(n10294), .ZN(n8416) );
  NAND2_X1 U10707 ( .A1(n8417), .A2(n7516), .ZN(P2_U3236) );
  INV_X1 U10708 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n8520) );
  XOR2_X1 U10709 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n8520), .Z(n8454) );
  INV_X1 U10710 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n8449) );
  XOR2_X1 U10711 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n8458) );
  INV_X1 U10712 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n8447) );
  INV_X1 U10713 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14392) );
  XOR2_X1 U10714 ( .A(n14392), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n8513) );
  INV_X1 U10715 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8445) );
  INV_X1 U10716 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8443) );
  INV_X1 U10717 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n8441) );
  XOR2_X1 U10718 ( .A(n8441), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n8511) );
  INV_X1 U10719 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8439) );
  INV_X1 U10720 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n13212) );
  XOR2_X1 U10721 ( .A(n8435), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n8503) );
  INV_X1 U10722 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n8433) );
  INV_X1 U10723 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8418) );
  INV_X1 U10724 ( .A(n8475), .ZN(n8474) );
  INV_X1 U10725 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n8424) );
  NOR2_X1 U10726 ( .A1(n8425), .A2(n8424), .ZN(n8427) );
  NOR2_X1 U10727 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8486), .ZN(n8426) );
  AND2_X1 U10728 ( .A1(n14805), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8428) );
  NOR2_X1 U10729 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n8429), .ZN(n8431) );
  XNOR2_X1 U10730 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8429), .ZN(n8493) );
  NOR2_X1 U10731 ( .A1(n8493), .A2(n8494), .ZN(n8430) );
  XOR2_X1 U10732 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n8467) );
  NOR2_X1 U10733 ( .A1(n8468), .A2(n8467), .ZN(n8432) );
  NAND2_X1 U10734 ( .A1(n8503), .A2(n8502), .ZN(n8434) );
  NAND2_X1 U10735 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n13212), .ZN(n8436) );
  OAI21_X1 U10736 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n13212), .A(n8436), .ZN(
        n8465) );
  NOR2_X1 U10737 ( .A1(n8466), .A2(n8465), .ZN(n8437) );
  XOR2_X1 U10738 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n8463) );
  NOR2_X1 U10739 ( .A1(n8464), .A2(n8463), .ZN(n8438) );
  NAND2_X1 U10740 ( .A1(n8511), .A2(n8510), .ZN(n8440) );
  XOR2_X1 U10741 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n8462) );
  NOR2_X1 U10742 ( .A1(n8461), .A2(n8462), .ZN(n8442) );
  AOI21_X2 U10743 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n8443), .A(n8442), .ZN(
        n8460) );
  XOR2_X1 U10744 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n8459) );
  NOR2_X1 U10745 ( .A1(n8460), .A2(n8459), .ZN(n8444) );
  NAND2_X1 U10746 ( .A1(n8513), .A2(n8512), .ZN(n8446) );
  OAI21_X2 U10747 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n8447), .A(n8446), .ZN(
        n8457) );
  NOR2_X1 U10748 ( .A1(n8458), .A2(n8457), .ZN(n8448) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8450) );
  NOR2_X1 U10750 ( .A1(n8451), .A2(n8450), .ZN(n8453) );
  XOR2_X1 U10751 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8451), .Z(n8455) );
  NOR2_X1 U10752 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n8455), .ZN(n8452) );
  NOR2_X1 U10753 ( .A1(n8453), .A2(n8452), .ZN(n8522) );
  XNOR2_X1 U10754 ( .A(n8454), .B(n8522), .ZN(n8517) );
  XOR2_X1 U10755 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8455), .Z(n8456) );
  XOR2_X1 U10756 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n8456), .Z(n14223) );
  XOR2_X1 U10757 ( .A(n8458), .B(n8457), .Z(n8516) );
  INV_X1 U10758 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14632) );
  INV_X1 U10759 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14619) );
  XOR2_X1 U10760 ( .A(n8460), .B(n8459), .Z(n14353) );
  INV_X1 U10761 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14605) );
  XOR2_X1 U10762 ( .A(n8462), .B(n8461), .Z(n14350) );
  XOR2_X1 U10763 ( .A(n8464), .B(n8463), .Z(n8509) );
  INV_X1 U10764 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8508) );
  XOR2_X1 U10765 ( .A(n8466), .B(n8465), .Z(n14212) );
  XOR2_X1 U10766 ( .A(n8468), .B(n8467), .Z(n8499) );
  OR2_X1 U10767 ( .A1(n14562), .A2(n8470), .ZN(n8485) );
  INV_X1 U10768 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8481) );
  XNOR2_X1 U10769 ( .A(n8472), .B(n8471), .ZN(n14179) );
  XNOR2_X1 U10770 ( .A(n8473), .B(n8474), .ZN(n8477) );
  NAND2_X1 U10771 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n8477), .ZN(n8479) );
  AOI21_X1 U10772 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n8476), .A(n8475), .ZN(
        n14974) );
  INV_X1 U10773 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n14973) );
  NOR2_X1 U10774 ( .A1(n14974), .A2(n14973), .ZN(n14983) );
  XOR2_X1 U10775 ( .A(n8477), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n14982) );
  NAND2_X1 U10776 ( .A1(n14983), .A2(n14982), .ZN(n8478) );
  NAND2_X1 U10777 ( .A1(n14179), .A2(n14180), .ZN(n8480) );
  NOR2_X1 U10778 ( .A1(n14179), .A2(n14180), .ZN(n14178) );
  XNOR2_X1 U10779 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n8482), .ZN(n14979) );
  NOR2_X1 U10780 ( .A1(n14978), .A2(n14979), .ZN(n8483) );
  INV_X1 U10781 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14980) );
  NAND2_X1 U10782 ( .A1(n14978), .A2(n14979), .ZN(n14977) );
  NAND2_X1 U10783 ( .A1(n14970), .A2(n14969), .ZN(n8484) );
  NAND2_X1 U10784 ( .A1(n8489), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8492) );
  XOR2_X1 U10785 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14805), .Z(n8491) );
  XOR2_X1 U10786 ( .A(n8491), .B(n8490), .Z(n14192) );
  NAND2_X1 U10787 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n8495), .ZN(n8497) );
  XOR2_X1 U10788 ( .A(n8494), .B(n8493), .Z(n14976) );
  INV_X1 U10789 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n12634) );
  NOR2_X1 U10790 ( .A1(n8499), .A2(n8498), .ZN(n8501) );
  NOR2_X1 U10791 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14203), .ZN(n8500) );
  XNOR2_X1 U10792 ( .A(n8503), .B(n8502), .ZN(n8505) );
  NAND2_X1 U10793 ( .A1(n8504), .A2(n8505), .ZN(n8506) );
  NAND2_X1 U10794 ( .A1(n14212), .A2(n14211), .ZN(n8507) );
  XNOR2_X1 U10795 ( .A(n8511), .B(n8510), .ZN(n14347) );
  INV_X1 U10796 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14590) );
  XNOR2_X1 U10797 ( .A(n8513), .B(n8512), .ZN(n14357) );
  NAND2_X1 U10798 ( .A1(n14358), .A2(n14357), .ZN(n8514) );
  NAND2_X1 U10799 ( .A1(n8518), .A2(n8517), .ZN(n8519) );
  AND2_X1 U10800 ( .A1(n8520), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n8521) );
  OAI22_X1 U10801 ( .A1(n8522), .A2(n8521), .B1(P3_ADDR_REG_18__SCAN_IN), .B2(
        n8520), .ZN(n8524) );
  XNOR2_X1 U10802 ( .A(n12684), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8523) );
  NOR2_X1 U10803 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n8532) );
  INV_X2 U10804 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9566) );
  NOR2_X1 U10805 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8543) );
  NOR2_X1 U10806 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8542) );
  NOR2_X1 U10807 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8541) );
  NOR2_X1 U10808 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8540) );
  NAND2_X1 U10809 ( .A1(n8579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8544) );
  MUX2_X1 U10810 ( .A(n8544), .B(P1_IR_REG_31__SCAN_IN), .S(n8573), .Z(n8545)
         );
  NAND2_X1 U10811 ( .A1(n8546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8547) );
  MUX2_X1 U10812 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8547), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8548) );
  INV_X1 U10813 ( .A(n8930), .ZN(n8552) );
  NOR2_X1 U10814 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n8557) );
  NOR2_X1 U10815 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8556) );
  NAND2_X1 U10816 ( .A1(n8559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8560) );
  MUX2_X1 U10817 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8560), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8561) );
  NAND2_X1 U10818 ( .A1(n8604), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8568) );
  NOR2_X2 U10819 ( .A1(n11714), .A2(n8563), .ZN(n8607) );
  NAND2_X1 U10820 ( .A1(n8607), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10821 ( .A1(n9739), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10822 ( .A1(n8606), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8565) );
  INV_X1 U10823 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8572) );
  NAND3_X1 U10824 ( .A1(n8574), .A2(n8573), .A3(n8572), .ZN(n8578) );
  NAND3_X1 U10825 ( .A1(n8574), .A2(n8573), .A3(P1_IR_REG_27__SCAN_IN), .ZN(
        n8576) );
  XNOR2_X1 U10826 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_27__SCAN_IN), .ZN(
        n8575) );
  NAND2_X1 U10827 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8581) );
  INV_X1 U10828 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8580) );
  MUX2_X1 U10829 ( .A(n8581), .B(P1_IR_REG_31__SCAN_IN), .S(n8580), .Z(n8584)
         );
  NAND2_X1 U10830 ( .A1(n8584), .A2(n8583), .ZN(n8855) );
  NAND2_X1 U10831 ( .A1(n8607), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U10832 ( .A1(n8604), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10833 ( .A1(n8606), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10834 ( .A1(n9739), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8587) );
  INV_X1 U10835 ( .A(SI_0_), .ZN(n8591) );
  INV_X1 U10836 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9378) );
  OAI21_X1 U10837 ( .B1(n6484), .B2(n8591), .A(n9378), .ZN(n8592) );
  AND2_X1 U10838 ( .A1(n8593), .A2(n8592), .ZN(n14174) );
  INV_X1 U10839 ( .A(n14032), .ZN(n11038) );
  NAND2_X1 U10840 ( .A1(n9528), .A2(n9533), .ZN(n9532) );
  NAND2_X1 U10841 ( .A1(n13431), .A2(n9158), .ZN(n8594) );
  NAND2_X1 U10842 ( .A1(n9532), .A2(n8594), .ZN(n9472) );
  NAND2_X1 U10843 ( .A1(n8604), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10844 ( .A1(n8606), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10845 ( .A1(n9739), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U10846 ( .A1(n8607), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8595) );
  INV_X1 U10847 ( .A(n9535), .ZN(n13667) );
  XNOR2_X1 U10848 ( .A(n8600), .B(n8599), .ZN(n11059) );
  OR2_X1 U10849 ( .A1(n9977), .A2(n8601), .ZN(n8602) );
  NAND2_X1 U10850 ( .A1(n13667), .A2(n14448), .ZN(n13447) );
  NAND2_X1 U10851 ( .A1(n9535), .A2(n14448), .ZN(n8603) );
  INV_X1 U10852 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10853 ( .A1(n11208), .A2(n8605), .ZN(n8611) );
  NAND2_X1 U10854 ( .A1(n8606), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U10855 ( .A1(n8607), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10856 ( .A1(n8612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8613) );
  XNOR2_X1 U10857 ( .A(n8613), .B(n8527), .ZN(n8873) );
  NOR2_X1 U10858 ( .A1(n8614), .A2(n8628), .ZN(n8615) );
  OR2_X1 U10859 ( .A1(n9804), .A2(n8615), .ZN(n14453) );
  INV_X1 U10861 ( .A(n8617), .ZN(n8618) );
  NAND2_X1 U10862 ( .A1(n8618), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U10863 ( .A1(n8620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10864 ( .A1(n8661), .A2(n13990), .ZN(n13428) );
  OR2_X1 U10865 ( .A1(n9153), .A2(n13428), .ZN(n8626) );
  NAND2_X1 U10866 ( .A1(n9805), .A2(n13990), .ZN(n13824) );
  INV_X1 U10867 ( .A(n13824), .ZN(n14507) );
  NAND2_X1 U10868 ( .A1(n14453), .A2(n14507), .ZN(n8641) );
  NAND2_X1 U10869 ( .A1(n9534), .A2(n14032), .ZN(n13438) );
  NAND2_X1 U10870 ( .A1(n13431), .A2(n13432), .ZN(n13436) );
  NAND2_X1 U10871 ( .A1(n13438), .A2(n13436), .ZN(n8627) );
  INV_X1 U10872 ( .A(n13431), .ZN(n9226) );
  NAND2_X1 U10873 ( .A1(n9226), .A2(n9158), .ZN(n13439) );
  AND2_X1 U10874 ( .A1(n8627), .A2(n13439), .ZN(n9474) );
  OAI21_X1 U10875 ( .B1(n8629), .B2(n13616), .A(n9812), .ZN(n8639) );
  NAND2_X1 U10876 ( .A1(n13928), .A2(n8661), .ZN(n8631) );
  INV_X1 U10877 ( .A(n13587), .ZN(n13604) );
  NAND2_X1 U10878 ( .A1(n10556), .A2(n13604), .ZN(n8630) );
  NAND2_X1 U10879 ( .A1(n8661), .A2(n10556), .ZN(n13597) );
  INV_X1 U10880 ( .A(n13597), .ZN(n8642) );
  INV_X1 U10881 ( .A(n6480), .ZN(n8848) );
  NAND2_X1 U10882 ( .A1(n13579), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U10883 ( .A1(n8606), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10884 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9741) );
  OAI21_X1 U10885 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9741), .ZN(n14420) );
  INV_X1 U10886 ( .A(n14420), .ZN(n8633) );
  NAND2_X1 U10887 ( .A1(n11208), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10888 ( .A1(n9739), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10889 ( .A1(n8642), .A2(n6480), .ZN(n14013) );
  OR2_X1 U10890 ( .A1(n13454), .A2(n14013), .ZN(n8638) );
  OAI21_X1 U10891 ( .B1(n9535), .B2(n14015), .A(n8638), .ZN(n14372) );
  AOI21_X1 U10892 ( .B1(n8639), .B2(n14411), .A(n14372), .ZN(n8640) );
  NAND2_X1 U10893 ( .A1(n8641), .A2(n8640), .ZN(n14458) );
  NAND2_X1 U10894 ( .A1(n13990), .A2(n13587), .ZN(n9164) );
  NAND2_X1 U10895 ( .A1(n8642), .A2(n9164), .ZN(n8645) );
  INV_X1 U10896 ( .A(n8818), .ZN(n8643) );
  NAND2_X1 U10897 ( .A1(n8645), .A2(n8644), .ZN(n9172) );
  NAND3_X1 U10898 ( .A1(n14170), .A2(P1_B_REG_SCAN_IN), .A3(n10994), .ZN(n8646) );
  INV_X1 U10899 ( .A(n8807), .ZN(n11044) );
  INV_X1 U10900 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U10901 ( .A1(n11044), .A2(n8813), .ZN(n8648) );
  INV_X1 U10902 ( .A(n8647), .ZN(n14168) );
  NAND2_X1 U10903 ( .A1(n14168), .A2(n10994), .ZN(n8810) );
  NAND2_X1 U10904 ( .A1(n8648), .A2(n8810), .ZN(n11041) );
  INV_X1 U10905 ( .A(n11041), .ZN(n14135) );
  NOR4_X1 U10906 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8652) );
  NOR4_X1 U10907 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8651) );
  NOR4_X1 U10908 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8650) );
  NOR4_X1 U10909 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8649) );
  AND4_X1 U10910 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n8658)
         );
  NOR2_X1 U10911 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .ZN(
        n8656) );
  NOR4_X1 U10912 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n8655) );
  NOR4_X1 U10913 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n8654) );
  NOR4_X1 U10914 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n8653) );
  AND4_X1 U10915 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), .ZN(n8657)
         );
  NAND2_X1 U10916 ( .A1(n8658), .A2(n8657), .ZN(n11043) );
  NOR2_X1 U10917 ( .A1(n11043), .A2(n11042), .ZN(n8659) );
  NAND2_X1 U10918 ( .A1(n14168), .A2(n14170), .ZN(n11045) );
  OAI21_X1 U10919 ( .B1(n8807), .B2(n8659), .A(n11045), .ZN(n9162) );
  NOR2_X1 U10920 ( .A1(n14135), .A2(n9162), .ZN(n8660) );
  NAND2_X1 U10921 ( .A1(n9170), .A2(n8660), .ZN(n13807) );
  INV_X1 U10922 ( .A(n8661), .ZN(n8662) );
  NAND2_X1 U10923 ( .A1(n8662), .A2(n13587), .ZN(n13596) );
  INV_X1 U10924 ( .A(n11048), .ZN(n8663) );
  OR2_X1 U10925 ( .A1(n8808), .A2(n9156), .ZN(n8817) );
  INV_X1 U10926 ( .A(n8817), .ZN(n9163) );
  MUX2_X1 U10927 ( .A(n14458), .B(P1_REG2_REG_3__SCAN_IN), .S(n6479), .Z(n8669) );
  INV_X1 U10928 ( .A(n14453), .ZN(n8664) );
  NAND2_X1 U10929 ( .A1(n13433), .A2(n13928), .ZN(n13598) );
  OR2_X1 U10930 ( .A1(n6479), .A2(n13598), .ZN(n13886) );
  NOR2_X1 U10931 ( .A1(n8664), .A2(n13886), .ZN(n8668) );
  NOR2_X1 U10932 ( .A1(n13432), .A2(n14032), .ZN(n9530) );
  AND2_X1 U10933 ( .A1(n9530), .A2(n14448), .ZN(n9479) );
  OAI211_X1 U10934 ( .C1(n9479), .C2(n6747), .A(n14429), .B(n14427), .ZN(
        n14455) );
  NOR2_X1 U10935 ( .A1(n14455), .A2(n14022), .ZN(n8667) );
  INV_X1 U10936 ( .A(n9165), .ZN(n11040) );
  NAND2_X1 U10937 ( .A1(n11040), .A2(n13604), .ZN(n8665) );
  OAI22_X1 U10938 ( .A1(n14422), .A2(n6747), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14421), .ZN(n8666) );
  NOR2_X1 U10939 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8672) );
  NOR2_X1 U10940 ( .A1(n8681), .A2(n11301), .ZN(n8679) );
  NOR2_X1 U10941 ( .A1(n8683), .A2(n11301), .ZN(n8684) );
  MUX2_X1 U10942 ( .A(n11301), .B(n8684), .S(P3_IR_REG_25__SCAN_IN), .Z(n8685)
         );
  INV_X1 U10943 ( .A(n8681), .ZN(n8686) );
  NAND2_X1 U10944 ( .A1(n8688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8690) );
  MUX2_X1 U10945 ( .A(n8690), .B(P3_IR_REG_31__SCAN_IN), .S(n8689), .Z(n8692)
         );
  INV_X1 U10946 ( .A(n8683), .ZN(n8691) );
  NAND2_X1 U10947 ( .A1(n6476), .A2(n8693), .ZN(n9368) );
  INV_X1 U10948 ( .A(n8695), .ZN(n8696) );
  AND2_X1 U10949 ( .A1(n7672), .A2(P1_U3086), .ZN(n10899) );
  INV_X2 U10950 ( .A(n10899), .ZN(n14165) );
  NAND2_X1 U10951 ( .A1(n8700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U10952 ( .A(n8701), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9733) );
  INV_X1 U10953 ( .A(n9733), .ZN(n8702) );
  OAI222_X1 U10954 ( .A1(n14166), .A2(n9732), .B1(n14165), .B2(n9731), .C1(
        P1_U3086), .C2(n8702), .ZN(P1_U3351) );
  OAI222_X1 U10955 ( .A1(n14166), .A2(n7600), .B1(n14165), .B2(n8601), .C1(
        P1_U3086), .C2(n11059), .ZN(P1_U3353) );
  NAND2_X1 U10956 ( .A1(n7672), .A2(n6473), .ZN(n12423) );
  NAND2_X1 U10957 ( .A1(n8735), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8703) );
  XNOR2_X1 U10958 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8780) );
  NAND2_X1 U10959 ( .A1(n8782), .A2(n8780), .ZN(n8705) );
  INV_X1 U10960 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10961 ( .A1(n8734), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10962 ( .A1(n8705), .A2(n8704), .ZN(n8787) );
  NAND2_X1 U10963 ( .A1(n8787), .A2(n8785), .ZN(n8707) );
  NAND2_X1 U10964 ( .A1(n8733), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10965 ( .A1(n8707), .A2(n8706), .ZN(n8753) );
  NAND2_X1 U10966 ( .A1(n8736), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U10967 ( .A1(n8759), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8709) );
  XNOR2_X1 U10968 ( .A(n8719), .B(n8718), .ZN(n10154) );
  NAND2_X2 U10969 ( .A1(n6802), .A2(P3_U3151), .ZN(n14186) );
  INV_X1 U10970 ( .A(SI_7_), .ZN(n8714) );
  NAND2_X1 U10971 ( .A1(n8710), .A2(n8711), .ZN(n8715) );
  NAND2_X1 U10972 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  INV_X1 U10973 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8712) );
  XNOR2_X1 U10974 ( .A(n8713), .B(n8712), .ZN(n9704) );
  OAI222_X1 U10975 ( .A1(n12423), .A2(n10154), .B1(n14186), .B2(n8714), .C1(
        n6473), .C2(n9704), .ZN(P3_U3288) );
  NOR2_X1 U10976 ( .A1(n8727), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9838) );
  INV_X1 U10977 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U10978 ( .A1(n9838), .A2(n9839), .ZN(n9841) );
  NAND2_X1 U10979 ( .A1(n9841), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8717) );
  XNOR2_X1 U10980 ( .A(n8717), .B(n8716), .ZN(n10098) );
  INV_X1 U10981 ( .A(SI_10_), .ZN(n8726) );
  INV_X1 U10982 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U10983 ( .A1(n8720), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U10984 ( .A1(n8722), .A2(n8721), .ZN(n8731) );
  INV_X1 U10985 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10986 ( .A1(n8723), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8724) );
  INV_X1 U10987 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U10988 ( .A(n8766), .B(n8765), .ZN(n10816) );
  OAI222_X1 U10989 ( .A1(P3_U3151), .A2(n10098), .B1(n14186), .B2(n8726), .C1(
        n12423), .C2(n10816), .ZN(P3_U3285) );
  NAND2_X1 U10990 ( .A1(n8727), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8728) );
  XNOR2_X1 U10991 ( .A(n8728), .B(P3_IR_REG_8__SCAN_IN), .ZN(n9849) );
  INV_X1 U10992 ( .A(n9849), .ZN(n10362) );
  INV_X1 U10993 ( .A(SI_8_), .ZN(n10365) );
  INV_X1 U10994 ( .A(n8729), .ZN(n8730) );
  XNOR2_X1 U10995 ( .A(n8731), .B(n8730), .ZN(n10361) );
  INV_X1 U10996 ( .A(n10361), .ZN(n8732) );
  OAI222_X1 U10997 ( .A1(n6473), .A2(n10362), .B1(n14186), .B2(n10365), .C1(
        n12423), .C2(n8732), .ZN(P3_U3287) );
  NOR2_X1 U10998 ( .A1(n6483), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12998) );
  INV_X2 U10999 ( .A(n12998), .ZN(n13010) );
  NAND2_X1 U11000 ( .A1(n6483), .A2(P2_U3088), .ZN(n13012) );
  INV_X1 U11001 ( .A(n13012), .ZN(n10901) );
  INV_X1 U11002 ( .A(n10901), .ZN(n10648) );
  OAI222_X1 U11003 ( .A1(n13010), .A2(n8733), .B1(n10648), .B2(n8761), .C1(
        n14545), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U11004 ( .A(n8939), .ZN(n12602) );
  OAI222_X1 U11005 ( .A1(n13010), .A2(n8734), .B1(n10648), .B2(n8601), .C1(
        n12602), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U11006 ( .A(n8937), .ZN(n12590) );
  OAI222_X1 U11007 ( .A1(n12590), .A2(P2_U3088), .B1(n10648), .B2(n8760), .C1(
        n8735), .C2(n13010), .ZN(P2_U3326) );
  OAI222_X1 U11008 ( .A1(n13010), .A2(n8736), .B1(n10648), .B2(n9731), .C1(
        n14556), .C2(P2_U3088), .ZN(P2_U3323) );
  NAND2_X1 U11009 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8738) );
  INV_X1 U11010 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U11011 ( .A(n8738), .B(P3_IR_REG_31__SCAN_IN), .S(n8737), .Z(n8741)
         );
  INV_X1 U11012 ( .A(n8739), .ZN(n8740) );
  OAI21_X1 U11013 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n9429) );
  INV_X1 U11014 ( .A(n9429), .ZN(n8745) );
  OAI222_X1 U11015 ( .A1(n9432), .A2(P3_U3151), .B1(n12423), .B2(n8745), .C1(
        n9431), .C2(n14186), .ZN(P3_U3294) );
  OR2_X1 U11016 ( .A1(n8710), .A2(n11301), .ZN(n8746) );
  XNOR2_X1 U11017 ( .A(n8746), .B(P3_IR_REG_6__SCAN_IN), .ZN(n9677) );
  INV_X1 U11018 ( .A(n9677), .ZN(n14796) );
  XNOR2_X1 U11019 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8747) );
  XNOR2_X1 U11020 ( .A(n8748), .B(n8747), .ZN(n10061) );
  INV_X1 U11021 ( .A(n10061), .ZN(n8749) );
  INV_X1 U11022 ( .A(SI_6_), .ZN(n10062) );
  OAI222_X1 U11023 ( .A1(n14796), .A2(n6473), .B1(n12423), .B2(n8749), .C1(
        n10062), .C2(n14186), .ZN(P3_U3289) );
  NAND2_X1 U11024 ( .A1(n8750), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8751) );
  XNOR2_X1 U11025 ( .A(n8751), .B(n8670), .ZN(n9277) );
  XNOR2_X1 U11026 ( .A(n8753), .B(n6774), .ZN(n10003) );
  INV_X1 U11027 ( .A(SI_4_), .ZN(n8754) );
  OAI222_X1 U11028 ( .A1(P3_U3151), .A2(n9277), .B1(n12423), .B2(n10003), .C1(
        n8754), .C2(n14186), .ZN(P3_U3291) );
  NOR2_X1 U11029 ( .A1(n8755), .A2(n14155), .ZN(n8756) );
  MUX2_X1 U11030 ( .A(n14155), .B(n8756), .S(P1_IR_REG_5__SCAN_IN), .Z(n8758)
         );
  OR2_X1 U11031 ( .A1(n8758), .A2(n8757), .ZN(n13691) );
  OAI222_X1 U11032 ( .A1(n14166), .A2(n9785), .B1(n14165), .B2(n9784), .C1(
        P1_U3086), .C2(n13691), .ZN(P1_U3350) );
  OAI222_X1 U11033 ( .A1(n13010), .A2(n8759), .B1(n10648), .B2(n9784), .C1(
        n14570), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U11034 ( .A1(n14166), .A2(n6991), .B1(n14165), .B2(n8760), .C1(
        P1_U3086), .C2(n8855), .ZN(P1_U3354) );
  OAI222_X1 U11035 ( .A1(n14166), .A2(n8762), .B1(n14165), .B2(n8761), .C1(
        P1_U3086), .C2(n8873), .ZN(P1_U3352) );
  OAI21_X1 U11036 ( .B1(n9841), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8764) );
  INV_X1 U11037 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8763) );
  XNOR2_X1 U11038 ( .A(n8764), .B(n8763), .ZN(n10217) );
  INV_X1 U11039 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11040 ( .A1(n8767), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8768) );
  XNOR2_X1 U11041 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8791) );
  XNOR2_X1 U11042 ( .A(n8792), .B(n8791), .ZN(n10921) );
  OAI222_X1 U11043 ( .A1(P3_U3151), .A2(n10217), .B1(n14186), .B2(n8769), .C1(
        n12423), .C2(n10921), .ZN(P3_U3284) );
  OR2_X1 U11044 ( .A1(n8757), .A2(n14155), .ZN(n8770) );
  XNOR2_X1 U11045 ( .A(n8770), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9916) );
  INV_X1 U11046 ( .A(n9916), .ZN(n8891) );
  OAI222_X1 U11047 ( .A1(n14166), .A2(n9919), .B1(n14165), .B2(n9915), .C1(
        P1_U3086), .C2(n8891), .ZN(P1_U3349) );
  OAI222_X1 U11048 ( .A1(n12614), .A2(P2_U3088), .B1(n10648), .B2(n9915), .C1(
        n8771), .C2(n13010), .ZN(P2_U3321) );
  INV_X1 U11049 ( .A(n8710), .ZN(n8775) );
  NAND2_X1 U11050 ( .A1(n8772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8773) );
  MUX2_X1 U11051 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8773), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8774) );
  NAND2_X1 U11052 ( .A1(n8775), .A2(n8774), .ZN(n9668) );
  XNOR2_X1 U11053 ( .A(n8777), .B(n7018), .ZN(n10017) );
  INV_X1 U11054 ( .A(SI_5_), .ZN(n8778) );
  OAI222_X1 U11055 ( .A1(n6473), .A2(n9668), .B1(n12423), .B2(n10017), .C1(
        n8778), .C2(n14186), .ZN(P3_U3290) );
  OR2_X1 U11056 ( .A1(n8739), .A2(n11301), .ZN(n8779) );
  INV_X1 U11057 ( .A(n9513), .ZN(n9141) );
  INV_X1 U11058 ( .A(n8780), .ZN(n8781) );
  XNOR2_X1 U11059 ( .A(n8782), .B(n8781), .ZN(n9512) );
  OAI222_X1 U11060 ( .A1(P3_U3151), .A2(n9141), .B1(n12423), .B2(n9512), .C1(
        n8783), .C2(n14186), .ZN(P3_U3293) );
  NAND2_X1 U11061 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6535), .ZN(n8784) );
  XNOR2_X1 U11062 ( .A(n8784), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9600) );
  INV_X1 U11063 ( .A(n9600), .ZN(n9241) );
  INV_X1 U11064 ( .A(n8785), .ZN(n8786) );
  XNOR2_X1 U11065 ( .A(n8787), .B(n8786), .ZN(n9599) );
  OAI222_X1 U11066 ( .A1(n6473), .A2(n9241), .B1(n12423), .B2(n9599), .C1(
        n8788), .C2(n14186), .ZN(P3_U3292) );
  OR2_X1 U11067 ( .A1(n8789), .A2(n11301), .ZN(n8790) );
  XNOR2_X1 U11068 ( .A(n8790), .B(P3_IR_REG_12__SCAN_IN), .ZN(n10537) );
  INV_X1 U11069 ( .A(n10537), .ZN(n10934) );
  XNOR2_X1 U11070 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9106) );
  INV_X1 U11071 ( .A(n9106), .ZN(n8793) );
  XNOR2_X1 U11072 ( .A(n9105), .B(n8793), .ZN(n10937) );
  INV_X1 U11073 ( .A(n10937), .ZN(n8794) );
  OAI222_X1 U11074 ( .A1(P3_U3151), .A2(n10934), .B1(n14186), .B2(n10935), 
        .C1(n12423), .C2(n8794), .ZN(P3_U3283) );
  INV_X1 U11075 ( .A(n9978), .ZN(n8806) );
  INV_X1 U11076 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11077 ( .A1(n8757), .A2(n8795), .ZN(n8814) );
  NAND2_X1 U11078 ( .A1(n8814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8796) );
  XNOR2_X1 U11079 ( .A(n8796), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9979) );
  INV_X1 U11080 ( .A(n14166), .ZN(n14157) );
  AOI22_X1 U11081 ( .A1(n9979), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14157), .ZN(n8797) );
  OAI21_X1 U11082 ( .B1(n8806), .B2(n14165), .A(n8797), .ZN(P1_U3348) );
  INV_X1 U11083 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8804) );
  XNOR2_X1 U11084 ( .A(n10597), .B(P3_B_REG_SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11085 ( .A1(n10851), .A2(n8798), .ZN(n8799) );
  NAND2_X1 U11086 ( .A1(n11031), .A2(n8804), .ZN(n8802) );
  INV_X1 U11087 ( .A(n6476), .ZN(n10898) );
  NAND2_X1 U11088 ( .A1(n10898), .A2(n10851), .ZN(n8801) );
  AND2_X1 U11089 ( .A1(n8802), .A2(n8801), .ZN(n12306) );
  NAND2_X1 U11090 ( .A1(n12306), .A2(n9015), .ZN(n8803) );
  OAI21_X1 U11091 ( .B1(n8804), .B2(n9015), .A(n8803), .ZN(P3_U3377) );
  OAI222_X1 U11092 ( .A1(n12631), .A2(P2_U3088), .B1(n10648), .B2(n8806), .C1(
        n8805), .C2(n13010), .ZN(P2_U3320) );
  NAND2_X1 U11093 ( .A1(n9163), .A2(n8807), .ZN(n14439) );
  INV_X1 U11094 ( .A(n8808), .ZN(n8812) );
  INV_X1 U11095 ( .A(n11045), .ZN(n8809) );
  AOI22_X1 U11096 ( .A1(n14439), .A2(n11042), .B1(n8812), .B2(n8809), .ZN(
        P1_U3446) );
  INV_X1 U11097 ( .A(n8810), .ZN(n8811) );
  AOI22_X1 U11098 ( .A1(n14439), .A2(n8813), .B1(n8812), .B2(n8811), .ZN(
        P1_U3445) );
  INV_X1 U11099 ( .A(n10187), .ZN(n8820) );
  NAND2_X1 U11100 ( .A1(n8822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U11101 ( .A(n8815), .B(P1_IR_REG_8__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U11102 ( .A1(n13709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n14157), .ZN(n8816) );
  OAI21_X1 U11103 ( .B1(n8820), .B2(n14165), .A(n8816), .ZN(P1_U3347) );
  NAND2_X1 U11104 ( .A1(n8818), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13645) );
  NAND2_X1 U11105 ( .A1(n8817), .A2(n13645), .ZN(n8847) );
  OR2_X1 U11106 ( .A1(n13597), .A2(n8818), .ZN(n8819) );
  NAND2_X1 U11107 ( .A1(n11132), .A2(n8819), .ZN(n8845) );
  INV_X1 U11108 ( .A(n14391), .ZN(n13746) );
  NOR2_X1 U11109 ( .A1(n13746), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11110 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8821) );
  INV_X1 U11111 ( .A(n8950), .ZN(n12640) );
  OAI222_X1 U11112 ( .A1(n13010), .A2(n8821), .B1(n10648), .B2(n8820), .C1(
        n12640), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U11113 ( .A(n10389), .ZN(n8827) );
  NOR2_X1 U11114 ( .A1(n8822), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8840) );
  OR2_X1 U11115 ( .A1(n8840), .A2(n14155), .ZN(n8824) );
  INV_X1 U11116 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8823) );
  OR2_X1 U11117 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  NAND2_X1 U11118 ( .A1(n8824), .A2(n8823), .ZN(n8829) );
  AOI22_X1 U11119 ( .A1(n13725), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14157), .ZN(n8826) );
  OAI21_X1 U11120 ( .B1(n8827), .B2(n14165), .A(n8826), .ZN(P1_U3346) );
  OAI222_X1 U11121 ( .A1(n13010), .A2(n8828), .B1(n10648), .B2(n8827), .C1(
        n8989), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U11122 ( .A(n10509), .ZN(n8837) );
  NAND2_X1 U11123 ( .A1(n8829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U11124 ( .A(n8830), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U11125 ( .A1(n10510), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14157), .ZN(n8831) );
  OAI21_X1 U11126 ( .B1(n8837), .B2(n14165), .A(n8831), .ZN(P1_U3345) );
  INV_X1 U11127 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U11128 ( .A1(n6938), .A2(P1_U4016), .ZN(n8832) );
  OAI21_X1 U11129 ( .B1(P1_U4016), .B2(n8833), .A(n8832), .ZN(P1_U3560) );
  INV_X1 U11130 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U11131 ( .A1(n8834), .A2(P2_U3947), .ZN(n8835) );
  OAI21_X1 U11132 ( .B1(n11450), .B2(P2_U3947), .A(n8835), .ZN(P2_U3562) );
  INV_X1 U11133 ( .A(n10432), .ZN(n8996) );
  INV_X1 U11134 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8836) );
  OAI222_X1 U11135 ( .A1(n8996), .A2(P2_U3088), .B1(n10648), .B2(n8837), .C1(
        n8836), .C2(n13010), .ZN(P2_U3317) );
  NAND2_X1 U11136 ( .A1(n12802), .A2(P2_U3947), .ZN(n8838) );
  OAI21_X1 U11137 ( .B1(n10481), .B2(P2_U3947), .A(n8838), .ZN(P2_U3551) );
  INV_X1 U11138 ( .A(n10573), .ZN(n8843) );
  NOR2_X1 U11139 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8839) );
  NAND2_X1 U11140 ( .A1(n8840), .A2(n8839), .ZN(n9568) );
  NAND2_X1 U11141 ( .A1(n9568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8841) );
  XNOR2_X1 U11142 ( .A(n8841), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10574) );
  INV_X1 U11143 ( .A(n10574), .ZN(n9550) );
  OAI222_X1 U11144 ( .A1(n14166), .A2(n8842), .B1(n14165), .B2(n8843), .C1(
        P1_U3086), .C2(n9550), .ZN(P1_U3344) );
  INV_X1 U11145 ( .A(n10435), .ZN(n12656) );
  OAI222_X1 U11146 ( .A1(n13010), .A2(n8844), .B1(n10648), .B2(n8843), .C1(
        n12656), .C2(P2_U3088), .ZN(P2_U3316) );
  INV_X1 U11147 ( .A(n8845), .ZN(n8846) );
  AND2_X1 U11148 ( .A1(n8847), .A2(n8846), .ZN(n8899) );
  INV_X1 U11149 ( .A(n8899), .ZN(n8849) );
  INV_X1 U11150 ( .A(n8855), .ZN(n13676) );
  XNOR2_X1 U11151 ( .A(n8855), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13669) );
  AND3_X1 U11152 ( .A1(n13669), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n13670) );
  AOI21_X1 U11153 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n13676), .A(n13670), .ZN(
        n11057) );
  INV_X1 U11154 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8850) );
  MUX2_X1 U11155 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8850), .S(n11059), .Z(
        n11056) );
  INV_X1 U11156 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n8851) );
  MUX2_X1 U11157 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n8851), .S(n8873), .Z(n8852)
         );
  AOI211_X1 U11158 ( .C1(n8853), .C2(n8852), .A(n8868), .B(n13737), .ZN(n8864)
         );
  NOR2_X1 U11159 ( .A1(n6480), .A2(n14163), .ZN(n8854) );
  AND2_X1 U11160 ( .A1(n8899), .A2(n8854), .ZN(n14387) );
  XNOR2_X1 U11161 ( .A(n8855), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n13679) );
  AND2_X1 U11162 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13678) );
  NAND2_X1 U11163 ( .A1(n13679), .A2(n13678), .ZN(n13677) );
  NAND2_X1 U11164 ( .A1(n13676), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11165 ( .A1(n13677), .A2(n8856), .ZN(n11051) );
  INV_X1 U11166 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U11167 ( .A(n8857), .B(P1_REG2_REG_2__SCAN_IN), .S(n11059), .Z(n8858) );
  AND2_X1 U11168 ( .A1(n11051), .A2(n8858), .ZN(n11052) );
  NOR2_X1 U11169 ( .A1(n11059), .A2(n8857), .ZN(n8861) );
  INV_X1 U11170 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n8859) );
  MUX2_X1 U11171 ( .A(n8859), .B(P1_REG2_REG_3__SCAN_IN), .S(n8873), .Z(n8860)
         );
  OAI21_X1 U11172 ( .B1(n11052), .B2(n8861), .A(n8860), .ZN(n8874) );
  INV_X1 U11173 ( .A(n8874), .ZN(n9409) );
  NOR3_X1 U11174 ( .A1(n11052), .A2(n8861), .A3(n8860), .ZN(n8862) );
  NOR3_X1 U11175 ( .A1(n13773), .A2(n9409), .A3(n8862), .ZN(n8863) );
  NOR2_X1 U11176 ( .A1(n8864), .A2(n8863), .ZN(n8867) );
  NOR2_X1 U11177 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8605), .ZN(n8865) );
  AOI21_X1 U11178 ( .B1(n13746), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n8865), .ZN(
        n8866) );
  OAI211_X1 U11179 ( .C1(n8873), .C2(n13772), .A(n8867), .B(n8866), .ZN(
        P1_U3246) );
  XNOR2_X1 U11180 ( .A(n9916), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n8872) );
  INV_X1 U11181 ( .A(n13691), .ZN(n13690) );
  INV_X1 U11182 ( .A(n8873), .ZN(n8869) );
  INV_X1 U11183 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8870) );
  MUX2_X1 U11184 ( .A(n8870), .B(P1_REG1_REG_4__SCAN_IN), .S(n9733), .Z(n9412)
         );
  NOR2_X1 U11185 ( .A1(n9413), .A2(n9412), .ZN(n9411) );
  AOI21_X1 U11186 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9733), .A(n9411), .ZN(
        n13684) );
  XNOR2_X1 U11187 ( .A(n13691), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n13685) );
  NAND2_X1 U11188 ( .A1(n13684), .A2(n13685), .ZN(n13683) );
  OAI21_X1 U11189 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13690), .A(n13683), .ZN(
        n8871) );
  NOR2_X1 U11190 ( .A1(n8871), .A2(n8872), .ZN(n8969) );
  AOI211_X1 U11191 ( .C1(n8872), .C2(n8871), .A(n13737), .B(n8969), .ZN(n8887)
         );
  OR2_X1 U11192 ( .A1(n8873), .A2(n8859), .ZN(n9406) );
  NAND2_X1 U11193 ( .A1(n8874), .A2(n9406), .ZN(n8877) );
  INV_X1 U11194 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8875) );
  MUX2_X1 U11195 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n8875), .S(n9733), .Z(n8876)
         );
  NAND2_X1 U11196 ( .A1(n8877), .A2(n8876), .ZN(n13694) );
  NAND2_X1 U11197 ( .A1(n9733), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13693) );
  NAND2_X1 U11198 ( .A1(n13694), .A2(n13693), .ZN(n8879) );
  INV_X1 U11199 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9818) );
  MUX2_X1 U11200 ( .A(n9818), .B(P1_REG2_REG_5__SCAN_IN), .S(n13691), .Z(n8878) );
  NAND2_X1 U11201 ( .A1(n8879), .A2(n8878), .ZN(n13696) );
  NAND2_X1 U11202 ( .A1(n13690), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U11203 ( .A1(n13696), .A2(n8884), .ZN(n8882) );
  INV_X1 U11204 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U11205 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n8880), .S(n9916), .Z(n8881)
         );
  NAND2_X1 U11206 ( .A1(n8882), .A2(n8881), .ZN(n8977) );
  MUX2_X1 U11207 ( .A(n8880), .B(P1_REG2_REG_6__SCAN_IN), .S(n9916), .Z(n8883)
         );
  NAND3_X1 U11208 ( .A1(n13696), .A2(n8884), .A3(n8883), .ZN(n8885) );
  AND3_X1 U11209 ( .A1(n14387), .A2(n8977), .A3(n8885), .ZN(n8886) );
  NOR2_X1 U11210 ( .A1(n8887), .A2(n8886), .ZN(n8890) );
  INV_X1 U11211 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U11212 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9931), .ZN(n8888) );
  AOI21_X1 U11213 ( .B1(n13746), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n8888), .ZN(
        n8889) );
  OAI211_X1 U11214 ( .C1(n8891), .C2(n13772), .A(n8890), .B(n8889), .ZN(
        P1_U3249) );
  INV_X1 U11215 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8893) );
  NOR2_X1 U11216 ( .A1(n14163), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8892) );
  OR2_X1 U11217 ( .A1(n6480), .A2(n8892), .ZN(n9404) );
  AOI21_X1 U11218 ( .B1(n14163), .B2(n8893), .A(n9404), .ZN(n8894) );
  INV_X1 U11219 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9405) );
  MUX2_X1 U11220 ( .A(n8894), .B(n9404), .S(P1_IR_REG_0__SCAN_IN), .Z(n8898)
         );
  INV_X1 U11221 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8895) );
  OAI22_X1 U11222 ( .A1(n14391), .A2(n6793), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8895), .ZN(n8897) );
  NOR3_X1 U11223 ( .A1(n13737), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9405), .ZN(
        n8896) );
  AOI211_X1 U11224 ( .C1(n8899), .C2(n8898), .A(n8897), .B(n8896), .ZN(n8900)
         );
  INV_X1 U11225 ( .A(n8900), .ZN(P1_U3243) );
  INV_X1 U11226 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U11227 ( .A1(n8903), .A2(n8901), .ZN(n12406) );
  NAND2_X4 U11228 ( .A1(n8905), .A2(n12419), .ZN(n11468) );
  INV_X1 U11229 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11230 ( .A1(n11433), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8911) );
  INV_X1 U11231 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9522) );
  OR2_X1 U11232 ( .A1(n9825), .A2(n9522), .ZN(n8910) );
  INV_X1 U11233 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8908) );
  INV_X1 U11234 ( .A(n9769), .ZN(n14892) );
  NAND2_X1 U11235 ( .A1(n14892), .A2(P3_U3897), .ZN(n8913) );
  OAI21_X1 U11236 ( .B1(P3_U3897), .B2(n13164), .A(n8913), .ZN(P3_U3493) );
  INV_X1 U11237 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n13251) );
  MUX2_X1 U11238 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n13251), .S(n8989), .Z(n8928) );
  INV_X1 U11239 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U11240 ( .A(n8939), .B(n8914), .ZN(n12606) );
  INV_X1 U11241 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8915) );
  XNOR2_X1 U11242 ( .A(n8937), .B(n8915), .ZN(n12594) );
  AND2_X1 U11243 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n12593) );
  NAND2_X1 U11244 ( .A1(n12594), .A2(n12593), .ZN(n12592) );
  NAND2_X1 U11245 ( .A1(n8937), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11246 ( .A1(n12592), .A2(n8916), .ZN(n12605) );
  NAND2_X1 U11247 ( .A1(n12606), .A2(n12605), .ZN(n12604) );
  NAND2_X1 U11248 ( .A1(n8939), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11249 ( .A1(n12604), .A2(n8917), .ZN(n14540) );
  XNOR2_X1 U11250 ( .A(n14545), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U11251 ( .A1(n14540), .A2(n14541), .ZN(n14539) );
  INV_X1 U11252 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8918) );
  OR2_X1 U11253 ( .A1(n14545), .A2(n8918), .ZN(n8919) );
  NAND2_X1 U11254 ( .A1(n14539), .A2(n8919), .ZN(n14554) );
  XNOR2_X1 U11255 ( .A(n14556), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n14555) );
  NAND2_X1 U11256 ( .A1(n14554), .A2(n14555), .ZN(n14553) );
  INV_X1 U11257 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8920) );
  OR2_X1 U11258 ( .A1(n14556), .A2(n8920), .ZN(n8921) );
  NAND2_X1 U11259 ( .A1(n14553), .A2(n8921), .ZN(n14568) );
  INV_X1 U11260 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14771) );
  MUX2_X1 U11261 ( .A(n14771), .B(P2_REG1_REG_5__SCAN_IN), .S(n14570), .Z(
        n14569) );
  NAND2_X1 U11262 ( .A1(n14568), .A2(n14569), .ZN(n14567) );
  INV_X1 U11263 ( .A(n14570), .ZN(n8944) );
  NAND2_X1 U11264 ( .A1(n8944), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11265 ( .A1(n14567), .A2(n8922), .ZN(n12620) );
  INV_X1 U11266 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14773) );
  MUX2_X1 U11267 ( .A(n14773), .B(P2_REG1_REG_6__SCAN_IN), .S(n12614), .Z(
        n12621) );
  NAND2_X1 U11268 ( .A1(n12620), .A2(n12621), .ZN(n12619) );
  OR2_X1 U11269 ( .A1(n12614), .A2(n14773), .ZN(n8923) );
  NAND2_X1 U11270 ( .A1(n12619), .A2(n8923), .ZN(n12629) );
  INV_X1 U11271 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9505) );
  MUX2_X1 U11272 ( .A(n9505), .B(P2_REG1_REG_7__SCAN_IN), .S(n12631), .Z(
        n12630) );
  NAND2_X1 U11273 ( .A1(n12629), .A2(n12630), .ZN(n12628) );
  OR2_X1 U11274 ( .A1(n12631), .A2(n9505), .ZN(n8924) );
  NAND2_X1 U11275 ( .A1(n12628), .A2(n8924), .ZN(n12643) );
  INV_X1 U11276 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14775) );
  MUX2_X1 U11277 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14775), .S(n8950), .Z(
        n12644) );
  NAND2_X1 U11278 ( .A1(n12643), .A2(n12644), .ZN(n12642) );
  NAND2_X1 U11279 ( .A1(n8950), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11280 ( .A1(n12642), .A2(n8925), .ZN(n8927) );
  OR2_X1 U11281 ( .A1(n8927), .A2(n8928), .ZN(n8991) );
  INV_X1 U11282 ( .A(n8991), .ZN(n8926) );
  AOI21_X1 U11283 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8961) );
  AOI21_X1 U11284 ( .B1(n9066), .B2(n8930), .A(n8929), .ZN(n8931) );
  OR2_X1 U11285 ( .A1(n8932), .A2(n8931), .ZN(n8935) );
  NOR2_X1 U11286 ( .A1(n8933), .A2(P2_U3088), .ZN(n12997) );
  NAND2_X1 U11287 ( .A1(n8935), .A2(n12997), .ZN(n8954) );
  INV_X1 U11288 ( .A(n13003), .ZN(n8955) );
  INV_X1 U11289 ( .A(n14665), .ZN(n14535) );
  AND2_X1 U11290 ( .A1(n8933), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11291 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9643) );
  OAI21_X1 U11292 ( .B1(n14661), .B2(n8989), .A(n9643), .ZN(n8959) );
  INV_X1 U11293 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8936) );
  XNOR2_X1 U11294 ( .A(n8939), .B(n8936), .ZN(n12609) );
  INV_X1 U11295 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10473) );
  XNOR2_X1 U11296 ( .A(n8937), .B(n10473), .ZN(n12597) );
  AND2_X1 U11297 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n12596) );
  NAND2_X1 U11298 ( .A1(n12597), .A2(n12596), .ZN(n12595) );
  NAND2_X1 U11299 ( .A1(n8937), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11300 ( .A1(n12595), .A2(n8938), .ZN(n12608) );
  NAND2_X1 U11301 ( .A1(n12609), .A2(n12608), .ZN(n12607) );
  NAND2_X1 U11302 ( .A1(n8939), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11303 ( .A1(n12607), .A2(n8940), .ZN(n14537) );
  XNOR2_X1 U11304 ( .A(n14545), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U11305 ( .A1(n14537), .A2(n14538), .ZN(n14536) );
  INV_X1 U11306 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8941) );
  OR2_X1 U11307 ( .A1(n14545), .A2(n8941), .ZN(n8942) );
  NAND2_X1 U11308 ( .A1(n14536), .A2(n8942), .ZN(n14550) );
  XNOR2_X1 U11309 ( .A(n14556), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U11310 ( .A1(n14550), .A2(n14551), .ZN(n14549) );
  OR2_X1 U11311 ( .A1(n14556), .A2(n7389), .ZN(n8943) );
  NAND2_X1 U11312 ( .A1(n14549), .A2(n8943), .ZN(n14564) );
  XNOR2_X1 U11313 ( .A(n14570), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U11314 ( .A1(n14564), .A2(n14565), .ZN(n14563) );
  NAND2_X1 U11315 ( .A1(n8944), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11316 ( .A1(n14563), .A2(n8945), .ZN(n12617) );
  INV_X1 U11317 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U11318 ( .A(n8946), .B(P2_REG2_REG_6__SCAN_IN), .S(n12614), .Z(
        n12618) );
  NAND2_X1 U11319 ( .A1(n12617), .A2(n12618), .ZN(n12616) );
  OR2_X1 U11320 ( .A1(n12614), .A2(n8946), .ZN(n8947) );
  NAND2_X1 U11321 ( .A1(n12616), .A2(n8947), .ZN(n12626) );
  MUX2_X1 U11322 ( .A(n8948), .B(P2_REG2_REG_7__SCAN_IN), .S(n12631), .Z(
        n12627) );
  NAND2_X1 U11323 ( .A1(n12626), .A2(n12627), .ZN(n12625) );
  INV_X1 U11324 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8948) );
  OR2_X1 U11325 ( .A1(n12631), .A2(n8948), .ZN(n8949) );
  NAND2_X1 U11326 ( .A1(n12625), .A2(n8949), .ZN(n12646) );
  INV_X1 U11327 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10700) );
  XNOR2_X1 U11328 ( .A(n8950), .B(n10700), .ZN(n12647) );
  NAND2_X1 U11329 ( .A1(n12646), .A2(n12647), .ZN(n12645) );
  NAND2_X1 U11330 ( .A1(n8950), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11331 ( .A1(n12645), .A2(n8951), .ZN(n8953) );
  INV_X1 U11332 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13210) );
  MUX2_X1 U11333 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13210), .S(n8989), .Z(n8952) );
  OR2_X1 U11334 ( .A1(n8953), .A2(n8952), .ZN(n8984) );
  NAND2_X1 U11335 ( .A1(n8953), .A2(n8952), .ZN(n8957) );
  INV_X1 U11336 ( .A(n8954), .ZN(n8956) );
  AOI21_X1 U11337 ( .B1(n8984), .B2(n8957), .A(n14637), .ZN(n8958) );
  AOI211_X1 U11338 ( .C1(n14535), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n8959), .B(
        n8958), .ZN(n8960) );
  OAI21_X1 U11339 ( .B1(n8961), .B2(n14633), .A(n8960), .ZN(P2_U3223) );
  INV_X1 U11340 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11341 ( .A1(n14657), .A2(n8962), .ZN(n8963) );
  OAI211_X1 U11342 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14633), .A(n8963), .B(
        n14661), .ZN(n8966) );
  INV_X1 U11343 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14765) );
  OAI22_X1 U11344 ( .A1(n14637), .A2(n8962), .B1(n14765), .B2(n14633), .ZN(
        n8965) );
  MUX2_X1 U11345 ( .A(n8966), .B(n8965), .S(n8964), .Z(n8968) );
  OAI22_X1 U11346 ( .A1(n14665), .A2(n14973), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7576), .ZN(n8967) );
  OR2_X1 U11347 ( .A1(n8968), .A2(n8967), .ZN(P2_U3214) );
  AOI21_X1 U11348 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9916), .A(n8969), .ZN(
        n8972) );
  INV_X1 U11349 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8970) );
  MUX2_X1 U11350 ( .A(n8970), .B(P1_REG1_REG_7__SCAN_IN), .S(n9979), .Z(n8971)
         );
  NOR2_X1 U11351 ( .A1(n8972), .A2(n8971), .ZN(n9194) );
  AOI211_X1 U11352 ( .C1(n8972), .C2(n8971), .A(n13737), .B(n9194), .ZN(n8982)
         );
  NAND2_X1 U11353 ( .A1(n9916), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U11354 ( .A1(n8977), .A2(n8976), .ZN(n8974) );
  INV_X1 U11355 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10000) );
  MUX2_X1 U11356 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10000), .S(n9979), .Z(n8973) );
  NAND2_X1 U11357 ( .A1(n8974), .A2(n8973), .ZN(n13707) );
  MUX2_X1 U11358 ( .A(n10000), .B(P1_REG2_REG_7__SCAN_IN), .S(n9979), .Z(n8975) );
  NAND3_X1 U11359 ( .A1(n8977), .A2(n8976), .A3(n8975), .ZN(n8978) );
  AND3_X1 U11360 ( .A1(n14387), .A2(n13707), .A3(n8978), .ZN(n8981) );
  NAND2_X1 U11361 ( .A1(n14383), .A2(n9979), .ZN(n8979) );
  NAND2_X1 U11362 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10116) );
  OAI211_X1 U11363 ( .C1(n14391), .C2(n8494), .A(n8979), .B(n10116), .ZN(n8980) );
  OR3_X1 U11364 ( .A1(n8982), .A2(n8981), .A3(n8980), .ZN(P1_U3250) );
  INV_X1 U11365 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10744) );
  MUX2_X1 U11366 ( .A(n10744), .B(P2_REG2_REG_10__SCAN_IN), .S(n10432), .Z(
        n8987) );
  NAND2_X1 U11367 ( .A1(n8989), .A2(n13210), .ZN(n8983) );
  NAND2_X1 U11368 ( .A1(n8984), .A2(n8983), .ZN(n8986) );
  OR2_X1 U11369 ( .A1(n8986), .A2(n8987), .ZN(n10415) );
  INV_X1 U11370 ( .A(n10415), .ZN(n8985) );
  AOI211_X1 U11371 ( .C1(n8987), .C2(n8986), .A(n8985), .B(n14637), .ZN(n8999)
         );
  INV_X1 U11372 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U11373 ( .A(n8988), .B(P2_REG1_REG_10__SCAN_IN), .S(n10432), .Z(
        n8994) );
  NAND2_X1 U11374 ( .A1(n8989), .A2(n13251), .ZN(n8990) );
  NAND2_X1 U11375 ( .A1(n8991), .A2(n8990), .ZN(n8993) );
  OR2_X1 U11376 ( .A1(n8993), .A2(n8994), .ZN(n10434) );
  INV_X1 U11377 ( .A(n10434), .ZN(n8992) );
  AOI211_X1 U11378 ( .C1(n8994), .C2(n8993), .A(n14633), .B(n8992), .ZN(n8998)
         );
  NAND2_X1 U11379 ( .A1(n14535), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U11380 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n9898) );
  OAI211_X1 U11381 ( .C1(n14661), .C2(n8996), .A(n8995), .B(n9898), .ZN(n8997)
         );
  OR3_X1 U11382 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(P2_U3224) );
  INV_X1 U11383 ( .A(n10790), .ZN(n9002) );
  NAND2_X1 U11384 ( .A1(n9000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9003) );
  XNOR2_X1 U11385 ( .A(n9003), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10791) );
  INV_X1 U11386 ( .A(n10791), .ZN(n9557) );
  OAI222_X1 U11387 ( .A1(n14165), .A2(n9002), .B1(n9557), .B2(P1_U3086), .C1(
        n9001), .C2(n14166), .ZN(P1_U3343) );
  OAI222_X1 U11388 ( .A1(n13010), .A2(n9107), .B1(n10648), .B2(n9002), .C1(
        P2_U3088), .C2(n14586), .ZN(P2_U3315) );
  INV_X1 U11389 ( .A(n10854), .ZN(n9008) );
  NAND2_X1 U11390 ( .A1(n9003), .A2(n9565), .ZN(n9004) );
  NAND2_X1 U11391 ( .A1(n9004), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U11392 ( .A1(n9005), .A2(n9566), .ZN(n9274) );
  OR2_X1 U11393 ( .A1(n9005), .A2(n9566), .ZN(n9006) );
  INV_X1 U11394 ( .A(n10855), .ZN(n9007) );
  OAI222_X1 U11395 ( .A1(n14165), .A2(n9008), .B1(n9007), .B2(P1_U3086), .C1(
        n9110), .C2(n14166), .ZN(P1_U3342) );
  OAI222_X1 U11396 ( .A1(n13010), .A2(n6767), .B1(n10648), .B2(n9008), .C1(
        P2_U3088), .C2(n14601), .ZN(P2_U3314) );
  INV_X1 U11397 ( .A(n12424), .ZN(n9022) );
  MUX2_X1 U11398 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9016), .Z(n9056) );
  XOR2_X1 U11399 ( .A(n9432), .B(n9056), .Z(n9060) );
  INV_X1 U11400 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9033) );
  XNOR2_X1 U11401 ( .A(n9060), .B(n6718), .ZN(n9042) );
  OR2_X1 U11402 ( .A1(n9020), .A2(n6473), .ZN(n10123) );
  NAND2_X1 U11403 ( .A1(n9347), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11404 ( .A1(n11613), .A2(n9020), .ZN(n9021) );
  AND2_X1 U11405 ( .A1(n11348), .A2(n9021), .ZN(n9028) );
  MUX2_X1 U11406 ( .A(n9037), .B(P3_U3897), .S(n9022), .Z(n12101) );
  INV_X1 U11407 ( .A(n9432), .ZN(n9058) );
  INV_X1 U11408 ( .A(n14788), .ZN(n12082) );
  INV_X1 U11409 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9027) );
  INV_X1 U11410 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9023) );
  NOR2_X1 U11411 ( .A1(n9023), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9188) );
  INV_X1 U11412 ( .A(n9188), .ZN(n9024) );
  OAI21_X1 U11413 ( .B1(n9432), .B2(n9188), .A(n6520), .ZN(n9026) );
  OR2_X1 U11414 ( .A1(n9026), .A2(n9027), .ZN(n9048) );
  INV_X1 U11415 ( .A(n9048), .ZN(n9025) );
  AOI21_X1 U11416 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9032) );
  INV_X1 U11417 ( .A(n9028), .ZN(n9030) );
  AOI22_X1 U11418 ( .A1(n14780), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9031) );
  OAI21_X1 U11419 ( .B1(n12082), .B2(n9032), .A(n9031), .ZN(n9040) );
  NAND2_X1 U11420 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n9033), .ZN(n9185) );
  INV_X1 U11421 ( .A(n9185), .ZN(n9034) );
  NAND2_X1 U11422 ( .A1(n8739), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9044) );
  OAI21_X1 U11423 ( .B1(n9432), .B2(n9034), .A(n9044), .ZN(n9035) );
  INV_X1 U11424 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9385) );
  OR2_X1 U11425 ( .A1(n9035), .A2(n9385), .ZN(n9045) );
  NAND2_X1 U11426 ( .A1(n9035), .A2(n9385), .ZN(n9038) );
  OR2_X1 U11427 ( .A1(n12424), .A2(n12069), .ZN(n9437) );
  INV_X1 U11428 ( .A(n9437), .ZN(n9036) );
  AOI21_X1 U11429 ( .B1(n9045), .B2(n9038), .A(n12109), .ZN(n9039) );
  AOI211_X1 U11430 ( .C1(n12101), .C2(n9058), .A(n9040), .B(n9039), .ZN(n9041)
         );
  OAI21_X1 U11431 ( .B1(n12113), .B2(n9042), .A(n9041), .ZN(P3_U3183) );
  INV_X1 U11432 ( .A(n12101), .ZN(n14797) );
  MUX2_X1 U11433 ( .A(n9043), .B(P3_REG2_REG_2__SCAN_IN), .S(n9513), .Z(n9047)
         );
  NAND2_X1 U11434 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U11435 ( .A1(n9046), .A2(n9047), .ZN(n9138) );
  OAI21_X1 U11436 ( .B1(n9047), .B2(n9046), .A(n9138), .ZN(n9055) );
  MUX2_X1 U11437 ( .A(n14951), .B(P3_REG1_REG_2__SCAN_IN), .S(n9513), .Z(n9050) );
  NAND2_X1 U11438 ( .A1(n9048), .A2(n6520), .ZN(n9049) );
  NAND2_X1 U11439 ( .A1(n9049), .A2(n9050), .ZN(n9143) );
  OAI21_X1 U11440 ( .B1(n9050), .B2(n9049), .A(n9143), .ZN(n9051) );
  AND2_X1 U11441 ( .A1(n14788), .A2(n9051), .ZN(n9054) );
  INV_X1 U11442 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9052) );
  OAI22_X1 U11443 ( .A1(n14804), .A2(n9052), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9522), .ZN(n9053) );
  AOI211_X1 U11444 ( .C1(n14801), .C2(n9055), .A(n9054), .B(n9053), .ZN(n9063)
         );
  INV_X1 U11445 ( .A(n9056), .ZN(n9057) );
  MUX2_X1 U11446 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12069), .Z(n9134) );
  XOR2_X1 U11447 ( .A(n9513), .B(n9134), .Z(n9135) );
  XNOR2_X1 U11448 ( .A(n9136), .B(n9135), .ZN(n9061) );
  NAND2_X1 U11449 ( .A1(n9061), .A2(n14792), .ZN(n9062) );
  OAI211_X1 U11450 ( .C1(n14797), .C2(n9141), .A(n9063), .B(n9062), .ZN(
        P3_U3184) );
  NOR2_X1 U11451 ( .A1(n9489), .A2(n9064), .ZN(n9065) );
  AND2_X1 U11452 ( .A1(n9065), .A2(n9491), .ZN(n9091) );
  INV_X1 U11453 ( .A(n9066), .ZN(n9069) );
  INV_X1 U11454 ( .A(n10289), .ZN(n9068) );
  AND3_X1 U11455 ( .A1(n14685), .A2(n9069), .A3(n14756), .ZN(n9070) );
  NAND2_X1 U11456 ( .A1(n9072), .A2(n9071), .ZN(n9074) );
  XNOR2_X1 U11457 ( .A(n9074), .B(n9073), .ZN(n9095) );
  NAND2_X1 U11458 ( .A1(n6487), .A2(n8271), .ZN(n9077) );
  OR2_X1 U11459 ( .A1(n9262), .A2(n10477), .ZN(n12453) );
  OAI21_X1 U11460 ( .B1(n12885), .B2(n9075), .A(n12453), .ZN(n9076) );
  NAND2_X1 U11461 ( .A1(n9095), .A2(n9077), .ZN(n9078) );
  NAND2_X1 U11462 ( .A1(n9097), .A2(n9078), .ZN(n9079) );
  XNOR2_X1 U11463 ( .A(n9262), .B(n8267), .ZN(n9117) );
  NAND2_X1 U11464 ( .A1(n6488), .A2(n8268), .ZN(n9118) );
  XNOR2_X1 U11465 ( .A(n9117), .B(n9118), .ZN(n9096) );
  INV_X1 U11466 ( .A(n9091), .ZN(n9081) );
  NAND2_X1 U11467 ( .A1(n9081), .A2(n9080), .ZN(n9085) );
  AND2_X1 U11468 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  NAND2_X1 U11469 ( .A1(n9085), .A2(n9084), .ZN(n9129) );
  NOR2_X1 U11470 ( .A1(n9129), .A2(P2_U3088), .ZN(n9182) );
  INV_X1 U11471 ( .A(n9182), .ZN(n12452) );
  AND2_X1 U11472 ( .A1(n14685), .A2(n9086), .ZN(n9087) );
  NAND2_X1 U11473 ( .A1(n9091), .A2(n9087), .ZN(n9088) );
  INV_X1 U11474 ( .A(n12569), .ZN(n12516) );
  INV_X1 U11475 ( .A(n9089), .ZN(n9090) );
  AND2_X1 U11476 ( .A1(n9091), .A2(n9090), .ZN(n12444) );
  NAND2_X1 U11477 ( .A1(n12880), .A2(n12587), .ZN(n9092) );
  OAI21_X1 U11478 ( .B1(n8378), .B2(n12773), .A(n9092), .ZN(n10306) );
  INV_X1 U11479 ( .A(n10306), .ZN(n9093) );
  OAI22_X1 U11480 ( .A1(n10309), .A2(n12516), .B1(n12429), .B2(n9093), .ZN(
        n9094) );
  AOI21_X1 U11481 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n12452), .A(n9094), .ZN(
        n9101) );
  OAI22_X1 U11482 ( .A1(n12476), .A2(n8378), .B1(n9095), .B2(n12571), .ZN(
        n9099) );
  INV_X1 U11483 ( .A(n9096), .ZN(n9098) );
  NAND3_X1 U11484 ( .A1(n9099), .A2(n9098), .A3(n9097), .ZN(n9100) );
  OAI211_X1 U11485 ( .C1(n12571), .C2(n9257), .A(n9101), .B(n9100), .ZN(
        P2_U3209) );
  NAND2_X1 U11486 ( .A1(n10711), .A2(n11009), .ZN(n9102) );
  NOR2_X1 U11487 ( .A1(n11008), .A2(n9102), .ZN(n11302) );
  NAND2_X1 U11488 ( .A1(n11302), .A2(n11303), .ZN(n11305) );
  NAND2_X1 U11489 ( .A1(n11305), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9103) );
  MUX2_X1 U11490 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9103), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9104) );
  NAND2_X1 U11491 ( .A1(n9104), .A2(n11332), .ZN(n12084) );
  XNOR2_X1 U11492 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n11298) );
  NAND2_X1 U11493 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  NAND2_X1 U11494 ( .A1(n9276), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9112) );
  XNOR2_X1 U11495 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n11284) );
  NAND2_X1 U11496 ( .A1(n11286), .A2(n11284), .ZN(n9115) );
  NAND2_X1 U11497 ( .A1(n9571), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9114) );
  AOI22_X1 U11498 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n9835), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9824), .ZN(n9214) );
  XOR2_X1 U11499 ( .A(n9215), .B(n9214), .Z(n11320) );
  INV_X1 U11500 ( .A(n11320), .ZN(n9116) );
  OAI222_X1 U11501 ( .A1(n6473), .A2(n12084), .B1(n14186), .B2(n11318), .C1(
        n12423), .C2(n9116), .ZN(P3_U3278) );
  INV_X1 U11502 ( .A(n9117), .ZN(n9119) );
  NAND2_X1 U11503 ( .A1(n9119), .A2(n9118), .ZN(n9124) );
  NAND2_X1 U11504 ( .A1(n9257), .A2(n9124), .ZN(n9128) );
  XNOR2_X1 U11505 ( .A(n14710), .B(n9262), .ZN(n9122) );
  INV_X1 U11506 ( .A(n9122), .ZN(n9299) );
  NAND2_X1 U11507 ( .A1(n6488), .A2(n12587), .ZN(n9121) );
  INV_X1 U11508 ( .A(n9121), .ZN(n9120) );
  NAND2_X1 U11509 ( .A1(n9299), .A2(n9120), .ZN(n9260) );
  NAND2_X1 U11510 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  NAND2_X1 U11511 ( .A1(n9260), .A2(n9123), .ZN(n9127) );
  INV_X1 U11512 ( .A(n9127), .ZN(n9125) );
  NAND2_X1 U11513 ( .A1(n9257), .A2(n9256), .ZN(n9305) );
  INV_X1 U11514 ( .A(n9305), .ZN(n9126) );
  AOI211_X1 U11515 ( .C1(n9128), .C2(n9127), .A(n12571), .B(n9126), .ZN(n9133)
         );
  NAND2_X1 U11516 ( .A1(n12444), .A2(n12882), .ZN(n12565) );
  INV_X1 U11517 ( .A(n12565), .ZN(n12492) );
  NAND2_X1 U11518 ( .A1(n12444), .A2(n12880), .ZN(n12561) );
  INV_X1 U11519 ( .A(n12561), .ZN(n12545) );
  AOI22_X1 U11520 ( .A1(n12492), .A2(n8268), .B1(n12545), .B2(n12586), .ZN(
        n9131) );
  AOI22_X1 U11521 ( .A1(n12569), .A2(n10785), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9130) );
  OAI211_X1 U11522 ( .C1(n12538), .C2(P2_REG3_REG_3__SCAN_IN), .A(n9131), .B(
        n9130), .ZN(n9132) );
  OR2_X1 U11523 ( .A1(n9133), .A2(n9132), .ZN(P2_U3190) );
  MUX2_X1 U11524 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12069), .Z(n9231) );
  XNOR2_X1 U11525 ( .A(n9231), .B(n9600), .ZN(n9233) );
  OAI22_X1 U11526 ( .A1(n9136), .A2(n9135), .B1(n9134), .B2(n9141), .ZN(n9234)
         );
  XOR2_X1 U11527 ( .A(n9233), .B(n9234), .Z(n9151) );
  NAND2_X1 U11528 ( .A1(n12101), .A2(n9600), .ZN(n9149) );
  INV_X1 U11529 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U11530 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9777), .ZN(n9612) );
  AOI21_X1 U11531 ( .B1(n14780), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n9612), .ZN(
        n9148) );
  NAND2_X1 U11532 ( .A1(n9141), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U11533 ( .A1(n9138), .A2(n9137), .ZN(n9235) );
  XNOR2_X1 U11534 ( .A(n9235), .B(n9600), .ZN(n9139) );
  NAND2_X1 U11535 ( .A1(P3_REG2_REG_3__SCAN_IN), .A2(n9139), .ZN(n9236) );
  OAI21_X1 U11536 ( .B1(n9139), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9236), .ZN(
        n9140) );
  NAND2_X1 U11537 ( .A1(n14801), .A2(n9140), .ZN(n9147) );
  NAND2_X1 U11538 ( .A1(n9141), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U11539 ( .A1(n9143), .A2(n9142), .ZN(n9242) );
  XNOR2_X1 U11540 ( .A(n9242), .B(n9600), .ZN(n9144) );
  NAND2_X1 U11541 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n9144), .ZN(n9243) );
  OAI21_X1 U11542 ( .B1(n9144), .B2(P3_REG1_REG_3__SCAN_IN), .A(n9243), .ZN(
        n9145) );
  NAND2_X1 U11543 ( .A1(n14788), .A2(n9145), .ZN(n9146) );
  AND4_X1 U11544 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n9150)
         );
  OAI21_X1 U11545 ( .B1(n9151), .B2(n12113), .A(n9150), .ZN(P3_U3185) );
  NAND2_X2 U11546 ( .A1(n9152), .A2(n13433), .ZN(n13063) );
  AOI22_X1 U11547 ( .A1(n14032), .A2(n13311), .B1(n9156), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9154) );
  AND2_X1 U11548 ( .A1(n9155), .A2(n9154), .ZN(n9399) );
  AOI22_X1 U11549 ( .A1(n14032), .A2(n9725), .B1(n9156), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9157) );
  NOR2_X1 U11550 ( .A1(n9399), .A2(n9398), .ZN(n9397) );
  AOI21_X1 U11551 ( .B1(n9399), .B2(n13022), .A(n9397), .ZN(n9224) );
  OR2_X1 U11552 ( .A1(n13431), .A2(n13062), .ZN(n9161) );
  NAND2_X1 U11553 ( .A1(n13432), .A2(n9725), .ZN(n9160) );
  NAND2_X1 U11554 ( .A1(n9161), .A2(n9160), .ZN(n9221) );
  XNOR2_X1 U11555 ( .A(n9222), .B(n9221), .ZN(n9223) );
  XOR2_X1 U11556 ( .A(n9224), .B(n9223), .Z(n9178) );
  OR2_X1 U11557 ( .A1(n11041), .A2(n9162), .ZN(n9171) );
  INV_X1 U11558 ( .A(n9171), .ZN(n9169) );
  NAND2_X1 U11559 ( .A1(n9163), .A2(n9169), .ZN(n9175) );
  INV_X1 U11560 ( .A(n9175), .ZN(n9168) );
  INV_X1 U11561 ( .A(n9164), .ZN(n9166) );
  AND2_X1 U11562 ( .A1(n14512), .A2(n13597), .ZN(n9167) );
  NAND2_X1 U11563 ( .A1(n9170), .A2(n9169), .ZN(n13332) );
  OR2_X1 U11564 ( .A1(n13332), .A2(n14013), .ZN(n13400) );
  INV_X1 U11565 ( .A(n13400), .ZN(n13420) );
  NAND2_X1 U11566 ( .A1(n11048), .A2(n9171), .ZN(n9174) );
  INV_X1 U11567 ( .A(n9172), .ZN(n9173) );
  NAND2_X1 U11568 ( .A1(n9174), .A2(n9173), .ZN(n9738) );
  OR2_X1 U11569 ( .A1(n9738), .A2(P1_U3086), .ZN(n11034) );
  AOI22_X1 U11570 ( .A1(n13667), .A2(n13420), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n11034), .ZN(n9177) );
  OR2_X1 U11571 ( .A1(n13332), .A2(n14015), .ZN(n13399) );
  INV_X1 U11572 ( .A(n13399), .ZN(n13419) );
  NAND2_X1 U11573 ( .A1(n14421), .A2(n9175), .ZN(n14364) );
  AOI22_X1 U11574 ( .A1(n6938), .A2(n13419), .B1(n14300), .B2(n13432), .ZN(
        n9176) );
  OAI211_X1 U11575 ( .C1(n9178), .C2(n13425), .A(n9177), .B(n9176), .ZN(
        P1_U3222) );
  INV_X1 U11576 ( .A(n8273), .ZN(n10469) );
  NOR2_X1 U11577 ( .A1(n12476), .A2(n10469), .ZN(n9181) );
  AND2_X1 U11578 ( .A1(n6488), .A2(n8273), .ZN(n9179) );
  OAI21_X1 U11579 ( .B1(n9179), .B2(n12571), .A(n12516), .ZN(n9180) );
  MUX2_X1 U11580 ( .A(n9181), .B(n9180), .S(n10477), .Z(n9184) );
  NAND2_X1 U11581 ( .A1(n12880), .A2(n8271), .ZN(n10292) );
  OAI22_X1 U11582 ( .A1(n9182), .A2(n7576), .B1(n12429), .B2(n10292), .ZN(
        n9183) );
  OR2_X1 U11583 ( .A1(n9184), .A2(n9183), .ZN(P2_U3204) );
  NOR3_X1 U11584 ( .A1(n14801), .A2(n14788), .A3(n14792), .ZN(n9192) );
  INV_X1 U11585 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9396) );
  OAI22_X1 U11586 ( .A1(n14804), .A2(n8476), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9396), .ZN(n9187) );
  NOR2_X1 U11587 ( .A1(n12109), .A2(n9185), .ZN(n9186) );
  AOI211_X1 U11588 ( .C1(n14788), .C2(n9188), .A(n9187), .B(n9186), .ZN(n9191)
         );
  MUX2_X1 U11589 ( .A(n9189), .B(n14797), .S(P3_IR_REG_0__SCAN_IN), .Z(n9190)
         );
  OAI211_X1 U11590 ( .C1(n9192), .C2(n6718), .A(n9191), .B(n9190), .ZN(
        P3_U3182) );
  INV_X1 U11591 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9193) );
  MUX2_X1 U11592 ( .A(n9193), .B(P1_REG1_REG_10__SCAN_IN), .S(n10510), .Z(
        n9198) );
  INV_X1 U11593 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9195) );
  MUX2_X1 U11594 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9195), .S(n13709), .Z(
        n13701) );
  INV_X1 U11595 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9196) );
  MUX2_X1 U11596 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9196), .S(n13725), .Z(
        n13716) );
  OAI21_X1 U11597 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n13725), .A(n13714), .ZN(
        n9197) );
  NOR2_X1 U11598 ( .A1(n9197), .A2(n9198), .ZN(n9419) );
  AOI211_X1 U11599 ( .C1(n9198), .C2(n9197), .A(n13737), .B(n9419), .ZN(n9213)
         );
  NAND2_X1 U11600 ( .A1(n9979), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U11601 ( .A1(n13707), .A2(n13706), .ZN(n9201) );
  INV_X1 U11602 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9199) );
  MUX2_X1 U11603 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9199), .S(n13709), .Z(n9200) );
  NAND2_X1 U11604 ( .A1(n9201), .A2(n9200), .ZN(n13722) );
  NAND2_X1 U11605 ( .A1(n13709), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13721) );
  NAND2_X1 U11606 ( .A1(n13722), .A2(n13721), .ZN(n9204) );
  INV_X1 U11607 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9202) );
  MUX2_X1 U11608 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9202), .S(n13725), .Z(n9203) );
  NAND2_X1 U11609 ( .A1(n9204), .A2(n9203), .ZN(n13724) );
  NAND2_X1 U11610 ( .A1(n13725), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9207) );
  INV_X1 U11611 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9205) );
  MUX2_X1 U11612 ( .A(n9205), .B(P1_REG2_REG_10__SCAN_IN), .S(n10510), .Z(
        n9206) );
  AOI21_X1 U11613 ( .B1(n13724), .B2(n9207), .A(n9206), .ZN(n9418) );
  NAND3_X1 U11614 ( .A1(n13724), .A2(n9207), .A3(n9206), .ZN(n9208) );
  NAND2_X1 U11615 ( .A1(n9208), .A2(n14387), .ZN(n9211) );
  AND2_X1 U11616 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10567) );
  AOI21_X1 U11617 ( .B1(n13746), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10567), 
        .ZN(n9210) );
  NAND2_X1 U11618 ( .A1(n14383), .A2(n10510), .ZN(n9209) );
  OAI211_X1 U11619 ( .C1(n9418), .C2(n9211), .A(n9210), .B(n9209), .ZN(n9212)
         );
  OR2_X1 U11620 ( .A1(n9213), .A2(n9212), .ZN(P1_U3253) );
  AOI22_X1 U11621 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10126), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7192), .ZN(n11329) );
  AOI22_X1 U11622 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10201), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n10203), .ZN(n9637) );
  XNOR2_X1 U11623 ( .A(n9636), .B(n9637), .ZN(n11347) );
  OAI222_X1 U11624 ( .A1(n12423), .A2(n11347), .B1(n14186), .B2(n9220), .C1(
        P3_U3151), .C2(n12091), .ZN(P3_U3276) );
  OAI22_X1 U11625 ( .A1(n9224), .A2(n9223), .B1(n9222), .B2(n9221), .ZN(n9721)
         );
  OAI22_X1 U11626 ( .A1(n9535), .A2(n13062), .B1(n14448), .B2(n13063), .ZN(
        n9717) );
  OAI22_X1 U11627 ( .A1(n9535), .A2(n13063), .B1(n14448), .B2(n13064), .ZN(
        n9225) );
  XNOR2_X1 U11628 ( .A(n9225), .B(n13022), .ZN(n9716) );
  XOR2_X1 U11629 ( .A(n9717), .B(n9716), .Z(n9720) );
  XOR2_X1 U11630 ( .A(n9721), .B(n9720), .Z(n9230) );
  INV_X1 U11631 ( .A(n14415), .ZN(n9810) );
  AOI22_X1 U11632 ( .A1(n9226), .A2(n13419), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n11034), .ZN(n9227) );
  OAI21_X1 U11633 ( .B1(n9810), .B2(n13400), .A(n9227), .ZN(n9228) );
  AOI21_X1 U11634 ( .B1(n14300), .B2(n9483), .A(n9228), .ZN(n9229) );
  OAI21_X1 U11635 ( .B1(n9230), .B2(n13425), .A(n9229), .ZN(P1_U3237) );
  MUX2_X1 U11636 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12069), .Z(n9278) );
  XNOR2_X1 U11637 ( .A(n9278), .B(n9277), .ZN(n9279) );
  INV_X1 U11638 ( .A(n9231), .ZN(n9232) );
  XOR2_X1 U11639 ( .A(n9279), .B(n9280), .Z(n9254) );
  INV_X1 U11640 ( .A(n9277), .ZN(n10004) );
  INV_X1 U11641 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U11642 ( .A1(n10004), .A2(n14863), .B1(P3_REG2_REG_4__SCAN_IN), 
        .B2(n9277), .ZN(n9239) );
  NAND2_X1 U11643 ( .A1(n9235), .A2(n9241), .ZN(n9237) );
  OAI21_X1 U11644 ( .B1(n9239), .B2(n9238), .A(n9287), .ZN(n9240) );
  NAND2_X1 U11645 ( .A1(n14801), .A2(n9240), .ZN(n9251) );
  INV_X1 U11646 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n14955) );
  AOI22_X1 U11647 ( .A1(n10004), .A2(n14955), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n9277), .ZN(n9246) );
  NAND2_X1 U11648 ( .A1(n9242), .A2(n9241), .ZN(n9244) );
  NAND2_X1 U11649 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  NAND2_X1 U11650 ( .A1(n9246), .A2(n9245), .ZN(n9285) );
  OAI21_X1 U11651 ( .B1(n9246), .B2(n9245), .A(n9285), .ZN(n9247) );
  NAND2_X1 U11652 ( .A1(n14788), .A2(n9247), .ZN(n9250) );
  NAND2_X1 U11653 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(n6473), .ZN(n10142) );
  INV_X1 U11654 ( .A(n10142), .ZN(n9248) );
  AOI21_X1 U11655 ( .B1(n14780), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n9248), .ZN(
        n9249) );
  NAND3_X1 U11656 ( .A1(n9251), .A2(n9250), .A3(n9249), .ZN(n9252) );
  AOI21_X1 U11657 ( .B1(n10004), .B2(n12101), .A(n9252), .ZN(n9253) );
  OAI21_X1 U11658 ( .B1(n9254), .B2(n12113), .A(n9253), .ZN(P3_U3186) );
  XNOR2_X1 U11659 ( .A(n9262), .B(n14717), .ZN(n9263) );
  INV_X1 U11660 ( .A(n9263), .ZN(n9255) );
  NAND2_X1 U11661 ( .A1(n6488), .A2(n12586), .ZN(n9259) );
  NAND2_X1 U11662 ( .A1(n9255), .A2(n9259), .ZN(n9258) );
  INV_X1 U11663 ( .A(n9258), .ZN(n9261) );
  XNOR2_X1 U11664 ( .A(n9263), .B(n9259), .ZN(n9306) );
  XNOR2_X1 U11666 ( .A(n9262), .B(n14727), .ZN(n9316) );
  NAND2_X1 U11667 ( .A1(n6488), .A2(n12585), .ZN(n9314) );
  XNOR2_X1 U11668 ( .A(n9316), .B(n9314), .ZN(n9264) );
  AOI22_X1 U11669 ( .A1(n12563), .A2(n12586), .B1(n12533), .B2(n9263), .ZN(
        n9265) );
  NOR2_X1 U11670 ( .A1(n9265), .A2(n9264), .ZN(n9272) );
  NAND2_X1 U11671 ( .A1(n9305), .A2(n9266), .ZN(n9304) );
  INV_X1 U11672 ( .A(n10338), .ZN(n9270) );
  OR2_X1 U11673 ( .A1(n12773), .A2(n10779), .ZN(n9267) );
  OAI21_X1 U11674 ( .B1(n9332), .B2(n12777), .A(n9267), .ZN(n10332) );
  AOI22_X1 U11675 ( .A1(n12444), .A2(n10332), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9269) );
  NAND2_X1 U11676 ( .A1(n12569), .A2(n14727), .ZN(n9268) );
  OAI211_X1 U11677 ( .C1(n12538), .C2(n9270), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U11678 ( .B1(n9272), .B2(n9304), .A(n9271), .ZN(n9273) );
  OAI21_X1 U11679 ( .B1(n9318), .B2(n12571), .A(n9273), .ZN(P2_U3199) );
  INV_X1 U11680 ( .A(n10969), .ZN(n9342) );
  NAND2_X1 U11681 ( .A1(n9274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9275) );
  XNOR2_X1 U11682 ( .A(n9275), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10970) );
  INV_X1 U11683 ( .A(n10970), .ZN(n10636) );
  OAI222_X1 U11684 ( .A1(n14165), .A2(n9342), .B1(n10636), .B2(P1_U3086), .C1(
        n9276), .C2(n14166), .ZN(P1_U3341) );
  OAI22_X1 U11685 ( .A1(n9280), .A2(n9279), .B1(n9278), .B2(n9277), .ZN(n9676)
         );
  INV_X1 U11686 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10035) );
  INV_X1 U11687 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9281) );
  MUX2_X1 U11688 ( .A(n10035), .B(n9281), .S(n12069), .Z(n9282) );
  INV_X1 U11689 ( .A(n9668), .ZN(n10018) );
  NAND2_X1 U11690 ( .A1(n9282), .A2(n10018), .ZN(n14790) );
  MUX2_X1 U11691 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12069), .Z(n9283) );
  NAND2_X1 U11692 ( .A1(n9283), .A2(n9668), .ZN(n9675) );
  NAND2_X1 U11693 ( .A1(n14790), .A2(n9675), .ZN(n9284) );
  XNOR2_X1 U11694 ( .A(n9676), .B(n9284), .ZN(n9296) );
  NAND2_X1 U11695 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n9286), .ZN(n9664) );
  OAI21_X1 U11696 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n9286), .A(n9664), .ZN(
        n9294) );
  NAND2_X1 U11697 ( .A1(P3_REG2_REG_5__SCAN_IN), .A2(n9288), .ZN(n9669) );
  OAI21_X1 U11698 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n9288), .A(n9669), .ZN(
        n9289) );
  NAND2_X1 U11699 ( .A1(n14801), .A2(n9289), .ZN(n9291) );
  NOR2_X1 U11700 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10010), .ZN(n10129) );
  INV_X1 U11701 ( .A(n10129), .ZN(n9290) );
  OAI211_X1 U11702 ( .C1(n14804), .C2(n8424), .A(n9291), .B(n9290), .ZN(n9293)
         );
  NOR2_X1 U11703 ( .A1(n14797), .A2(n9668), .ZN(n9292) );
  AOI211_X1 U11704 ( .C1(n14788), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9295)
         );
  OAI21_X1 U11705 ( .B1(n9296), .B2(n12113), .A(n9295), .ZN(P3_U3187) );
  NAND2_X1 U11706 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14560) );
  INV_X1 U11707 ( .A(n14560), .ZN(n9297) );
  AOI21_X1 U11708 ( .B1(n12569), .B2(n14717), .A(n9297), .ZN(n9298) );
  OAI21_X1 U11709 ( .B1(n12561), .B2(n10266), .A(n9298), .ZN(n9303) );
  INV_X1 U11710 ( .A(n9306), .ZN(n9300) );
  NAND3_X1 U11711 ( .A1(n12563), .A2(n9300), .A3(n9299), .ZN(n9301) );
  AOI21_X1 U11712 ( .B1(n9301), .B2(n12565), .A(n10265), .ZN(n9302) );
  AOI211_X1 U11713 ( .C1(n12558), .C2(n10269), .A(n9303), .B(n9302), .ZN(n9309) );
  OAI21_X1 U11714 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(n9307) );
  NAND2_X1 U11715 ( .A1(n9307), .A2(n12533), .ZN(n9308) );
  NAND2_X1 U11716 ( .A1(n9309), .A2(n9308), .ZN(P2_U3202) );
  XNOR2_X1 U11717 ( .A(n14737), .B(n11762), .ZN(n9310) );
  AND2_X1 U11718 ( .A1(n6488), .A2(n12584), .ZN(n9311) );
  NAND2_X1 U11719 ( .A1(n9310), .A2(n9311), .ZN(n9333) );
  INV_X1 U11720 ( .A(n9310), .ZN(n9331) );
  INV_X1 U11721 ( .A(n9311), .ZN(n9312) );
  NAND2_X1 U11722 ( .A1(n9331), .A2(n9312), .ZN(n9313) );
  NAND2_X1 U11723 ( .A1(n9333), .A2(n9313), .ZN(n9323) );
  INV_X1 U11724 ( .A(n9314), .ZN(n9315) );
  OR2_X1 U11725 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  NAND2_X1 U11726 ( .A1(n9318), .A2(n9317), .ZN(n9322) );
  INV_X1 U11727 ( .A(n9322), .ZN(n9320) );
  INV_X1 U11728 ( .A(n9334), .ZN(n9321) );
  AOI211_X1 U11729 ( .C1(n9323), .C2(n9322), .A(n12571), .B(n9321), .ZN(n9329)
         );
  INV_X1 U11730 ( .A(n9324), .ZN(n10283) );
  NAND2_X1 U11731 ( .A1(n12880), .A2(n12583), .ZN(n9325) );
  OAI21_X1 U11732 ( .B1(n10266), .B2(n12773), .A(n9325), .ZN(n10279) );
  AOI22_X1 U11733 ( .A1(n12444), .A2(n10279), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9327) );
  NAND2_X1 U11734 ( .A1(n12569), .A2(n14737), .ZN(n9326) );
  OAI211_X1 U11735 ( .C1(n12538), .C2(n10283), .A(n9327), .B(n9326), .ZN(n9328) );
  OR2_X1 U11736 ( .A1(n9329), .A2(n9328), .ZN(P2_U3211) );
  XNOR2_X1 U11737 ( .A(n9501), .B(n11762), .ZN(n9574) );
  NAND2_X1 U11738 ( .A1(n6488), .A2(n12583), .ZN(n9572) );
  XNOR2_X1 U11739 ( .A(n9574), .B(n9572), .ZN(n9335) );
  INV_X1 U11740 ( .A(n9335), .ZN(n9330) );
  AOI21_X1 U11741 ( .B1(n9334), .B2(n9330), .A(n12571), .ZN(n9337) );
  NOR3_X1 U11742 ( .A1(n12476), .A2(n9332), .A3(n9331), .ZN(n9336) );
  OAI21_X1 U11743 ( .B1(n9337), .B2(n9336), .A(n9575), .ZN(n9341) );
  AOI22_X1 U11744 ( .A1(n12882), .A2(n12584), .B1(n12880), .B2(n12582), .ZN(
        n9497) );
  OAI22_X1 U11745 ( .A1(n12429), .A2(n9497), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9338), .ZN(n9339) );
  AOI21_X1 U11746 ( .B1(n14670), .B2(n12558), .A(n9339), .ZN(n9340) );
  OAI211_X1 U11747 ( .C1(n14674), .C2(n12516), .A(n9341), .B(n9340), .ZN(
        P2_U3185) );
  OAI222_X1 U11748 ( .A1(n13010), .A2(n9343), .B1(n10648), .B2(n9342), .C1(
        P2_U3088), .C2(n14611), .ZN(P2_U3313) );
  INV_X1 U11749 ( .A(n9344), .ZN(n9345) );
  NAND2_X1 U11750 ( .A1(n9345), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9346) );
  MUX2_X1 U11751 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9346), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9348) );
  NAND2_X1 U11752 ( .A1(n11499), .A2(n9639), .ZN(n9350) );
  NAND2_X1 U11753 ( .A1(n12091), .A2(n11499), .ZN(n9349) );
  NAND2_X1 U11754 ( .A1(n11656), .A2(n9350), .ZN(n12307) );
  OAI211_X1 U11755 ( .C1(n11656), .C2(n9350), .A(n9349), .B(n12307), .ZN(n9765) );
  NAND2_X1 U11756 ( .A1(n10898), .A2(n10597), .ZN(n9351) );
  NAND2_X1 U11757 ( .A1(n12306), .A2(n12405), .ZN(n9621) );
  INV_X1 U11758 ( .A(n9621), .ZN(n9365) );
  NOR2_X1 U11759 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n9356) );
  NOR4_X1 U11760 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9355) );
  NOR4_X1 U11761 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9354) );
  NOR4_X1 U11762 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9353) );
  NAND4_X1 U11763 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n9362)
         );
  NOR4_X1 U11764 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9360) );
  NOR4_X1 U11765 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9359) );
  NOR4_X1 U11766 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9358) );
  NOR4_X1 U11767 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9357) );
  NAND4_X1 U11768 ( .A1(n9360), .A2(n9359), .A3(n9358), .A4(n9357), .ZN(n9361)
         );
  NOR2_X1 U11769 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  NAND2_X1 U11770 ( .A1(n9365), .A2(n9618), .ZN(n9461) );
  INV_X1 U11771 ( .A(n9618), .ZN(n9366) );
  NOR2_X1 U11772 ( .A1(n12306), .A2(n9366), .ZN(n9367) );
  NAND2_X1 U11773 ( .A1(n9367), .A2(n12313), .ZN(n9458) );
  INV_X1 U11774 ( .A(n9458), .ZN(n9371) );
  NAND2_X1 U11775 ( .A1(n12100), .A2(n11804), .ZN(n12308) );
  NAND2_X1 U11776 ( .A1(n11499), .A2(n9622), .ZN(n11650) );
  OR2_X1 U11777 ( .A1(n12308), .A2(n11650), .ZN(n9459) );
  NAND2_X1 U11778 ( .A1(n12091), .A2(n9639), .ZN(n12309) );
  NAND2_X1 U11779 ( .A1(n12309), .A2(n11613), .ZN(n9617) );
  OAI211_X1 U11780 ( .C1(n9371), .C2(n9459), .A(n9368), .B(n9617), .ZN(n9369)
         );
  AOI21_X1 U11781 ( .B1(n9765), .B2(n9461), .A(n9369), .ZN(n9372) );
  INV_X1 U11782 ( .A(n12309), .ZN(n9764) );
  NAND2_X1 U11783 ( .A1(n9619), .A2(n9764), .ZN(n9436) );
  NOR2_X1 U11784 ( .A1(n9436), .A2(n12310), .ZN(n9462) );
  INV_X1 U11785 ( .A(n9462), .ZN(n9370) );
  OAI22_X1 U11786 ( .A1(n9372), .A2(P3_U3151), .B1(n9371), .B2(n9370), .ZN(
        n9593) );
  NOR2_X1 U11787 ( .A1(n9593), .A2(n12404), .ZN(n9523) );
  INV_X1 U11788 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9633) );
  OR2_X1 U11789 ( .A1(n11468), .A2(n9633), .ZN(n9374) );
  OR2_X1 U11790 ( .A1(n9825), .A2(n9396), .ZN(n9373) );
  INV_X1 U11791 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U11792 ( .A1(n11433), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9376) );
  XNOR2_X1 U11793 ( .A(n9378), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9379) );
  MUX2_X1 U11794 ( .A(n9379), .B(SI_0_), .S(n6802), .Z(n12425) );
  MUX2_X1 U11795 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12425), .S(n11348), .Z(n9448)
         );
  AND2_X1 U11796 ( .A1(n14889), .A2(n9635), .ZN(n11503) );
  NOR2_X1 U11797 ( .A1(n14888), .A2(n11503), .ZN(n11626) );
  INV_X1 U11798 ( .A(n11626), .ZN(n9394) );
  NAND2_X1 U11799 ( .A1(n9765), .A2(n14886), .ZN(n9467) );
  OR2_X1 U11800 ( .A1(n9458), .A2(n9459), .ZN(n9380) );
  OAI21_X1 U11801 ( .B1(n9461), .B2(n9467), .A(n9380), .ZN(n9381) );
  NAND2_X1 U11802 ( .A1(n9619), .A2(n14916), .ZN(n9382) );
  NAND2_X1 U11803 ( .A1(n11433), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9389) );
  INV_X1 U11804 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n14903) );
  OR2_X1 U11805 ( .A1(n9825), .A2(n14903), .ZN(n9388) );
  INV_X1 U11806 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9386) );
  INV_X1 U11807 ( .A(n12030), .ZN(n14870) );
  NAND2_X1 U11808 ( .A1(n11348), .A2(n9437), .ZN(n9391) );
  OR2_X1 U11809 ( .A1(n14867), .A2(n9436), .ZN(n9392) );
  OAI22_X1 U11810 ( .A1(n11994), .A2(n9635), .B1(n14870), .B2(n11988), .ZN(
        n9393) );
  AOI21_X1 U11811 ( .B1(n9394), .B2(n11984), .A(n9393), .ZN(n9395) );
  OAI21_X1 U11812 ( .B1(n9523), .B2(n9396), .A(n9395), .ZN(P3_U3172) );
  INV_X1 U11813 ( .A(n13678), .ZN(n9401) );
  AOI21_X1 U11814 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(n11037) );
  INV_X1 U11815 ( .A(n11037), .ZN(n9400) );
  MUX2_X1 U11816 ( .A(n9401), .B(n9400), .S(n14163), .Z(n9402) );
  NOR2_X1 U11817 ( .A1(n9402), .A2(n6480), .ZN(n9403) );
  AOI211_X1 U11818 ( .C1(n9405), .C2(n9404), .A(n13668), .B(n9403), .ZN(n11063) );
  INV_X1 U11819 ( .A(n11063), .ZN(n9417) );
  MUX2_X1 U11820 ( .A(n8875), .B(P1_REG2_REG_4__SCAN_IN), .S(n9733), .Z(n9407)
         );
  NAND2_X1 U11821 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  OAI211_X1 U11822 ( .C1(n9409), .C2(n9408), .A(n14387), .B(n13694), .ZN(n9410) );
  NAND2_X1 U11823 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9747) );
  OAI211_X1 U11824 ( .C1(n14391), .C2(n7129), .A(n9410), .B(n9747), .ZN(n9415)
         );
  AOI211_X1 U11825 ( .C1(n9413), .C2(n9412), .A(n9411), .B(n13737), .ZN(n9414)
         );
  AOI211_X1 U11826 ( .C1(n14383), .C2(n9733), .A(n9415), .B(n9414), .ZN(n9416)
         );
  NAND2_X1 U11827 ( .A1(n9417), .A2(n9416), .ZN(P1_U3247) );
  AOI21_X1 U11828 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10510), .A(n9418), .ZN(
        n9547) );
  INV_X1 U11829 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9549) );
  MUX2_X1 U11830 ( .A(n9549), .B(P1_REG2_REG_11__SCAN_IN), .S(n10574), .Z(
        n9546) );
  XNOR2_X1 U11831 ( .A(n9547), .B(n9546), .ZN(n9428) );
  INV_X1 U11832 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9420) );
  MUX2_X1 U11833 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9420), .S(n10574), .Z(
        n9421) );
  OAI21_X1 U11834 ( .B1(n9422), .B2(n9421), .A(n9553), .ZN(n9423) );
  NAND2_X1 U11835 ( .A1(n9423), .A2(n14386), .ZN(n9427) );
  NAND2_X1 U11836 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14304)
         );
  INV_X1 U11837 ( .A(n14304), .ZN(n9425) );
  NOR2_X1 U11838 ( .A1(n13772), .A2(n9550), .ZN(n9424) );
  AOI211_X1 U11839 ( .C1(n13746), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9425), .B(
        n9424), .ZN(n9426) );
  OAI211_X1 U11840 ( .C1(n13773), .C2(n9428), .A(n9427), .B(n9426), .ZN(
        P1_U3254) );
  AND2_X2 U11841 ( .A1(n11348), .A2(n7672), .ZN(n11453) );
  OR2_X1 U11842 ( .A1(n10155), .A2(n9431), .ZN(n9434) );
  OR2_X1 U11843 ( .A1(n11348), .A2(n9432), .ZN(n9433) );
  INV_X1 U11844 ( .A(n14887), .ZN(n9446) );
  INV_X1 U11845 ( .A(n14889), .ZN(n9439) );
  INV_X1 U11846 ( .A(n9436), .ZN(n9438) );
  NAND2_X1 U11847 ( .A1(n9438), .A2(n14890), .ZN(n11659) );
  OAI22_X1 U11848 ( .A1(n9439), .A2(n12009), .B1(n9769), .B2(n11988), .ZN(
        n9440) );
  AOI21_X1 U11849 ( .B1(n9446), .B2(n12017), .A(n9440), .ZN(n9456) );
  INV_X1 U11850 ( .A(n11650), .ZN(n9441) );
  NAND2_X1 U11851 ( .A1(n12405), .A2(n9441), .ZN(n9443) );
  OAI21_X1 U11852 ( .B1(n12091), .B2(n9466), .A(n9639), .ZN(n9442) );
  AND2_X4 U11853 ( .A1(n9443), .A2(n9442), .ZN(n11892) );
  OR2_X1 U11854 ( .A1(n12030), .A2(n14887), .ZN(n11501) );
  NAND3_X1 U11855 ( .A1(n12030), .A2(n9446), .A3(n11892), .ZN(n9447) );
  AND2_X1 U11856 ( .A1(n9510), .A2(n9447), .ZN(n9453) );
  NAND2_X1 U11857 ( .A1(n14889), .A2(n9448), .ZN(n14895) );
  NAND2_X1 U11858 ( .A1(n12030), .A2(n14887), .ZN(n11507) );
  INV_X1 U11859 ( .A(n14895), .ZN(n9449) );
  AOI21_X1 U11860 ( .B1(n9760), .B2(n11844), .A(n9449), .ZN(n9450) );
  INV_X1 U11861 ( .A(n14888), .ZN(n9451) );
  NAND2_X1 U11862 ( .A1(n11507), .A2(n11501), .ZN(n14894) );
  NAND3_X1 U11863 ( .A1(n9451), .A2(n14894), .A3(n6828), .ZN(n9452) );
  OAI211_X1 U11864 ( .C1(n9453), .C2(n14895), .A(n9511), .B(n9452), .ZN(n9454)
         );
  NAND2_X1 U11865 ( .A1(n9454), .A2(n11984), .ZN(n9455) );
  OAI211_X1 U11866 ( .C1(n9523), .C2(n14903), .A(n9456), .B(n9455), .ZN(
        P3_U3162) );
  INV_X1 U11867 ( .A(n9765), .ZN(n9457) );
  OAI22_X1 U11868 ( .A1(n9461), .A2(n9459), .B1(n9458), .B2(n9457), .ZN(n9460)
         );
  NAND2_X1 U11869 ( .A1(n9460), .A2(n9619), .ZN(n9465) );
  INV_X1 U11870 ( .A(n9461), .ZN(n9463) );
  NAND2_X1 U11871 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  NAND2_X1 U11872 ( .A1(n9622), .A2(n9466), .ZN(n11655) );
  AOI21_X1 U11873 ( .B1(n14873), .B2(n9467), .A(n11626), .ZN(n9468) );
  AOI21_X1 U11874 ( .B1(n14891), .B2(n12030), .A(n9468), .ZN(n9629) );
  OAI21_X1 U11875 ( .B1(n9635), .B2(n14886), .A(n9629), .ZN(n12387) );
  NAND2_X1 U11876 ( .A1(n12387), .A2(n14948), .ZN(n9469) );
  OAI21_X1 U11877 ( .B1(n9375), .B2(n14948), .A(n9469), .ZN(P3_U3390) );
  OAI21_X1 U11878 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n14451) );
  INV_X1 U11879 ( .A(n14451), .ZN(n9486) );
  OAI21_X1 U11880 ( .B1(n13610), .B2(n9474), .A(n9473), .ZN(n9476) );
  OAI22_X1 U11881 ( .A1(n9810), .A2(n14013), .B1(n13431), .B2(n14015), .ZN(
        n9475) );
  AOI21_X1 U11882 ( .B1(n9476), .B2(n14411), .A(n9475), .ZN(n9477) );
  OAI21_X1 U11883 ( .B1(n9486), .B2(n13824), .A(n9477), .ZN(n14449) );
  NAND2_X1 U11884 ( .A1(n14449), .A2(n14419), .ZN(n9485) );
  INV_X1 U11885 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9478) );
  OAI22_X1 U11886 ( .A1(n14419), .A2(n8857), .B1(n9478), .B2(n14421), .ZN(
        n9482) );
  INV_X1 U11887 ( .A(n9479), .ZN(n9480) );
  OAI211_X1 U11888 ( .C1(n14448), .C2(n9530), .A(n9480), .B(n14429), .ZN(
        n14447) );
  NOR2_X1 U11889 ( .A1(n14447), .A2(n14022), .ZN(n9481) );
  AOI211_X1 U11890 ( .C1(n14033), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9484)
         );
  OAI211_X1 U11891 ( .C1(n9486), .C2(n13886), .A(n9485), .B(n9484), .ZN(
        P1_U3291) );
  NOR2_X1 U11892 ( .A1(n9488), .A2(n9487), .ZN(n9490) );
  AND2_X1 U11893 ( .A1(n14685), .A2(n9489), .ZN(n14686) );
  OAI21_X1 U11894 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n14676) );
  INV_X1 U11895 ( .A(n14676), .ZN(n9503) );
  XNOR2_X1 U11896 ( .A(n9496), .B(n9495), .ZN(n9499) );
  INV_X1 U11897 ( .A(n9497), .ZN(n9498) );
  AOI21_X1 U11898 ( .B1(n9499), .B2(n12879), .A(n9498), .ZN(n14679) );
  INV_X1 U11899 ( .A(n10281), .ZN(n9500) );
  AOI211_X1 U11900 ( .C1(n9501), .C2(n9500), .A(n12865), .B(n10702), .ZN(
        n14668) );
  AOI21_X1 U11901 ( .B1(n14738), .B2(n9501), .A(n14668), .ZN(n9502) );
  OAI211_X1 U11902 ( .C1(n9503), .C2(n14720), .A(n14679), .B(n9502), .ZN(n9507) );
  NAND2_X1 U11903 ( .A1(n9507), .A2(n14779), .ZN(n9504) );
  OAI21_X1 U11904 ( .B1(n14779), .B2(n9505), .A(n9504), .ZN(P2_U3506) );
  INV_X1 U11905 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U11906 ( .A1(n9507), .A2(n14764), .ZN(n9508) );
  OAI21_X1 U11907 ( .B1(n14764), .B2(n9509), .A(n9508), .ZN(P2_U3451) );
  NAND2_X1 U11908 ( .A1(n9511), .A2(n9510), .ZN(n9598) );
  NAND2_X1 U11909 ( .A1(n11453), .A2(n9512), .ZN(n9516) );
  OR2_X1 U11910 ( .A1(n10155), .A2(SI_2_), .ZN(n9515) );
  OR2_X1 U11911 ( .A1(n11348), .A2(n9513), .ZN(n9514) );
  XNOR2_X1 U11912 ( .A(n9761), .B(n11892), .ZN(n9594) );
  XNOR2_X1 U11913 ( .A(n9594), .B(n9769), .ZN(n9597) );
  XOR2_X1 U11914 ( .A(n9598), .B(n9597), .Z(n9527) );
  INV_X2 U11915 ( .A(n9828), .ZN(n11465) );
  NAND2_X1 U11916 ( .A1(n11465), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9521) );
  INV_X1 U11917 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9517) );
  OR2_X1 U11918 ( .A1(n9605), .A2(n9517), .ZN(n9520) );
  OR2_X1 U11919 ( .A1(n9825), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9519) );
  INV_X1 U11920 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9776) );
  INV_X1 U11921 ( .A(n14853), .ZN(n14868) );
  OAI22_X1 U11922 ( .A1(n14870), .A2(n12009), .B1(n14868), .B2(n11988), .ZN(
        n9525) );
  NOR2_X1 U11923 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  AOI211_X1 U11924 ( .C1(n9761), .C2(n12017), .A(n9525), .B(n9524), .ZN(n9526)
         );
  OAI21_X1 U11925 ( .B1(n12019), .B2(n9527), .A(n9526), .ZN(P3_U3177) );
  INV_X1 U11926 ( .A(n9528), .ZN(n13609) );
  AND2_X1 U11927 ( .A1(n13432), .A2(n14032), .ZN(n9529) );
  NOR2_X1 U11928 ( .A1(n9530), .A2(n9529), .ZN(n9539) );
  XNOR2_X1 U11929 ( .A(n9539), .B(n9226), .ZN(n9531) );
  MUX2_X1 U11930 ( .A(n13609), .B(n9531), .S(n9534), .Z(n9538) );
  OAI21_X1 U11931 ( .B1(n9528), .B2(n9533), .A(n9532), .ZN(n14445) );
  OAI22_X1 U11932 ( .A1(n9535), .A2(n14013), .B1(n9534), .B2(n14015), .ZN(
        n9536) );
  AOI21_X1 U11933 ( .B1(n14445), .B2(n14507), .A(n9536), .ZN(n9537) );
  OAI21_X1 U11934 ( .B1(n14501), .B2(n9538), .A(n9537), .ZN(n14443) );
  INV_X1 U11935 ( .A(n14443), .ZN(n9544) );
  INV_X1 U11936 ( .A(n13886), .ZN(n14407) );
  NAND2_X1 U11937 ( .A1(n9539), .A2(n14429), .ZN(n14442) );
  AOI22_X1 U11938 ( .A1(n6479), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14400), .ZN(n9541) );
  NAND2_X1 U11939 ( .A1(n14033), .A2(n13432), .ZN(n9540) );
  OAI211_X1 U11940 ( .C1(n14442), .C2(n14022), .A(n9541), .B(n9540), .ZN(n9542) );
  AOI21_X1 U11941 ( .B1(n14445), .B2(n14407), .A(n9542), .ZN(n9543) );
  OAI21_X1 U11942 ( .B1(n9544), .B2(n6479), .A(n9543), .ZN(P1_U3292) );
  INV_X1 U11943 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9545) );
  AOI22_X1 U11944 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9557), .B1(n10791), 
        .B2(n9545), .ZN(n9552) );
  OR2_X1 U11945 ( .A1(n9547), .A2(n9546), .ZN(n9548) );
  OAI21_X1 U11946 ( .B1(n9550), .B2(n9549), .A(n9548), .ZN(n9551) );
  NOR2_X1 U11947 ( .A1(n9552), .A2(n9551), .ZN(n9872) );
  AOI21_X1 U11948 ( .B1(n9552), .B2(n9551), .A(n9872), .ZN(n9561) );
  INV_X1 U11949 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U11950 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n10791), .B1(n9557), 
        .B2(n14220), .ZN(n9555) );
  OAI21_X1 U11951 ( .B1(n9555), .B2(n9554), .A(n9866), .ZN(n9559) );
  AOI22_X1 U11952 ( .A1(n13746), .A2(P1_ADDR_REG_12__SCAN_IN), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(P1_U3086), .ZN(n9556) );
  OAI21_X1 U11953 ( .B1(n9557), .B2(n13772), .A(n9556), .ZN(n9558) );
  AOI21_X1 U11954 ( .B1(n9559), .B2(n14386), .A(n9558), .ZN(n9560) );
  OAI21_X1 U11955 ( .B1(n9561), .B2(n13773), .A(n9560), .ZN(P1_U3255) );
  INV_X1 U11956 ( .A(n11066), .ZN(n9570) );
  OAI222_X1 U11957 ( .A1(n10445), .A2(P2_U3088), .B1(n10648), .B2(n9570), .C1(
        n9562), .C2(n13010), .ZN(P2_U3312) );
  INV_X1 U11958 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9563) );
  NAND4_X1 U11959 ( .A1(n9566), .A2(n9565), .A3(n9564), .A4(n9563), .ZN(n9567)
         );
  OAI21_X1 U11960 ( .B1(n9568), .B2(n9567), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9569) );
  XNOR2_X1 U11961 ( .A(n9569), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14384) );
  INV_X1 U11962 ( .A(n14384), .ZN(n10628) );
  OAI222_X1 U11963 ( .A1(n14166), .A2(n9571), .B1(n14165), .B2(n9570), .C1(
        P1_U3086), .C2(n10628), .ZN(P1_U3340) );
  INV_X1 U11964 ( .A(n9572), .ZN(n9573) );
  XNOR2_X1 U11965 ( .A(n10705), .B(n11743), .ZN(n9577) );
  NAND2_X1 U11966 ( .A1(n6488), .A2(n12582), .ZN(n9578) );
  NAND2_X1 U11967 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  NAND2_X1 U11968 ( .A1(n9583), .A2(n9576), .ZN(n9580) );
  INV_X1 U11969 ( .A(n9577), .ZN(n9585) );
  INV_X1 U11970 ( .A(n9578), .ZN(n9579) );
  NAND2_X1 U11971 ( .A1(n9585), .A2(n9579), .ZN(n9581) );
  INV_X1 U11972 ( .A(n9580), .ZN(n9582) );
  NAND2_X1 U11973 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  AOI22_X1 U11974 ( .A1(n9640), .A2(n9585), .B1(n9584), .B2(n9583), .ZN(n9592)
         );
  AOI22_X1 U11975 ( .A1(n12545), .A2(n12581), .B1(n12558), .B2(n9586), .ZN(
        n9587) );
  NAND2_X1 U11976 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n12639) );
  OAI211_X1 U11977 ( .C1(n9588), .C2(n12565), .A(n9587), .B(n12639), .ZN(n9589) );
  AOI21_X1 U11978 ( .B1(n10705), .B2(n12569), .A(n9589), .ZN(n9591) );
  NAND3_X1 U11979 ( .A1(n9640), .A2(n12563), .A3(n12582), .ZN(n9590) );
  OAI211_X1 U11980 ( .C1(n9592), .C2(n12571), .A(n9591), .B(n9590), .ZN(
        P2_U3193) );
  INV_X1 U11981 ( .A(n9594), .ZN(n9595) );
  AND2_X1 U11982 ( .A1(n9595), .A2(n9769), .ZN(n9596) );
  OR2_X1 U11983 ( .A1(n11348), .A2(n9600), .ZN(n9601) );
  OAI211_X1 U11984 ( .C1(n10155), .C2(SI_3_), .A(n9602), .B(n9601), .ZN(n9762)
         );
  XNOR2_X1 U11985 ( .A(n11892), .B(n9762), .ZN(n10052) );
  XNOR2_X1 U11986 ( .A(n10052), .B(n14853), .ZN(n9603) );
  NAND2_X1 U11987 ( .A1(n9604), .A2(n9603), .ZN(n10055) );
  OAI211_X1 U11988 ( .C1(n9604), .C2(n9603), .A(n10055), .B(n11984), .ZN(n9616) );
  INV_X1 U11989 ( .A(n9762), .ZN(n14917) );
  NAND2_X1 U11990 ( .A1(n11465), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9611) );
  INV_X1 U11991 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9606) );
  OR2_X1 U11992 ( .A1(n9605), .A2(n9606), .ZN(n9610) );
  NOR2_X1 U11993 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n10011) );
  AND2_X1 U11994 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9607) );
  NOR2_X1 U11995 ( .A1(n10011), .A2(n9607), .ZN(n14859) );
  OR2_X1 U11996 ( .A1(n11400), .A2(n14859), .ZN(n9609) );
  OR2_X1 U11997 ( .A1(n11468), .A2(n14863), .ZN(n9608) );
  AND4_X2 U11998 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9608), .ZN(n10131)
         );
  AOI21_X1 U11999 ( .B1(n12029), .B2(n12013), .A(n9612), .ZN(n9613) );
  OAI21_X1 U12000 ( .B1(n9769), .B2(n12009), .A(n9613), .ZN(n9614) );
  AOI21_X1 U12001 ( .B1(n14917), .B2(n12017), .A(n9614), .ZN(n9615) );
  OAI211_X1 U12002 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12003), .A(n9616), .B(
        n9615), .ZN(P3_U3158) );
  AND3_X1 U12003 ( .A1(n9619), .A2(n9618), .A3(n9617), .ZN(n9620) );
  NAND2_X1 U12004 ( .A1(n11804), .A2(n9622), .ZN(n9623) );
  AND2_X1 U12005 ( .A1(n9766), .A2(n12310), .ZN(n12315) );
  INV_X1 U12006 ( .A(n12315), .ZN(n9624) );
  OR2_X1 U12007 ( .A1(n12306), .A2(n9624), .ZN(n9625) );
  OAI21_X1 U12008 ( .B1(n12405), .B2(n12315), .A(n9625), .ZN(n9626) );
  INV_X1 U12009 ( .A(n9626), .ZN(n9627) );
  NAND2_X1 U12010 ( .A1(n12317), .A2(n9627), .ZN(n9631) );
  INV_X1 U12011 ( .A(n9631), .ZN(n9628) );
  NAND2_X1 U12012 ( .A1(n9628), .A2(n14901), .ZN(n12117) );
  OR2_X1 U12013 ( .A1(n12117), .A2(n14886), .ZN(n12252) );
  INV_X1 U12014 ( .A(n9629), .ZN(n9630) );
  AOI21_X1 U12015 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n14884), .A(n9630), .ZN(
        n9632) );
  MUX2_X1 U12016 ( .A(n9633), .B(n9632), .S(n14228), .Z(n9634) );
  OAI21_X1 U12017 ( .B1(n9635), .B2(n12252), .A(n9634), .ZN(P3_U3233) );
  XNOR2_X1 U12018 ( .A(n9755), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11360) );
  INV_X1 U12019 ( .A(n11360), .ZN(n9638) );
  OAI222_X1 U12020 ( .A1(P3_U3151), .A2(n9639), .B1(n12423), .B2(n9638), .C1(
        n11361), .C2(n14186), .ZN(P3_U3275) );
  XNOR2_X1 U12021 ( .A(n10324), .B(n11762), .ZN(n9901) );
  NOR2_X1 U12022 ( .A1(n12885), .A2(n10738), .ZN(n9903) );
  XNOR2_X1 U12023 ( .A(n9901), .B(n9903), .ZN(n9641) );
  OAI21_X1 U12024 ( .B1(n9640), .B2(n9641), .A(n9902), .ZN(n9642) );
  NAND2_X1 U12025 ( .A1(n9642), .A2(n12533), .ZN(n9646) );
  AOI22_X1 U12026 ( .A1(n12882), .A2(n12582), .B1(n12880), .B2(n12580), .ZN(
        n9650) );
  OAI21_X1 U12027 ( .B1(n12429), .B2(n9650), .A(n9643), .ZN(n9644) );
  AOI21_X1 U12028 ( .B1(n10322), .B2(n12558), .A(n9644), .ZN(n9645) );
  OAI211_X1 U12029 ( .C1(n10324), .C2(n12516), .A(n9646), .B(n9645), .ZN(
        P2_U3203) );
  XNOR2_X1 U12030 ( .A(n9647), .B(n9648), .ZN(n10330) );
  AOI21_X1 U12031 ( .B1(n9649), .B2(n9648), .A(n12774), .ZN(n9653) );
  INV_X1 U12032 ( .A(n9650), .ZN(n9651) );
  AOI21_X1 U12033 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n10325) );
  AOI21_X1 U12034 ( .B1(n10701), .B2(n9655), .A(n12865), .ZN(n9654) );
  AND2_X1 U12035 ( .A1(n9654), .A2(n10745), .ZN(n10328) );
  AOI21_X1 U12036 ( .B1(n14738), .B2(n9655), .A(n10328), .ZN(n9656) );
  OAI211_X1 U12037 ( .C1(n10330), .C2(n14720), .A(n10325), .B(n9656), .ZN(
        n9658) );
  NAND2_X1 U12038 ( .A1(n9658), .A2(n14779), .ZN(n9657) );
  OAI21_X1 U12039 ( .B1(n14779), .B2(n13251), .A(n9657), .ZN(P2_U3508) );
  INV_X1 U12040 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12041 ( .A1(n9658), .A2(n14764), .ZN(n9659) );
  OAI21_X1 U12042 ( .B1(n14764), .B2(n9660), .A(n9659), .ZN(P2_U3457) );
  INV_X1 U12043 ( .A(n11070), .ZN(n9753) );
  NAND2_X1 U12044 ( .A1(n9661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9662) );
  XNOR2_X1 U12045 ( .A(n9662), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13736) );
  INV_X1 U12046 ( .A(n13736), .ZN(n10640) );
  OAI222_X1 U12047 ( .A1(n14165), .A2(n9753), .B1(n10640), .B2(P1_U3086), .C1(
        n6812), .C2(n14166), .ZN(P1_U3339) );
  INV_X1 U12048 ( .A(n9704), .ZN(n10156) );
  INV_X1 U12049 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n14958) );
  MUX2_X1 U12050 ( .A(n14958), .B(P3_REG1_REG_6__SCAN_IN), .S(n9677), .Z(
        n14785) );
  NAND2_X1 U12051 ( .A1(n9668), .A2(n9663), .ZN(n9665) );
  NAND2_X1 U12052 ( .A1(n9665), .A2(n9664), .ZN(n14786) );
  NAND2_X1 U12053 ( .A1(n14785), .A2(n14786), .ZN(n14784) );
  XNOR2_X1 U12054 ( .A(n10156), .B(n9698), .ZN(n9666) );
  NAND2_X1 U12055 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n9666), .ZN(n9699) );
  OAI21_X1 U12056 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n9666), .A(n9699), .ZN(
        n9691) );
  INV_X1 U12057 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n14845) );
  AOI22_X1 U12058 ( .A1(n9677), .A2(n14845), .B1(P3_REG2_REG_6__SCAN_IN), .B2(
        n14796), .ZN(n14783) );
  NAND2_X1 U12059 ( .A1(n9668), .A2(n9667), .ZN(n9670) );
  NAND2_X1 U12060 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(n9671), .ZN(n9705) );
  OAI21_X1 U12061 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n9671), .A(n9705), .ZN(
        n9672) );
  NAND2_X1 U12062 ( .A1(n9672), .A2(n14801), .ZN(n9674) );
  AND2_X1 U12063 ( .A1(n6473), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10234) );
  AOI21_X1 U12064 ( .B1(n14780), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10234), .ZN(
        n9673) );
  OAI211_X1 U12065 ( .C1(n14797), .C2(n9704), .A(n9674), .B(n9673), .ZN(n9690)
         );
  NAND2_X1 U12066 ( .A1(n9676), .A2(n9675), .ZN(n14791) );
  MUX2_X1 U12067 ( .A(n14845), .B(n14958), .S(n12069), .Z(n9678) );
  NAND2_X1 U12068 ( .A1(n9678), .A2(n9677), .ZN(n9681) );
  INV_X1 U12069 ( .A(n9678), .ZN(n9679) );
  NAND2_X1 U12070 ( .A1(n9679), .A2(n14796), .ZN(n9680) );
  NAND2_X1 U12071 ( .A1(n9681), .A2(n9680), .ZN(n14789) );
  INV_X1 U12072 ( .A(n9681), .ZN(n9687) );
  INV_X1 U12073 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10072) );
  INV_X1 U12074 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U12075 ( .A(n10072), .B(n9682), .S(n12069), .Z(n9683) );
  NAND2_X1 U12076 ( .A1(n9683), .A2(n10156), .ZN(n9693) );
  INV_X1 U12077 ( .A(n9683), .ZN(n9684) );
  NAND2_X1 U12078 ( .A1(n9684), .A2(n9704), .ZN(n9685) );
  AND2_X1 U12079 ( .A1(n9693), .A2(n9685), .ZN(n9686) );
  OR3_X1 U12080 ( .A1(n14794), .A2(n9687), .A3(n9686), .ZN(n9688) );
  AOI21_X1 U12081 ( .B1(n9694), .B2(n9688), .A(n12113), .ZN(n9689) );
  AOI211_X1 U12082 ( .C1(n14788), .C2(n9691), .A(n9690), .B(n9689), .ZN(n9692)
         );
  INV_X1 U12083 ( .A(n9692), .ZN(P3_U3189) );
  MUX2_X1 U12084 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12069), .Z(n9837) );
  XNOR2_X1 U12085 ( .A(n9837), .B(n9849), .ZN(n9695) );
  OAI21_X1 U12086 ( .B1(n9696), .B2(n9695), .A(n9836), .ZN(n9697) );
  NAND2_X1 U12087 ( .A1(n9697), .A2(n14792), .ZN(n9715) );
  INV_X1 U12088 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U12089 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10362), .B1(n9849), .B2(
        n14961), .ZN(n9702) );
  NAND2_X1 U12090 ( .A1(n9704), .A2(n9698), .ZN(n9700) );
  NAND2_X1 U12091 ( .A1(n9702), .A2(n9701), .ZN(n9845) );
  OAI21_X1 U12092 ( .B1(n9702), .B2(n9701), .A(n9845), .ZN(n9713) );
  INV_X1 U12093 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U12094 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10362), .B1(n9849), .B2(
        n9848), .ZN(n9708) );
  NAND2_X1 U12095 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  OAI21_X1 U12096 ( .B1(n9708), .B2(n9707), .A(n9847), .ZN(n9709) );
  NAND2_X1 U12097 ( .A1(n9709), .A2(n14801), .ZN(n9711) );
  NOR2_X1 U12098 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10163), .ZN(n10460) );
  AOI21_X1 U12099 ( .B1(n14780), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10460), .ZN(
        n9710) );
  OAI211_X1 U12100 ( .C1(n14797), .C2(n10362), .A(n9711), .B(n9710), .ZN(n9712) );
  AOI21_X1 U12101 ( .B1(n14788), .B2(n9713), .A(n9712), .ZN(n9714) );
  NAND2_X1 U12102 ( .A1(n9715), .A2(n9714), .ZN(P3_U3190) );
  INV_X1 U12103 ( .A(n9716), .ZN(n9719) );
  INV_X1 U12104 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U12105 ( .A1(n14415), .A2(n9725), .ZN(n9723) );
  NAND2_X1 U12106 ( .A1(n14363), .A2(n13311), .ZN(n9722) );
  NAND2_X1 U12107 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  XNOR2_X1 U12108 ( .A(n9724), .B(n13022), .ZN(n9727) );
  AND2_X1 U12109 ( .A1(n14363), .A2(n9725), .ZN(n9726) );
  AOI21_X1 U12110 ( .B1(n14415), .B2(n13313), .A(n9726), .ZN(n9728) );
  XNOR2_X1 U12111 ( .A(n9727), .B(n9728), .ZN(n14368) );
  NAND2_X1 U12112 ( .A1(n14369), .A2(n14368), .ZN(n14367) );
  OR2_X1 U12113 ( .A1(n9977), .A2(n9731), .ZN(n9736) );
  OR2_X1 U12114 ( .A1(n13574), .A2(n9732), .ZN(n9735) );
  INV_X2 U12115 ( .A(n11132), .ZN(n11102) );
  NAND2_X1 U12116 ( .A1(n11102), .A2(n9733), .ZN(n9734) );
  OAI22_X1 U12117 ( .A1(n13454), .A2(n13062), .B1(n14461), .B2(n13063), .ZN(
        n9781) );
  OAI22_X1 U12118 ( .A1(n13454), .A2(n13063), .B1(n14461), .B2(n13064), .ZN(
        n9737) );
  XNOR2_X1 U12119 ( .A(n9737), .B(n13022), .ZN(n9782) );
  XOR2_X1 U12120 ( .A(n9783), .B(n9782), .Z(n9751) );
  NAND2_X1 U12121 ( .A1(n9739), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9746) );
  INV_X1 U12122 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9740) );
  NOR2_X1 U12123 ( .A1(n9741), .A2(n9740), .ZN(n9793) );
  AND2_X1 U12124 ( .A1(n9741), .A2(n9740), .ZN(n9742) );
  NOR2_X1 U12125 ( .A1(n9793), .A2(n9742), .ZN(n9807) );
  NAND2_X1 U12126 ( .A1(n11208), .A2(n9807), .ZN(n9745) );
  NAND2_X1 U12127 ( .A1(n8606), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U12128 ( .A1(n13579), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9743) );
  NAND4_X1 U12129 ( .A1(n9746), .A2(n9745), .A3(n9744), .A4(n9743), .ZN(n14414) );
  AOI22_X1 U12130 ( .A1(n13420), .A2(n14414), .B1(n13419), .B2(n14415), .ZN(
        n9748) );
  OAI211_X1 U12131 ( .C1(n14420), .C2(n14376), .A(n9748), .B(n9747), .ZN(n9749) );
  AOI21_X1 U12132 ( .B1(n14300), .B2(n13608), .A(n9749), .ZN(n9750) );
  OAI21_X1 U12133 ( .B1(n9751), .B2(n13425), .A(n9750), .ZN(P1_U3230) );
  INV_X1 U12134 ( .A(n14643), .ZN(n9754) );
  OAI222_X1 U12135 ( .A1(P2_U3088), .A2(n9754), .B1(n10648), .B2(n9753), .C1(
        n9752), .C2(n13010), .ZN(P2_U3311) );
  NAND2_X1 U12136 ( .A1(n9755), .A2(n10481), .ZN(n9758) );
  NAND2_X1 U12137 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9756), .ZN(n9757) );
  AOI22_X1 U12138 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n10646), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n7231), .ZN(n9858) );
  XNOR2_X1 U12139 ( .A(n9859), .B(n7032), .ZN(n11371) );
  INV_X1 U12140 ( .A(n11371), .ZN(n9759) );
  INV_X1 U12141 ( .A(SI_21_), .ZN(n11372) );
  OAI222_X1 U12142 ( .A1(n12423), .A2(n9759), .B1(n14186), .B2(n11372), .C1(
        n6473), .C2(n11499), .ZN(P3_U3274) );
  INV_X1 U12143 ( .A(n9761), .ZN(n14880) );
  NAND2_X1 U12144 ( .A1(n14892), .A2(n14880), .ZN(n11509) );
  NAND2_X1 U12145 ( .A1(n9769), .A2(n9761), .ZN(n11508) );
  AND2_X1 U12146 ( .A1(n11509), .A2(n11508), .ZN(n14872) );
  NAND2_X1 U12147 ( .A1(n14866), .A2(n14872), .ZN(n14865) );
  OR2_X2 U12148 ( .A1(n14853), .A2(n9762), .ZN(n14847) );
  NAND2_X1 U12149 ( .A1(n14853), .A2(n9762), .ZN(n11516) );
  INV_X1 U12150 ( .A(n9771), .ZN(n11629) );
  OAI21_X1 U12151 ( .B1(n9763), .B2(n11629), .A(n14848), .ZN(n14918) );
  INV_X1 U12152 ( .A(n14918), .ZN(n9780) );
  NOR2_X1 U12153 ( .A1(n14901), .A2(n11499), .ZN(n14881) );
  NAND2_X1 U12154 ( .A1(n14228), .A2(n14881), .ZN(n14904) );
  NAND3_X1 U12155 ( .A1(n9765), .A2(n9764), .A3(n14886), .ZN(n9767) );
  OAI22_X1 U12156 ( .A1(n9769), .A2(n14869), .B1(n10131), .B2(n14867), .ZN(
        n9775) );
  NAND2_X1 U12157 ( .A1(n14894), .A2(n14895), .ZN(n14893) );
  NAND2_X1 U12158 ( .A1(n14893), .A2(n14871), .ZN(n9768) );
  NAND2_X1 U12159 ( .A1(n9769), .A2(n14880), .ZN(n9770) );
  OAI211_X1 U12160 ( .C1(n9772), .C2(n9771), .A(n10028), .B(n14896), .ZN(n9773) );
  INV_X1 U12161 ( .A(n9773), .ZN(n9774) );
  AOI211_X1 U12162 ( .C1(n14878), .C2(n14918), .A(n9775), .B(n9774), .ZN(
        n14920) );
  MUX2_X1 U12163 ( .A(n9776), .B(n14920), .S(n14228), .Z(n9779) );
  AOI22_X1 U12164 ( .A1(n14231), .A2(n14917), .B1(n14884), .B2(n9777), .ZN(
        n9778) );
  OAI211_X1 U12165 ( .C1(n9780), .C2(n14904), .A(n9779), .B(n9778), .ZN(
        P3_U3230) );
  NAND2_X1 U12166 ( .A1(n14414), .A2(n9725), .ZN(n9789) );
  OR2_X1 U12167 ( .A1(n9977), .A2(n9784), .ZN(n9787) );
  OR2_X1 U12168 ( .A1(n13574), .A2(n9785), .ZN(n9786) );
  NAND2_X1 U12169 ( .A1(n14468), .A2(n13311), .ZN(n9788) );
  NAND2_X1 U12170 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  XNOR2_X1 U12171 ( .A(n9790), .B(n7528), .ZN(n9911) );
  AND2_X1 U12172 ( .A1(n14468), .A2(n9725), .ZN(n9791) );
  AOI21_X1 U12173 ( .B1(n14414), .B2(n13313), .A(n9791), .ZN(n9910) );
  XNOR2_X1 U12174 ( .A(n9911), .B(n9910), .ZN(n9792) );
  XNOR2_X1 U12175 ( .A(n9909), .B(n9792), .ZN(n9803) );
  NAND2_X1 U12176 ( .A1(n9793), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9923) );
  OR2_X1 U12177 ( .A1(n9793), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9794) );
  AND2_X1 U12178 ( .A1(n9923), .A2(n9794), .ZN(n14401) );
  NAND2_X1 U12179 ( .A1(n11208), .A2(n14401), .ZN(n9799) );
  INV_X2 U12180 ( .A(n11138), .ZN(n13580) );
  NAND2_X1 U12181 ( .A1(n13580), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U12182 ( .A1(n8606), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U12183 ( .A1(n11209), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9796) );
  NAND4_X1 U12184 ( .A1(n9799), .A2(n9798), .A3(n9797), .A4(n9796), .ZN(n13665) );
  AOI22_X1 U12185 ( .A1(n13666), .A2(n14416), .B1(n14413), .B2(n13665), .ZN(
        n9815) );
  NAND2_X1 U12186 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13687) );
  INV_X1 U12187 ( .A(n14376), .ZN(n13403) );
  NAND2_X1 U12188 ( .A1(n13403), .A2(n9807), .ZN(n9800) );
  OAI211_X1 U12189 ( .C1(n9815), .C2(n13332), .A(n13687), .B(n9800), .ZN(n9801) );
  AOI21_X1 U12190 ( .B1(n14300), .B2(n14468), .A(n9801), .ZN(n9802) );
  OAI21_X1 U12191 ( .B1(n9803), .B2(n13425), .A(n9802), .ZN(P1_U3227) );
  INV_X1 U12192 ( .A(n14468), .ZN(n9973) );
  INV_X1 U12193 ( .A(n13611), .ZN(n9985) );
  XNOR2_X1 U12194 ( .A(n9985), .B(n9975), .ZN(n14470) );
  INV_X1 U12195 ( .A(n9805), .ZN(n9806) );
  AOI211_X1 U12196 ( .C1(n14468), .C2(n14428), .A(n14076), .B(n14405), .ZN(
        n14467) );
  INV_X1 U12197 ( .A(n9807), .ZN(n9808) );
  OAI22_X1 U12198 ( .A1(n14422), .A2(n9973), .B1(n9808), .B2(n14421), .ZN(
        n9809) );
  AOI21_X1 U12199 ( .B1(n14467), .B2(n14432), .A(n9809), .ZN(n9820) );
  NAND2_X1 U12200 ( .A1(n9810), .A2(n14363), .ZN(n9811) );
  NAND2_X1 U12201 ( .A1(n13666), .A2(n14461), .ZN(n9813) );
  NAND2_X1 U12202 ( .A1(n13454), .A2(n13608), .ZN(n9814) );
  XNOR2_X1 U12203 ( .A(n9986), .B(n13611), .ZN(n9816) );
  OAI21_X1 U12204 ( .B1(n9816), .B2(n14501), .A(n9815), .ZN(n14466) );
  INV_X1 U12205 ( .A(n14466), .ZN(n9817) );
  MUX2_X1 U12206 ( .A(n9818), .B(n9817), .S(n14419), .Z(n9819) );
  OAI211_X1 U12207 ( .C1(n14470), .C2(n14025), .A(n9820), .B(n9819), .ZN(
        P1_U3288) );
  INV_X1 U12208 ( .A(n11078), .ZN(n9834) );
  NAND2_X1 U12209 ( .A1(n9821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9822) );
  MUX2_X1 U12210 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9822), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9823) );
  INV_X1 U12211 ( .A(n13752), .ZN(n13748) );
  OAI222_X1 U12212 ( .A1(n14165), .A2(n9834), .B1(n13748), .B2(P1_U3086), .C1(
        n9824), .C2(n14166), .ZN(P1_U3338) );
  INV_X1 U12213 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U12214 ( .A1(n10011), .A2(n10010), .ZN(n10022) );
  NAND2_X1 U12215 ( .A1(n10373), .A2(n10372), .ZN(n10613) );
  NAND2_X1 U12216 ( .A1(n10953), .A2(n10952), .ZN(n11278) );
  NOR2_X2 U12217 ( .A1(n11292), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n11312) );
  AND2_X2 U12218 ( .A1(n11312), .A2(n11933), .ZN(n11322) );
  AND2_X2 U12219 ( .A1(n11322), .A2(n13126), .ZN(n11341) );
  NAND2_X1 U12220 ( .A1(n11340), .A2(n11341), .ZN(n11353) );
  NOR2_X2 U12221 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n11353), .ZN(n11365) );
  INV_X1 U12222 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U12223 ( .A1(n11365), .A2(n11960), .ZN(n11376) );
  OR2_X2 U12224 ( .A1(n11376), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n11387) );
  NOR2_X2 U12225 ( .A1(n11387), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11398) );
  INV_X1 U12226 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n11875) );
  AND2_X2 U12227 ( .A1(n11398), .A2(n11875), .ZN(n11411) );
  NAND2_X1 U12228 ( .A1(n11411), .A2(n11952), .ZN(n11422) );
  OR2_X2 U12229 ( .A1(n11422), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n11435) );
  NOR2_X2 U12230 ( .A1(n11435), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11437) );
  INV_X1 U12231 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U12232 ( .A1(n11437), .A2(n9826), .ZN(n11254) );
  INV_X1 U12233 ( .A(n11254), .ZN(n9827) );
  INV_X1 U12234 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U12235 ( .A1(n9827), .A2(n11895), .ZN(n12116) );
  NAND2_X1 U12236 ( .A1(n6804), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9832) );
  INV_X1 U12237 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12319) );
  OR2_X1 U12238 ( .A1(n9828), .A2(n12319), .ZN(n9831) );
  INV_X1 U12239 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9829) );
  OR2_X1 U12240 ( .A1(n11468), .A2(n9829), .ZN(n9830) );
  NAND4_X1 U12241 ( .A1(n11472), .A2(n9832), .A3(n9831), .A4(n9830), .ZN(
        n11897) );
  NAND2_X1 U12242 ( .A1(n11897), .A2(P3_U3897), .ZN(n9833) );
  OAI21_X1 U12243 ( .B1(P3_U3897), .B2(n13128), .A(n9833), .ZN(P3_U3520) );
  INV_X1 U12244 ( .A(n12670), .ZN(n10450) );
  OAI222_X1 U12245 ( .A1(n13010), .A2(n9835), .B1(n10648), .B2(n9834), .C1(
        P2_U3088), .C2(n10450), .ZN(P2_U3310) );
  OAI21_X1 U12246 ( .B1(n9837), .B2(n10362), .A(n9836), .ZN(n9953) );
  MUX2_X1 U12247 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12069), .Z(n9843) );
  OR2_X1 U12248 ( .A1(n9838), .A2(n11301), .ZN(n9840) );
  MUX2_X1 U12249 ( .A(n9840), .B(P3_IR_REG_31__SCAN_IN), .S(n9839), .Z(n9842)
         );
  NAND2_X1 U12250 ( .A1(n9842), .A2(n9841), .ZN(n14185) );
  NAND2_X1 U12251 ( .A1(n9843), .A2(n14185), .ZN(n9952) );
  NAND2_X1 U12252 ( .A1(n6637), .A2(n9952), .ZN(n9844) );
  XNOR2_X1 U12253 ( .A(n9953), .B(n9844), .ZN(n9857) );
  INV_X1 U12254 ( .A(n14185), .ZN(n10602) );
  XNOR2_X1 U12255 ( .A(n10602), .B(n9954), .ZN(n9846) );
  NAND2_X1 U12256 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n9846), .ZN(n9955) );
  OAI21_X1 U12257 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n9846), .A(n9955), .ZN(
        n9855) );
  NAND2_X1 U12258 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n9850), .ZN(n9961) );
  OAI21_X1 U12259 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n9850), .A(n9961), .ZN(
        n9851) );
  NAND2_X1 U12260 ( .A1(n9851), .A2(n14801), .ZN(n9853) );
  AND2_X1 U12261 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n10620) );
  AOI21_X1 U12262 ( .B1(n14780), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10620), .ZN(
        n9852) );
  OAI211_X1 U12263 ( .C1(n14797), .C2(n14185), .A(n9853), .B(n9852), .ZN(n9854) );
  AOI21_X1 U12264 ( .B1(n14788), .B2(n9855), .A(n9854), .ZN(n9856) );
  OAI21_X1 U12265 ( .B1(n9857), .B2(n12113), .A(n9856), .ZN(P3_U3191) );
  INV_X1 U12266 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11785) );
  INV_X1 U12267 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U12268 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11785), .B2(n9861), .ZN(n10121) );
  XNOR2_X1 U12269 ( .A(n10122), .B(n10121), .ZN(n11382) );
  INV_X1 U12270 ( .A(n11382), .ZN(n9863) );
  INV_X1 U12271 ( .A(n12423), .ZN(n14205) );
  OAI22_X1 U12272 ( .A1(n11804), .A2(P3_U3151), .B1(SI_22_), .B2(n14186), .ZN(
        n9862) );
  AOI21_X1 U12273 ( .B1(n9863), .B2(n14205), .A(n9862), .ZN(P3_U3273) );
  INV_X1 U12274 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n13223) );
  NOR2_X1 U12275 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13223), .ZN(n9864) );
  AOI21_X1 U12276 ( .B1(n13746), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9864), .ZN(
        n9865) );
  INV_X1 U12277 ( .A(n9865), .ZN(n9871) );
  OAI21_X1 U12278 ( .B1(n10791), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9866), .ZN(
        n9869) );
  INV_X1 U12279 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9867) );
  MUX2_X1 U12280 ( .A(n9867), .B(P1_REG1_REG_13__SCAN_IN), .S(n10855), .Z(
        n9868) );
  NOR2_X1 U12281 ( .A1(n9869), .A2(n9868), .ZN(n9943) );
  AOI211_X1 U12282 ( .C1(n9869), .C2(n9868), .A(n9943), .B(n13737), .ZN(n9870)
         );
  AOI211_X1 U12283 ( .C1(n14383), .C2(n10855), .A(n9871), .B(n9870), .ZN(n9879) );
  NOR2_X1 U12284 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n10791), .ZN(n9873) );
  NOR2_X1 U12285 ( .A1(n9873), .A2(n9872), .ZN(n9877) );
  INV_X1 U12286 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U12287 ( .A(n9874), .B(P1_REG2_REG_13__SCAN_IN), .S(n10855), .Z(
        n9875) );
  INV_X1 U12288 ( .A(n9875), .ZN(n9876) );
  NAND2_X1 U12289 ( .A1(n9876), .A2(n9877), .ZN(n9937) );
  OAI211_X1 U12290 ( .C1(n9877), .C2(n9876), .A(n14387), .B(n9937), .ZN(n9878)
         );
  NAND2_X1 U12291 ( .A1(n9879), .A2(n9878), .ZN(P1_U3256) );
  INV_X1 U12292 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U12293 ( .A1(n11465), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9886) );
  INV_X1 U12294 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9880) );
  OR2_X1 U12295 ( .A1(n11466), .A2(n9880), .ZN(n9885) );
  INV_X1 U12296 ( .A(n11437), .ZN(n9881) );
  NAND2_X1 U12297 ( .A1(n9881), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9882) );
  AND2_X1 U12298 ( .A1(n11254), .A2(n9882), .ZN(n11859) );
  OR2_X1 U12299 ( .A1(n9825), .A2(n11859), .ZN(n9884) );
  INV_X1 U12300 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n11706) );
  OR2_X1 U12301 ( .A1(n11468), .A2(n11706), .ZN(n9883) );
  NAND2_X1 U12302 ( .A1(n11998), .A2(P3_U3897), .ZN(n9887) );
  OAI21_X1 U12303 ( .B1(P3_U3897), .B2(n13246), .A(n9887), .ZN(P3_U3518) );
  INV_X1 U12304 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9897) );
  XNOR2_X1 U12305 ( .A(n9888), .B(n9889), .ZN(n10316) );
  XNOR2_X1 U12306 ( .A(n9890), .B(n9889), .ZN(n9892) );
  NAND2_X1 U12307 ( .A1(n12880), .A2(n12578), .ZN(n9891) );
  OAI21_X1 U12308 ( .B1(n10040), .B2(n12773), .A(n9891), .ZN(n10044) );
  AOI21_X1 U12309 ( .B1(n9892), .B2(n12879), .A(n10044), .ZN(n10321) );
  INV_X1 U12310 ( .A(n9893), .ZN(n10746) );
  AOI211_X1 U12311 ( .C1(n9894), .C2(n10746), .A(n12865), .B(n10766), .ZN(
        n10319) );
  AOI21_X1 U12312 ( .B1(n14738), .B2(n9894), .A(n10319), .ZN(n9895) );
  OAI211_X1 U12313 ( .C1(n10316), .C2(n14720), .A(n10321), .B(n9895), .ZN(
        n12976) );
  NAND2_X1 U12314 ( .A1(n12976), .A2(n14764), .ZN(n9896) );
  OAI21_X1 U12315 ( .B1(n14764), .B2(n9897), .A(n9896), .ZN(P2_U3463) );
  AOI22_X1 U12316 ( .A1(n12545), .A2(n12579), .B1(n12558), .B2(n10742), .ZN(
        n9899) );
  OAI211_X1 U12317 ( .C1(n10738), .C2(n12565), .A(n9899), .B(n9898), .ZN(n9907) );
  XNOR2_X1 U12318 ( .A(n10750), .B(n11762), .ZN(n10041) );
  AND2_X1 U12319 ( .A1(n6488), .A2(n12580), .ZN(n9900) );
  NAND2_X1 U12320 ( .A1(n10041), .A2(n9900), .ZN(n10043) );
  OAI21_X1 U12321 ( .B1(n10041), .B2(n9900), .A(n10043), .ZN(n9905) );
  AOI211_X1 U12322 ( .C1(n9905), .C2(n9904), .A(n12571), .B(n6628), .ZN(n9906)
         );
  AOI211_X1 U12323 ( .C1(n10750), .C2(n12569), .A(n9907), .B(n9906), .ZN(n9908) );
  INV_X1 U12324 ( .A(n9908), .ZN(P2_U3189) );
  INV_X1 U12325 ( .A(n9911), .ZN(n9914) );
  INV_X1 U12326 ( .A(n9910), .ZN(n9913) );
  AOI21_X2 U12327 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n10112) );
  OR2_X1 U12328 ( .A1(n9915), .A2(n9977), .ZN(n9918) );
  NAND2_X1 U12329 ( .A1(n11102), .A2(n9916), .ZN(n9917) );
  AOI22_X1 U12330 ( .A1(n13665), .A2(n9725), .B1(n13311), .B2(n13464), .ZN(
        n9920) );
  XNOR2_X1 U12331 ( .A(n9920), .B(n13022), .ZN(n10109) );
  AND2_X1 U12332 ( .A1(n13464), .A2(n9725), .ZN(n9921) );
  AOI21_X1 U12333 ( .B1(n13665), .B2(n13313), .A(n9921), .ZN(n10110) );
  XNOR2_X1 U12334 ( .A(n10109), .B(n10110), .ZN(n10111) );
  XNOR2_X1 U12335 ( .A(n10112), .B(n10111), .ZN(n9936) );
  NAND2_X1 U12336 ( .A1(n14414), .A2(n14416), .ZN(n9930) );
  NAND2_X1 U12337 ( .A1(n13580), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9928) );
  INV_X1 U12338 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12339 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  AND2_X1 U12340 ( .A1(n9992), .A2(n9924), .ZN(n10114) );
  NAND2_X1 U12341 ( .A1(n11208), .A2(n10114), .ZN(n9927) );
  NAND2_X1 U12342 ( .A1(n8606), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12343 ( .A1(n11209), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9925) );
  NAND4_X1 U12344 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n13664) );
  NAND2_X1 U12345 ( .A1(n13664), .A2(n14413), .ZN(n9929) );
  NAND2_X1 U12346 ( .A1(n9930), .A2(n9929), .ZN(n14398) );
  INV_X1 U12347 ( .A(n14401), .ZN(n9932) );
  OAI22_X1 U12348 ( .A1(n14376), .A2(n9932), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9931), .ZN(n9934) );
  INV_X1 U12349 ( .A(n14300), .ZN(n13393) );
  NOR2_X1 U12350 ( .A1(n13393), .A2(n14475), .ZN(n9933) );
  AOI211_X1 U12351 ( .C1(n14373), .C2(n14398), .A(n9934), .B(n9933), .ZN(n9935) );
  OAI21_X1 U12352 ( .B1(n9936), .B2(n13425), .A(n9935), .ZN(P1_U3239) );
  NAND2_X1 U12353 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10855), .ZN(n9938) );
  NAND2_X1 U12354 ( .A1(n9938), .A2(n9937), .ZN(n9941) );
  INV_X1 U12355 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9939) );
  MUX2_X1 U12356 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9939), .S(n10970), .Z(
        n9940) );
  NAND2_X1 U12357 ( .A1(n9940), .A2(n9941), .ZN(n10635) );
  OAI211_X1 U12358 ( .C1(n9941), .C2(n9940), .A(n14387), .B(n10635), .ZN(n9951) );
  INV_X1 U12359 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U12360 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9942), .S(n10970), .Z(
        n9945) );
  OAI21_X1 U12361 ( .B1(n9945), .B2(n9944), .A(n10627), .ZN(n9949) );
  NAND2_X1 U12362 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14294)
         );
  INV_X1 U12363 ( .A(n14294), .ZN(n9946) );
  AOI21_X1 U12364 ( .B1(n13746), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9946), .ZN(
        n9947) );
  OAI21_X1 U12365 ( .B1(n10636), .B2(n13772), .A(n9947), .ZN(n9948) );
  AOI21_X1 U12366 ( .B1(n9949), .B2(n14386), .A(n9948), .ZN(n9950) );
  NAND2_X1 U12367 ( .A1(n9951), .A2(n9950), .ZN(P1_U3257) );
  MUX2_X1 U12368 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12069), .Z(n10092) );
  XNOR2_X1 U12369 ( .A(n10092), .B(n10098), .ZN(n10093) );
  XOR2_X1 U12370 ( .A(n10093), .B(n10094), .Z(n9972) );
  INV_X1 U12371 ( .A(n10098), .ZN(n10817) );
  INV_X1 U12372 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U12373 ( .A1(n10817), .A2(n14966), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n10098), .ZN(n9958) );
  NAND2_X1 U12374 ( .A1(n14185), .A2(n9954), .ZN(n9956) );
  NAND2_X1 U12375 ( .A1(n9956), .A2(n9955), .ZN(n9957) );
  OAI21_X1 U12376 ( .B1(n9958), .B2(n9957), .A(n10095), .ZN(n9970) );
  INV_X1 U12377 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U12378 ( .A1(n10817), .A2(n9959), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n10098), .ZN(n9964) );
  NAND2_X1 U12379 ( .A1(n14185), .A2(n9960), .ZN(n9962) );
  OAI21_X1 U12380 ( .B1(n9964), .B2(n9963), .A(n10099), .ZN(n9965) );
  NAND2_X1 U12381 ( .A1(n9965), .A2(n14801), .ZN(n9968) );
  INV_X1 U12382 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U12383 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9966), .ZN(n10831) );
  AOI21_X1 U12384 ( .B1(n14780), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n10831), 
        .ZN(n9967) );
  OAI211_X1 U12385 ( .C1(n14797), .C2(n10098), .A(n9968), .B(n9967), .ZN(n9969) );
  AOI21_X1 U12386 ( .B1(n14788), .B2(n9970), .A(n9969), .ZN(n9971) );
  OAI21_X1 U12387 ( .B1(n9972), .B2(n12113), .A(n9971), .ZN(P3_U3192) );
  INV_X1 U12388 ( .A(n14414), .ZN(n9987) );
  AND2_X1 U12389 ( .A1(n9987), .A2(n9973), .ZN(n9974) );
  OR2_X1 U12390 ( .A1(n13665), .A2(n13464), .ZN(n9976) );
  NAND2_X1 U12391 ( .A1(n9978), .A2(n13595), .ZN(n9981) );
  AOI22_X1 U12392 ( .A1(n13594), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11102), 
        .B2(n9979), .ZN(n9980) );
  NAND2_X1 U12393 ( .A1(n9981), .A2(n9980), .ZN(n14484) );
  XNOR2_X1 U12394 ( .A(n13664), .B(n14484), .ZN(n13613) );
  XNOR2_X1 U12395 ( .A(n10194), .B(n13613), .ZN(n14486) );
  INV_X1 U12396 ( .A(n9982), .ZN(n14404) );
  NAND2_X1 U12397 ( .A1(n9982), .A2(n10192), .ZN(n10195) );
  INV_X1 U12398 ( .A(n10195), .ZN(n10196) );
  AOI211_X1 U12399 ( .C1(n14484), .C2(n14404), .A(n14076), .B(n10196), .ZN(
        n14483) );
  INV_X1 U12400 ( .A(n10114), .ZN(n9983) );
  OAI22_X1 U12401 ( .A1(n14422), .A2(n10192), .B1(n9983), .B2(n14421), .ZN(
        n9984) );
  AOI21_X1 U12402 ( .B1(n14483), .B2(n14432), .A(n9984), .ZN(n10002) );
  NAND2_X1 U12403 ( .A1(n9987), .A2(n14468), .ZN(n9988) );
  INV_X1 U12404 ( .A(n13665), .ZN(n9989) );
  NAND2_X1 U12405 ( .A1(n9989), .A2(n13464), .ZN(n9990) );
  INV_X1 U12406 ( .A(n13613), .ZN(n10193) );
  XNOR2_X1 U12407 ( .A(n10184), .B(n10193), .ZN(n9998) );
  NAND2_X1 U12408 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  AND2_X1 U12409 ( .A1(n10179), .A2(n9993), .ZN(n10357) );
  NAND2_X1 U12410 ( .A1(n11208), .A2(n10357), .ZN(n9997) );
  NAND2_X1 U12411 ( .A1(n13580), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U12412 ( .A1(n8606), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U12413 ( .A1(n11209), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9994) );
  NAND4_X1 U12414 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n13663) );
  AOI22_X1 U12415 ( .A1(n14416), .A2(n13665), .B1(n13663), .B2(n14413), .ZN(
        n10117) );
  OAI21_X1 U12416 ( .B1(n9998), .B2(n14501), .A(n10117), .ZN(n14482) );
  INV_X1 U12417 ( .A(n14482), .ZN(n9999) );
  MUX2_X1 U12418 ( .A(n10000), .B(n9999), .S(n14419), .Z(n10001) );
  OAI211_X1 U12419 ( .C1(n14486), .C2(n14025), .A(n10002), .B(n10001), .ZN(
        P1_U3286) );
  NAND2_X1 U12420 ( .A1(n14848), .A2(n14847), .ZN(n10008) );
  OR2_X1 U12421 ( .A1(n11454), .A2(SI_4_), .ZN(n10006) );
  OR2_X1 U12422 ( .A1(n11348), .A2(n10004), .ZN(n10005) );
  NAND2_X1 U12423 ( .A1(n10131), .A2(n10146), .ZN(n11520) );
  INV_X1 U12424 ( .A(n10146), .ZN(n14858) );
  INV_X1 U12425 ( .A(n14852), .ZN(n11518) );
  NAND2_X1 U12426 ( .A1(n11465), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10016) );
  INV_X1 U12427 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10009) );
  OR2_X1 U12428 ( .A1(n11466), .A2(n10009), .ZN(n10015) );
  OR2_X1 U12429 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  AND2_X1 U12430 ( .A1(n10022), .A2(n10012), .ZN(n10132) );
  OR2_X1 U12431 ( .A1(n11400), .A2(n10132), .ZN(n10014) );
  OR2_X1 U12432 ( .A1(n11468), .A2(n10035), .ZN(n10013) );
  AND4_X2 U12433 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n14833) );
  NAND2_X1 U12434 ( .A1(n11464), .A2(n10017), .ZN(n10021) );
  OR2_X1 U12435 ( .A1(n11454), .A2(SI_5_), .ZN(n10020) );
  OR2_X1 U12436 ( .A1(n11348), .A2(n10018), .ZN(n10019) );
  NAND2_X1 U12437 ( .A1(n14833), .A2(n10135), .ZN(n11524) );
  INV_X1 U12438 ( .A(n10135), .ZN(n10149) );
  NAND2_X1 U12439 ( .A1(n14854), .A2(n10149), .ZN(n11528) );
  XNOR2_X1 U12440 ( .A(n10160), .B(n11623), .ZN(n14927) );
  INV_X1 U12441 ( .A(n14927), .ZN(n10039) );
  NAND2_X1 U12442 ( .A1(n11465), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12443 ( .A1(n10022), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10023) );
  AND2_X1 U12444 ( .A1(n10070), .A2(n10023), .ZN(n14842) );
  OR2_X1 U12445 ( .A1(n11400), .A2(n14842), .ZN(n10025) );
  OR2_X1 U12446 ( .A1(n11468), .A2(n14845), .ZN(n10024) );
  INV_X1 U12447 ( .A(n12028), .ZN(n10236) );
  OAI22_X1 U12448 ( .A1(n10236), .A2(n14867), .B1(n10131), .B2(n14869), .ZN(
        n10034) );
  NAND2_X1 U12449 ( .A1(n14851), .A2(n14852), .ZN(n10030) );
  NAND2_X1 U12450 ( .A1(n12029), .A2(n10146), .ZN(n10029) );
  NAND2_X1 U12451 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NAND2_X1 U12452 ( .A1(n10031), .A2(n11623), .ZN(n10032) );
  AOI21_X1 U12453 ( .B1(n10151), .B2(n10032), .A(n14873), .ZN(n10033) );
  AOI211_X1 U12454 ( .C1(n14927), .C2(n14878), .A(n10034), .B(n10033), .ZN(
        n14924) );
  MUX2_X1 U12455 ( .A(n10035), .B(n14924), .S(n14228), .Z(n10038) );
  AND2_X1 U12456 ( .A1(n10135), .A2(n14916), .ZN(n14926) );
  INV_X1 U12457 ( .A(n10132), .ZN(n10036) );
  AOI22_X1 U12458 ( .A1(n14861), .A2(n14926), .B1(n14884), .B2(n10036), .ZN(
        n10037) );
  OAI211_X1 U12459 ( .C1(n10039), .C2(n14904), .A(n10038), .B(n10037), .ZN(
        P3_U3228) );
  NOR2_X1 U12460 ( .A1(n12476), .A2(n10040), .ZN(n10042) );
  AOI22_X1 U12461 ( .A1(n6628), .A2(n12533), .B1(n10042), .B2(n10041), .ZN(
        n10051) );
  NAND2_X1 U12462 ( .A1(n6488), .A2(n12579), .ZN(n10081) );
  NOR2_X1 U12463 ( .A1(n10315), .A2(n12516), .ZN(n10048) );
  INV_X1 U12464 ( .A(n10313), .ZN(n10046) );
  NAND2_X1 U12465 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12655)
         );
  NAND2_X1 U12466 ( .A1(n12444), .A2(n10044), .ZN(n10045) );
  OAI211_X1 U12467 ( .C1(n12538), .C2(n10046), .A(n12655), .B(n10045), .ZN(
        n10047) );
  AOI211_X1 U12468 ( .C1(n10086), .C2(n12533), .A(n10048), .B(n10047), .ZN(
        n10049) );
  OAI21_X1 U12469 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(P2_U3208) );
  INV_X1 U12470 ( .A(n10052), .ZN(n10053) );
  NAND2_X1 U12471 ( .A1(n10053), .A2(n14853), .ZN(n10054) );
  NAND2_X1 U12472 ( .A1(n10055), .A2(n10054), .ZN(n10140) );
  XNOR2_X1 U12473 ( .A(n10146), .B(n6828), .ZN(n10056) );
  XNOR2_X1 U12474 ( .A(n10056), .B(n10131), .ZN(n10141) );
  NAND2_X1 U12475 ( .A1(n10056), .A2(n10131), .ZN(n10057) );
  XNOR2_X1 U12476 ( .A(n10135), .B(n11892), .ZN(n10058) );
  XNOR2_X1 U12477 ( .A(n10058), .B(n14833), .ZN(n10127) );
  INV_X1 U12478 ( .A(n10058), .ZN(n10059) );
  NAND2_X1 U12479 ( .A1(n10059), .A2(n14833), .ZN(n10060) );
  NAND2_X1 U12480 ( .A1(n11464), .A2(n10061), .ZN(n10065) );
  OR2_X1 U12481 ( .A1(n10155), .A2(n10062), .ZN(n10064) );
  OR2_X1 U12482 ( .A1(n11348), .A2(n14796), .ZN(n10063) );
  XNOR2_X1 U12483 ( .A(n14841), .B(n11844), .ZN(n10231) );
  XNOR2_X1 U12484 ( .A(n10231), .B(n12028), .ZN(n10066) );
  AOI21_X1 U12485 ( .B1(n10067), .B2(n10066), .A(n12019), .ZN(n10068) );
  NAND2_X1 U12486 ( .A1(n10068), .A2(n10232), .ZN(n10080) );
  INV_X1 U12487 ( .A(n14841), .ZN(n10152) );
  NAND2_X1 U12488 ( .A1(n11433), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10076) );
  INV_X1 U12489 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n10069) );
  OR2_X1 U12490 ( .A1(n11466), .A2(n10069), .ZN(n10075) );
  AND2_X1 U12491 ( .A1(n10070), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10071) );
  NOR2_X1 U12492 ( .A1(n10164), .A2(n10071), .ZN(n10240) );
  OR2_X1 U12493 ( .A1(n9825), .A2(n10240), .ZN(n10074) );
  OR2_X1 U12494 ( .A1(n11468), .A2(n10072), .ZN(n10073) );
  NAND2_X1 U12495 ( .A1(n14854), .A2(n11999), .ZN(n10077) );
  NAND2_X1 U12496 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14802) );
  OAI211_X1 U12497 ( .C1(n14832), .C2(n11988), .A(n10077), .B(n14802), .ZN(
        n10078) );
  AOI21_X1 U12498 ( .B1(n10152), .B2(n12017), .A(n10078), .ZN(n10079) );
  OAI211_X1 U12499 ( .C1(n14842), .C2(n12015), .A(n10080), .B(n10079), .ZN(
        P3_U3179) );
  INV_X1 U12500 ( .A(n10081), .ZN(n10082) );
  XNOR2_X1 U12501 ( .A(n10768), .B(n11762), .ZN(n10243) );
  NAND2_X1 U12502 ( .A1(n6488), .A2(n12578), .ZN(n10241) );
  XNOR2_X1 U12503 ( .A(n10243), .B(n10241), .ZN(n10084) );
  AOI22_X1 U12504 ( .A1(n12492), .A2(n12579), .B1(n12558), .B2(n10767), .ZN(
        n10083) );
  NAND2_X1 U12505 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14588)
         );
  OAI211_X1 U12506 ( .C1(n10759), .C2(n12561), .A(n10083), .B(n14588), .ZN(
        n10088) );
  AOI22_X1 U12507 ( .A1(n6525), .A2(n12533), .B1(n12563), .B2(n12579), .ZN(
        n10085) );
  NOR3_X1 U12508 ( .A1(n10086), .A2(n10085), .A3(n10084), .ZN(n10087) );
  AOI211_X1 U12509 ( .C1(n10768), .C2(n12569), .A(n10088), .B(n10087), .ZN(
        n10089) );
  OAI21_X1 U12510 ( .B1(n10242), .B2(n12571), .A(n10089), .ZN(P2_U3196) );
  INV_X1 U12511 ( .A(n11090), .ZN(n10125) );
  NAND2_X1 U12512 ( .A1(n10090), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U12513 ( .A(n10091), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13767) );
  INV_X1 U12514 ( .A(n13767), .ZN(n13760) );
  OAI222_X1 U12515 ( .A1(n14165), .A2(n10125), .B1(n13760), .B2(P1_U3086), 
        .C1(n7192), .C2(n14166), .ZN(P1_U3337) );
  MUX2_X1 U12516 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12069), .Z(n10204) );
  XNOR2_X1 U12517 ( .A(n10204), .B(n10922), .ZN(n10206) );
  XOR2_X1 U12518 ( .A(n10206), .B(n10207), .Z(n10108) );
  NAND2_X1 U12519 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10098), .ZN(n10096) );
  XNOR2_X1 U12520 ( .A(n10216), .B(n10922), .ZN(n10097) );
  NAND2_X1 U12521 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10097), .ZN(n10218) );
  OAI21_X1 U12522 ( .B1(n10097), .B2(P3_REG1_REG_11__SCAN_IN), .A(n10218), 
        .ZN(n10106) );
  NAND2_X1 U12523 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n10098), .ZN(n10100) );
  NAND2_X1 U12524 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n10101), .ZN(n10212) );
  OAI21_X1 U12525 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n10101), .A(n10212), 
        .ZN(n10102) );
  NAND2_X1 U12526 ( .A1(n10102), .A2(n14801), .ZN(n10104) );
  AND2_X1 U12527 ( .A1(n6473), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11002) );
  AOI21_X1 U12528 ( .B1(n14780), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11002), 
        .ZN(n10103) );
  OAI211_X1 U12529 ( .C1(n14797), .C2(n10217), .A(n10104), .B(n10103), .ZN(
        n10105) );
  AOI21_X1 U12530 ( .B1(n14788), .B2(n10106), .A(n10105), .ZN(n10107) );
  OAI21_X1 U12531 ( .B1(n10108), .B2(n12113), .A(n10107), .ZN(P3_U3193) );
  AOI22_X1 U12532 ( .A1(n13664), .A2(n13313), .B1(n9725), .B2(n14484), .ZN(
        n10348) );
  AOI22_X1 U12533 ( .A1(n13664), .A2(n9725), .B1(n13311), .B2(n14484), .ZN(
        n10113) );
  XNOR2_X1 U12534 ( .A(n10113), .B(n13022), .ZN(n10349) );
  XOR2_X1 U12535 ( .A(n10348), .B(n10349), .Z(n10350) );
  XNOR2_X1 U12536 ( .A(n10351), .B(n10350), .ZN(n10120) );
  NAND2_X1 U12537 ( .A1(n13403), .A2(n10114), .ZN(n10115) );
  OAI211_X1 U12538 ( .C1(n10117), .C2(n13332), .A(n10116), .B(n10115), .ZN(
        n10118) );
  AOI21_X1 U12539 ( .B1(n14300), .B2(n14484), .A(n10118), .ZN(n10119) );
  OAI21_X1 U12540 ( .B1(n10120), .B2(n13425), .A(n10119), .ZN(P1_U3213) );
  INV_X1 U12541 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10904) );
  INV_X1 U12542 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U12543 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n10904), .B2(n11143), .ZN(n10594) );
  XNOR2_X1 U12544 ( .A(n10595), .B(n10594), .ZN(n11393) );
  NAND2_X1 U12545 ( .A1(n11393), .A2(n14205), .ZN(n10124) );
  OAI211_X1 U12546 ( .C1(n11394), .C2(n14186), .A(n10124), .B(n10123), .ZN(
        P3_U3272) );
  OAI222_X1 U12547 ( .A1(n13010), .A2(n10126), .B1(n10648), .B2(n10125), .C1(
        P2_U3088), .C2(n14660), .ZN(P2_U3309) );
  XOR2_X1 U12548 ( .A(n10128), .B(n10127), .Z(n10137) );
  AOI21_X1 U12549 ( .B1(n12013), .B2(n12028), .A(n10129), .ZN(n10130) );
  OAI21_X1 U12550 ( .B1(n10131), .B2(n12009), .A(n10130), .ZN(n10134) );
  NOR2_X1 U12551 ( .A1(n12015), .A2(n10132), .ZN(n10133) );
  AOI211_X1 U12552 ( .C1(n10135), .C2(n12017), .A(n10134), .B(n10133), .ZN(
        n10136) );
  OAI21_X1 U12553 ( .B1(n10137), .B2(n12019), .A(n10136), .ZN(P3_U3167) );
  INV_X1 U12554 ( .A(n10138), .ZN(n10139) );
  AOI21_X1 U12555 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10148) );
  NAND2_X1 U12556 ( .A1(n11999), .A2(n14853), .ZN(n10143) );
  OAI211_X1 U12557 ( .C1(n14833), .C2(n11988), .A(n10143), .B(n10142), .ZN(
        n10145) );
  NOR2_X1 U12558 ( .A1(n12015), .A2(n14859), .ZN(n10144) );
  AOI211_X1 U12559 ( .C1(n10146), .C2(n12017), .A(n10145), .B(n10144), .ZN(
        n10147) );
  OAI21_X1 U12560 ( .B1(n10148), .B2(n12019), .A(n10147), .ZN(P3_U3170) );
  NAND2_X1 U12561 ( .A1(n14833), .A2(n10149), .ZN(n10150) );
  OR2_X2 U12562 ( .A1(n12028), .A2(n14841), .ZN(n11532) );
  NAND2_X1 U12563 ( .A1(n12028), .A2(n14841), .ZN(n11530) );
  NAND2_X1 U12564 ( .A1(n14837), .A2(n14836), .ZN(n14835) );
  NAND2_X1 U12565 ( .A1(n12028), .A2(n10152), .ZN(n10153) );
  NAND2_X1 U12566 ( .A1(n14835), .A2(n10153), .ZN(n10367) );
  OR2_X1 U12567 ( .A1(n11454), .A2(SI_7_), .ZN(n10158) );
  OR2_X1 U12568 ( .A1(n11348), .A2(n10156), .ZN(n10157) );
  NAND2_X1 U12569 ( .A1(n14832), .A2(n10368), .ZN(n11533) );
  NAND2_X1 U12570 ( .A1(n11533), .A2(n11534), .ZN(n10366) );
  XNOR2_X1 U12571 ( .A(n10367), .B(n10366), .ZN(n10172) );
  INV_X1 U12572 ( .A(n14836), .ZN(n11630) );
  INV_X1 U12573 ( .A(n10366), .ZN(n11625) );
  OAI21_X1 U12574 ( .B1(n10161), .B2(n11625), .A(n10360), .ZN(n14934) );
  NAND2_X1 U12575 ( .A1(n11433), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10169) );
  INV_X1 U12576 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n10162) );
  OR2_X1 U12577 ( .A1(n11466), .A2(n10162), .ZN(n10168) );
  NOR2_X1 U12578 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  OR2_X1 U12579 ( .A1(n10373), .A2(n10165), .ZN(n10384) );
  INV_X1 U12580 ( .A(n10384), .ZN(n10466) );
  OR2_X1 U12581 ( .A1(n11400), .A2(n10466), .ZN(n10167) );
  OR2_X1 U12582 ( .A1(n11468), .A2(n9848), .ZN(n10166) );
  OAI22_X1 U12583 ( .A1(n10236), .A2(n14869), .B1(n14819), .B2(n14867), .ZN(
        n10170) );
  AOI21_X1 U12584 ( .B1(n14934), .B2(n14878), .A(n10170), .ZN(n10171) );
  OAI21_X1 U12585 ( .B1(n10172), .B2(n14873), .A(n10171), .ZN(n14932) );
  INV_X1 U12586 ( .A(n14932), .ZN(n10177) );
  INV_X1 U12587 ( .A(n14904), .ZN(n11708) );
  INV_X1 U12588 ( .A(n10240), .ZN(n10173) );
  AOI22_X1 U12589 ( .A1(n14861), .A2(n14933), .B1(n14884), .B2(n10173), .ZN(
        n10174) );
  OAI21_X1 U12590 ( .B1(n10072), .B2(n14228), .A(n10174), .ZN(n10175) );
  AOI21_X1 U12591 ( .B1(n14934), .B2(n11708), .A(n10175), .ZN(n10176) );
  OAI21_X1 U12592 ( .B1(n10177), .B2(n14908), .A(n10176), .ZN(P3_U3226) );
  NOR2_X1 U12593 ( .A1(n10400), .A2(n7524), .ZN(n10502) );
  NAND2_X1 U12594 ( .A1(n11208), .A2(n10502), .ZN(n10183) );
  NAND2_X1 U12595 ( .A1(n13580), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U12596 ( .A1(n11209), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U12597 ( .A1(n8606), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10180) );
  NAND4_X1 U12598 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n13662) );
  NAND2_X1 U12599 ( .A1(n10192), .A2(n13664), .ZN(n10185) );
  NAND2_X1 U12600 ( .A1(n10187), .A2(n13595), .ZN(n10189) );
  AOI22_X1 U12601 ( .A1(n13594), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11102), 
        .B2(n13709), .ZN(n10188) );
  XNOR2_X1 U12602 ( .A(n13472), .B(n13663), .ZN(n13614) );
  XOR2_X1 U12603 ( .A(n10392), .B(n13614), .Z(n10190) );
  AOI222_X1 U12604 ( .A1(n13664), .A2(n14416), .B1(n13662), .B2(n14413), .C1(
        n14411), .C2(n10190), .ZN(n14491) );
  INV_X1 U12605 ( .A(n14491), .ZN(n10191) );
  AOI21_X1 U12606 ( .B1(n10357), .B2(n14400), .A(n10191), .ZN(n10200) );
  INV_X1 U12607 ( .A(n13664), .ZN(n10355) );
  XNOR2_X1 U12608 ( .A(n10397), .B(n13614), .ZN(n14494) );
  INV_X1 U12609 ( .A(n13472), .ZN(n14492) );
  OAI211_X1 U12610 ( .C1(n10196), .C2(n14492), .A(n14429), .B(n10399), .ZN(
        n14490) );
  AOI22_X1 U12611 ( .A1(n14033), .A2(n13472), .B1(n6479), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n10197) );
  OAI21_X1 U12612 ( .B1(n14490), .B2(n14022), .A(n10197), .ZN(n10198) );
  AOI21_X1 U12613 ( .B1(n14494), .B2(n14433), .A(n10198), .ZN(n10199) );
  OAI21_X1 U12614 ( .B1(n10200), .B2(n6479), .A(n10199), .ZN(P1_U3285) );
  INV_X1 U12615 ( .A(n11101), .ZN(n10202) );
  OAI222_X1 U12616 ( .A1(n12679), .A2(P2_U3088), .B1(n10648), .B2(n10202), 
        .C1(n10201), .C2(n13010), .ZN(P2_U3308) );
  OAI222_X1 U12617 ( .A1(n14166), .A2(n10203), .B1(n14165), .B2(n10202), .C1(
        P1_U3086), .C2(n13990), .ZN(P1_U3336) );
  INV_X1 U12618 ( .A(n10204), .ZN(n10205) );
  MUX2_X1 U12619 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12069), .Z(n10534) );
  XNOR2_X1 U12620 ( .A(n10534), .B(n10537), .ZN(n10208) );
  OAI211_X1 U12621 ( .C1(n10209), .C2(n10208), .A(n10535), .B(n14792), .ZN(
        n10230) );
  INV_X1 U12622 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U12623 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n10934), .B1(n10537), 
        .B2(n10210), .ZN(n10215) );
  NAND2_X1 U12624 ( .A1(n10217), .A2(n10211), .ZN(n10213) );
  OAI21_X1 U12625 ( .B1(n10215), .B2(n10214), .A(n10540), .ZN(n10228) );
  NAND2_X1 U12626 ( .A1(n10217), .A2(n10216), .ZN(n10219) );
  INV_X1 U12627 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n10220) );
  MUX2_X1 U12628 ( .A(n10220), .B(P3_REG1_REG_12__SCAN_IN), .S(n10537), .Z(
        n10221) );
  NAND2_X1 U12629 ( .A1(n10221), .A2(n10222), .ZN(n10546) );
  OAI21_X1 U12630 ( .B1(n10222), .B2(n10221), .A(n10546), .ZN(n10223) );
  NAND2_X1 U12631 ( .A1(n10223), .A2(n14788), .ZN(n10226) );
  INV_X1 U12632 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12633 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10224), .ZN(n11915) );
  AOI21_X1 U12634 ( .B1(n14780), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11915), 
        .ZN(n10225) );
  OAI211_X1 U12635 ( .C1(n14797), .C2(n10934), .A(n10226), .B(n10225), .ZN(
        n10227) );
  AOI21_X1 U12636 ( .B1(n14801), .B2(n10228), .A(n10227), .ZN(n10229) );
  NAND2_X1 U12637 ( .A1(n10230), .A2(n10229), .ZN(P3_U3194) );
  XNOR2_X1 U12638 ( .A(n10366), .B(n11892), .ZN(n10454) );
  OAI211_X1 U12639 ( .C1(n10233), .C2(n10454), .A(n10457), .B(n11984), .ZN(
        n10239) );
  INV_X1 U12640 ( .A(n14819), .ZN(n12026) );
  AOI21_X1 U12641 ( .B1(n12026), .B2(n12013), .A(n10234), .ZN(n10235) );
  OAI21_X1 U12642 ( .B1(n10236), .B2(n12009), .A(n10235), .ZN(n10237) );
  AOI21_X1 U12643 ( .B1(n10368), .B2(n12017), .A(n10237), .ZN(n10238) );
  OAI211_X1 U12644 ( .C1(n10240), .C2(n12015), .A(n10239), .B(n10238), .ZN(
        P3_U3153) );
  INV_X1 U12645 ( .A(n10241), .ZN(n10244) );
  XNOR2_X1 U12646 ( .A(n14270), .B(n11743), .ZN(n10246) );
  AND2_X1 U12647 ( .A1(n6487), .A2(n8326), .ZN(n10245) );
  NAND2_X1 U12648 ( .A1(n10246), .A2(n10245), .ZN(n10248) );
  OAI21_X1 U12649 ( .B1(n10246), .B2(n10245), .A(n10248), .ZN(n10487) );
  NOR2_X1 U12650 ( .A1(n12476), .A2(n10759), .ZN(n10247) );
  AOI22_X1 U12651 ( .A1(n10485), .A2(n12533), .B1(n10247), .B2(n10246), .ZN(
        n10257) );
  XNOR2_X1 U12652 ( .A(n10687), .B(n11743), .ZN(n11717) );
  NAND2_X1 U12653 ( .A1(n6488), .A2(n12577), .ZN(n11716) );
  XNOR2_X1 U12654 ( .A(n11717), .B(n11716), .ZN(n10250) );
  INV_X1 U12655 ( .A(n10250), .ZN(n10256) );
  INV_X1 U12656 ( .A(n10248), .ZN(n10249) );
  NAND2_X1 U12657 ( .A1(n6633), .A2(n12533), .ZN(n10255) );
  NAND2_X1 U12658 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14617)
         );
  OAI21_X1 U12659 ( .B1(n12561), .B2(n11719), .A(n14617), .ZN(n10253) );
  OAI22_X1 U12660 ( .A1(n12565), .A2(n10759), .B1(n12538), .B2(n10685), .ZN(
        n10252) );
  AOI211_X1 U12661 ( .C1(n10687), .C2(n12569), .A(n10253), .B(n10252), .ZN(
        n10254) );
  OAI211_X1 U12662 ( .C1(n10257), .C2(n10256), .A(n10255), .B(n10254), .ZN(
        P2_U3187) );
  XNOR2_X1 U12663 ( .A(n10258), .B(n10259), .ZN(n14721) );
  AOI21_X1 U12664 ( .B1(n10782), .B2(n14717), .A(n12865), .ZN(n10260) );
  AND2_X1 U12665 ( .A1(n10260), .A2(n10334), .ZN(n14719) );
  NAND3_X1 U12666 ( .A1(n10778), .A2(n10262), .A3(n10261), .ZN(n10263) );
  NAND2_X1 U12667 ( .A1(n10264), .A2(n10263), .ZN(n10268) );
  OAI22_X1 U12668 ( .A1(n10266), .A2(n12777), .B1(n10265), .B2(n12773), .ZN(
        n10267) );
  AOI21_X1 U12669 ( .B1(n10268), .B2(n12879), .A(n10267), .ZN(n14724) );
  NOR2_X1 U12670 ( .A1(n14724), .A2(n12858), .ZN(n10272) );
  AOI22_X1 U12671 ( .A1(n12858), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n10269), 
        .B2(n14669), .ZN(n10270) );
  OAI21_X1 U12672 ( .B1(n14673), .B2(n6738), .A(n10270), .ZN(n10271) );
  AOI211_X1 U12673 ( .C1(n14667), .C2(n14719), .A(n10272), .B(n10271), .ZN(
        n10273) );
  OAI21_X1 U12674 ( .B1(n12893), .B2(n14721), .A(n10273), .ZN(P2_U3261) );
  OAI21_X1 U12675 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(n14744) );
  INV_X1 U12676 ( .A(n14744), .ZN(n14741) );
  XNOR2_X1 U12677 ( .A(n10278), .B(n10277), .ZN(n10280) );
  AOI21_X1 U12678 ( .B1(n10280), .B2(n12879), .A(n10279), .ZN(n14735) );
  MUX2_X1 U12679 ( .A(n8946), .B(n14735), .S(n12889), .Z(n10287) );
  INV_X1 U12680 ( .A(n10337), .ZN(n10282) );
  AOI211_X1 U12681 ( .C1(n14737), .C2(n10282), .A(n12865), .B(n10281), .ZN(
        n14736) );
  OAI22_X1 U12682 ( .A1(n14673), .A2(n10284), .B1(n12886), .B2(n10283), .ZN(
        n10285) );
  AOI21_X1 U12683 ( .B1(n14667), .B2(n14736), .A(n10285), .ZN(n10286) );
  OAI211_X1 U12684 ( .C1(n14741), .C2(n12893), .A(n10287), .B(n10286), .ZN(
        P2_U3259) );
  AOI21_X1 U12685 ( .B1(n10288), .B2(n12889), .A(n14667), .ZN(n10299) );
  NAND2_X1 U12686 ( .A1(n10289), .A2(n10477), .ZN(n14689) );
  INV_X1 U12687 ( .A(n14691), .ZN(n10291) );
  NAND2_X1 U12688 ( .A1(n6485), .A2(n12774), .ZN(n10290) );
  NAND2_X1 U12689 ( .A1(n10291), .A2(n10290), .ZN(n10293) );
  AND2_X1 U12690 ( .A1(n10293), .A2(n10292), .ZN(n14690) );
  OAI22_X1 U12691 ( .A1(n14680), .A2(n14690), .B1(n7576), .B2(n12886), .ZN(
        n10297) );
  INV_X1 U12692 ( .A(n10294), .ZN(n10295) );
  NAND2_X1 U12693 ( .A1(n12889), .A2(n10295), .ZN(n12854) );
  NOR2_X1 U12694 ( .A1(n12854), .A2(n14691), .ZN(n10296) );
  AOI211_X1 U12695 ( .C1(n14680), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10297), .B(
        n10296), .ZN(n10298) );
  OAI21_X1 U12696 ( .B1(n10299), .B2(n14689), .A(n10298), .ZN(P2_U3265) );
  XNOR2_X1 U12697 ( .A(n10300), .B(n10305), .ZN(n14705) );
  NAND2_X1 U12698 ( .A1(n8267), .A2(n10475), .ZN(n10301) );
  NAND2_X1 U12699 ( .A1(n10301), .A2(n12971), .ZN(n10302) );
  NOR2_X1 U12700 ( .A1(n10783), .A2(n10302), .ZN(n14703) );
  OAI21_X1 U12701 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(n10307) );
  AOI21_X1 U12702 ( .B1(n10307), .B2(n12879), .A(n10306), .ZN(n14701) );
  NOR2_X1 U12703 ( .A1(n12858), .A2(n14701), .ZN(n10311) );
  AOI22_X1 U12704 ( .A1(n12858), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14669), .ZN(n10308) );
  OAI21_X1 U12705 ( .B1(n14673), .B2(n10309), .A(n10308), .ZN(n10310) );
  AOI211_X1 U12706 ( .C1(n14703), .C2(n14667), .A(n10311), .B(n10310), .ZN(
        n10312) );
  OAI21_X1 U12707 ( .B1(n12893), .B2(n14705), .A(n10312), .ZN(P2_U3263) );
  AOI22_X1 U12708 ( .A1(n12858), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10313), 
        .B2(n14669), .ZN(n10314) );
  OAI21_X1 U12709 ( .B1(n14673), .B2(n10315), .A(n10314), .ZN(n10318) );
  NOR2_X1 U12710 ( .A1(n10316), .A2(n12893), .ZN(n10317) );
  AOI211_X1 U12711 ( .C1(n10319), .C2(n14667), .A(n10318), .B(n10317), .ZN(
        n10320) );
  OAI21_X1 U12712 ( .B1(n14680), .B2(n10321), .A(n10320), .ZN(P2_U3254) );
  AOI22_X1 U12713 ( .A1(n14680), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10322), 
        .B2(n14669), .ZN(n10323) );
  OAI21_X1 U12714 ( .B1(n14673), .B2(n10324), .A(n10323), .ZN(n10327) );
  NOR2_X1 U12715 ( .A1(n10325), .A2(n12858), .ZN(n10326) );
  AOI211_X1 U12716 ( .C1(n10328), .C2(n14667), .A(n10327), .B(n10326), .ZN(
        n10329) );
  OAI21_X1 U12717 ( .B1(n12893), .B2(n10330), .A(n10329), .ZN(P2_U3256) );
  XOR2_X1 U12718 ( .A(n10341), .B(n10331), .Z(n10333) );
  AOI21_X1 U12719 ( .B1(n10333), .B2(n12879), .A(n10332), .ZN(n14730) );
  NAND2_X1 U12720 ( .A1(n10334), .A2(n14727), .ZN(n10335) );
  NAND2_X1 U12721 ( .A1(n10335), .A2(n12971), .ZN(n10336) );
  NOR2_X1 U12722 ( .A1(n10337), .A2(n10336), .ZN(n14726) );
  AOI22_X1 U12723 ( .A1(n12858), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n10338), 
        .B2(n14669), .ZN(n10339) );
  OAI21_X1 U12724 ( .B1(n14673), .B2(n10340), .A(n10339), .ZN(n10345) );
  INV_X1 U12725 ( .A(n10341), .ZN(n10342) );
  XNOR2_X1 U12726 ( .A(n10343), .B(n10342), .ZN(n14729) );
  NOR2_X1 U12727 ( .A1(n12893), .A2(n14729), .ZN(n10344) );
  AOI211_X1 U12728 ( .C1(n14726), .C2(n14667), .A(n10345), .B(n10344), .ZN(
        n10346) );
  OAI21_X1 U12729 ( .B1(n14680), .B2(n14730), .A(n10346), .ZN(P2_U3260) );
  AOI22_X1 U12730 ( .A1(n13472), .A2(n9725), .B1(n13663), .B2(n13313), .ZN(
        n10491) );
  AOI22_X1 U12731 ( .A1(n13472), .A2(n13311), .B1(n13663), .B2(n9725), .ZN(
        n10347) );
  XNOR2_X1 U12732 ( .A(n10347), .B(n13022), .ZN(n10492) );
  XOR2_X1 U12733 ( .A(n10491), .B(n10492), .Z(n10353) );
  OAI21_X1 U12734 ( .B1(n10353), .B2(n10352), .A(n10499), .ZN(n10354) );
  NAND2_X1 U12735 ( .A1(n10354), .A2(n14366), .ZN(n10359) );
  AND2_X1 U12736 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n13704) );
  OAI22_X1 U12737 ( .A1(n10565), .A2(n13400), .B1(n10355), .B2(n13399), .ZN(
        n10356) );
  AOI211_X1 U12738 ( .C1(n10357), .C2(n13403), .A(n13704), .B(n10356), .ZN(
        n10358) );
  OAI211_X1 U12739 ( .C1(n14492), .C2(n13393), .A(n10359), .B(n10358), .ZN(
        P1_U3221) );
  OR2_X1 U12740 ( .A1(n11348), .A2(n10362), .ZN(n10363) );
  OAI211_X1 U12741 ( .C1(n11454), .C2(n10365), .A(n10364), .B(n10363), .ZN(
        n10463) );
  NAND2_X1 U12742 ( .A1(n14819), .A2(n10463), .ZN(n11539) );
  INV_X1 U12743 ( .A(n10463), .ZN(n10940) );
  NAND2_X1 U12744 ( .A1(n12026), .A2(n10940), .ZN(n11540) );
  XNOR2_X1 U12745 ( .A(n10918), .B(n6676), .ZN(n10383) );
  NAND2_X1 U12746 ( .A1(n10367), .A2(n10366), .ZN(n10370) );
  NAND2_X1 U12747 ( .A1(n12027), .A2(n10368), .ZN(n10369) );
  OAI21_X1 U12748 ( .B1(n6632), .B2(n6676), .A(n10942), .ZN(n10381) );
  NAND2_X1 U12749 ( .A1(n11465), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n10379) );
  INV_X1 U12750 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n10371) );
  OR2_X1 U12751 ( .A1(n11466), .A2(n10371), .ZN(n10378) );
  OR2_X1 U12752 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  AND2_X1 U12753 ( .A1(n10613), .A2(n10374), .ZN(n14823) );
  OR2_X1 U12754 ( .A1(n11400), .A2(n14823), .ZN(n10377) );
  INV_X1 U12755 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10375) );
  OR2_X1 U12756 ( .A1(n11468), .A2(n10375), .ZN(n10376) );
  OAI22_X1 U12757 ( .A1(n14832), .A2(n14869), .B1(n10919), .B2(n14867), .ZN(
        n10380) );
  AOI21_X1 U12758 ( .B1(n10381), .B2(n14896), .A(n10380), .ZN(n10382) );
  OAI21_X1 U12759 ( .B1(n14900), .B2(n10383), .A(n10382), .ZN(n14935) );
  INV_X1 U12760 ( .A(n14935), .ZN(n10388) );
  INV_X1 U12761 ( .A(n10383), .ZN(n14938) );
  NOR2_X1 U12762 ( .A1(n10940), .A2(n14886), .ZN(n14936) );
  AOI22_X1 U12763 ( .A1(n14861), .A2(n14936), .B1(n14884), .B2(n10384), .ZN(
        n10385) );
  OAI21_X1 U12764 ( .B1(n9848), .B2(n14228), .A(n10385), .ZN(n10386) );
  AOI21_X1 U12765 ( .B1(n14938), .B2(n11708), .A(n10386), .ZN(n10387) );
  OAI21_X1 U12766 ( .B1(n10388), .B2(n14908), .A(n10387), .ZN(P3_U3225) );
  NAND2_X1 U12767 ( .A1(n10389), .A2(n13595), .ZN(n10391) );
  AOI22_X1 U12768 ( .A1(n13594), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11102), 
        .B2(n13725), .ZN(n10390) );
  NAND2_X1 U12769 ( .A1(n10392), .A2(n13614), .ZN(n10394) );
  NAND2_X1 U12770 ( .A1(n14492), .A2(n13663), .ZN(n10393) );
  INV_X1 U12771 ( .A(n10508), .ZN(n10395) );
  AOI21_X1 U12772 ( .B1(n13617), .B2(n10396), .A(n10395), .ZN(n14502) );
  OR2_X1 U12773 ( .A1(n6479), .A2(n14501), .ZN(n13962) );
  XOR2_X1 U12774 ( .A(n10516), .B(n13617), .Z(n14504) );
  INV_X1 U12775 ( .A(n14504), .ZN(n14508) );
  NAND2_X1 U12776 ( .A1(n14508), .A2(n14433), .ZN(n10413) );
  INV_X1 U12777 ( .A(n10524), .ZN(n10398) );
  AOI211_X1 U12778 ( .C1(n14498), .C2(n10399), .A(n14076), .B(n10398), .ZN(
        n14496) );
  NAND2_X1 U12779 ( .A1(n14498), .A2(n14033), .ZN(n10410) );
  AOI22_X1 U12780 ( .A1(n6479), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10502), .B2(
        n14400), .ZN(n10409) );
  NAND2_X1 U12781 ( .A1(n13663), .A2(n14416), .ZN(n10407) );
  OR2_X1 U12782 ( .A1(n10400), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U12783 ( .A1(n10400), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10518) );
  AND2_X1 U12784 ( .A1(n10401), .A2(n10518), .ZN(n10568) );
  NAND2_X1 U12785 ( .A1(n11208), .A2(n10568), .ZN(n10405) );
  NAND2_X1 U12786 ( .A1(n13580), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U12787 ( .A1(n11209), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U12788 ( .A1(n8606), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10402) );
  NAND4_X1 U12789 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n13661) );
  NAND2_X1 U12790 ( .A1(n13661), .A2(n14413), .ZN(n10406) );
  NAND2_X1 U12791 ( .A1(n10407), .A2(n10406), .ZN(n14497) );
  NAND2_X1 U12792 ( .A1(n14497), .A2(n14419), .ZN(n10408) );
  NAND3_X1 U12793 ( .A1(n10410), .A2(n10409), .A3(n10408), .ZN(n10411) );
  AOI21_X1 U12794 ( .B1(n14496), .B2(n14432), .A(n10411), .ZN(n10412) );
  OAI211_X1 U12795 ( .C1(n14502), .C2(n13962), .A(n10413), .B(n10412), .ZN(
        P1_U3284) );
  INV_X1 U12796 ( .A(n14611), .ZN(n10443) );
  NAND2_X1 U12797 ( .A1(n10432), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10414) );
  AND2_X1 U12798 ( .A1(n10415), .A2(n10414), .ZN(n12653) );
  INV_X1 U12799 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10416) );
  MUX2_X1 U12800 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10416), .S(n10435), .Z(
        n12652) );
  NAND2_X1 U12801 ( .A1(n12653), .A2(n12652), .ZN(n12651) );
  OR2_X1 U12802 ( .A1(n10435), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10417) );
  NAND2_X1 U12803 ( .A1(n12651), .A2(n10417), .ZN(n14577) );
  INV_X1 U12804 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10418) );
  OR2_X1 U12805 ( .A1(n14586), .A2(n10418), .ZN(n10419) );
  NAND2_X1 U12806 ( .A1(n14586), .A2(n10418), .ZN(n10420) );
  AND2_X1 U12807 ( .A1(n10419), .A2(n10420), .ZN(n14578) );
  NAND2_X1 U12808 ( .A1(n14577), .A2(n14578), .ZN(n14576) );
  NAND2_X1 U12809 ( .A1(n14576), .A2(n10420), .ZN(n14592) );
  INV_X1 U12810 ( .A(n14601), .ZN(n10440) );
  INV_X1 U12811 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U12812 ( .A1(n10440), .A2(n10421), .ZN(n10423) );
  NAND2_X1 U12813 ( .A1(n14601), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10422) );
  AND2_X1 U12814 ( .A1(n10423), .A2(n10422), .ZN(n14591) );
  NAND2_X1 U12815 ( .A1(n10440), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10424) );
  NAND2_X1 U12816 ( .A1(n14593), .A2(n10424), .ZN(n10425) );
  XNOR2_X1 U12817 ( .A(n10425), .B(n14611), .ZN(n14607) );
  AND2_X1 U12818 ( .A1(n14607), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14606) );
  AOI21_X1 U12819 ( .B1(n10443), .B2(n10425), .A(n14606), .ZN(n10426) );
  NOR2_X1 U12820 ( .A1(n10426), .A2(n10445), .ZN(n10427) );
  INV_X1 U12821 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14621) );
  XNOR2_X1 U12822 ( .A(n10426), .B(n10445), .ZN(n14622) );
  NOR2_X1 U12823 ( .A1(n14621), .A2(n14622), .ZN(n14620) );
  NOR2_X1 U12824 ( .A1(n10427), .A2(n14620), .ZN(n14640) );
  NAND2_X1 U12825 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14643), .ZN(n10428) );
  OAI21_X1 U12826 ( .B1(n14643), .B2(P2_REG2_REG_16__SCAN_IN), .A(n10428), 
        .ZN(n14639) );
  NOR2_X1 U12827 ( .A1(n14640), .A2(n14639), .ZN(n14638) );
  AOI21_X1 U12828 ( .B1(n14643), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14638), 
        .ZN(n10431) );
  NAND2_X1 U12829 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n12670), .ZN(n10429) );
  OAI21_X1 U12830 ( .B1(n12670), .B2(P2_REG2_REG_17__SCAN_IN), .A(n10429), 
        .ZN(n10430) );
  NOR2_X1 U12831 ( .A1(n10431), .A2(n10430), .ZN(n12664) );
  AOI211_X1 U12832 ( .C1(n10431), .C2(n10430), .A(n12664), .B(n14637), .ZN(
        n10453) );
  INV_X1 U12833 ( .A(n10445), .ZN(n14629) );
  NAND2_X1 U12834 ( .A1(n10432), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U12835 ( .A1(n10434), .A2(n10433), .ZN(n12660) );
  INV_X1 U12836 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n13181) );
  MUX2_X1 U12837 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13181), .S(n10435), .Z(
        n12659) );
  NAND2_X1 U12838 ( .A1(n12660), .A2(n12659), .ZN(n12658) );
  NAND2_X1 U12839 ( .A1(n10435), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10436) );
  AND2_X1 U12840 ( .A1(n12658), .A2(n10436), .ZN(n14581) );
  OR2_X1 U12841 ( .A1(n14586), .A2(n14281), .ZN(n10437) );
  INV_X1 U12842 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U12843 ( .A1(n14586), .A2(n14281), .ZN(n10438) );
  AND2_X1 U12844 ( .A1(n10437), .A2(n10438), .ZN(n14582) );
  NAND2_X1 U12845 ( .A1(n14581), .A2(n14582), .ZN(n14580) );
  NAND2_X1 U12846 ( .A1(n14580), .A2(n10438), .ZN(n14596) );
  INV_X1 U12847 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10439) );
  MUX2_X1 U12848 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10439), .S(n14601), .Z(
        n14595) );
  NAND2_X1 U12849 ( .A1(n10440), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U12850 ( .A1(n14597), .A2(n10441), .ZN(n14610) );
  NAND2_X1 U12851 ( .A1(n14611), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10442) );
  OAI21_X1 U12852 ( .B1(n14611), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10442), 
        .ZN(n14609) );
  AND2_X1 U12853 ( .A1(n14610), .A2(n14609), .ZN(n14612) );
  AOI21_X1 U12854 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n10443), .A(n14612), 
        .ZN(n10444) );
  INV_X1 U12855 ( .A(n10444), .ZN(n10446) );
  XOR2_X1 U12856 ( .A(n10445), .B(n10444), .Z(n14623) );
  AND2_X1 U12857 ( .A1(n14623), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n14624) );
  AOI21_X1 U12858 ( .B1(n14629), .B2(n10446), .A(n14624), .ZN(n14636) );
  XNOR2_X1 U12859 ( .A(n14643), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14635) );
  NOR2_X1 U12860 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  AOI21_X1 U12861 ( .B1(n14643), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14634), 
        .ZN(n10448) );
  XNOR2_X1 U12862 ( .A(n12670), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10447) );
  NOR2_X1 U12863 ( .A1(n10448), .A2(n10447), .ZN(n12669) );
  AOI211_X1 U12864 ( .C1(n10448), .C2(n10447), .A(n12669), .B(n14633), .ZN(
        n10452) );
  NAND2_X1 U12865 ( .A1(n14535), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U12866 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12496)
         );
  OAI211_X1 U12867 ( .C1(n10450), .C2(n14661), .A(n10449), .B(n12496), .ZN(
        n10451) );
  OR3_X1 U12868 ( .A1(n10453), .A2(n10452), .A3(n10451), .ZN(P2_U3231) );
  INV_X1 U12869 ( .A(n10454), .ZN(n10455) );
  NAND2_X1 U12870 ( .A1(n10455), .A2(n12027), .ZN(n10456) );
  NAND2_X1 U12871 ( .A1(n10457), .A2(n10456), .ZN(n10459) );
  XNOR2_X1 U12872 ( .A(n11892), .B(n10463), .ZN(n10606) );
  XNOR2_X1 U12873 ( .A(n10606), .B(n14819), .ZN(n10458) );
  NAND2_X1 U12874 ( .A1(n10459), .A2(n10458), .ZN(n10609) );
  OAI211_X1 U12875 ( .C1(n10459), .C2(n10458), .A(n10609), .B(n11984), .ZN(
        n10465) );
  AOI21_X1 U12876 ( .B1(n14809), .B2(n12013), .A(n10460), .ZN(n10461) );
  OAI21_X1 U12877 ( .B1(n14832), .B2(n12009), .A(n10461), .ZN(n10462) );
  AOI21_X1 U12878 ( .B1(n10463), .B2(n12017), .A(n10462), .ZN(n10464) );
  OAI211_X1 U12879 ( .C1(n10466), .C2(n12015), .A(n10465), .B(n10464), .ZN(
        P3_U3161) );
  OAI21_X1 U12880 ( .B1(n8380), .B2(n10468), .A(n10467), .ZN(n10472) );
  OAI22_X1 U12881 ( .A1(n8269), .A2(n12777), .B1(n10469), .B2(n12773), .ZN(
        n10471) );
  XNOR2_X1 U12882 ( .A(n8380), .B(n12456), .ZN(n10478) );
  INV_X1 U12883 ( .A(n10478), .ZN(n14698) );
  NOR2_X1 U12884 ( .A1(n14698), .A2(n6485), .ZN(n10470) );
  AOI211_X1 U12885 ( .C1(n12879), .C2(n10472), .A(n10471), .B(n10470), .ZN(
        n14697) );
  INV_X1 U12886 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n12589) );
  OAI22_X1 U12887 ( .A1(n12889), .A2(n10473), .B1(n12589), .B2(n12886), .ZN(
        n10474) );
  AOI21_X1 U12888 ( .B1(n12896), .B2(n14695), .A(n10474), .ZN(n10480) );
  INV_X1 U12889 ( .A(n12854), .ZN(n10772) );
  INV_X1 U12890 ( .A(n10475), .ZN(n10476) );
  AOI211_X1 U12891 ( .C1(n10477), .C2(n14695), .A(n10476), .B(n12865), .ZN(
        n14694) );
  AOI22_X1 U12892 ( .A1(n10772), .A2(n10478), .B1(n14667), .B2(n14694), .ZN(
        n10479) );
  OAI211_X1 U12893 ( .C1(n14680), .C2(n14697), .A(n10480), .B(n10479), .ZN(
        P2_U3264) );
  INV_X1 U12894 ( .A(n11113), .ZN(n10554) );
  OAI222_X1 U12895 ( .A1(n14165), .A2(n10554), .B1(n14166), .B2(n10481), .C1(
        P1_U3086), .C2(n13587), .ZN(P1_U3335) );
  OAI22_X1 U12896 ( .A1(n10483), .A2(n12777), .B1(n10482), .B2(n12773), .ZN(
        n10663) );
  AOI22_X1 U12897 ( .A1(n12444), .A2(n10663), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10484) );
  OAI21_X1 U12898 ( .B1(n10669), .B2(n12538), .A(n10484), .ZN(n10489) );
  AOI211_X1 U12899 ( .C1(n10487), .C2(n10486), .A(n12571), .B(n10485), .ZN(
        n10488) );
  AOI211_X1 U12900 ( .C1(n10671), .C2(n12569), .A(n10489), .B(n10488), .ZN(
        n10490) );
  INV_X1 U12901 ( .A(n10490), .ZN(P2_U3206) );
  NAND2_X1 U12902 ( .A1(n10492), .A2(n10491), .ZN(n10497) );
  AND2_X1 U12903 ( .A1(n10499), .A2(n10497), .ZN(n10501) );
  NAND2_X1 U12904 ( .A1(n14498), .A2(n13311), .ZN(n10494) );
  NAND2_X1 U12905 ( .A1(n13662), .A2(n9725), .ZN(n10493) );
  NAND2_X1 U12906 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  XNOR2_X1 U12907 ( .A(n10495), .B(n13022), .ZN(n10557) );
  AND2_X1 U12908 ( .A1(n13662), .A2(n13313), .ZN(n10496) );
  AOI21_X1 U12909 ( .B1(n14498), .B2(n9725), .A(n10496), .ZN(n10560) );
  XNOR2_X1 U12910 ( .A(n10557), .B(n10560), .ZN(n10500) );
  AND2_X1 U12911 ( .A1(n10500), .A2(n10497), .ZN(n10498) );
  OAI211_X1 U12912 ( .C1(n10501), .C2(n10500), .A(n14366), .B(n10558), .ZN(
        n10506) );
  INV_X1 U12913 ( .A(n10502), .ZN(n10503) );
  NAND2_X1 U12914 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13718) );
  OAI21_X1 U12915 ( .B1(n14376), .B2(n10503), .A(n13718), .ZN(n10504) );
  AOI21_X1 U12916 ( .B1(n14497), .B2(n14373), .A(n10504), .ZN(n10505) );
  OAI211_X1 U12917 ( .C1(n7109), .C2(n13393), .A(n10506), .B(n10505), .ZN(
        P1_U3231) );
  NAND2_X1 U12918 ( .A1(n14498), .A2(n10565), .ZN(n10507) );
  NAND2_X1 U12919 ( .A1(n10509), .A2(n13595), .ZN(n10512) );
  AOI22_X1 U12920 ( .A1(n13594), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11102), 
        .B2(n10510), .ZN(n10511) );
  XNOR2_X1 U12921 ( .A(n13482), .B(n13661), .ZN(n13619) );
  INV_X1 U12922 ( .A(n13619), .ZN(n10513) );
  AOI21_X1 U12923 ( .B1(n10514), .B2(n10513), .A(n14501), .ZN(n10515) );
  AOI22_X1 U12924 ( .A1(n10515), .A2(n10572), .B1(n14416), .B2(n13662), .ZN(
        n14511) );
  XNOR2_X1 U12925 ( .A(n10586), .B(n13619), .ZN(n14516) );
  NAND2_X1 U12926 ( .A1(n14516), .A2(n14433), .ZN(n10530) );
  NAND2_X1 U12927 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NAND2_X1 U12928 ( .A1(n10578), .A2(n10519), .ZN(n14306) );
  INV_X1 U12929 ( .A(n14306), .ZN(n10589) );
  NAND2_X1 U12930 ( .A1(n11208), .A2(n10589), .ZN(n10523) );
  NAND2_X1 U12931 ( .A1(n13580), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U12932 ( .A1(n8606), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U12933 ( .A1(n11209), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10520) );
  NAND4_X1 U12934 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n13660) );
  AOI211_X1 U12935 ( .C1(n13482), .C2(n10524), .A(n14076), .B(n10588), .ZN(
        n10525) );
  AOI21_X1 U12936 ( .B1(n14413), .B2(n13660), .A(n10525), .ZN(n14510) );
  INV_X1 U12937 ( .A(n14510), .ZN(n10528) );
  INV_X1 U12938 ( .A(n13482), .ZN(n14513) );
  AOI22_X1 U12939 ( .A1(n6479), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n10568), 
        .B2(n14400), .ZN(n10526) );
  OAI21_X1 U12940 ( .B1(n14513), .B2(n14422), .A(n10526), .ZN(n10527) );
  AOI21_X1 U12941 ( .B1(n10528), .B2(n14432), .A(n10527), .ZN(n10529) );
  OAI211_X1 U12942 ( .C1(n6479), .C2(n14511), .A(n10530), .B(n10529), .ZN(
        P1_U3283) );
  MUX2_X1 U12943 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12069), .Z(n10708) );
  NAND2_X1 U12944 ( .A1(n10531), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10532) );
  MUX2_X1 U12945 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10532), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n10533) );
  NAND2_X1 U12946 ( .A1(n10533), .A2(n11008), .ZN(n14191) );
  XNOR2_X1 U12947 ( .A(n10708), .B(n14191), .ZN(n10539) );
  INV_X1 U12948 ( .A(n10534), .ZN(n10536) );
  OAI21_X1 U12949 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(n10538) );
  AOI21_X1 U12950 ( .B1(n10539), .B2(n10538), .A(n10709), .ZN(n10552) );
  NAND2_X1 U12951 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n10934), .ZN(n10541) );
  NAND2_X1 U12952 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n10542), .ZN(n10723) );
  OAI21_X1 U12953 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n10542), .A(n10723), 
        .ZN(n10545) );
  AND2_X1 U12954 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11973) );
  AOI21_X1 U12955 ( .B1(n14780), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11973), 
        .ZN(n10543) );
  OAI21_X1 U12956 ( .B1(n14797), .B2(n14191), .A(n10543), .ZN(n10544) );
  AOI21_X1 U12957 ( .B1(n10545), .B2(n14801), .A(n10544), .ZN(n10551) );
  NAND2_X1 U12958 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10934), .ZN(n10547) );
  NAND2_X1 U12959 ( .A1(n10547), .A2(n10546), .ZN(n10717) );
  XNOR2_X1 U12960 ( .A(n10717), .B(n11268), .ZN(n10548) );
  NAND2_X1 U12961 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n10548), .ZN(n10718) );
  OAI21_X1 U12962 ( .B1(n10548), .B2(P3_REG1_REG_13__SCAN_IN), .A(n10718), 
        .ZN(n10549) );
  NAND2_X1 U12963 ( .A1(n10549), .A2(n14788), .ZN(n10550) );
  OAI211_X1 U12964 ( .C1(n10552), .C2(n12113), .A(n10551), .B(n10550), .ZN(
        P3_U3195) );
  OAI222_X1 U12965 ( .A1(P2_U3088), .A2(n10555), .B1(n10648), .B2(n10554), 
        .C1(n10553), .C2(n13010), .ZN(P2_U3307) );
  INV_X1 U12966 ( .A(n11121), .ZN(n10647) );
  INV_X1 U12967 ( .A(n10556), .ZN(n13605) );
  OAI222_X1 U12968 ( .A1(n14165), .A2(n10647), .B1(n13605), .B2(P1_U3086), 
        .C1(n7231), .C2(n14166), .ZN(P1_U3334) );
  INV_X1 U12969 ( .A(n10557), .ZN(n10559) );
  NAND2_X1 U12970 ( .A1(n13482), .A2(n13311), .ZN(n10562) );
  NAND2_X1 U12971 ( .A1(n13661), .A2(n9725), .ZN(n10561) );
  NAND2_X1 U12972 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  XNOR2_X1 U12973 ( .A(n10563), .B(n13022), .ZN(n10873) );
  AND2_X1 U12974 ( .A1(n13661), .A2(n13313), .ZN(n10564) );
  AOI21_X1 U12975 ( .B1(n13482), .B2(n9725), .A(n10564), .ZN(n10872) );
  XNOR2_X1 U12976 ( .A(n10873), .B(n10872), .ZN(n10875) );
  XNOR2_X1 U12977 ( .A(n10876), .B(n10875), .ZN(n10571) );
  INV_X1 U12978 ( .A(n13660), .ZN(n10803) );
  OAI22_X1 U12979 ( .A1(n10803), .A2(n13400), .B1(n10565), .B2(n13399), .ZN(
        n10566) );
  AOI211_X1 U12980 ( .C1(n13403), .C2(n10568), .A(n10567), .B(n10566), .ZN(
        n10570) );
  NAND2_X1 U12981 ( .A1(n13482), .A2(n14300), .ZN(n10569) );
  OAI211_X1 U12982 ( .C1(n10571), .C2(n13425), .A(n10570), .B(n10569), .ZN(
        P1_U3217) );
  INV_X1 U12983 ( .A(n13661), .ZN(n10584) );
  NAND2_X1 U12984 ( .A1(n10573), .A2(n13595), .ZN(n10576) );
  AOI22_X1 U12985 ( .A1(n13594), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11102), 
        .B2(n10574), .ZN(n10575) );
  XNOR2_X1 U12986 ( .A(n14301), .B(n13660), .ZN(n13620) );
  XNOR2_X1 U12987 ( .A(n10794), .B(n10805), .ZN(n10585) );
  AND2_X1 U12988 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  NOR2_X1 U12989 ( .A1(n10796), .A2(n10579), .ZN(n10887) );
  NAND2_X1 U12990 ( .A1(n11208), .A2(n10887), .ZN(n10583) );
  NAND2_X1 U12991 ( .A1(n13580), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U12992 ( .A1(n8606), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U12993 ( .A1(n11209), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10580) );
  NAND4_X1 U12994 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(
        n13659) );
  INV_X1 U12995 ( .A(n13659), .ZN(n10853) );
  OAI22_X1 U12996 ( .A1(n10584), .A2(n14015), .B1(n10853), .B2(n14013), .ZN(
        n14303) );
  AOI21_X1 U12997 ( .B1(n10585), .B2(n14411), .A(n14303), .ZN(n14330) );
  XNOR2_X1 U12998 ( .A(n10806), .B(n10805), .ZN(n14333) );
  INV_X1 U12999 ( .A(n10807), .ZN(n10587) );
  OAI211_X1 U13000 ( .C1(n14331), .C2(n10588), .A(n10587), .B(n14429), .ZN(
        n14329) );
  AOI22_X1 U13001 ( .A1(n6479), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10589), 
        .B2(n14400), .ZN(n10591) );
  NAND2_X1 U13002 ( .A1(n14301), .A2(n14033), .ZN(n10590) );
  OAI211_X1 U13003 ( .C1(n14329), .C2(n14022), .A(n10591), .B(n10590), .ZN(
        n10592) );
  AOI21_X1 U13004 ( .B1(n14333), .B2(n14433), .A(n10592), .ZN(n10593) );
  OAI21_X1 U13005 ( .B1(n6479), .B2(n14330), .A(n10593), .ZN(P1_U3282) );
  XOR2_X1 U13006 ( .A(n11156), .B(n10845), .Z(n11406) );
  INV_X1 U13007 ( .A(SI_24_), .ZN(n11407) );
  OAI22_X1 U13008 ( .A1(n10597), .A2(n6473), .B1(n11407), .B2(n14186), .ZN(
        n10598) );
  AOI21_X1 U13009 ( .B1(n11406), .B2(n14205), .A(n10598), .ZN(n10599) );
  INV_X1 U13010 ( .A(n10599), .ZN(P3_U3271) );
  XNOR2_X1 U13011 ( .A(n10601), .B(n10600), .ZN(n14182) );
  NAND2_X1 U13012 ( .A1(n11464), .A2(n14182), .ZN(n10605) );
  OR2_X1 U13013 ( .A1(n11348), .A2(n10602), .ZN(n10604) );
  OR2_X1 U13014 ( .A1(n11454), .A2(SI_9_), .ZN(n10603) );
  XNOR2_X1 U13015 ( .A(n10943), .B(n6828), .ZN(n10813) );
  XNOR2_X1 U13016 ( .A(n10813), .B(n10919), .ZN(n10612) );
  INV_X1 U13017 ( .A(n10606), .ZN(n10607) );
  OR2_X1 U13018 ( .A1(n10607), .A2(n14819), .ZN(n10608) );
  NAND2_X1 U13019 ( .A1(n10609), .A2(n10608), .ZN(n10611) );
  OR2_X2 U13020 ( .A1(n10611), .A2(n10612), .ZN(n10815) );
  INV_X1 U13021 ( .A(n10815), .ZN(n10610) );
  AOI21_X1 U13022 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10625) );
  NAND2_X1 U13023 ( .A1(n11465), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n10619) );
  NAND2_X1 U13024 ( .A1(n10613), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13025 ( .A1(n10823), .A2(n10614), .ZN(n14810) );
  INV_X1 U13026 ( .A(n14810), .ZN(n10836) );
  OR2_X1 U13027 ( .A1(n11400), .A2(n10836), .ZN(n10618) );
  INV_X1 U13028 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n10615) );
  OR2_X1 U13029 ( .A1(n11466), .A2(n10615), .ZN(n10617) );
  OR2_X1 U13030 ( .A1(n11468), .A2(n9959), .ZN(n10616) );
  AOI21_X1 U13031 ( .B1(n14237), .B2(n12013), .A(n10620), .ZN(n10621) );
  OAI21_X1 U13032 ( .B1(n14819), .B2(n12009), .A(n10621), .ZN(n10623) );
  NOR2_X1 U13033 ( .A1(n12015), .A2(n14823), .ZN(n10622) );
  AOI211_X1 U13034 ( .C1(n10943), .C2(n12017), .A(n10623), .B(n10622), .ZN(
        n10624) );
  OAI21_X1 U13035 ( .B1(n10625), .B2(n12019), .A(n10624), .ZN(P3_U3171) );
  INV_X1 U13036 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13037 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13349)
         );
  OAI21_X1 U13038 ( .B1(n14391), .B2(n10626), .A(n13349), .ZN(n10634) );
  NAND2_X1 U13039 ( .A1(n10628), .A2(n10629), .ZN(n10630) );
  INV_X1 U13040 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U13041 ( .A1(n14382), .A2(n14381), .ZN(n14380) );
  NAND2_X1 U13042 ( .A1(n10630), .A2(n14380), .ZN(n10632) );
  XNOR2_X1 U13043 ( .A(n13736), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10631) );
  NOR2_X1 U13044 ( .A1(n10631), .A2(n10632), .ZN(n13735) );
  AOI211_X1 U13045 ( .C1(n10632), .C2(n10631), .A(n13735), .B(n13737), .ZN(
        n10633) );
  AOI211_X1 U13046 ( .C1(n14383), .C2(n13736), .A(n10634), .B(n10633), .ZN(
        n10645) );
  OAI21_X1 U13047 ( .B1(n9939), .B2(n10636), .A(n10635), .ZN(n10637) );
  NOR2_X1 U13048 ( .A1(n14384), .A2(n10637), .ZN(n10638) );
  XNOR2_X1 U13049 ( .A(n14384), .B(n10637), .ZN(n14378) );
  NOR2_X1 U13050 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14378), .ZN(n14377) );
  NOR2_X1 U13051 ( .A1(n10638), .A2(n14377), .ZN(n10643) );
  INV_X1 U13052 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10641) );
  NAND2_X1 U13053 ( .A1(n13736), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13731) );
  INV_X1 U13054 ( .A(n13731), .ZN(n10639) );
  AOI21_X1 U13055 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n10642) );
  NAND2_X1 U13056 ( .A1(n10642), .A2(n10643), .ZN(n13730) );
  OAI211_X1 U13057 ( .C1(n10643), .C2(n10642), .A(n14387), .B(n13730), .ZN(
        n10644) );
  NAND2_X1 U13058 ( .A1(n10645), .A2(n10644), .ZN(P1_U3259) );
  OAI222_X1 U13059 ( .A1(P2_U3088), .A2(n10649), .B1(n10648), .B2(n10647), 
        .C1(n10646), .C2(n13010), .ZN(P2_U3306) );
  XNOR2_X1 U13060 ( .A(n10650), .B(n7292), .ZN(n10840) );
  INV_X1 U13061 ( .A(n10840), .ZN(n10661) );
  XNOR2_X1 U13062 ( .A(n10652), .B(n10651), .ZN(n10653) );
  NOR2_X1 U13063 ( .A1(n10653), .A2(n12774), .ZN(n10838) );
  AND2_X1 U13064 ( .A1(n12882), .A2(n12577), .ZN(n10654) );
  AOI21_X1 U13065 ( .B1(n12862), .B2(n12880), .A(n10654), .ZN(n11776) );
  INV_X1 U13066 ( .A(n11776), .ZN(n10655) );
  OAI21_X1 U13067 ( .B1(n10838), .B2(n10655), .A(n12889), .ZN(n10660) );
  OAI22_X1 U13068 ( .A1(n12889), .A2(n14621), .B1(n11774), .B2(n12886), .ZN(
        n10658) );
  INV_X1 U13069 ( .A(n10656), .ZN(n12876) );
  OAI211_X1 U13070 ( .C1(n11718), .C2(n10683), .A(n12876), .B(n12971), .ZN(
        n10837) );
  NOR2_X1 U13071 ( .A1(n10837), .A2(n12811), .ZN(n10657) );
  AOI211_X1 U13072 ( .C1(n12896), .C2(n11779), .A(n10658), .B(n10657), .ZN(
        n10659) );
  OAI211_X1 U13073 ( .C1(n10661), .C2(n12893), .A(n10660), .B(n10659), .ZN(
        P2_U3250) );
  XOR2_X1 U13074 ( .A(n10662), .B(n10666), .Z(n10665) );
  INV_X1 U13075 ( .A(n10663), .ZN(n10664) );
  OAI21_X1 U13076 ( .B1(n10665), .B2(n12774), .A(n10664), .ZN(n14271) );
  INV_X1 U13077 ( .A(n14271), .ZN(n10675) );
  XNOR2_X1 U13078 ( .A(n10667), .B(n10666), .ZN(n14273) );
  INV_X1 U13079 ( .A(n10765), .ZN(n10668) );
  OAI211_X1 U13080 ( .C1(n10668), .C2(n14270), .A(n12971), .B(n10680), .ZN(
        n14269) );
  OAI22_X1 U13081 ( .A1(n12889), .A2(n10421), .B1(n10669), .B2(n12886), .ZN(
        n10670) );
  AOI21_X1 U13082 ( .B1(n10671), .B2(n12896), .A(n10670), .ZN(n10672) );
  OAI21_X1 U13083 ( .B1(n14269), .B2(n12811), .A(n10672), .ZN(n10673) );
  AOI21_X1 U13084 ( .B1(n14273), .B2(n14677), .A(n10673), .ZN(n10674) );
  OAI21_X1 U13085 ( .B1(n10675), .B2(n14680), .A(n10674), .ZN(P2_U3252) );
  XNOR2_X1 U13086 ( .A(n10676), .B(n10679), .ZN(n10677) );
  OAI222_X1 U13087 ( .A1(n12777), .A2(n11719), .B1(n12773), .B2(n10759), .C1(
        n12774), .C2(n10677), .ZN(n14265) );
  INV_X1 U13088 ( .A(n14265), .ZN(n10691) );
  XOR2_X1 U13089 ( .A(n10678), .B(n10679), .Z(n14267) );
  NAND2_X1 U13090 ( .A1(n10687), .A2(n10680), .ZN(n10681) );
  NAND2_X1 U13091 ( .A1(n10681), .A2(n12971), .ZN(n10682) );
  OR2_X1 U13092 ( .A1(n10683), .A2(n10682), .ZN(n14263) );
  NAND2_X1 U13093 ( .A1(n14680), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10684) );
  OAI21_X1 U13094 ( .B1(n12886), .B2(n10685), .A(n10684), .ZN(n10686) );
  AOI21_X1 U13095 ( .B1(n10687), .B2(n12896), .A(n10686), .ZN(n10688) );
  OAI21_X1 U13096 ( .B1(n14263), .B2(n12811), .A(n10688), .ZN(n10689) );
  AOI21_X1 U13097 ( .B1(n14267), .B2(n14677), .A(n10689), .ZN(n10690) );
  OAI21_X1 U13098 ( .B1(n10691), .B2(n14680), .A(n10690), .ZN(P2_U3251) );
  NAND2_X1 U13099 ( .A1(n10692), .A2(n10694), .ZN(n10693) );
  NAND2_X1 U13100 ( .A1(n7195), .A2(n10693), .ZN(n14747) );
  AOI22_X1 U13101 ( .A1(n12880), .A2(n12581), .B1(n12882), .B2(n12583), .ZN(
        n10698) );
  XNOR2_X1 U13102 ( .A(n10695), .B(n10694), .ZN(n10696) );
  NAND2_X1 U13103 ( .A1(n10696), .A2(n12879), .ZN(n10697) );
  OAI211_X1 U13104 ( .C1(n14747), .C2(n6485), .A(n10698), .B(n10697), .ZN(
        n14750) );
  NAND2_X1 U13105 ( .A1(n14750), .A2(n12889), .ZN(n10707) );
  OAI22_X1 U13106 ( .A1(n12889), .A2(n10700), .B1(n10699), .B2(n12886), .ZN(
        n10704) );
  OAI211_X1 U13107 ( .C1(n10702), .C2(n14749), .A(n12971), .B(n10701), .ZN(
        n14748) );
  NOR2_X1 U13108 ( .A1(n12811), .A2(n14748), .ZN(n10703) );
  AOI211_X1 U13109 ( .C1(n12896), .C2(n10705), .A(n10704), .B(n10703), .ZN(
        n10706) );
  OAI211_X1 U13110 ( .C1(n14747), .C2(n12854), .A(n10707), .B(n10706), .ZN(
        P2_U3257) );
  INV_X1 U13111 ( .A(n10708), .ZN(n10710) );
  NAND2_X1 U13112 ( .A1(n11008), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10712) );
  XNOR2_X1 U13113 ( .A(n10712), .B(n10711), .ZN(n14196) );
  NAND2_X1 U13114 ( .A1(n14196), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n11018) );
  OR2_X1 U13115 ( .A1(n14196), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n10713) );
  AND2_X1 U13116 ( .A1(n11018), .A2(n10713), .ZN(n10725) );
  NAND2_X1 U13117 ( .A1(n14196), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11021) );
  OR2_X1 U13118 ( .A1(n14196), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10714) );
  AND2_X1 U13119 ( .A1(n11021), .A2(n10714), .ZN(n10721) );
  MUX2_X1 U13120 ( .A(n10725), .B(n10721), .S(n12069), .Z(n10715) );
  OAI211_X1 U13121 ( .C1(n10716), .C2(n10715), .A(n11012), .B(n14792), .ZN(
        n10734) );
  NAND2_X1 U13122 ( .A1(n14191), .A2(n10717), .ZN(n10719) );
  NAND2_X1 U13123 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  NAND2_X1 U13124 ( .A1(n10720), .A2(n10721), .ZN(n11020) );
  OAI21_X1 U13125 ( .B1(n10721), .B2(n10720), .A(n11020), .ZN(n10732) );
  NAND2_X1 U13126 ( .A1(n14191), .A2(n10722), .ZN(n10724) );
  OAI21_X1 U13127 ( .B1(n10726), .B2(n10725), .A(n11017), .ZN(n10727) );
  NAND2_X1 U13128 ( .A1(n10727), .A2(n14801), .ZN(n10730) );
  INV_X1 U13129 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n10728) );
  NOR2_X1 U13130 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10728), .ZN(n11866) );
  AOI21_X1 U13131 ( .B1(n14780), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11866), 
        .ZN(n10729) );
  OAI211_X1 U13132 ( .C1(n14797), .C2(n14196), .A(n10730), .B(n10729), .ZN(
        n10731) );
  AOI21_X1 U13133 ( .B1(n14788), .B2(n10732), .A(n10731), .ZN(n10733) );
  NAND2_X1 U13134 ( .A1(n10734), .A2(n10733), .ZN(P3_U3196) );
  XNOR2_X1 U13135 ( .A(n10735), .B(n10736), .ZN(n14754) );
  XNOR2_X1 U13136 ( .A(n10737), .B(n10736), .ZN(n10740) );
  OAI22_X1 U13137 ( .A1(n10758), .A2(n12777), .B1(n12773), .B2(n10738), .ZN(
        n10739) );
  AOI21_X1 U13138 ( .B1(n10740), .B2(n12879), .A(n10739), .ZN(n10741) );
  OAI21_X1 U13139 ( .B1(n14754), .B2(n6485), .A(n10741), .ZN(n14758) );
  NAND2_X1 U13140 ( .A1(n14758), .A2(n12889), .ZN(n10752) );
  INV_X1 U13141 ( .A(n10742), .ZN(n10743) );
  OAI22_X1 U13142 ( .A1(n12889), .A2(n10744), .B1(n10743), .B2(n12886), .ZN(
        n10749) );
  INV_X1 U13143 ( .A(n10750), .ZN(n14757) );
  INV_X1 U13144 ( .A(n10745), .ZN(n10747) );
  OAI211_X1 U13145 ( .C1(n14757), .C2(n10747), .A(n10746), .B(n12971), .ZN(
        n14755) );
  NOR2_X1 U13146 ( .A1(n14755), .A2(n12811), .ZN(n10748) );
  AOI211_X1 U13147 ( .C1(n12896), .C2(n10750), .A(n10749), .B(n10748), .ZN(
        n10751) );
  OAI211_X1 U13148 ( .C1(n14754), .C2(n12854), .A(n10752), .B(n10751), .ZN(
        P2_U3255) );
  XNOR2_X1 U13149 ( .A(n10753), .B(n10754), .ZN(n14278) );
  NAND2_X1 U13150 ( .A1(n14278), .A2(n14745), .ZN(n10764) );
  NOR2_X1 U13151 ( .A1(n10755), .A2(n10754), .ZN(n10757) );
  OR3_X1 U13152 ( .A1(n10757), .A2(n10756), .A3(n12774), .ZN(n10762) );
  OAI22_X1 U13153 ( .A1(n10759), .A2(n12777), .B1(n10758), .B2(n12773), .ZN(
        n10760) );
  INV_X1 U13154 ( .A(n10760), .ZN(n10761) );
  AND2_X1 U13155 ( .A1(n10762), .A2(n10761), .ZN(n10763) );
  AND2_X1 U13156 ( .A1(n10764), .A2(n10763), .ZN(n14280) );
  OAI211_X1 U13157 ( .C1(n10766), .C2(n14276), .A(n12971), .B(n10765), .ZN(
        n14275) );
  AOI22_X1 U13158 ( .A1(n14680), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10767), 
        .B2(n14669), .ZN(n10770) );
  NAND2_X1 U13159 ( .A1(n12896), .A2(n10768), .ZN(n10769) );
  OAI211_X1 U13160 ( .C1(n14275), .C2(n12811), .A(n10770), .B(n10769), .ZN(
        n10771) );
  AOI21_X1 U13161 ( .B1(n14278), .B2(n10772), .A(n10771), .ZN(n10773) );
  OAI21_X1 U13162 ( .B1(n14280), .B2(n14680), .A(n10773), .ZN(P2_U3253) );
  XNOR2_X1 U13163 ( .A(n10774), .B(n10775), .ZN(n14713) );
  OR2_X1 U13164 ( .A1(n10776), .A2(n10775), .ZN(n10777) );
  AOI21_X1 U13165 ( .B1(n10778), .B2(n10777), .A(n12774), .ZN(n10781) );
  OAI22_X1 U13166 ( .A1(n10779), .A2(n12777), .B1(n8269), .B2(n12773), .ZN(
        n10780) );
  OR2_X1 U13167 ( .A1(n10781), .A2(n10780), .ZN(n14712) );
  OAI211_X1 U13168 ( .C1(n14710), .C2(n10783), .A(n12971), .B(n10782), .ZN(
        n14709) );
  AOI22_X1 U13169 ( .A1(n12858), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n14669), 
        .B2(n10784), .ZN(n10787) );
  NAND2_X1 U13170 ( .A1(n12896), .A2(n10785), .ZN(n10786) );
  OAI211_X1 U13171 ( .C1(n12811), .C2(n14709), .A(n10787), .B(n10786), .ZN(
        n10788) );
  AOI21_X1 U13172 ( .B1(n12889), .B2(n14712), .A(n10788), .ZN(n10789) );
  OAI21_X1 U13173 ( .B1(n14713), .B2(n12893), .A(n10789), .ZN(P2_U3262) );
  NAND2_X1 U13174 ( .A1(n10790), .A2(n13595), .ZN(n10793) );
  AOI22_X1 U13175 ( .A1(n13594), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11102), 
        .B2(n10791), .ZN(n10792) );
  XNOR2_X1 U13176 ( .A(n13490), .B(n13659), .ZN(n13622) );
  OR2_X1 U13177 ( .A1(n14301), .A2(n10803), .ZN(n10795) );
  XOR2_X1 U13178 ( .A(n13622), .B(n10852), .Z(n10802) );
  NOR2_X1 U13179 ( .A1(n10796), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10797) );
  NAND2_X1 U13180 ( .A1(n11208), .A2(n7525), .ZN(n10801) );
  NAND2_X1 U13181 ( .A1(n13580), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10800) );
  NAND2_X1 U13182 ( .A1(n11209), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13183 ( .A1(n8606), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13184 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n13658) );
  OAI22_X1 U13185 ( .A1(n10803), .A2(n14015), .B1(n10973), .B2(n14013), .ZN(
        n10890) );
  AOI21_X1 U13186 ( .B1(n10802), .B2(n14411), .A(n10890), .ZN(n14215) );
  XNOR2_X1 U13187 ( .A(n10859), .B(n13622), .ZN(n14218) );
  OAI21_X1 U13188 ( .B1(n10807), .B2(n14216), .A(n14429), .ZN(n10808) );
  OR2_X1 U13189 ( .A1(n10867), .A2(n10808), .ZN(n14214) );
  AOI22_X1 U13190 ( .A1(n6479), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n10887), 
        .B2(n14400), .ZN(n10810) );
  NAND2_X1 U13191 ( .A1(n13490), .A2(n14033), .ZN(n10809) );
  OAI211_X1 U13192 ( .C1(n14214), .C2(n14022), .A(n10810), .B(n10809), .ZN(
        n10811) );
  AOI21_X1 U13193 ( .B1(n14218), .B2(n14433), .A(n10811), .ZN(n10812) );
  OAI21_X1 U13194 ( .B1(n6479), .B2(n14215), .A(n10812), .ZN(P1_U3281) );
  NAND2_X1 U13195 ( .A1(n10813), .A2(n10919), .ZN(n10814) );
  OR2_X1 U13196 ( .A1(n11454), .A2(SI_10_), .ZN(n10819) );
  OR2_X1 U13197 ( .A1(n11348), .A2(n10817), .ZN(n10818) );
  XNOR2_X1 U13198 ( .A(n10945), .B(n11892), .ZN(n10996) );
  XNOR2_X1 U13199 ( .A(n10996), .B(n14818), .ZN(n10821) );
  OAI211_X1 U13200 ( .C1(n10822), .C2(n10821), .A(n10999), .B(n11984), .ZN(
        n10835) );
  NAND2_X1 U13201 ( .A1(n11465), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13202 ( .A1(n10823), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10824) );
  AND2_X1 U13203 ( .A1(n10928), .A2(n10824), .ZN(n14238) );
  OR2_X1 U13204 ( .A1(n11400), .A2(n14238), .ZN(n10829) );
  INV_X1 U13205 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10825) );
  OR2_X1 U13206 ( .A1(n11468), .A2(n10825), .ZN(n10828) );
  INV_X1 U13207 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n10826) );
  OR2_X1 U13208 ( .A1(n11466), .A2(n10826), .ZN(n10827) );
  NAND4_X1 U13209 ( .A1(n10830), .A2(n10829), .A3(n10828), .A4(n10827), .ZN(
        n14807) );
  AOI21_X1 U13210 ( .B1(n12013), .B2(n14807), .A(n10831), .ZN(n10832) );
  OAI21_X1 U13211 ( .B1(n10919), .B2(n12009), .A(n10832), .ZN(n10833) );
  AOI21_X1 U13212 ( .B1(n10945), .B2(n12017), .A(n10833), .ZN(n10834) );
  OAI211_X1 U13213 ( .C1(n10836), .C2(n12015), .A(n10835), .B(n10834), .ZN(
        P3_U3157) );
  INV_X1 U13214 ( .A(n14720), .ZN(n14274) );
  OAI211_X1 U13215 ( .C1(n11718), .C2(n14756), .A(n10837), .B(n11776), .ZN(
        n10839) );
  AOI211_X1 U13216 ( .C1(n14274), .C2(n10840), .A(n10839), .B(n10838), .ZN(
        n10843) );
  NAND2_X1 U13217 ( .A1(n14777), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10841) );
  OAI21_X1 U13218 ( .B1(n10843), .B2(n14777), .A(n10841), .ZN(P2_U3514) );
  NAND2_X1 U13219 ( .A1(n14762), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10842) );
  OAI21_X1 U13220 ( .B1(n10843), .B2(n14762), .A(n10842), .ZN(P2_U3475) );
  NAND2_X1 U13221 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n10844), .ZN(n10847) );
  NAND2_X1 U13222 ( .A1(n10845), .A2(n11156), .ZN(n10846) );
  AOI22_X1 U13223 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13011), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n14172), .ZN(n10848) );
  INV_X1 U13224 ( .A(n10848), .ZN(n10849) );
  XNOR2_X1 U13225 ( .A(n10894), .B(n10849), .ZN(n11417) );
  INV_X1 U13226 ( .A(n11417), .ZN(n10850) );
  OAI222_X1 U13227 ( .A1(n6473), .A2(n10851), .B1(n14186), .B2(n11418), .C1(
        n12423), .C2(n10850), .ZN(P3_U3270) );
  NAND2_X1 U13228 ( .A1(n10854), .A2(n13595), .ZN(n10857) );
  AOI22_X1 U13229 ( .A1(n13594), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10855), 
        .B2(n11102), .ZN(n10856) );
  XNOR2_X1 U13230 ( .A(n13499), .B(n10973), .ZN(n13624) );
  INV_X1 U13231 ( .A(n13624), .ZN(n10965) );
  XNOR2_X1 U13232 ( .A(n10966), .B(n10965), .ZN(n14322) );
  XNOR2_X1 U13233 ( .A(n10974), .B(n13624), .ZN(n14328) );
  NAND2_X1 U13234 ( .A1(n14328), .A2(n14433), .ZN(n10871) );
  NAND2_X1 U13235 ( .A1(n8606), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U13236 ( .A1(n10860), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10977) );
  OR2_X1 U13237 ( .A1(n10860), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U13238 ( .A1(n10977), .A2(n10861), .ZN(n14296) );
  INV_X1 U13239 ( .A(n14296), .ZN(n10985) );
  NAND2_X1 U13240 ( .A1(n11208), .A2(n10985), .ZN(n10864) );
  NAND2_X1 U13241 ( .A1(n13580), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13242 ( .A1(n11209), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10862) );
  INV_X1 U13243 ( .A(n14016), .ZN(n13657) );
  AOI22_X1 U13244 ( .A1(n13657), .A2(n14413), .B1(n14416), .B2(n13659), .ZN(
        n14323) );
  AOI22_X1 U13245 ( .A1(n6479), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7525), .B2(
        n14400), .ZN(n10866) );
  OAI21_X1 U13246 ( .B1(n14323), .B2(n6479), .A(n10866), .ZN(n10869) );
  OAI211_X1 U13247 ( .C1(n10867), .C2(n14325), .A(n14429), .B(n10987), .ZN(
        n14324) );
  NOR2_X1 U13248 ( .A1(n14324), .A2(n14022), .ZN(n10868) );
  AOI211_X1 U13249 ( .C1(n14033), .C2(n13499), .A(n10869), .B(n10868), .ZN(
        n10870) );
  OAI211_X1 U13250 ( .C1(n14322), .C2(n13962), .A(n10871), .B(n10870), .ZN(
        P1_U3280) );
  INV_X1 U13251 ( .A(n10872), .ZN(n10874) );
  AOI22_X1 U13252 ( .A1(n14301), .A2(n9725), .B1(n13313), .B2(n13660), .ZN(
        n10878) );
  AOI22_X1 U13253 ( .A1(n14301), .A2(n13311), .B1(n9725), .B2(n13660), .ZN(
        n10877) );
  XNOR2_X1 U13254 ( .A(n10877), .B(n13022), .ZN(n10879) );
  XOR2_X1 U13255 ( .A(n10878), .B(n10879), .Z(n14299) );
  NAND2_X1 U13256 ( .A1(n10879), .A2(n10878), .ZN(n10884) );
  AND2_X1 U13257 ( .A1(n14297), .A2(n10884), .ZN(n10886) );
  NAND2_X1 U13258 ( .A1(n13490), .A2(n13311), .ZN(n10881) );
  NAND2_X1 U13259 ( .A1(n13659), .A2(n9725), .ZN(n10880) );
  NAND2_X1 U13260 ( .A1(n10881), .A2(n10880), .ZN(n10882) );
  XNOR2_X1 U13261 ( .A(n10882), .B(n13022), .ZN(n10907) );
  AND2_X1 U13262 ( .A1(n13659), .A2(n13313), .ZN(n10883) );
  AOI21_X1 U13263 ( .B1(n13490), .B2(n9725), .A(n10883), .ZN(n10910) );
  XNOR2_X1 U13264 ( .A(n10907), .B(n10910), .ZN(n10885) );
  NAND3_X1 U13265 ( .A1(n14297), .A2(n10885), .A3(n10884), .ZN(n10908) );
  OAI211_X1 U13266 ( .C1(n10886), .C2(n10885), .A(n14366), .B(n10908), .ZN(
        n10892) );
  INV_X1 U13267 ( .A(n10887), .ZN(n10888) );
  OAI22_X1 U13268 ( .A1(n14376), .A2(n10888), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10577), .ZN(n10889) );
  AOI21_X1 U13269 ( .B1(n10890), .B2(n14373), .A(n10889), .ZN(n10891) );
  OAI211_X1 U13270 ( .C1(n14216), .C2(n13393), .A(n10892), .B(n10891), .ZN(
        P1_U3224) );
  NAND2_X1 U13271 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13011), .ZN(n10893) );
  AOI22_X1 U13272 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13006), .B2(n7241), .ZN(n10895) );
  INV_X1 U13273 ( .A(n10895), .ZN(n10896) );
  XNOR2_X1 U13274 ( .A(n11247), .B(n10896), .ZN(n11429) );
  INV_X1 U13275 ( .A(n11429), .ZN(n10897) );
  OAI222_X1 U13276 ( .A1(P3_U3151), .A2(n10898), .B1(n14186), .B2(n11430), 
        .C1(n12423), .C2(n10897), .ZN(P3_U3269) );
  NAND2_X1 U13277 ( .A1(n11142), .A2(n10899), .ZN(n10900) );
  OAI211_X1 U13278 ( .C1(n11143), .C2(n14166), .A(n10900), .B(n13645), .ZN(
        P1_U3332) );
  NAND2_X1 U13279 ( .A1(n11142), .A2(n10901), .ZN(n10903) );
  OAI211_X1 U13280 ( .C1(n10904), .C2(n13010), .A(n10903), .B(n10902), .ZN(
        P2_U3304) );
  INV_X1 U13281 ( .A(n11155), .ZN(n10995) );
  AOI22_X1 U13282 ( .A1(n10905), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n12998), .ZN(n10906) );
  OAI21_X1 U13283 ( .B1(n10995), .B2(n13012), .A(n10906), .ZN(P2_U3303) );
  INV_X1 U13284 ( .A(n10907), .ZN(n10909) );
  OAI21_X1 U13285 ( .B1(n10910), .B2(n10909), .A(n10908), .ZN(n13021) );
  AND2_X1 U13286 ( .A1(n13658), .A2(n13313), .ZN(n10911) );
  AOI21_X1 U13287 ( .B1(n13499), .B2(n9725), .A(n10911), .ZN(n13016) );
  AOI22_X1 U13288 ( .A1(n13499), .A2(n13311), .B1(n9725), .B2(n13658), .ZN(
        n10912) );
  XNOR2_X1 U13289 ( .A(n10912), .B(n13022), .ZN(n13017) );
  XOR2_X1 U13290 ( .A(n13016), .B(n13017), .Z(n13020) );
  XNOR2_X1 U13291 ( .A(n13021), .B(n13020), .ZN(n10916) );
  AOI22_X1 U13292 ( .A1(n13403), .A2(n7525), .B1(P1_REG3_REG_13__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10913) );
  OAI21_X1 U13293 ( .B1(n14323), .B2(n13332), .A(n10913), .ZN(n10914) );
  AOI21_X1 U13294 ( .B1(n13499), .B2(n14300), .A(n10914), .ZN(n10915) );
  OAI21_X1 U13295 ( .B1(n10916), .B2(n13425), .A(n10915), .ZN(P1_U3234) );
  NAND2_X1 U13296 ( .A1(n14228), .A2(n14878), .ZN(n10917) );
  INV_X1 U13297 ( .A(n10943), .ZN(n14827) );
  NAND2_X1 U13298 ( .A1(n14809), .A2(n14827), .ZN(n11544) );
  NAND2_X1 U13299 ( .A1(n10919), .A2(n10943), .ZN(n11543) );
  NAND2_X1 U13300 ( .A1(n14818), .A2(n10945), .ZN(n11547) );
  INV_X1 U13301 ( .A(n10945), .ZN(n14815) );
  NAND2_X1 U13302 ( .A1(n14237), .A2(n14815), .ZN(n11548) );
  NAND2_X1 U13303 ( .A1(n11547), .A2(n11548), .ZN(n14814) );
  AND2_X2 U13304 ( .A1(n14811), .A2(n11548), .ZN(n14241) );
  OR2_X1 U13305 ( .A1(n11454), .A2(SI_11_), .ZN(n10924) );
  OR2_X1 U13306 ( .A1(n11348), .A2(n10922), .ZN(n10923) );
  NAND2_X1 U13307 ( .A1(n11913), .A2(n11005), .ZN(n11552) );
  INV_X1 U13308 ( .A(n11005), .ZN(n14242) );
  NAND2_X1 U13309 ( .A1(n14807), .A2(n14242), .ZN(n11553) );
  NAND2_X1 U13310 ( .A1(n11552), .A2(n11553), .ZN(n11632) );
  NAND2_X1 U13311 ( .A1(n11465), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n10933) );
  INV_X1 U13312 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n10927) );
  OR2_X1 U13313 ( .A1(n11466), .A2(n10927), .ZN(n10932) );
  OR2_X1 U13314 ( .A1(n11468), .A2(n10210), .ZN(n10931) );
  AND2_X1 U13315 ( .A1(n10928), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U13316 ( .A1(n10953), .A2(n10929), .ZN(n11917) );
  OR2_X1 U13317 ( .A1(n11400), .A2(n11917), .ZN(n10930) );
  NAND4_X1 U13318 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n14235) );
  OAI22_X1 U13319 ( .A1(n11454), .A2(n10935), .B1(n11348), .B2(n10934), .ZN(
        n10936) );
  INV_X1 U13320 ( .A(n10936), .ZN(n10939) );
  NAND2_X1 U13321 ( .A1(n14235), .A2(n11812), .ZN(n11557) );
  NAND2_X1 U13322 ( .A1(n11556), .A2(n11557), .ZN(n11633) );
  INV_X1 U13323 ( .A(n11633), .ZN(n11264) );
  XNOR2_X1 U13324 ( .A(n11265), .B(n11264), .ZN(n14252) );
  INV_X1 U13325 ( .A(n14252), .ZN(n10964) );
  NAND2_X1 U13326 ( .A1(n14819), .A2(n10940), .ZN(n10941) );
  NAND2_X1 U13327 ( .A1(n11543), .A2(n11544), .ZN(n11538) );
  NAND2_X1 U13328 ( .A1(n14809), .A2(n10943), .ZN(n10944) );
  NAND2_X1 U13329 ( .A1(n14821), .A2(n10944), .ZN(n14806) );
  NAND2_X1 U13330 ( .A1(n14806), .A2(n14814), .ZN(n10947) );
  NAND2_X1 U13331 ( .A1(n14237), .A2(n10945), .ZN(n10946) );
  NAND2_X1 U13332 ( .A1(n10947), .A2(n10946), .ZN(n14234) );
  AND2_X1 U13333 ( .A1(n14807), .A2(n11005), .ZN(n10948) );
  NAND2_X1 U13334 ( .A1(n10950), .A2(n11633), .ZN(n11662) );
  OAI211_X1 U13335 ( .C1(n10950), .C2(n11633), .A(n11662), .B(n14896), .ZN(
        n10960) );
  NAND2_X1 U13336 ( .A1(n11433), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n10958) );
  INV_X1 U13337 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n10951) );
  OR2_X1 U13338 ( .A1(n11466), .A2(n10951), .ZN(n10957) );
  OR2_X1 U13339 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  AND2_X1 U13340 ( .A1(n10954), .A2(n11278), .ZN(n12300) );
  OR2_X1 U13341 ( .A1(n11400), .A2(n12300), .ZN(n10956) );
  INV_X1 U13342 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12301) );
  OR2_X1 U13343 ( .A1(n11468), .A2(n12301), .ZN(n10955) );
  NAND4_X1 U13344 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n12282) );
  AOI22_X1 U13345 ( .A1(n14890), .A2(n14807), .B1(n12282), .B2(n14891), .ZN(
        n10959) );
  NAND2_X1 U13346 ( .A1(n10960), .A2(n10959), .ZN(n14250) );
  NAND2_X1 U13347 ( .A1(n14250), .A2(n14228), .ZN(n10963) );
  NOR2_X1 U13348 ( .A1(n11812), .A2(n14886), .ZN(n14251) );
  OAI22_X1 U13349 ( .A1(n14228), .A2(n10210), .B1(n11917), .B2(n14902), .ZN(
        n10961) );
  AOI21_X1 U13350 ( .B1(n14861), .B2(n14251), .A(n10961), .ZN(n10962) );
  OAI211_X1 U13351 ( .C1(n12305), .C2(n10964), .A(n10963), .B(n10962), .ZN(
        P3_U3221) );
  NAND2_X1 U13352 ( .A1(n10966), .A2(n10965), .ZN(n10968) );
  OR2_X1 U13353 ( .A1(n13499), .A2(n10973), .ZN(n10967) );
  NAND2_X1 U13354 ( .A1(n10968), .A2(n10967), .ZN(n11064) );
  NAND2_X1 U13355 ( .A1(n10969), .A2(n13595), .ZN(n10972) );
  AOI22_X1 U13356 ( .A1(n10970), .A2(n11102), .B1(n13594), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10971) );
  XNOR2_X1 U13357 ( .A(n14291), .B(n14016), .ZN(n13504) );
  XNOR2_X1 U13358 ( .A(n11064), .B(n13504), .ZN(n14321) );
  INV_X1 U13359 ( .A(n14321), .ZN(n10993) );
  NOR2_X1 U13360 ( .A1(n10975), .A2(n13504), .ZN(n14318) );
  INV_X1 U13361 ( .A(n11218), .ZN(n14317) );
  OR3_X1 U13362 ( .A1(n14318), .A2(n14317), .A3(n14025), .ZN(n10992) );
  NAND2_X1 U13363 ( .A1(n8606), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13364 ( .A1(n11209), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n10981) );
  INV_X1 U13365 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13366 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  AND2_X1 U13367 ( .A1(n11083), .A2(n10978), .ZN(n14019) );
  NAND2_X1 U13368 ( .A1(n11208), .A2(n14019), .ZN(n10980) );
  NAND2_X1 U13369 ( .A1(n13580), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10979) );
  OR2_X1 U13370 ( .A1(n14001), .A2(n14013), .ZN(n10984) );
  NAND2_X1 U13371 ( .A1(n13658), .A2(n14416), .ZN(n10983) );
  NAND2_X1 U13372 ( .A1(n10984), .A2(n10983), .ZN(n14293) );
  INV_X1 U13373 ( .A(n14293), .ZN(n14313) );
  AOI22_X1 U13374 ( .A1(n6479), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10985), 
        .B2(n14400), .ZN(n10986) );
  OAI21_X1 U13375 ( .B1(n14313), .B2(n6479), .A(n10986), .ZN(n10990) );
  AOI21_X1 U13376 ( .B1(n10987), .B2(n14291), .A(n14076), .ZN(n10988) );
  NAND2_X1 U13377 ( .A1(n10988), .A2(n14012), .ZN(n14314) );
  NOR2_X1 U13378 ( .A1(n14314), .A2(n14022), .ZN(n10989) );
  AOI211_X1 U13379 ( .C1(n14033), .C2(n14291), .A(n10990), .B(n10989), .ZN(
        n10991) );
  OAI211_X1 U13380 ( .C1(n10993), .C2(n13962), .A(n10992), .B(n10991), .ZN(
        P1_U3279) );
  OAI222_X1 U13381 ( .A1(n14166), .A2(n11156), .B1(n14165), .B2(n10995), .C1(
        P1_U3086), .C2(n10994), .ZN(P1_U3331) );
  INV_X1 U13382 ( .A(n10996), .ZN(n10997) );
  OR2_X1 U13383 ( .A1(n10997), .A2(n14818), .ZN(n10998) );
  NAND2_X1 U13384 ( .A1(n11809), .A2(n11810), .ZN(n11000) );
  XNOR2_X1 U13385 ( .A(n11000), .B(n11913), .ZN(n11007) );
  NOR2_X1 U13386 ( .A1(n14818), .A2(n12009), .ZN(n11001) );
  AOI211_X1 U13387 ( .C1(n12013), .C2(n14235), .A(n11002), .B(n11001), .ZN(
        n11003) );
  OAI21_X1 U13388 ( .B1(n12015), .B2(n14238), .A(n11003), .ZN(n11004) );
  AOI21_X1 U13389 ( .B1(n11005), .B2(n12017), .A(n11004), .ZN(n11006) );
  OAI21_X1 U13390 ( .B1(n11007), .B2(n12019), .A(n11006), .ZN(P3_U3176) );
  OAI21_X1 U13391 ( .B1(n11008), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n11010) );
  XNOR2_X1 U13392 ( .A(n11010), .B(n11009), .ZN(n14199) );
  MUX2_X1 U13393 ( .A(n11018), .B(n11021), .S(n12069), .Z(n11011) );
  XOR2_X1 U13394 ( .A(n14199), .B(n12047), .Z(n11015) );
  INV_X1 U13395 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12273) );
  INV_X1 U13396 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n11013) );
  MUX2_X1 U13397 ( .A(n12273), .B(n11013), .S(n12069), .Z(n11014) );
  NAND2_X1 U13398 ( .A1(n11015), .A2(n11014), .ZN(n12046) );
  OAI21_X1 U13399 ( .B1(n11015), .B2(n11014), .A(n12046), .ZN(n11016) );
  INV_X1 U13400 ( .A(n11016), .ZN(n11030) );
  NAND2_X1 U13401 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(n11019), .ZN(n12033) );
  OAI21_X1 U13402 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n11019), .A(n12033), 
        .ZN(n11028) );
  NAND2_X1 U13403 ( .A1(n12101), .A2(n6882), .ZN(n11026) );
  AND2_X1 U13404 ( .A1(n6473), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12012) );
  AOI21_X1 U13405 ( .B1(n14780), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12012), 
        .ZN(n11025) );
  NAND2_X1 U13406 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n11022), .ZN(n12038) );
  OAI21_X1 U13407 ( .B1(n11022), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12038), 
        .ZN(n11023) );
  NAND2_X1 U13408 ( .A1(n14788), .A2(n11023), .ZN(n11024) );
  NAND3_X1 U13409 ( .A1(n11026), .A2(n11025), .A3(n11024), .ZN(n11027) );
  AOI21_X1 U13410 ( .B1(n11028), .B2(n14801), .A(n11027), .ZN(n11029) );
  OAI21_X1 U13411 ( .B1(n11030), .B2(n12113), .A(n11029), .ZN(P3_U3197) );
  AND2_X1 U13412 ( .A1(n11032), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13413 ( .A1(n11032), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13414 ( .A1(n11032), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13415 ( .A1(n11032), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13416 ( .A1(n11032), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13417 ( .A1(n11032), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13418 ( .A1(n11032), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13419 ( .A1(n11032), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13420 ( .A1(n11032), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13421 ( .A1(n11032), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13422 ( .A1(n11032), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13423 ( .A1(n11032), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13424 ( .A1(n11032), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13425 ( .A1(n11032), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13426 ( .A1(n11032), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13427 ( .A1(n11032), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13428 ( .A1(n11032), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13429 ( .A1(n11032), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13430 ( .A1(n11032), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13431 ( .A1(n11032), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13432 ( .A1(n11032), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13433 ( .A1(n11032), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13434 ( .A1(n11032), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13435 ( .A1(n11032), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13436 ( .A1(n11032), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13437 ( .A1(n11032), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13438 ( .A1(n11032), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13439 ( .A1(n11032), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13440 ( .A1(n11032), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13441 ( .A1(n11032), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  OAI222_X1 U13442 ( .A1(P2_U3088), .A2(n11033), .B1(n13012), .B2(n11715), 
        .C1(n11447), .C2(n13010), .ZN(P2_U3297) );
  AOI22_X1 U13443 ( .A1(n9226), .A2(n13420), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n11034), .ZN(n11036) );
  NAND2_X1 U13444 ( .A1(n14300), .A2(n14032), .ZN(n11035) );
  OAI211_X1 U13445 ( .C1(n11037), .C2(n13425), .A(n11036), .B(n11035), .ZN(
        P1_U3232) );
  NOR2_X1 U13446 ( .A1(n13431), .A2(n14013), .ZN(n14035) );
  OR2_X1 U13447 ( .A1(n13596), .A2(n13990), .ZN(n14503) );
  NAND2_X1 U13448 ( .A1(n6938), .A2(n11038), .ZN(n13434) );
  AND2_X1 U13449 ( .A1(n13438), .A2(n13434), .ZN(n14029) );
  AOI21_X1 U13450 ( .B1(n14316), .B2(n14501), .A(n14029), .ZN(n11039) );
  AOI211_X1 U13451 ( .C1(n11040), .C2(n14032), .A(n14035), .B(n11039), .ZN(
        n14441) );
  NAND2_X1 U13452 ( .A1(n11044), .A2(n11042), .ZN(n11046) );
  AOI22_X1 U13453 ( .A1(n11046), .A2(n11045), .B1(n11044), .B2(n11043), .ZN(
        n11047) );
  NAND2_X1 U13454 ( .A1(n14532), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11050) );
  OAI21_X1 U13455 ( .B1(n14441), .B2(n14532), .A(n11050), .ZN(P1_U3528) );
  INV_X1 U13456 ( .A(n11051), .ZN(n11054) );
  MUX2_X1 U13457 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n8857), .S(n11059), .Z(
        n11053) );
  AOI211_X1 U13458 ( .C1(n11054), .C2(n11053), .A(n11052), .B(n13773), .ZN(
        n11062) );
  AOI211_X1 U13459 ( .C1(n11057), .C2(n11056), .A(n11055), .B(n13737), .ZN(
        n11061) );
  AOI22_X1 U13460 ( .A1(n13746), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n11058) );
  OAI21_X1 U13461 ( .B1(n11059), .B2(n13772), .A(n11058), .ZN(n11060) );
  OR4_X1 U13462 ( .A1(n11063), .A2(n11062), .A3(n11061), .A4(n11060), .ZN(
        P1_U3245) );
  NAND2_X1 U13463 ( .A1(n11064), .A2(n7255), .ZN(n11065) );
  OR2_X1 U13464 ( .A1(n14291), .A2(n14016), .ZN(n13505) );
  NAND2_X1 U13465 ( .A1(n11066), .A2(n13595), .ZN(n11068) );
  AOI22_X1 U13466 ( .A1(n13594), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11102), 
        .B2(n14384), .ZN(n11067) );
  NAND2_X1 U13467 ( .A1(n14307), .A2(n14001), .ZN(n13508) );
  NAND2_X1 U13468 ( .A1(n14011), .A2(n14024), .ZN(n11069) );
  NAND2_X1 U13469 ( .A1(n11070), .A2(n13595), .ZN(n11072) );
  AOI22_X1 U13470 ( .A1(n13594), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11102), 
        .B2(n13736), .ZN(n11071) );
  NAND2_X1 U13471 ( .A1(n13579), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13472 ( .A1(n8606), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11075) );
  XNOR2_X1 U13473 ( .A(n11083), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U13474 ( .A1(n11208), .A2(n14005), .ZN(n11074) );
  NAND2_X1 U13475 ( .A1(n13580), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11073) );
  XNOR2_X1 U13476 ( .A(n14132), .B(n13655), .ZN(n13626) );
  INV_X1 U13477 ( .A(n13626), .ZN(n13999) );
  OR2_X1 U13478 ( .A1(n14008), .A2(n13655), .ZN(n11077) );
  NAND2_X1 U13479 ( .A1(n11078), .A2(n13595), .ZN(n11080) );
  AOI22_X1 U13480 ( .A1(n13594), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11102), 
        .B2(n13752), .ZN(n11079) );
  NAND2_X1 U13481 ( .A1(n13580), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11088) );
  INV_X1 U13482 ( .A(n11083), .ZN(n11081) );
  AOI21_X1 U13483 ( .B1(n11081), .B2(P1_REG3_REG_16__SCAN_IN), .A(
        P1_REG3_REG_17__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U13484 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n11082) );
  OR2_X1 U13485 ( .A1(n11084), .A2(n11093), .ZN(n13364) );
  INV_X1 U13486 ( .A(n13364), .ZN(n13989) );
  NAND2_X1 U13487 ( .A1(n11208), .A2(n13989), .ZN(n11087) );
  NAND2_X1 U13488 ( .A1(n8606), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U13489 ( .A1(n13579), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U13490 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n13966) );
  OR2_X1 U13491 ( .A1(n14126), .A2(n13966), .ZN(n11219) );
  NAND2_X1 U13492 ( .A1(n14126), .A2(n13966), .ZN(n11220) );
  NAND2_X1 U13493 ( .A1(n11219), .A2(n11220), .ZN(n13977) );
  INV_X1 U13494 ( .A(n13977), .ZN(n13980) );
  INV_X1 U13495 ( .A(n13966), .ZN(n14002) );
  OR2_X1 U13496 ( .A1(n14126), .A2(n14002), .ZN(n11089) );
  NAND2_X1 U13497 ( .A1(n11090), .A2(n13595), .ZN(n11092) );
  AOI22_X1 U13498 ( .A1(n13594), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11102), 
        .B2(n13767), .ZN(n11091) );
  NAND2_X1 U13499 ( .A1(n11093), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11107) );
  OR2_X1 U13500 ( .A1(n11093), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11094) );
  AND2_X1 U13501 ( .A1(n11107), .A2(n11094), .ZN(n13971) );
  NAND2_X1 U13502 ( .A1(n11208), .A2(n13971), .ZN(n11098) );
  NAND2_X1 U13503 ( .A1(n13580), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13504 ( .A1(n13579), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U13505 ( .A1(n8606), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11095) );
  NAND4_X1 U13506 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n13654) );
  OR2_X1 U13507 ( .A1(n13972), .A2(n13654), .ZN(n11222) );
  NAND2_X1 U13508 ( .A1(n13972), .A2(n13654), .ZN(n11221) );
  NAND2_X1 U13509 ( .A1(n11222), .A2(n11221), .ZN(n13967) );
  NAND2_X1 U13510 ( .A1(n13963), .A2(n13967), .ZN(n11100) );
  INV_X1 U13511 ( .A(n13654), .ZN(n13982) );
  OR2_X1 U13512 ( .A1(n13972), .A2(n13982), .ZN(n11099) );
  NAND2_X1 U13513 ( .A1(n11100), .A2(n11099), .ZN(n13951) );
  NAND2_X1 U13514 ( .A1(n11101), .A2(n13595), .ZN(n11104) );
  AOI22_X1 U13515 ( .A1(n13594), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13928), 
        .B2(n11102), .ZN(n11103) );
  NAND2_X1 U13516 ( .A1(n13579), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11106) );
  NAND2_X1 U13517 ( .A1(n8606), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U13518 ( .A1(n11106), .A2(n11105), .ZN(n11110) );
  INV_X1 U13519 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U13520 ( .A1(n11107), .A2(n13130), .ZN(n11108) );
  NAND2_X1 U13521 ( .A1(n11116), .A2(n11108), .ZN(n13954) );
  INV_X1 U13522 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13765) );
  OAI22_X1 U13523 ( .A1(n13954), .A2(n11153), .B1(n11138), .B2(n13765), .ZN(
        n11109) );
  XNOR2_X1 U13524 ( .A(n14116), .B(n13965), .ZN(n13950) );
  INV_X1 U13525 ( .A(n13950), .ZN(n11112) );
  INV_X1 U13526 ( .A(n13965), .ZN(n13401) );
  NAND2_X1 U13527 ( .A1(n14116), .A2(n13401), .ZN(n11111) );
  NAND2_X1 U13528 ( .A1(n11113), .A2(n13595), .ZN(n11115) );
  OR2_X1 U13529 ( .A1(n13574), .A2(n10481), .ZN(n11114) );
  INV_X1 U13530 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U13531 ( .A1(n11116), .A2(n13379), .ZN(n11117) );
  NAND2_X1 U13532 ( .A1(n11125), .A2(n11117), .ZN(n13942) );
  AOI22_X1 U13533 ( .A1(n13579), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n8606), 
        .B2(P1_REG0_REG_20__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U13534 ( .A1(n9739), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11118) );
  OAI211_X1 U13535 ( .C1(n13942), .C2(n11153), .A(n11119), .B(n11118), .ZN(
        n13653) );
  INV_X1 U13536 ( .A(n13653), .ZN(n13531) );
  NAND2_X1 U13537 ( .A1(n14108), .A2(n13653), .ZN(n11120) );
  NAND2_X1 U13538 ( .A1(n11121), .A2(n13595), .ZN(n11123) );
  OR2_X1 U13539 ( .A1(n13574), .A2(n7231), .ZN(n11122) );
  INV_X1 U13540 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n11129) );
  INV_X1 U13541 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n11124) );
  AND2_X1 U13542 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  NOR2_X1 U13543 ( .A1(n11133), .A2(n11126), .ZN(n13926) );
  NAND2_X1 U13544 ( .A1(n13926), .A2(n11208), .ZN(n11128) );
  AOI22_X1 U13545 ( .A1(n8606), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n13580), 
        .B2(P1_REG1_REG_21__SCAN_IN), .ZN(n11127) );
  OAI211_X1 U13546 ( .C1(n9795), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n13652) );
  INV_X1 U13547 ( .A(n13652), .ZN(n13387) );
  XNOR2_X1 U13548 ( .A(n13923), .B(n13387), .ZN(n13921) );
  INV_X1 U13549 ( .A(n13921), .ZN(n13919) );
  NAND2_X1 U13550 ( .A1(n11130), .A2(n7672), .ZN(n11131) );
  XNOR2_X1 U13551 ( .A(n11131), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14173) );
  NOR2_X1 U13552 ( .A1(n11133), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11134) );
  OR2_X1 U13553 ( .A1(n11146), .A2(n11134), .ZN(n13911) );
  INV_X1 U13554 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U13555 ( .A1(n13579), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U13556 ( .A1(n8606), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11135) );
  OAI211_X1 U13557 ( .C1(n11138), .C2(n11137), .A(n11136), .B(n11135), .ZN(
        n11139) );
  INV_X1 U13558 ( .A(n11139), .ZN(n11140) );
  XNOR2_X1 U13559 ( .A(n13915), .B(n13651), .ZN(n13907) );
  INV_X1 U13560 ( .A(n13651), .ZN(n11228) );
  NAND2_X1 U13561 ( .A1(n14094), .A2(n11228), .ZN(n11141) );
  NAND2_X1 U13562 ( .A1(n11142), .A2(n13595), .ZN(n11145) );
  OR2_X1 U13563 ( .A1(n13574), .A2(n11143), .ZN(n11144) );
  OR2_X1 U13564 ( .A1(n11146), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U13565 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n11146), .ZN(n11160) );
  NAND2_X1 U13566 ( .A1(n11147), .A2(n11160), .ZN(n13893) );
  INV_X1 U13567 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U13568 ( .A1(n13579), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U13569 ( .A1(n9739), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11148) );
  OAI211_X1 U13570 ( .C1(n13584), .C2(n11150), .A(n11149), .B(n11148), .ZN(
        n11151) );
  INV_X1 U13571 ( .A(n11151), .ZN(n11152) );
  XNOR2_X1 U13572 ( .A(n14087), .B(n13388), .ZN(n13890) );
  INV_X1 U13573 ( .A(n13890), .ZN(n13898) );
  NAND2_X1 U13574 ( .A1(n13899), .A2(n13898), .ZN(n13897) );
  NAND2_X1 U13575 ( .A1(n14087), .A2(n13388), .ZN(n11154) );
  NAND2_X1 U13576 ( .A1(n11155), .A2(n13595), .ZN(n11158) );
  OR2_X1 U13577 ( .A1(n13574), .A2(n11156), .ZN(n11157) );
  INV_X1 U13578 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11161) );
  INV_X1 U13579 ( .A(n11160), .ZN(n11159) );
  NAND2_X1 U13580 ( .A1(n11159), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11170) );
  INV_X1 U13581 ( .A(n11170), .ZN(n11169) );
  AOI21_X1 U13582 ( .B1(n11161), .B2(n11160), .A(n11169), .ZN(n13882) );
  NAND2_X1 U13583 ( .A1(n11208), .A2(n13882), .ZN(n11165) );
  NAND2_X1 U13584 ( .A1(n9739), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U13585 ( .A1(n13579), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U13586 ( .A1(n8606), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11162) );
  NAND4_X1 U13587 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n13858) );
  XNOR2_X1 U13588 ( .A(n14083), .B(n13340), .ZN(n13871) );
  OR2_X1 U13589 ( .A1(n13340), .A2(n14083), .ZN(n11166) );
  NAND2_X1 U13590 ( .A1(n13009), .A2(n13595), .ZN(n11168) );
  OR2_X1 U13591 ( .A1(n13574), .A2(n14172), .ZN(n11167) );
  INV_X1 U13592 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13339) );
  NAND2_X1 U13593 ( .A1(n11169), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11179) );
  INV_X1 U13594 ( .A(n11179), .ZN(n11178) );
  AOI21_X1 U13595 ( .B1(n13339), .B2(n11170), .A(n11178), .ZN(n13338) );
  NAND2_X1 U13596 ( .A1(n11208), .A2(n13338), .ZN(n11174) );
  NAND2_X1 U13597 ( .A1(n9739), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U13598 ( .A1(n13579), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U13599 ( .A1(n8606), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11171) );
  NAND4_X1 U13600 ( .A1(n11174), .A2(n11173), .A3(n11172), .A4(n11171), .ZN(
        n13875) );
  NAND2_X1 U13601 ( .A1(n14074), .A2(n13875), .ZN(n11233) );
  OR2_X1 U13602 ( .A1(n14074), .A2(n13875), .ZN(n11175) );
  INV_X1 U13603 ( .A(n13875), .ZN(n13372) );
  NAND2_X1 U13604 ( .A1(n14074), .A2(n13372), .ZN(n13831) );
  NAND2_X1 U13605 ( .A1(n13005), .A2(n13595), .ZN(n11177) );
  OR2_X1 U13606 ( .A1(n13574), .A2(n7241), .ZN(n11176) );
  INV_X1 U13607 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U13608 ( .A1(n11178), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11189) );
  INV_X1 U13609 ( .A(n11189), .ZN(n11190) );
  AOI21_X1 U13610 ( .B1(n13408), .B2(n11179), .A(n11190), .ZN(n13842) );
  NAND2_X1 U13611 ( .A1(n11208), .A2(n13842), .ZN(n11183) );
  NAND2_X1 U13612 ( .A1(n9739), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U13613 ( .A1(n13579), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U13614 ( .A1(n8606), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11180) );
  NAND4_X1 U13615 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n13859) );
  INV_X1 U13616 ( .A(n13859), .ZN(n13341) );
  NAND2_X1 U13617 ( .A1(n13839), .A2(n13341), .ZN(n11186) );
  OR2_X1 U13618 ( .A1(n13839), .A2(n13341), .ZN(n11184) );
  NAND2_X1 U13619 ( .A1(n13001), .A2(n13595), .ZN(n11188) );
  OR2_X1 U13620 ( .A1(n13574), .A2(n14162), .ZN(n11187) );
  NAND2_X1 U13621 ( .A1(n9739), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11195) );
  INV_X1 U13622 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U13623 ( .A1(n13112), .A2(n11189), .ZN(n11191) );
  NAND2_X1 U13624 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n11190), .ZN(n11207) );
  NAND2_X1 U13625 ( .A1(n11208), .A2(n13825), .ZN(n11194) );
  NAND2_X1 U13626 ( .A1(n8606), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13627 ( .A1(n13579), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11192) );
  NAND4_X1 U13628 ( .A1(n11195), .A2(n11194), .A3(n11193), .A4(n11192), .ZN(
        n13835) );
  NAND2_X1 U13629 ( .A1(n14063), .A2(n13321), .ZN(n11197) );
  OR2_X1 U13630 ( .A1(n14063), .A2(n13321), .ZN(n11196) );
  NAND2_X1 U13631 ( .A1(n11246), .A2(n13595), .ZN(n11199) );
  OR2_X1 U13632 ( .A1(n13574), .A2(n11442), .ZN(n11198) );
  XNOR2_X1 U13633 ( .A(n11207), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U13634 ( .A1(n11208), .A2(n13318), .ZN(n11203) );
  NAND2_X1 U13635 ( .A1(n9739), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U13636 ( .A1(n8606), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U13637 ( .A1(n13579), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11200) );
  NAND4_X1 U13638 ( .A1(n11203), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n13798) );
  INV_X1 U13639 ( .A(n13798), .ZN(n11204) );
  NAND2_X1 U13640 ( .A1(n14058), .A2(n11204), .ZN(n13793) );
  OR2_X1 U13641 ( .A1(n14058), .A2(n11204), .ZN(n11205) );
  INV_X1 U13642 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13319) );
  NOR2_X1 U13643 ( .A1(n11207), .A2(n13319), .ZN(n13805) );
  NAND2_X1 U13644 ( .A1(n11208), .A2(n13805), .ZN(n11213) );
  NAND2_X1 U13645 ( .A1(n9739), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U13646 ( .A1(n11209), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U13647 ( .A1(n8606), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11210) );
  NAND4_X1 U13648 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n13650) );
  NAND2_X1 U13649 ( .A1(n13650), .A2(n14413), .ZN(n11215) );
  NAND2_X1 U13650 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  INV_X1 U13651 ( .A(n11219), .ZN(n13520) );
  INV_X1 U13652 ( .A(n11221), .ZN(n11223) );
  NAND2_X1 U13653 ( .A1(n11225), .A2(n11224), .ZN(n13933) );
  INV_X1 U13654 ( .A(n13939), .ZN(n11226) );
  OR2_X2 U13655 ( .A1(n13933), .A2(n11226), .ZN(n13934) );
  INV_X1 U13656 ( .A(n13923), .ZN(n14101) );
  NAND2_X1 U13657 ( .A1(n14101), .A2(n13387), .ZN(n11227) );
  NAND2_X1 U13658 ( .A1(n13896), .A2(n13388), .ZN(n11231) );
  NOR2_X1 U13659 ( .A1(n13896), .A2(n13388), .ZN(n11230) );
  INV_X1 U13660 ( .A(n14083), .ZN(n13884) );
  NAND2_X1 U13661 ( .A1(n13884), .A2(n13340), .ZN(n11232) );
  INV_X1 U13662 ( .A(n13852), .ZN(n13854) );
  INV_X1 U13663 ( .A(n13838), .ZN(n13832) );
  NAND2_X1 U13664 ( .A1(n13837), .A2(n13832), .ZN(n11235) );
  NAND2_X1 U13665 ( .A1(n13839), .A2(n13859), .ZN(n11234) );
  NAND2_X1 U13666 ( .A1(n11235), .A2(n11234), .ZN(n13816) );
  INV_X1 U13667 ( .A(n14063), .ZN(n13827) );
  NAND2_X1 U13668 ( .A1(n13827), .A2(n13321), .ZN(n11236) );
  INV_X1 U13669 ( .A(n13631), .ZN(n11237) );
  NAND2_X1 U13670 ( .A1(n11238), .A2(n13631), .ZN(n11239) );
  INV_X1 U13671 ( .A(n14058), .ZN(n11243) );
  INV_X1 U13672 ( .A(n14126), .ZN(n13979) );
  NAND2_X1 U13673 ( .A1(n14003), .A2(n13979), .ZN(n13986) );
  OR2_X2 U13674 ( .A1(n13972), .A2(n13986), .ZN(n13969) );
  INV_X1 U13675 ( .A(n14074), .ZN(n13855) );
  OR2_X1 U13676 ( .A1(n11243), .A2(n6527), .ZN(n11240) );
  AND3_X1 U13677 ( .A1(n13808), .A2(n11240), .A3(n14429), .ZN(n14057) );
  NAND2_X1 U13678 ( .A1(n14057), .A2(n14432), .ZN(n11242) );
  AOI22_X1 U13679 ( .A1(n6479), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13318), 
        .B2(n14400), .ZN(n11241) );
  OAI211_X1 U13680 ( .C1(n11243), .C2(n14422), .A(n11242), .B(n11241), .ZN(
        n11244) );
  AOI21_X1 U13681 ( .B1(n14056), .B2(n14433), .A(n11244), .ZN(n11245) );
  OAI21_X1 U13682 ( .B1(n6479), .B2(n14060), .A(n11245), .ZN(P1_U3265) );
  INV_X1 U13683 ( .A(n11246), .ZN(n13000) );
  OAI222_X1 U13684 ( .A1(n14166), .A2(n11442), .B1(n14165), .B2(n13000), .C1(
        P1_U3086), .C2(n6480), .ZN(P1_U3327) );
  NAND2_X1 U13685 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13002), .ZN(n11249) );
  NOR2_X1 U13686 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n7241), .ZN(n11248) );
  AOI22_X1 U13687 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11443), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11442), .ZN(n11250) );
  XNOR2_X1 U13688 ( .A(n11444), .B(n11250), .ZN(n12420) );
  NAND2_X1 U13689 ( .A1(n12420), .A2(n11453), .ZN(n11252) );
  OR2_X1 U13690 ( .A1(n11454), .A2(n12421), .ZN(n11251) );
  NAND2_X1 U13691 ( .A1(n11465), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n11259) );
  INV_X1 U13692 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n11253) );
  OR2_X1 U13693 ( .A1(n11466), .A2(n11253), .ZN(n11258) );
  NAND2_X1 U13694 ( .A1(n11254), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n11255) );
  OR2_X1 U13695 ( .A1(n11400), .A2(n12129), .ZN(n11257) );
  INV_X1 U13696 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12130) );
  OR2_X1 U13697 ( .A1(n11468), .A2(n12130), .ZN(n11256) );
  NAND2_X1 U13698 ( .A1(n12321), .A2(n11795), .ZN(n11483) );
  AOI22_X1 U13699 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13002), .B2(n14162), .ZN(n11260) );
  INV_X1 U13700 ( .A(SI_27_), .ZN(n11712) );
  NAND2_X1 U13701 ( .A1(n12325), .A2(n12124), .ZN(n12131) );
  AND2_X1 U13702 ( .A1(n11483), .A2(n12131), .ZN(n11481) );
  NAND2_X1 U13703 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  XNOR2_X1 U13704 ( .A(n11267), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n14188) );
  OAI22_X1 U13705 ( .A1(n11454), .A2(SI_13_), .B1(n11268), .B2(n11348), .ZN(
        n11269) );
  INV_X1 U13706 ( .A(n11269), .ZN(n11270) );
  NAND2_X1 U13707 ( .A1(n11271), .A2(n11270), .ZN(n11971) );
  OR2_X1 U13708 ( .A1(n11971), .A2(n12282), .ZN(n11562) );
  INV_X1 U13709 ( .A(n11562), .ZN(n11272) );
  NAND2_X1 U13710 ( .A1(n11971), .A2(n12282), .ZN(n11561) );
  XNOR2_X1 U13711 ( .A(n11273), .B(n6629), .ZN(n14194) );
  OAI22_X1 U13712 ( .A1(n11454), .A2(n7053), .B1(n11348), .B2(n14196), .ZN(
        n11274) );
  INV_X1 U13713 ( .A(n11274), .ZN(n11275) );
  NAND2_X1 U13714 ( .A1(n11276), .A2(n11275), .ZN(n12378) );
  NAND2_X1 U13715 ( .A1(n11433), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11283) );
  INV_X1 U13716 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11277) );
  OR2_X1 U13717 ( .A1(n11466), .A2(n11277), .ZN(n11282) );
  NAND2_X1 U13718 ( .A1(n11278), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11279) );
  AND2_X1 U13719 ( .A1(n11292), .A2(n11279), .ZN(n12286) );
  OR2_X1 U13720 ( .A1(n11400), .A2(n12286), .ZN(n11281) );
  INV_X1 U13721 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12287) );
  OR2_X1 U13722 ( .A1(n11468), .A2(n12287), .ZN(n11280) );
  OR2_X1 U13723 ( .A1(n12378), .A2(n12010), .ZN(n11567) );
  NAND2_X1 U13724 ( .A1(n12378), .A2(n12010), .ZN(n11566) );
  NAND2_X1 U13725 ( .A1(n11567), .A2(n11566), .ZN(n12290) );
  INV_X1 U13726 ( .A(n11284), .ZN(n11285) );
  XNOR2_X1 U13727 ( .A(n11286), .B(n11285), .ZN(n14197) );
  NAND2_X1 U13728 ( .A1(n14197), .A2(n11464), .ZN(n11290) );
  OAI22_X1 U13729 ( .A1(n11454), .A2(n11287), .B1(n11348), .B2(n14199), .ZN(
        n11288) );
  INV_X1 U13730 ( .A(n11288), .ZN(n11289) );
  NAND2_X1 U13731 ( .A1(n11465), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n11297) );
  INV_X1 U13732 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11291) );
  OR2_X1 U13733 ( .A1(n11466), .A2(n11291), .ZN(n11296) );
  AND2_X1 U13734 ( .A1(n11292), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n11293) );
  NOR2_X1 U13735 ( .A1(n11312), .A2(n11293), .ZN(n12272) );
  OR2_X1 U13736 ( .A1(n11400), .A2(n12272), .ZN(n11295) );
  OR2_X1 U13737 ( .A1(n11468), .A2(n12273), .ZN(n11294) );
  NAND4_X1 U13738 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n12283) );
  INV_X1 U13739 ( .A(n12283), .ZN(n11934) );
  OR2_X1 U13740 ( .A1(n12374), .A2(n11934), .ZN(n11570) );
  NAND2_X1 U13741 ( .A1(n12374), .A2(n11934), .ZN(n11575) );
  NAND2_X1 U13742 ( .A1(n12277), .A2(n12276), .ZN(n12275) );
  NAND2_X1 U13743 ( .A1(n12275), .A2(n11575), .ZN(n12265) );
  INV_X1 U13744 ( .A(n11298), .ZN(n11299) );
  XNOR2_X1 U13745 ( .A(n11300), .B(n11299), .ZN(n14200) );
  NAND2_X1 U13746 ( .A1(n14200), .A2(n11464), .ZN(n11310) );
  OR2_X1 U13747 ( .A1(n11302), .A2(n11301), .ZN(n11304) );
  MUX2_X1 U13748 ( .A(n11304), .B(P3_IR_REG_31__SCAN_IN), .S(n11303), .Z(
        n11306) );
  NAND2_X1 U13749 ( .A1(n11306), .A2(n11305), .ZN(n14202) );
  OAI22_X1 U13750 ( .A1(n11454), .A2(n11307), .B1(n11348), .B2(n14202), .ZN(
        n11308) );
  INV_X1 U13751 ( .A(n11308), .ZN(n11309) );
  NAND2_X1 U13752 ( .A1(n11310), .A2(n11309), .ZN(n12370) );
  NAND2_X1 U13753 ( .A1(n11465), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n11317) );
  INV_X1 U13754 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n11311) );
  OR2_X1 U13755 ( .A1(n11466), .A2(n11311), .ZN(n11316) );
  NOR2_X1 U13756 ( .A1(n11312), .A2(n11933), .ZN(n11313) );
  OR2_X1 U13757 ( .A1(n11400), .A2(n6519), .ZN(n11315) );
  INV_X1 U13758 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12262) );
  OR2_X1 U13759 ( .A1(n11468), .A2(n12262), .ZN(n11314) );
  OR2_X1 U13760 ( .A1(n12370), .A2(n11929), .ZN(n11577) );
  NAND2_X1 U13761 ( .A1(n12370), .A2(n11929), .ZN(n11576) );
  NAND2_X1 U13762 ( .A1(n11577), .A2(n11576), .ZN(n11666) );
  OAI22_X1 U13763 ( .A1(n11454), .A2(n11318), .B1(n11348), .B2(n12084), .ZN(
        n11319) );
  AOI21_X1 U13764 ( .B1(n11320), .B2(n11464), .A(n11319), .ZN(n12253) );
  NAND2_X1 U13765 ( .A1(n11433), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n11327) );
  INV_X1 U13766 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n11321) );
  OR2_X1 U13767 ( .A1(n11466), .A2(n11321), .ZN(n11326) );
  NOR2_X1 U13768 ( .A1(n11322), .A2(n13126), .ZN(n11323) );
  NOR2_X1 U13769 ( .A1(n11341), .A2(n11323), .ZN(n12254) );
  OR2_X1 U13770 ( .A1(n11400), .A2(n12254), .ZN(n11325) );
  INV_X1 U13771 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12255) );
  OR2_X1 U13772 ( .A1(n11468), .A2(n12255), .ZN(n11324) );
  NAND4_X1 U13773 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n12260) );
  NAND2_X1 U13774 ( .A1(n12253), .A2(n12260), .ZN(n11489) );
  INV_X1 U13775 ( .A(n12253), .ZN(n12366) );
  INV_X1 U13776 ( .A(n12260), .ZN(n11328) );
  NAND2_X1 U13777 ( .A1(n12366), .A2(n11328), .ZN(n11496) );
  NAND2_X1 U13778 ( .A1(n11489), .A2(n11496), .ZN(n11669) );
  INV_X1 U13779 ( .A(n11329), .ZN(n11330) );
  XNOR2_X1 U13780 ( .A(n11331), .B(n11330), .ZN(n14206) );
  NAND2_X1 U13781 ( .A1(n14206), .A2(n11464), .ZN(n11338) );
  INV_X1 U13782 ( .A(SI_18_), .ZN(n11335) );
  NAND2_X1 U13783 ( .A1(n11332), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n11334) );
  INV_X1 U13784 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n11333) );
  XNOR2_X1 U13785 ( .A(n11334), .B(n11333), .ZN(n14208) );
  OAI22_X1 U13786 ( .A1(n11454), .A2(n11335), .B1(n11348), .B2(n14208), .ZN(
        n11336) );
  INV_X1 U13787 ( .A(n11336), .ZN(n11337) );
  NAND2_X1 U13788 ( .A1(n11465), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n11346) );
  INV_X1 U13789 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n11339) );
  OR2_X1 U13790 ( .A1(n11466), .A2(n11339), .ZN(n11345) );
  OR2_X1 U13791 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  AND2_X1 U13792 ( .A1(n11342), .A2(n11353), .ZN(n12240) );
  OR2_X1 U13793 ( .A1(n12240), .A2(n11400), .ZN(n11344) );
  INV_X1 U13794 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13209) );
  OR2_X1 U13795 ( .A1(n11468), .A2(n13209), .ZN(n11343) );
  NAND2_X1 U13796 ( .A1(n12362), .A2(n12224), .ZN(n11491) );
  NAND2_X1 U13797 ( .A1(n11347), .A2(n11464), .ZN(n11351) );
  OAI22_X1 U13798 ( .A1(n11454), .A2(SI_19_), .B1(n12100), .B2(n11348), .ZN(
        n11349) );
  INV_X1 U13799 ( .A(n11349), .ZN(n11350) );
  NAND2_X1 U13800 ( .A1(n11351), .A2(n11350), .ZN(n11888) );
  NAND2_X1 U13801 ( .A1(n11465), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n11358) );
  INV_X1 U13802 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n11352) );
  OR2_X1 U13803 ( .A1(n11466), .A2(n11352), .ZN(n11357) );
  AND2_X1 U13804 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n11353), .ZN(n11354) );
  NOR2_X1 U13805 ( .A1(n11365), .A2(n11354), .ZN(n12229) );
  OR2_X1 U13806 ( .A1(n11400), .A2(n12229), .ZN(n11356) );
  INV_X1 U13807 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12230) );
  OR2_X1 U13808 ( .A1(n11468), .A2(n12230), .ZN(n11355) );
  NAND4_X1 U13809 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n12238) );
  NAND2_X1 U13810 ( .A1(n11888), .A2(n12238), .ZN(n11621) );
  INV_X1 U13811 ( .A(n11621), .ZN(n11359) );
  OR2_X1 U13812 ( .A1(n11888), .A2(n12238), .ZN(n11622) );
  NAND2_X1 U13813 ( .A1(n11360), .A2(n11464), .ZN(n11363) );
  NAND2_X1 U13814 ( .A1(n11433), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n11370) );
  INV_X1 U13815 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n11364) );
  OR2_X1 U13816 ( .A1(n11466), .A2(n11364), .ZN(n11369) );
  OR2_X1 U13817 ( .A1(n11365), .A2(n11960), .ZN(n11366) );
  AND2_X1 U13818 ( .A1(n11366), .A2(n11376), .ZN(n12215) );
  OR2_X1 U13819 ( .A1(n11400), .A2(n12215), .ZN(n11368) );
  INV_X1 U13820 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12216) );
  OR2_X1 U13821 ( .A1(n11468), .A2(n12216), .ZN(n11367) );
  NAND4_X1 U13822 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n12025) );
  XNOR2_X1 U13823 ( .A(n12354), .B(n12025), .ZN(n12218) );
  INV_X1 U13824 ( .A(n12218), .ZN(n11674) );
  INV_X1 U13825 ( .A(n12354), .ZN(n11966) );
  NAND2_X1 U13826 ( .A1(n11966), .A2(n12025), .ZN(n11488) );
  NAND2_X1 U13827 ( .A1(n12217), .A2(n11488), .ZN(n12200) );
  OR2_X1 U13828 ( .A1(n11454), .A2(n11372), .ZN(n11373) );
  NAND2_X1 U13829 ( .A1(n11465), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n11381) );
  INV_X1 U13830 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n11375) );
  OR2_X1 U13831 ( .A1(n11466), .A2(n11375), .ZN(n11380) );
  NAND2_X1 U13832 ( .A1(n11376), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n11377) );
  AND2_X1 U13833 ( .A1(n11387), .A2(n11377), .ZN(n12207) );
  OR2_X1 U13834 ( .A1(n11400), .A2(n12207), .ZN(n11379) );
  INV_X1 U13835 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12208) );
  OR2_X1 U13836 ( .A1(n11468), .A2(n12208), .ZN(n11378) );
  NAND2_X1 U13837 ( .A1(n12351), .A2(n11961), .ZN(n11588) );
  NAND2_X1 U13838 ( .A1(n11465), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n11392) );
  INV_X1 U13839 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n11386) );
  OR2_X1 U13840 ( .A1(n11466), .A2(n11386), .ZN(n11391) );
  INV_X1 U13841 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12194) );
  OR2_X1 U13842 ( .A1(n11468), .A2(n12194), .ZN(n11390) );
  AND2_X1 U13843 ( .A1(n11387), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11388) );
  NOR2_X1 U13844 ( .A1(n11398), .A2(n11388), .ZN(n12193) );
  OR2_X1 U13845 ( .A1(n11400), .A2(n12193), .ZN(n11389) );
  NAND4_X1 U13846 ( .A1(n11392), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(
        n12178) );
  NAND2_X1 U13847 ( .A1(n12346), .A2(n12206), .ZN(n11485) );
  OR2_X1 U13848 ( .A1(n11454), .A2(n11394), .ZN(n11395) );
  NAND2_X1 U13849 ( .A1(n11465), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n11404) );
  INV_X1 U13850 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n11397) );
  OR2_X1 U13851 ( .A1(n11466), .A2(n11397), .ZN(n11403) );
  NOR2_X1 U13852 ( .A1(n11398), .A2(n11875), .ZN(n11399) );
  NOR2_X1 U13853 ( .A1(n11411), .A2(n11399), .ZN(n12183) );
  OR2_X1 U13854 ( .A1(n11400), .A2(n12183), .ZN(n11402) );
  INV_X1 U13855 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12184) );
  OR2_X1 U13856 ( .A1(n11468), .A2(n12184), .ZN(n11401) );
  NAND2_X1 U13857 ( .A1(n11845), .A2(n12191), .ZN(n12164) );
  NAND2_X1 U13858 ( .A1(n12341), .A2(n12156), .ZN(n11405) );
  NAND2_X1 U13859 ( .A1(n12164), .A2(n11405), .ZN(n11678) );
  OR2_X1 U13860 ( .A1(n11454), .A2(n11407), .ZN(n11408) );
  NAND2_X1 U13861 ( .A1(n11433), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n11416) );
  INV_X1 U13862 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n11410) );
  OR2_X1 U13863 ( .A1(n11466), .A2(n11410), .ZN(n11415) );
  OR2_X1 U13864 ( .A1(n11411), .A2(n11952), .ZN(n11412) );
  AND2_X1 U13865 ( .A1(n11422), .A2(n11412), .ZN(n12159) );
  OR2_X1 U13866 ( .A1(n9825), .A2(n12159), .ZN(n11414) );
  INV_X1 U13867 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12160) );
  OR2_X1 U13868 ( .A1(n11468), .A2(n12160), .ZN(n11413) );
  NAND4_X1 U13869 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n12177) );
  XNOR2_X1 U13870 ( .A(n12337), .B(n12177), .ZN(n12163) );
  AND2_X1 U13871 ( .A1(n12163), .A2(n12164), .ZN(n11599) );
  NAND2_X1 U13872 ( .A1(n11433), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n11427) );
  INV_X1 U13873 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n11421) );
  OR2_X1 U13874 ( .A1(n11466), .A2(n11421), .ZN(n11426) );
  NAND2_X1 U13875 ( .A1(n11422), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n11423) );
  AND2_X1 U13876 ( .A1(n11435), .A2(n11423), .ZN(n12145) );
  OR2_X1 U13877 ( .A1(n9825), .A2(n12145), .ZN(n11425) );
  INV_X1 U13878 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12146) );
  OR2_X1 U13879 ( .A1(n11468), .A2(n12146), .ZN(n11424) );
  NAND2_X1 U13880 ( .A1(n12333), .A2(n12155), .ZN(n11600) );
  NAND2_X1 U13881 ( .A1(n12337), .A2(n12140), .ZN(n12147) );
  NAND2_X1 U13882 ( .A1(n11429), .A2(n11464), .ZN(n11432) );
  NAND2_X1 U13883 ( .A1(n11465), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n11441) );
  INV_X1 U13884 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n11434) );
  OR2_X1 U13885 ( .A1(n11466), .A2(n11434), .ZN(n11440) );
  AND2_X1 U13886 ( .A1(n11435), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11436) );
  NOR2_X1 U13887 ( .A1(n11437), .A2(n11436), .ZN(n12002) );
  OR2_X1 U13888 ( .A1(n9825), .A2(n12002), .ZN(n11439) );
  INV_X1 U13889 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n11689) );
  OR2_X1 U13890 ( .A1(n11468), .A2(n11689), .ZN(n11438) );
  NOR2_X1 U13891 ( .A1(n12329), .A2(n12141), .ZN(n11612) );
  NAND2_X1 U13892 ( .A1(n12329), .A2(n12141), .ZN(n11602) );
  OR2_X1 U13893 ( .A1(n12325), .A2(n12124), .ZN(n11608) );
  INV_X1 U13894 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14160) );
  INV_X1 U13895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U13896 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14160), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n12995), .ZN(n11449) );
  NOR2_X1 U13897 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n11442), .ZN(n11445) );
  OAI22_X1 U13898 ( .A1(n11445), .A2(n11444), .B1(P2_DATAO_REG_28__SCAN_IN), 
        .B2(n11443), .ZN(n11448) );
  XOR2_X1 U13899 ( .A(n11449), .B(n11448), .Z(n12416) );
  NOR2_X1 U13900 ( .A1(n11454), .A2(n12417), .ZN(n11446) );
  AOI21_X1 U13901 ( .B1(n12416), .B2(n11464), .A(n11446), .ZN(n11475) );
  NAND2_X1 U13902 ( .A1(n11475), .A2(n11897), .ZN(n11620) );
  INV_X1 U13903 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13573) );
  OAI22_X1 U13904 ( .A1(n13573), .A2(n11447), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U13905 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14160), .B1(n11449), 
        .B2(n11448), .ZN(n11462) );
  INV_X1 U13906 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U13907 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n11451), .B2(n11450), .ZN(n11452) );
  INV_X1 U13908 ( .A(SI_31_), .ZN(n12408) );
  OR2_X1 U13909 ( .A1(n11454), .A2(n12408), .ZN(n11455) );
  NAND2_X1 U13910 ( .A1(n11456), .A2(n11455), .ZN(n14245) );
  NAND2_X1 U13911 ( .A1(n11465), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11460) );
  INV_X1 U13912 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11457) );
  OR2_X1 U13913 ( .A1(n11466), .A2(n11457), .ZN(n11459) );
  INV_X1 U13914 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n14227) );
  OR2_X1 U13915 ( .A1(n11468), .A2(n14227), .ZN(n11458) );
  NAND4_X1 U13916 ( .A1(n11472), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n14225) );
  INV_X1 U13917 ( .A(n14225), .ZN(n11477) );
  XNOR2_X1 U13918 ( .A(n11462), .B(n11461), .ZN(n12413) );
  INV_X1 U13919 ( .A(SI_30_), .ZN(n12414) );
  NOR2_X1 U13920 ( .A1(n11454), .A2(n12414), .ZN(n11463) );
  AOI21_X1 U13921 ( .B1(n12413), .B2(n11464), .A(n11463), .ZN(n11478) );
  INV_X1 U13922 ( .A(n11478), .ZN(n14248) );
  NAND2_X1 U13923 ( .A1(n11465), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n11471) );
  INV_X1 U13924 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14260) );
  OR2_X1 U13925 ( .A1(n11466), .A2(n14260), .ZN(n11470) );
  INV_X1 U13926 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n11467) );
  OR2_X1 U13927 ( .A1(n11468), .A2(n11467), .ZN(n11469) );
  NAND4_X1 U13928 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n12021) );
  INV_X1 U13929 ( .A(n12021), .ZN(n11473) );
  NAND2_X1 U13930 ( .A1(n14248), .A2(n11473), .ZN(n11474) );
  OAI21_X1 U13931 ( .B1(n14245), .B2(n11477), .A(n11474), .ZN(n11647) );
  INV_X1 U13932 ( .A(n11475), .ZN(n11805) );
  INV_X1 U13933 ( .A(n11897), .ZN(n12125) );
  NAND2_X1 U13934 ( .A1(n11805), .A2(n12125), .ZN(n11619) );
  OAI21_X1 U13935 ( .B1(n11478), .B2(n14225), .A(n11619), .ZN(n11476) );
  AND2_X1 U13936 ( .A1(n11478), .A2(n12021), .ZN(n11646) );
  INV_X1 U13937 ( .A(n11481), .ZN(n11482) );
  OAI21_X1 U13938 ( .B1(n11482), .B2(n12310), .A(n11484), .ZN(n11614) );
  NOR2_X1 U13939 ( .A1(n12023), .A2(n11613), .ZN(n11607) );
  XNOR2_X1 U13940 ( .A(n12147), .B(n11613), .ZN(n11598) );
  MUX2_X1 U13941 ( .A(n11486), .B(n11485), .S(n12310), .Z(n11593) );
  NAND2_X1 U13942 ( .A1(n11486), .A2(n11485), .ZN(n12189) );
  INV_X1 U13943 ( .A(n12189), .ZN(n12195) );
  INV_X1 U13944 ( .A(n12025), .ZN(n12225) );
  NAND2_X1 U13945 ( .A1(n12354), .A2(n12225), .ZN(n11487) );
  MUX2_X1 U13946 ( .A(n11488), .B(n11487), .S(n12310), .Z(n11587) );
  NAND3_X1 U13947 ( .A1(n11622), .A2(n11491), .A3(n12310), .ZN(n11495) );
  INV_X1 U13948 ( .A(n11489), .ZN(n11490) );
  NAND2_X1 U13949 ( .A1(n11491), .A2(n11490), .ZN(n11493) );
  AND3_X1 U13950 ( .A1(n11493), .A2(n11613), .A3(n11492), .ZN(n11494) );
  NAND2_X1 U13951 ( .A1(n11494), .A2(n11621), .ZN(n11498) );
  AND2_X1 U13952 ( .A1(n11495), .A2(n11498), .ZN(n11585) );
  INV_X1 U13953 ( .A(n11496), .ZN(n11497) );
  NAND2_X1 U13954 ( .A1(n11498), .A2(n11497), .ZN(n11582) );
  AOI21_X1 U13955 ( .B1(n11503), .B2(n11656), .A(n11499), .ZN(n11500) );
  NOR2_X1 U13956 ( .A1(n11500), .A2(n14888), .ZN(n11502) );
  MUX2_X1 U13957 ( .A(n11613), .B(n11502), .S(n11501), .Z(n11515) );
  INV_X1 U13958 ( .A(n14894), .ZN(n11505) );
  INV_X1 U13959 ( .A(n11503), .ZN(n11504) );
  NAND3_X1 U13960 ( .A1(n11505), .A2(n11613), .A3(n11504), .ZN(n11506) );
  OAI211_X1 U13961 ( .C1(n11613), .C2(n11507), .A(n11506), .B(n7410), .ZN(
        n11514) );
  NAND2_X1 U13962 ( .A1(n11508), .A2(n14847), .ZN(n11511) );
  NAND2_X1 U13963 ( .A1(n11516), .A2(n11509), .ZN(n11510) );
  MUX2_X1 U13964 ( .A(n11511), .B(n11510), .S(n11613), .Z(n11512) );
  INV_X1 U13965 ( .A(n11512), .ZN(n11513) );
  OAI21_X1 U13966 ( .B1(n11515), .B2(n11514), .A(n11513), .ZN(n11519) );
  MUX2_X1 U13967 ( .A(n11516), .B(n14847), .S(n11613), .Z(n11517) );
  NAND3_X1 U13968 ( .A1(n11519), .A2(n11518), .A3(n11517), .ZN(n11523) );
  MUX2_X1 U13969 ( .A(n11521), .B(n11520), .S(n12310), .Z(n11522) );
  NAND3_X1 U13970 ( .A1(n11523), .A2(n11623), .A3(n11522), .ZN(n11527) );
  NAND2_X1 U13971 ( .A1(n11524), .A2(n11532), .ZN(n11525) );
  NAND2_X1 U13972 ( .A1(n11525), .A2(n11613), .ZN(n11526) );
  NAND2_X1 U13973 ( .A1(n11527), .A2(n11526), .ZN(n11531) );
  AOI21_X1 U13974 ( .B1(n11530), .B2(n11528), .A(n11613), .ZN(n11529) );
  AOI21_X1 U13975 ( .B1(n11531), .B2(n11530), .A(n11529), .ZN(n11537) );
  OAI21_X1 U13976 ( .B1(n11613), .B2(n11532), .A(n11625), .ZN(n11536) );
  MUX2_X1 U13977 ( .A(n11534), .B(n11533), .S(n11613), .Z(n11535) );
  OAI211_X1 U13978 ( .C1(n11537), .C2(n11536), .A(n11624), .B(n11535), .ZN(
        n11542) );
  MUX2_X1 U13979 ( .A(n11540), .B(n11539), .S(n12310), .Z(n11541) );
  NAND3_X1 U13980 ( .A1(n11542), .A2(n14826), .A3(n11541), .ZN(n11546) );
  MUX2_X1 U13981 ( .A(n11544), .B(n11543), .S(n11613), .Z(n11545) );
  NAND2_X1 U13982 ( .A1(n11546), .A2(n11545), .ZN(n11551) );
  MUX2_X1 U13983 ( .A(n11548), .B(n11547), .S(n11613), .Z(n11549) );
  NAND2_X1 U13984 ( .A1(n10926), .A2(n11549), .ZN(n11550) );
  AOI21_X1 U13985 ( .B1(n11551), .B2(n10920), .A(n11550), .ZN(n11560) );
  NAND2_X1 U13986 ( .A1(n11552), .A2(n11556), .ZN(n11555) );
  NAND2_X1 U13987 ( .A1(n11557), .A2(n11553), .ZN(n11554) );
  MUX2_X1 U13988 ( .A(n11555), .B(n11554), .S(n11613), .Z(n11559) );
  NAND2_X1 U13989 ( .A1(n11562), .A2(n11561), .ZN(n12295) );
  INV_X1 U13990 ( .A(n12295), .ZN(n11636) );
  MUX2_X1 U13991 ( .A(n11557), .B(n11556), .S(n11613), .Z(n11558) );
  OAI211_X1 U13992 ( .C1(n11560), .C2(n11559), .A(n11636), .B(n11558), .ZN(
        n11564) );
  MUX2_X1 U13993 ( .A(n11562), .B(n11561), .S(n11613), .Z(n11563) );
  NAND2_X1 U13994 ( .A1(n11564), .A2(n11563), .ZN(n11565) );
  INV_X1 U13995 ( .A(n12290), .ZN(n11637) );
  NAND2_X1 U13996 ( .A1(n11565), .A2(n11637), .ZN(n11569) );
  MUX2_X1 U13997 ( .A(n11567), .B(n11566), .S(n12310), .Z(n11568) );
  NAND3_X1 U13998 ( .A1(n11569), .A2(n12276), .A3(n11568), .ZN(n11574) );
  NAND2_X1 U13999 ( .A1(n11577), .A2(n11570), .ZN(n11571) );
  NAND2_X1 U14000 ( .A1(n11571), .A2(n12310), .ZN(n11573) );
  INV_X1 U14001 ( .A(n11576), .ZN(n11572) );
  AOI21_X1 U14002 ( .B1(n11574), .B2(n11573), .A(n11572), .ZN(n11579) );
  AOI21_X1 U14003 ( .B1(n11576), .B2(n11575), .A(n12310), .ZN(n11578) );
  OAI22_X1 U14004 ( .A1(n11579), .A2(n11578), .B1(n11577), .B2(n12310), .ZN(
        n11580) );
  NAND2_X1 U14005 ( .A1(n11580), .A2(n12250), .ZN(n11581) );
  AOI21_X1 U14006 ( .B1(n11582), .B2(n11581), .A(n12237), .ZN(n11584) );
  MUX2_X1 U14007 ( .A(n11622), .B(n11621), .S(n12310), .Z(n11583) );
  OAI211_X1 U14008 ( .C1(n11585), .C2(n11584), .A(n12218), .B(n11583), .ZN(
        n11586) );
  NAND3_X1 U14009 ( .A1(n11587), .A2(n11586), .A3(n12204), .ZN(n11591) );
  MUX2_X1 U14010 ( .A(n11589), .B(n11588), .S(n11613), .Z(n11590) );
  NAND3_X1 U14011 ( .A1(n12195), .A2(n11591), .A3(n11590), .ZN(n11592) );
  NAND3_X1 U14012 ( .A1(n11593), .A2(n12174), .A3(n11592), .ZN(n11595) );
  NAND3_X1 U14013 ( .A1(n12341), .A2(n12156), .A3(n11613), .ZN(n11594) );
  NAND2_X1 U14014 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  NAND2_X1 U14015 ( .A1(n12163), .A2(n11596), .ZN(n11597) );
  OAI211_X1 U14016 ( .C1(n11599), .C2(n11598), .A(n12138), .B(n11597), .ZN(
        n11605) );
  MUX2_X1 U14017 ( .A(n11601), .B(n11600), .S(n12310), .Z(n11604) );
  INV_X1 U14018 ( .A(n11602), .ZN(n11603) );
  AOI21_X1 U14019 ( .B1(n11605), .B2(n11604), .A(n11683), .ZN(n11606) );
  AOI21_X1 U14020 ( .B1(n11607), .B2(n12329), .A(n11606), .ZN(n11610) );
  INV_X1 U14021 ( .A(n11701), .ZN(n11696) );
  INV_X1 U14022 ( .A(n11608), .ZN(n11609) );
  AOI22_X1 U14023 ( .A1(n11610), .A2(n11696), .B1(n11609), .B2(n12310), .ZN(
        n11611) );
  INV_X1 U14024 ( .A(n11620), .ZN(n11615) );
  AOI211_X1 U14025 ( .C1(n11616), .C2(n11619), .A(n11646), .B(n11615), .ZN(
        n11618) );
  OAI21_X1 U14026 ( .B1(n11618), .B2(n11647), .A(n11645), .ZN(n11652) );
  INV_X1 U14027 ( .A(n11652), .ZN(n11651) );
  INV_X1 U14028 ( .A(n12232), .ZN(n11640) );
  INV_X1 U14029 ( .A(n12276), .ZN(n11639) );
  NAND4_X1 U14030 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11628) );
  NOR4_X1 U14031 ( .A1(n11628), .A2(n14852), .A3(n11627), .A4(n14894), .ZN(
        n11631) );
  NAND4_X1 U14032 ( .A1(n11631), .A2(n14826), .A3(n11630), .A4(n11629), .ZN(
        n11634) );
  NOR4_X1 U14033 ( .A1(n11634), .A2(n11633), .A3(n14814), .A4(n11632), .ZN(
        n11635) );
  NAND4_X1 U14034 ( .A1(n12250), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11638) );
  NOR4_X1 U14035 ( .A1(n11640), .A2(n11666), .A3(n11639), .A4(n11638), .ZN(
        n11641) );
  NAND4_X1 U14036 ( .A1(n12204), .A2(n12218), .A3(n12242), .A4(n11641), .ZN(
        n11642) );
  NOR4_X1 U14037 ( .A1(n11678), .A2(n12189), .A3(n11683), .A4(n11642), .ZN(
        n11643) );
  AND4_X1 U14038 ( .A1(n12138), .A2(n11696), .A3(n11643), .A4(n12163), .ZN(
        n11644) );
  XNOR2_X1 U14039 ( .A(n11648), .B(n12100), .ZN(n11649) );
  OAI22_X1 U14040 ( .A1(n11651), .A2(n14901), .B1(n11650), .B2(n11649), .ZN(
        n11654) );
  INV_X1 U14041 ( .A(P3_B_REG_SCAN_IN), .ZN(n11799) );
  AOI21_X1 U14042 ( .B1(n11657), .B2(n11656), .A(n11799), .ZN(n11658) );
  OAI21_X1 U14043 ( .B1(n11659), .B2(n12092), .A(n11658), .ZN(n11660) );
  INV_X1 U14044 ( .A(n11812), .ZN(n11919) );
  NAND2_X1 U14045 ( .A1(n14235), .A2(n11919), .ZN(n11661) );
  NAND2_X1 U14046 ( .A1(n11662), .A2(n11661), .ZN(n12296) );
  NAND2_X1 U14047 ( .A1(n12296), .A2(n12295), .ZN(n12294) );
  INV_X1 U14048 ( .A(n12282), .ZN(n11967) );
  OR2_X1 U14049 ( .A1(n11971), .A2(n11967), .ZN(n11663) );
  NAND2_X1 U14050 ( .A1(n12294), .A2(n11663), .ZN(n12281) );
  NAND2_X1 U14051 ( .A1(n12378), .A2(n12297), .ZN(n11664) );
  OR2_X1 U14052 ( .A1(n12374), .A2(n12283), .ZN(n11665) );
  NAND2_X1 U14053 ( .A1(n12259), .A2(n11666), .ZN(n11668) );
  NAND2_X1 U14054 ( .A1(n12370), .A2(n12270), .ZN(n11667) );
  NAND2_X1 U14055 ( .A1(n11668), .A2(n11667), .ZN(n12246) );
  NAND2_X1 U14056 ( .A1(n12246), .A2(n11669), .ZN(n11671) );
  NAND2_X1 U14057 ( .A1(n12366), .A2(n12260), .ZN(n11670) );
  OR2_X1 U14058 ( .A1(n12362), .A2(n12247), .ZN(n11672) );
  INV_X1 U14059 ( .A(n11888), .ZN(n12358) );
  NAND2_X1 U14060 ( .A1(n12358), .A2(n12238), .ZN(n11673) );
  NAND2_X1 U14061 ( .A1(n12227), .A2(n11673), .ZN(n12212) );
  NAND2_X1 U14062 ( .A1(n12354), .A2(n12025), .ZN(n11675) );
  OR2_X1 U14063 ( .A1(n12351), .A2(n12213), .ZN(n12188) );
  INV_X1 U14064 ( .A(n12346), .ZN(n11676) );
  NAND2_X1 U14065 ( .A1(n11676), .A2(n12206), .ZN(n11677) );
  AND2_X1 U14066 ( .A1(n12188), .A2(n11677), .ZN(n12170) );
  AND2_X1 U14067 ( .A1(n12170), .A2(n11678), .ZN(n11679) );
  NAND2_X1 U14068 ( .A1(n12346), .A2(n12178), .ZN(n12171) );
  NAND2_X1 U14069 ( .A1(n12341), .A2(n12191), .ZN(n11680) );
  NAND2_X1 U14070 ( .A1(n12181), .A2(n11680), .ZN(n12153) );
  INV_X1 U14071 ( .A(n12163), .ZN(n11681) );
  NAND2_X1 U14072 ( .A1(n12337), .A2(n12177), .ZN(n11789) );
  NAND2_X1 U14073 ( .A1(n12333), .A2(n12024), .ZN(n11695) );
  NAND2_X1 U14074 ( .A1(n12143), .A2(n11695), .ZN(n11682) );
  XNOR2_X1 U14075 ( .A(n11682), .B(n11683), .ZN(n11687) );
  XNOR2_X1 U14076 ( .A(n11684), .B(n11683), .ZN(n12330) );
  OAI22_X1 U14077 ( .A1(n12155), .A2(n14869), .B1(n12124), .B2(n14867), .ZN(
        n11685) );
  OAI22_X1 U14078 ( .A1(n14228), .A2(n11689), .B1(n12002), .B2(n14902), .ZN(
        n11690) );
  AOI21_X1 U14079 ( .B1(n12329), .B2(n14231), .A(n11690), .ZN(n11692) );
  NAND2_X1 U14080 ( .A1(n12330), .A2(n11708), .ZN(n11691) );
  OAI211_X1 U14081 ( .C1(n12332), .C2(n14908), .A(n11692), .B(n11691), .ZN(
        P3_U3207) );
  OAI21_X1 U14082 ( .B1(n11693), .B2(n11696), .A(n12132), .ZN(n12326) );
  OAI22_X1 U14083 ( .A1(n12141), .A2(n14869), .B1(n11795), .B2(n14867), .ZN(
        n11705) );
  NAND2_X1 U14084 ( .A1(n12329), .A2(n12023), .ZN(n11694) );
  AND2_X1 U14085 ( .A1(n11695), .A2(n11694), .ZN(n11702) );
  AND2_X1 U14086 ( .A1(n12143), .A2(n11702), .ZN(n11698) );
  OR2_X1 U14087 ( .A1(n12329), .A2(n12023), .ZN(n11699) );
  NAND2_X1 U14088 ( .A1(n11699), .A2(n11696), .ZN(n11697) );
  AND2_X1 U14089 ( .A1(n12148), .A2(n11700), .ZN(n11793) );
  NAND2_X1 U14090 ( .A1(n12137), .A2(n11793), .ZN(n11703) );
  NAND2_X1 U14091 ( .A1(n11703), .A2(n11787), .ZN(n11704) );
  OAI22_X1 U14092 ( .A1(n14228), .A2(n11706), .B1(n11859), .B2(n14902), .ZN(
        n11707) );
  AOI21_X1 U14093 ( .B1(n12325), .B2(n14231), .A(n11707), .ZN(n11710) );
  NAND2_X1 U14094 ( .A1(n12326), .A2(n11708), .ZN(n11709) );
  OAI211_X1 U14095 ( .C1(n12328), .C2(n14908), .A(n11710), .B(n11709), .ZN(
        P3_U3206) );
  INV_X1 U14096 ( .A(n11711), .ZN(n11713) );
  OAI222_X1 U14097 ( .A1(n6473), .A2(n12069), .B1(n12423), .B2(n11713), .C1(
        n11712), .C2(n14186), .ZN(P3_U3268) );
  OAI222_X1 U14098 ( .A1(n14165), .A2(n11715), .B1(n11714), .B2(P1_U3086), 
        .C1(n13573), .C2(n14166), .ZN(P1_U3325) );
  XNOR2_X1 U14099 ( .A(n12946), .B(n11762), .ZN(n11736) );
  NAND2_X1 U14100 ( .A1(n12817), .A2(n6488), .ZN(n11737) );
  NOR2_X1 U14101 ( .A1(n12525), .A2(n12885), .ZN(n11733) );
  XNOR2_X1 U14102 ( .A(n12837), .B(n11762), .ZN(n11730) );
  NOR2_X1 U14103 ( .A1(n12498), .A2(n12885), .ZN(n11722) );
  XNOR2_X1 U14104 ( .A(n12495), .B(n11762), .ZN(n11721) );
  INV_X1 U14105 ( .A(n11721), .ZN(n12500) );
  XNOR2_X1 U14106 ( .A(n11721), .B(n11722), .ZN(n12487) );
  OAI21_X1 U14107 ( .B1(n11722), .B2(n12500), .A(n12486), .ZN(n11723) );
  XNOR2_X1 U14108 ( .A(n12966), .B(n11762), .ZN(n11726) );
  NAND2_X1 U14109 ( .A1(n12881), .A2(n6488), .ZN(n11724) );
  XNOR2_X1 U14110 ( .A(n11726), .B(n11724), .ZN(n12501) );
  INV_X1 U14111 ( .A(n11724), .ZN(n11725) );
  XNOR2_X1 U14112 ( .A(n12853), .B(n11743), .ZN(n12441) );
  NOR2_X1 U14113 ( .A1(n12443), .A2(n12885), .ZN(n11728) );
  NAND2_X1 U14114 ( .A1(n12441), .A2(n11728), .ZN(n11731) );
  OAI21_X1 U14115 ( .B1(n12441), .B2(n11728), .A(n11731), .ZN(n12549) );
  INV_X1 U14116 ( .A(n12549), .ZN(n11729) );
  XNOR2_X1 U14117 ( .A(n11730), .B(n11733), .ZN(n12450) );
  XNOR2_X1 U14118 ( .A(n12951), .B(n11762), .ZN(n12523) );
  AND2_X1 U14119 ( .A1(n12802), .A2(n6487), .ZN(n11735) );
  NOR2_X1 U14120 ( .A1(n12523), .A2(n11735), .ZN(n11734) );
  NAND2_X1 U14121 ( .A1(n12523), .A2(n11735), .ZN(n12520) );
  XNOR2_X1 U14122 ( .A(n11736), .B(n11737), .ZN(n12463) );
  XNOR2_X1 U14123 ( .A(n12796), .B(n11762), .ZN(n11739) );
  AND2_X1 U14124 ( .A1(n6968), .A2(n6488), .ZN(n11738) );
  INV_X1 U14125 ( .A(n11739), .ZN(n11740) );
  NAND2_X1 U14126 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  XNOR2_X1 U14127 ( .A(n12783), .B(n11743), .ZN(n11744) );
  XNOR2_X1 U14128 ( .A(n12766), .B(n11743), .ZN(n11747) );
  AND2_X1 U14129 ( .A1(n6488), .A2(n12746), .ZN(n11748) );
  NAND2_X1 U14130 ( .A1(n11747), .A2(n11748), .ZN(n12472) );
  NAND2_X1 U14131 ( .A1(n11745), .A2(n11744), .ZN(n12470) );
  NAND3_X1 U14132 ( .A1(n12471), .A2(n12472), .A3(n12470), .ZN(n11751) );
  XNOR2_X1 U14133 ( .A(n12926), .B(n11762), .ZN(n12562) );
  AND2_X1 U14134 ( .A1(n6488), .A2(n12758), .ZN(n11746) );
  NAND2_X1 U14135 ( .A1(n12562), .A2(n11746), .ZN(n11752) );
  OAI21_X1 U14136 ( .B1(n12562), .B2(n11746), .A(n11752), .ZN(n12475) );
  INV_X1 U14137 ( .A(n11747), .ZN(n12477) );
  INV_X1 U14138 ( .A(n11748), .ZN(n11749) );
  NOR2_X1 U14139 ( .A1(n12475), .A2(n12473), .ZN(n11750) );
  XNOR2_X1 U14140 ( .A(n12734), .B(n9262), .ZN(n11756) );
  NAND2_X1 U14141 ( .A1(n6487), .A2(n12747), .ZN(n11755) );
  XNOR2_X1 U14142 ( .A(n11756), .B(n11755), .ZN(n12564) );
  INV_X1 U14143 ( .A(n11752), .ZN(n11753) );
  NOR2_X1 U14144 ( .A1(n12564), .A2(n11753), .ZN(n11754) );
  NAND2_X1 U14145 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  XNOR2_X1 U14146 ( .A(n12915), .B(n11762), .ZN(n11759) );
  AND2_X1 U14147 ( .A1(n6488), .A2(n12576), .ZN(n11758) );
  NAND2_X1 U14148 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  OAI21_X1 U14149 ( .B1(n11759), .B2(n11758), .A(n11760), .ZN(n12426) );
  NAND2_X1 U14150 ( .A1(n6488), .A2(n12575), .ZN(n11761) );
  XNOR2_X1 U14151 ( .A(n11762), .B(n11761), .ZN(n11763) );
  XNOR2_X1 U14152 ( .A(n12909), .B(n11763), .ZN(n11764) );
  XNOR2_X1 U14153 ( .A(n11765), .B(n11764), .ZN(n11771) );
  INV_X1 U14154 ( .A(n11766), .ZN(n12699) );
  OAI22_X1 U14155 ( .A1(n11767), .A2(n12777), .B1(n12773), .B2(n12729), .ZN(
        n12696) );
  AOI22_X1 U14156 ( .A1(n12444), .A2(n12696), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11768) );
  OAI21_X1 U14157 ( .B1(n12699), .B2(n12538), .A(n11768), .ZN(n11769) );
  AOI21_X1 U14158 ( .B1(n12909), .B2(n12569), .A(n11769), .ZN(n11770) );
  OAI21_X1 U14159 ( .B1(n11771), .B2(n12571), .A(n11770), .ZN(P2_U3192) );
  INV_X1 U14160 ( .A(n11772), .ZN(n11773) );
  AOI22_X1 U14161 ( .A1(n11773), .A2(n12533), .B1(n12563), .B2(n12883), .ZN(
        n11781) );
  NOR2_X1 U14162 ( .A1(n12538), .A2(n11774), .ZN(n11778) );
  OAI22_X1 U14163 ( .A1(n12429), .A2(n11776), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11775), .ZN(n11777) );
  AOI211_X1 U14164 ( .C1(n11779), .C2(n12569), .A(n11778), .B(n11777), .ZN(
        n11780) );
  OAI21_X1 U14165 ( .B1(n11782), .B2(n11781), .A(n11780), .ZN(P2_U3213) );
  INV_X1 U14166 ( .A(n11783), .ZN(n11784) );
  OAI222_X1 U14167 ( .A1(n13010), .A2(n11785), .B1(n13012), .B2(n11784), .C1(
        P2_U3088), .C2(n6489), .ZN(P2_U3305) );
  INV_X1 U14168 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n11807) );
  OR2_X1 U14169 ( .A1(n12325), .A2(n11998), .ZN(n11792) );
  INV_X1 U14170 ( .A(n11787), .ZN(n11788) );
  AND2_X1 U14171 ( .A1(n11789), .A2(n11791), .ZN(n11790) );
  INV_X1 U14172 ( .A(n12133), .ZN(n11794) );
  INV_X1 U14173 ( .A(n11795), .ZN(n12022) );
  NAND2_X1 U14174 ( .A1(n12321), .A2(n12022), .ZN(n11796) );
  NAND2_X1 U14175 ( .A1(n12127), .A2(n11796), .ZN(n11797) );
  XNOR2_X1 U14176 ( .A(n11797), .B(n11803), .ZN(n11798) );
  NAND2_X1 U14177 ( .A1(n11798), .A2(n14896), .ZN(n11802) );
  NOR2_X1 U14178 ( .A1(n12424), .A2(n11799), .ZN(n11800) );
  NOR2_X1 U14179 ( .A1(n14867), .A2(n11800), .ZN(n14224) );
  AOI22_X1 U14180 ( .A1(n14224), .A2(n12021), .B1(n12022), .B2(n14890), .ZN(
        n11801) );
  NAND2_X1 U14181 ( .A1(n11802), .A2(n11801), .ZN(n12115) );
  NAND2_X1 U14182 ( .A1(n11805), .A2(n14916), .ZN(n12118) );
  INV_X1 U14183 ( .A(n11808), .ZN(P3_U3456) );
  XNOR2_X1 U14184 ( .A(n12325), .B(n11892), .ZN(n11889) );
  XNOR2_X1 U14185 ( .A(n11889), .B(n11998), .ZN(n11890) );
  NAND2_X1 U14186 ( .A1(n11809), .A2(n14807), .ZN(n11811) );
  XNOR2_X1 U14187 ( .A(n11812), .B(n6828), .ZN(n11814) );
  XNOR2_X1 U14188 ( .A(n11814), .B(n14235), .ZN(n11912) );
  INV_X1 U14189 ( .A(n11814), .ZN(n11816) );
  INV_X1 U14190 ( .A(n14235), .ZN(n11815) );
  NAND2_X1 U14191 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  XNOR2_X1 U14192 ( .A(n11971), .B(n11892), .ZN(n11968) );
  AND2_X1 U14193 ( .A1(n11968), .A2(n11967), .ZN(n11818) );
  XNOR2_X1 U14194 ( .A(n12378), .B(n6828), .ZN(n11819) );
  XNOR2_X1 U14195 ( .A(n11819), .B(n12297), .ZN(n11863) );
  NAND2_X1 U14196 ( .A1(n11864), .A2(n11863), .ZN(n11822) );
  INV_X1 U14197 ( .A(n11819), .ZN(n11820) );
  NAND2_X1 U14198 ( .A1(n11820), .A2(n12297), .ZN(n11821) );
  NAND2_X1 U14199 ( .A1(n11822), .A2(n11821), .ZN(n12008) );
  XNOR2_X1 U14200 ( .A(n12374), .B(n6828), .ZN(n11823) );
  XNOR2_X1 U14201 ( .A(n11823), .B(n12283), .ZN(n12007) );
  NAND2_X1 U14202 ( .A1(n12008), .A2(n12007), .ZN(n11826) );
  INV_X1 U14203 ( .A(n11823), .ZN(n11824) );
  NAND2_X1 U14204 ( .A1(n11824), .A2(n12283), .ZN(n11825) );
  XNOR2_X1 U14205 ( .A(n12370), .B(n11892), .ZN(n11930) );
  AND2_X1 U14206 ( .A1(n11930), .A2(n12270), .ZN(n11827) );
  INV_X1 U14207 ( .A(n11930), .ZN(n11828) );
  NAND2_X1 U14208 ( .A1(n11828), .A2(n11929), .ZN(n11829) );
  XNOR2_X1 U14209 ( .A(n12253), .B(n6828), .ZN(n11832) );
  XNOR2_X1 U14210 ( .A(n11832), .B(n12260), .ZN(n11940) );
  NAND2_X1 U14211 ( .A1(n11831), .A2(n11830), .ZN(n11942) );
  NAND2_X1 U14212 ( .A1(n11832), .A2(n12260), .ZN(n11833) );
  NAND2_X1 U14213 ( .A1(n11942), .A2(n11833), .ZN(n11987) );
  XNOR2_X1 U14214 ( .A(n12362), .B(n6828), .ZN(n11834) );
  XNOR2_X1 U14215 ( .A(n11834), .B(n12247), .ZN(n11986) );
  NAND2_X1 U14216 ( .A1(n11987), .A2(n11986), .ZN(n11985) );
  INV_X1 U14217 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U14218 ( .A1(n11835), .A2(n12247), .ZN(n11836) );
  NAND2_X1 U14219 ( .A1(n11985), .A2(n11836), .ZN(n11883) );
  XNOR2_X1 U14220 ( .A(n11888), .B(n11892), .ZN(n11837) );
  XNOR2_X1 U14221 ( .A(n11837), .B(n12238), .ZN(n11882) );
  NAND2_X1 U14222 ( .A1(n11883), .A2(n11882), .ZN(n11881) );
  INV_X1 U14223 ( .A(n11837), .ZN(n11838) );
  NAND2_X1 U14224 ( .A1(n11838), .A2(n12238), .ZN(n11839) );
  XNOR2_X1 U14225 ( .A(n12354), .B(n6828), .ZN(n11840) );
  XNOR2_X1 U14226 ( .A(n11840), .B(n12025), .ZN(n11958) );
  INV_X1 U14227 ( .A(n11840), .ZN(n11841) );
  NAND2_X1 U14228 ( .A1(n11841), .A2(n12025), .ZN(n11842) );
  XNOR2_X1 U14229 ( .A(n12351), .B(n6828), .ZN(n11843) );
  XNOR2_X1 U14230 ( .A(n11843), .B(n11961), .ZN(n11903) );
  XNOR2_X1 U14231 ( .A(n12346), .B(n11892), .ZN(n11871) );
  XNOR2_X1 U14232 ( .A(n12337), .B(n6828), .ZN(n11951) );
  XNOR2_X1 U14233 ( .A(n11845), .B(n6828), .ZN(n11949) );
  INV_X1 U14234 ( .A(n11949), .ZN(n11846) );
  OAI22_X1 U14235 ( .A1(n11951), .A2(n12140), .B1(n12156), .B2(n11846), .ZN(
        n11851) );
  AOI21_X1 U14236 ( .B1(n11871), .B2(n12178), .A(n11851), .ZN(n11853) );
  OR2_X1 U14237 ( .A1(n11871), .A2(n12178), .ZN(n11850) );
  NAND3_X1 U14238 ( .A1(n11846), .A2(n12156), .A3(n12140), .ZN(n11849) );
  OAI21_X1 U14239 ( .B1(n11949), .B2(n12191), .A(n12177), .ZN(n11847) );
  NAND2_X1 U14240 ( .A1(n11951), .A2(n11847), .ZN(n11848) );
  OAI211_X1 U14241 ( .C1(n11851), .C2(n11850), .A(n11849), .B(n11848), .ZN(
        n11852) );
  XNOR2_X1 U14242 ( .A(n12333), .B(n11892), .ZN(n11854) );
  XNOR2_X1 U14243 ( .A(n11854), .B(n12024), .ZN(n11923) );
  XNOR2_X1 U14244 ( .A(n12329), .B(n11892), .ZN(n11855) );
  XNOR2_X1 U14245 ( .A(n11855), .B(n12141), .ZN(n11997) );
  INV_X1 U14246 ( .A(n11855), .ZN(n11856) );
  XOR2_X1 U14247 ( .A(n11890), .B(n11891), .Z(n11862) );
  AOI22_X1 U14248 ( .A1(n11999), .A2(n12023), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(n6473), .ZN(n11858) );
  NAND2_X1 U14249 ( .A1(n12022), .A2(n12013), .ZN(n11857) );
  OAI211_X1 U14250 ( .C1(n12003), .C2(n11859), .A(n11858), .B(n11857), .ZN(
        n11860) );
  AOI21_X1 U14251 ( .B1(n12325), .B2(n12017), .A(n11860), .ZN(n11861) );
  OAI21_X1 U14252 ( .B1(n11862), .B2(n12019), .A(n11861), .ZN(P3_U3154) );
  XNOR2_X1 U14253 ( .A(n11864), .B(n11863), .ZN(n11870) );
  NOR2_X1 U14254 ( .A1(n11934), .A2(n11988), .ZN(n11865) );
  AOI211_X1 U14255 ( .C1(n11999), .C2(n12282), .A(n11866), .B(n11865), .ZN(
        n11867) );
  OAI21_X1 U14256 ( .B1(n12003), .B2(n12286), .A(n11867), .ZN(n11868) );
  AOI21_X1 U14257 ( .B1(n12378), .B2(n12017), .A(n11868), .ZN(n11869) );
  OAI21_X1 U14258 ( .B1(n11870), .B2(n12019), .A(n11869), .ZN(P3_U3155) );
  INV_X1 U14259 ( .A(n11871), .ZN(n11872) );
  AND2_X1 U14260 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  XNOR2_X1 U14261 ( .A(n11950), .B(n12156), .ZN(n11880) );
  OAI22_X1 U14262 ( .A1(n12140), .A2(n11988), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11875), .ZN(n11876) );
  AOI21_X1 U14263 ( .B1(n11999), .B2(n12178), .A(n11876), .ZN(n11877) );
  OAI21_X1 U14264 ( .B1(n12003), .B2(n12183), .A(n11877), .ZN(n11878) );
  AOI21_X1 U14265 ( .B1(n12341), .B2(n12017), .A(n11878), .ZN(n11879) );
  OAI21_X1 U14266 ( .B1(n11880), .B2(n12019), .A(n11879), .ZN(P3_U3156) );
  OAI211_X1 U14267 ( .C1(n11883), .C2(n11882), .A(n11881), .B(n11984), .ZN(
        n11887) );
  NAND2_X1 U14268 ( .A1(n6473), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12102) );
  OAI21_X1 U14269 ( .B1(n12225), .B2(n11988), .A(n12102), .ZN(n11885) );
  NOR2_X1 U14270 ( .A1(n12015), .A2(n12229), .ZN(n11884) );
  AOI211_X1 U14271 ( .C1(n11999), .C2(n12247), .A(n11885), .B(n11884), .ZN(
        n11886) );
  OAI211_X1 U14272 ( .C1(n11994), .C2(n11888), .A(n11887), .B(n11886), .ZN(
        P3_U3159) );
  OAI22_X1 U14273 ( .A1(n11891), .A2(n11890), .B1(n11889), .B2(n11998), .ZN(
        n11894) );
  XNOR2_X1 U14274 ( .A(n12133), .B(n11892), .ZN(n11893) );
  XNOR2_X1 U14275 ( .A(n11894), .B(n11893), .ZN(n11901) );
  OAI22_X1 U14276 ( .A1(n12124), .A2(n12009), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11895), .ZN(n11896) );
  AOI21_X1 U14277 ( .B1(n12013), .B2(n11897), .A(n11896), .ZN(n11898) );
  OAI21_X1 U14278 ( .B1(n12015), .B2(n12129), .A(n11898), .ZN(n11899) );
  AOI21_X1 U14279 ( .B1(n12321), .B2(n12017), .A(n11899), .ZN(n11900) );
  OAI21_X1 U14280 ( .B1(n11901), .B2(n12019), .A(n11900), .ZN(P3_U3160) );
  AOI21_X1 U14281 ( .B1(n11903), .B2(n11902), .A(n6562), .ZN(n11908) );
  AOI22_X1 U14282 ( .A1(n12013), .A2(n12178), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11905) );
  NAND2_X1 U14283 ( .A1(n11999), .A2(n12025), .ZN(n11904) );
  OAI211_X1 U14284 ( .C1(n12003), .C2(n12207), .A(n11905), .B(n11904), .ZN(
        n11906) );
  AOI21_X1 U14285 ( .B1(n12351), .B2(n12017), .A(n11906), .ZN(n11907) );
  OAI21_X1 U14286 ( .B1(n11908), .B2(n12019), .A(n11907), .ZN(P3_U3163) );
  INV_X1 U14287 ( .A(n11909), .ZN(n11910) );
  AOI21_X1 U14288 ( .B1(n11912), .B2(n11911), .A(n11910), .ZN(n11921) );
  NOR2_X1 U14289 ( .A1(n11913), .A2(n12009), .ZN(n11914) );
  AOI211_X1 U14290 ( .C1(n12013), .C2(n12282), .A(n11915), .B(n11914), .ZN(
        n11916) );
  OAI21_X1 U14291 ( .B1(n12015), .B2(n11917), .A(n11916), .ZN(n11918) );
  AOI21_X1 U14292 ( .B1(n11919), .B2(n12017), .A(n11918), .ZN(n11920) );
  OAI21_X1 U14293 ( .B1(n11921), .B2(n12019), .A(n11920), .ZN(P3_U3164) );
  XOR2_X1 U14294 ( .A(n11923), .B(n11922), .Z(n11928) );
  AOI22_X1 U14295 ( .A1(n12013), .A2(n12023), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11925) );
  NAND2_X1 U14296 ( .A1(n11999), .A2(n12177), .ZN(n11924) );
  OAI211_X1 U14297 ( .C1(n12003), .C2(n12145), .A(n11925), .B(n11924), .ZN(
        n11926) );
  AOI21_X1 U14298 ( .B1(n12333), .B2(n12017), .A(n11926), .ZN(n11927) );
  OAI21_X1 U14299 ( .B1(n11928), .B2(n12019), .A(n11927), .ZN(P3_U3165) );
  XNOR2_X1 U14300 ( .A(n11930), .B(n11929), .ZN(n11931) );
  XNOR2_X1 U14301 ( .A(n11932), .B(n11931), .ZN(n11939) );
  NOR2_X1 U14302 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11933), .ZN(n12043) );
  NOR2_X1 U14303 ( .A1(n11934), .A2(n12009), .ZN(n11935) );
  AOI211_X1 U14304 ( .C1(n12013), .C2(n12260), .A(n12043), .B(n11935), .ZN(
        n11936) );
  OAI21_X1 U14305 ( .B1(n12015), .B2(n6519), .A(n11936), .ZN(n11937) );
  AOI21_X1 U14306 ( .B1(n12370), .B2(n12017), .A(n11937), .ZN(n11938) );
  OAI21_X1 U14307 ( .B1(n11939), .B2(n12019), .A(n11938), .ZN(P3_U3166) );
  AOI21_X1 U14308 ( .B1(n11941), .B2(n11940), .A(n12019), .ZN(n11943) );
  NAND2_X1 U14309 ( .A1(n11943), .A2(n11942), .ZN(n11947) );
  NAND2_X1 U14310 ( .A1(n6473), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12059) );
  OAI21_X1 U14311 ( .B1(n12224), .B2(n11988), .A(n12059), .ZN(n11945) );
  NOR2_X1 U14312 ( .A1(n12015), .A2(n12254), .ZN(n11944) );
  AOI211_X1 U14313 ( .C1(n11999), .C2(n12270), .A(n11945), .B(n11944), .ZN(
        n11946) );
  OAI211_X1 U14314 ( .C1(n12253), .C2(n11994), .A(n11947), .B(n11946), .ZN(
        P3_U3168) );
  OAI22_X1 U14315 ( .A1(n12155), .A2(n11988), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11952), .ZN(n11953) );
  AOI21_X1 U14316 ( .B1(n11999), .B2(n12191), .A(n11953), .ZN(n11954) );
  OAI21_X1 U14317 ( .B1(n12015), .B2(n12159), .A(n11954), .ZN(n11955) );
  AOI21_X1 U14318 ( .B1(n12337), .B2(n12017), .A(n11955), .ZN(n11956) );
  OAI211_X1 U14319 ( .C1(n11959), .C2(n11958), .A(n11957), .B(n11984), .ZN(
        n11965) );
  OAI22_X1 U14320 ( .A1(n11961), .A2(n11988), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11960), .ZN(n11963) );
  NOR2_X1 U14321 ( .A1(n12003), .A2(n12215), .ZN(n11962) );
  AOI211_X1 U14322 ( .C1(n11999), .C2(n12238), .A(n11963), .B(n11962), .ZN(
        n11964) );
  OAI211_X1 U14323 ( .C1(n11966), .C2(n11994), .A(n11965), .B(n11964), .ZN(
        P3_U3173) );
  XNOR2_X1 U14324 ( .A(n11968), .B(n11967), .ZN(n11969) );
  XNOR2_X1 U14325 ( .A(n11970), .B(n11969), .ZN(n11977) );
  INV_X1 U14326 ( .A(n11971), .ZN(n12383) );
  NOR2_X1 U14327 ( .A1(n12010), .A2(n11988), .ZN(n11972) );
  AOI211_X1 U14328 ( .C1(n11999), .C2(n14235), .A(n11973), .B(n11972), .ZN(
        n11974) );
  OAI21_X1 U14329 ( .B1(n12015), .B2(n12300), .A(n11974), .ZN(n11975) );
  AOI21_X1 U14330 ( .B1(n12383), .B2(n12017), .A(n11975), .ZN(n11976) );
  OAI21_X1 U14331 ( .B1(n11977), .B2(n12019), .A(n11976), .ZN(P3_U3174) );
  XNOR2_X1 U14332 ( .A(n11978), .B(n12178), .ZN(n11983) );
  AOI22_X1 U14333 ( .A1(n12013), .A2(n12191), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(n6473), .ZN(n11980) );
  NAND2_X1 U14334 ( .A1(n12213), .A2(n11999), .ZN(n11979) );
  OAI211_X1 U14335 ( .C1(n12003), .C2(n12193), .A(n11980), .B(n11979), .ZN(
        n11981) );
  AOI21_X1 U14336 ( .B1(n12346), .B2(n12017), .A(n11981), .ZN(n11982) );
  OAI21_X1 U14337 ( .B1(n11983), .B2(n12019), .A(n11982), .ZN(P3_U3175) );
  INV_X1 U14338 ( .A(n12362), .ZN(n11995) );
  OAI211_X1 U14339 ( .C1(n11987), .C2(n11986), .A(n11985), .B(n11984), .ZN(
        n11993) );
  INV_X1 U14340 ( .A(n12238), .ZN(n11989) );
  NAND2_X1 U14341 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12080)
         );
  OAI21_X1 U14342 ( .B1(n11989), .B2(n11988), .A(n12080), .ZN(n11991) );
  NOR2_X1 U14343 ( .A1(n12003), .A2(n12240), .ZN(n11990) );
  AOI211_X1 U14344 ( .C1(n11999), .C2(n12260), .A(n11991), .B(n11990), .ZN(
        n11992) );
  OAI211_X1 U14345 ( .C1(n11995), .C2(n11994), .A(n11993), .B(n11992), .ZN(
        P3_U3178) );
  XOR2_X1 U14346 ( .A(n11997), .B(n11996), .Z(n12006) );
  AOI22_X1 U14347 ( .A1(n11998), .A2(n12013), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12001) );
  NAND2_X1 U14348 ( .A1(n12024), .A2(n11999), .ZN(n12000) );
  OAI211_X1 U14349 ( .C1(n12003), .C2(n12002), .A(n12001), .B(n12000), .ZN(
        n12004) );
  AOI21_X1 U14350 ( .B1(n12329), .B2(n12017), .A(n12004), .ZN(n12005) );
  OAI21_X1 U14351 ( .B1(n12006), .B2(n12019), .A(n12005), .ZN(P3_U3180) );
  XNOR2_X1 U14352 ( .A(n12008), .B(n12007), .ZN(n12020) );
  NOR2_X1 U14353 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  AOI211_X1 U14354 ( .C1(n12013), .C2(n12270), .A(n12012), .B(n12011), .ZN(
        n12014) );
  OAI21_X1 U14355 ( .B1(n12015), .B2(n12272), .A(n12014), .ZN(n12016) );
  AOI21_X1 U14356 ( .B1(n12374), .B2(n12017), .A(n12016), .ZN(n12018) );
  OAI21_X1 U14357 ( .B1(n12020), .B2(n12019), .A(n12018), .ZN(P3_U3181) );
  MUX2_X1 U14358 ( .A(n14225), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12031), .Z(
        P3_U3522) );
  MUX2_X1 U14359 ( .A(n12021), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12031), .Z(
        P3_U3521) );
  MUX2_X1 U14360 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12022), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14361 ( .A(n12023), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12031), .Z(
        P3_U3517) );
  MUX2_X1 U14362 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12024), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14363 ( .A(n12177), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12031), .Z(
        P3_U3515) );
  MUX2_X1 U14364 ( .A(n12191), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12031), .Z(
        P3_U3514) );
  MUX2_X1 U14365 ( .A(n12178), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12031), .Z(
        P3_U3513) );
  MUX2_X1 U14366 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12213), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14367 ( .A(n12025), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12031), .Z(
        P3_U3511) );
  MUX2_X1 U14368 ( .A(n12238), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12031), .Z(
        P3_U3510) );
  MUX2_X1 U14369 ( .A(n12247), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12031), .Z(
        P3_U3509) );
  MUX2_X1 U14370 ( .A(n12260), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12031), .Z(
        P3_U3508) );
  MUX2_X1 U14371 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12270), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14372 ( .A(n12283), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12031), .Z(
        P3_U3506) );
  MUX2_X1 U14373 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12297), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14374 ( .A(n12282), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12031), .Z(
        P3_U3504) );
  MUX2_X1 U14375 ( .A(n14235), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12031), .Z(
        P3_U3503) );
  MUX2_X1 U14376 ( .A(n14807), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12031), .Z(
        P3_U3502) );
  MUX2_X1 U14377 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14237), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14378 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n14809), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14379 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12026), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14380 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12027), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14381 ( .A(n12028), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12031), .Z(
        P3_U3497) );
  MUX2_X1 U14382 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n14854), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14383 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12029), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14384 ( .A(n14853), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12031), .Z(
        P3_U3494) );
  MUX2_X1 U14385 ( .A(n12030), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12031), .Z(
        P3_U3492) );
  MUX2_X1 U14386 ( .A(n14889), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12031), .Z(
        P3_U3491) );
  INV_X1 U14387 ( .A(n14202), .ZN(n12055) );
  AOI22_X1 U14388 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14202), .B1(n12055), 
        .B2(n12262), .ZN(n12036) );
  NAND2_X1 U14389 ( .A1(n14199), .A2(n12032), .ZN(n12034) );
  OAI21_X1 U14390 ( .B1(n12036), .B2(n12035), .A(n12054), .ZN(n12052) );
  NAND2_X1 U14391 ( .A1(n14199), .A2(n12037), .ZN(n12039) );
  NAND2_X1 U14392 ( .A1(n12039), .A2(n12038), .ZN(n12041) );
  XNOR2_X1 U14393 ( .A(n12055), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U14394 ( .A1(n12040), .A2(n12041), .ZN(n12056) );
  OAI21_X1 U14395 ( .B1(n12041), .B2(n12040), .A(n12056), .ZN(n12042) );
  NAND2_X1 U14396 ( .A1(n12042), .A2(n14788), .ZN(n12045) );
  AOI21_X1 U14397 ( .B1(n14780), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12043), 
        .ZN(n12044) );
  OAI211_X1 U14398 ( .C1(n14797), .C2(n14202), .A(n12045), .B(n12044), .ZN(
        n12051) );
  MUX2_X1 U14399 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12069), .Z(n12062) );
  XNOR2_X1 U14400 ( .A(n12062), .B(n14202), .ZN(n12049) );
  OAI21_X1 U14401 ( .B1(n12047), .B2(n14199), .A(n12046), .ZN(n12048) );
  NOR2_X1 U14402 ( .A1(n12048), .A2(n12049), .ZN(n12061) );
  AOI211_X1 U14403 ( .C1(n12049), .C2(n12048), .A(n12113), .B(n12061), .ZN(
        n12050) );
  AOI211_X1 U14404 ( .C1(n14801), .C2(n12052), .A(n12051), .B(n12050), .ZN(
        n12053) );
  INV_X1 U14405 ( .A(n12053), .ZN(P3_U3198) );
  XNOR2_X1 U14406 ( .A(n12085), .B(n12255), .ZN(n12068) );
  NAND2_X1 U14407 ( .A1(n14202), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12057) );
  XOR2_X1 U14408 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12075), .Z(n12060) );
  NAND2_X1 U14409 ( .A1(n14780), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12058) );
  OAI211_X1 U14410 ( .C1(n12082), .C2(n12060), .A(n12059), .B(n12058), .ZN(
        n12066) );
  MUX2_X1 U14411 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12069), .Z(n12071) );
  XNOR2_X1 U14412 ( .A(n12071), .B(n12084), .ZN(n12063) );
  NOR2_X1 U14413 ( .A1(n12064), .A2(n12063), .ZN(n12070) );
  AOI211_X1 U14414 ( .C1(n12064), .C2(n12063), .A(n12113), .B(n12070), .ZN(
        n12065) );
  AOI211_X1 U14415 ( .C1(n12101), .C2(n6888), .A(n12066), .B(n12065), .ZN(
        n12067) );
  OAI21_X1 U14416 ( .B1(n12068), .B2(n12109), .A(n12067), .ZN(P3_U3199) );
  MUX2_X1 U14417 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12069), .Z(n12073) );
  AOI21_X1 U14418 ( .B1(n12071), .B2(n12084), .A(n12070), .ZN(n12094) );
  AOI21_X1 U14419 ( .B1(n12073), .B2(n12072), .A(n12093), .ZN(n12090) );
  INV_X1 U14420 ( .A(n14208), .ZN(n12105) );
  INV_X1 U14421 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12074) );
  XNOR2_X1 U14422 ( .A(n14208), .B(n12074), .ZN(n12096) );
  NAND2_X1 U14423 ( .A1(n12075), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U14424 ( .A1(n12076), .A2(n12084), .ZN(n12077) );
  NAND2_X1 U14425 ( .A1(n12078), .A2(n12077), .ZN(n12097) );
  XOR2_X1 U14426 ( .A(n12096), .B(n12097), .Z(n12081) );
  NAND2_X1 U14427 ( .A1(n14780), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U14428 ( .C1(n12082), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12088) );
  XNOR2_X1 U14429 ( .A(n14208), .B(P3_REG2_REG_18__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U14430 ( .A1(n12085), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12084), 
        .B2(n12083), .ZN(n12107) );
  XOR2_X1 U14431 ( .A(n12106), .B(n12107), .Z(n12086) );
  NOR2_X1 U14432 ( .A1(n12086), .A2(n12109), .ZN(n12087) );
  AOI211_X1 U14433 ( .C1(n12101), .C2(n12105), .A(n12088), .B(n12087), .ZN(
        n12089) );
  OAI21_X1 U14434 ( .B1(n12090), .B2(n12113), .A(n12089), .ZN(P3_U3200) );
  XNOR2_X1 U14435 ( .A(n12091), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12098) );
  XNOR2_X1 U14436 ( .A(n12091), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12108) );
  MUX2_X1 U14437 ( .A(n12098), .B(n12108), .S(n12092), .Z(n12095) );
  AOI22_X1 U14438 ( .A1(n12097), .A2(n12096), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n14208), .ZN(n12099) );
  XNOR2_X1 U14439 ( .A(n12099), .B(n12098), .ZN(n12111) );
  NAND2_X1 U14440 ( .A1(n12101), .A2(n12100), .ZN(n12103) );
  OAI211_X1 U14441 ( .C1(n12104), .C2(n14804), .A(n12103), .B(n12102), .ZN(
        n12110) );
  OAI21_X1 U14442 ( .B1(n12114), .B2(n12113), .A(n12112), .ZN(P3_U3201) );
  NAND2_X1 U14443 ( .A1(n12115), .A2(n14228), .ZN(n12121) );
  NOR2_X1 U14444 ( .A1(n14902), .A2(n12116), .ZN(n14226) );
  NOR2_X1 U14445 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  AOI211_X1 U14446 ( .C1(n14908), .C2(P3_REG2_REG_29__SCAN_IN), .A(n14226), 
        .B(n12119), .ZN(n12120) );
  OAI211_X1 U14447 ( .C1(n12122), .C2(n12305), .A(n12121), .B(n12120), .ZN(
        P3_U3204) );
  AOI21_X1 U14448 ( .B1(n12123), .B2(n12133), .A(n14873), .ZN(n12128) );
  OAI22_X1 U14449 ( .A1(n12125), .A2(n14867), .B1(n12124), .B2(n14869), .ZN(
        n12126) );
  AOI21_X1 U14450 ( .B1(n12128), .B2(n12127), .A(n12126), .ZN(n12323) );
  OAI22_X1 U14451 ( .A1(n14228), .A2(n12130), .B1(n12129), .B2(n14902), .ZN(
        n12135) );
  NOR2_X1 U14452 ( .A1(n12324), .A2(n12305), .ZN(n12134) );
  OAI21_X1 U14453 ( .B1(n14908), .B2(n12323), .A(n12136), .ZN(P3_U3205) );
  INV_X1 U14454 ( .A(n12137), .ZN(n12139) );
  AOI21_X1 U14455 ( .B1(n12139), .B2(n12138), .A(n14873), .ZN(n12144) );
  OAI22_X1 U14456 ( .A1(n12141), .A2(n14867), .B1(n12140), .B2(n14869), .ZN(
        n12142) );
  AOI21_X1 U14457 ( .B1(n12144), .B2(n12143), .A(n12142), .ZN(n12335) );
  OAI22_X1 U14458 ( .A1(n14228), .A2(n12146), .B1(n12145), .B2(n14902), .ZN(
        n12151) );
  NAND2_X1 U14459 ( .A1(n12161), .A2(n12147), .ZN(n12149) );
  XNOR2_X1 U14460 ( .A(n12149), .B(n12148), .ZN(n12336) );
  NOR2_X1 U14461 ( .A1(n12336), .A2(n12305), .ZN(n12150) );
  AOI211_X1 U14462 ( .C1(n14231), .C2(n12333), .A(n12151), .B(n12150), .ZN(
        n12152) );
  OAI21_X1 U14463 ( .B1(n12335), .B2(n14908), .A(n12152), .ZN(P3_U3208) );
  INV_X1 U14464 ( .A(n12153), .ZN(n12154) );
  AOI21_X1 U14465 ( .B1(n12154), .B2(n12163), .A(n14873), .ZN(n12158) );
  OAI22_X1 U14466 ( .A1(n12156), .A2(n14869), .B1(n12155), .B2(n14867), .ZN(
        n12157) );
  AOI21_X1 U14467 ( .B1(n12158), .B2(n11786), .A(n12157), .ZN(n12339) );
  OAI22_X1 U14468 ( .A1(n14228), .A2(n12160), .B1(n12159), .B2(n14902), .ZN(
        n12168) );
  INV_X1 U14469 ( .A(n12161), .ZN(n12166) );
  AOI21_X1 U14470 ( .B1(n12162), .B2(n12164), .A(n12163), .ZN(n12165) );
  NOR2_X1 U14471 ( .A1(n12166), .A2(n12165), .ZN(n12340) );
  NOR2_X1 U14472 ( .A1(n12340), .A2(n12305), .ZN(n12167) );
  AOI211_X1 U14473 ( .C1(n14231), .C2(n12337), .A(n12168), .B(n12167), .ZN(
        n12169) );
  OAI21_X1 U14474 ( .B1(n14908), .B2(n12339), .A(n12169), .ZN(P3_U3209) );
  NAND2_X1 U14475 ( .A1(n12201), .A2(n12170), .ZN(n12172) );
  AND2_X1 U14476 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  AOI21_X1 U14477 ( .B1(n12173), .B2(n12174), .A(n14873), .ZN(n12182) );
  OR2_X1 U14478 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  NAND2_X1 U14479 ( .A1(n12162), .A2(n12176), .ZN(n12345) );
  AOI22_X1 U14480 ( .A1(n14890), .A2(n12178), .B1(n12177), .B2(n14891), .ZN(
        n12179) );
  OAI21_X1 U14481 ( .B1(n12345), .B2(n14900), .A(n12179), .ZN(n12180) );
  AOI21_X1 U14482 ( .B1(n12182), .B2(n12181), .A(n12180), .ZN(n12343) );
  OAI22_X1 U14483 ( .A1(n14228), .A2(n12184), .B1(n12183), .B2(n14902), .ZN(
        n12185) );
  AOI21_X1 U14484 ( .B1(n12341), .B2(n14231), .A(n12185), .ZN(n12187) );
  OR2_X1 U14485 ( .A1(n14904), .A2(n12345), .ZN(n12186) );
  OAI211_X1 U14486 ( .C1(n12343), .C2(n14908), .A(n12187), .B(n12186), .ZN(
        P3_U3210) );
  NAND2_X1 U14487 ( .A1(n12201), .A2(n12188), .ZN(n12190) );
  XNOR2_X1 U14488 ( .A(n12190), .B(n12189), .ZN(n12192) );
  AOI222_X1 U14489 ( .A1(n12192), .A2(n14896), .B1(n12191), .B2(n14891), .C1(
        n12213), .C2(n14890), .ZN(n12348) );
  OAI22_X1 U14490 ( .A1(n14228), .A2(n12194), .B1(n12193), .B2(n14902), .ZN(
        n12198) );
  XNOR2_X1 U14491 ( .A(n12196), .B(n12195), .ZN(n12349) );
  NOR2_X1 U14492 ( .A1(n12349), .A2(n12305), .ZN(n12197) );
  AOI211_X1 U14493 ( .C1(n14231), .C2(n12346), .A(n12198), .B(n12197), .ZN(
        n12199) );
  OAI21_X1 U14494 ( .B1(n12348), .B2(n14908), .A(n12199), .ZN(P3_U3211) );
  XNOR2_X1 U14495 ( .A(n12200), .B(n12204), .ZN(n12353) );
  INV_X1 U14496 ( .A(n12201), .ZN(n12202) );
  AOI21_X1 U14497 ( .B1(n12204), .B2(n12203), .A(n12202), .ZN(n12205) );
  OAI222_X1 U14498 ( .A1(n14869), .A2(n12225), .B1(n14867), .B2(n12206), .C1(
        n12205), .C2(n14873), .ZN(n12350) );
  NAND2_X1 U14499 ( .A1(n12350), .A2(n14228), .ZN(n12211) );
  OAI22_X1 U14500 ( .A1(n14228), .A2(n12208), .B1(n12207), .B2(n14902), .ZN(
        n12209) );
  AOI21_X1 U14501 ( .B1(n12351), .B2(n14231), .A(n12209), .ZN(n12210) );
  OAI211_X1 U14502 ( .C1(n12305), .C2(n12353), .A(n12211), .B(n12210), .ZN(
        P3_U3212) );
  XNOR2_X1 U14503 ( .A(n12212), .B(n12218), .ZN(n12214) );
  AOI222_X1 U14504 ( .A1(n12214), .A2(n14896), .B1(n12213), .B2(n14891), .C1(
        n12238), .C2(n14890), .ZN(n12356) );
  OAI22_X1 U14505 ( .A1(n14228), .A2(n12216), .B1(n12215), .B2(n14902), .ZN(
        n12221) );
  OAI21_X1 U14506 ( .B1(n12219), .B2(n12218), .A(n12217), .ZN(n12357) );
  NOR2_X1 U14507 ( .A1(n12357), .A2(n12305), .ZN(n12220) );
  AOI211_X1 U14508 ( .C1(n14231), .C2(n12354), .A(n12221), .B(n12220), .ZN(
        n12222) );
  OAI21_X1 U14509 ( .B1(n12356), .B2(n14908), .A(n12222), .ZN(P3_U3213) );
  AOI21_X1 U14510 ( .B1(n12223), .B2(n12232), .A(n14873), .ZN(n12228) );
  OAI22_X1 U14511 ( .A1(n12225), .A2(n14867), .B1(n12224), .B2(n14869), .ZN(
        n12226) );
  AOI21_X1 U14512 ( .B1(n12228), .B2(n12227), .A(n12226), .ZN(n12360) );
  OAI22_X1 U14513 ( .A1(n14228), .A2(n12230), .B1(n12229), .B2(n14902), .ZN(
        n12234) );
  XNOR2_X1 U14514 ( .A(n12231), .B(n12232), .ZN(n12361) );
  NOR2_X1 U14515 ( .A1(n12361), .A2(n12305), .ZN(n12233) );
  AOI211_X1 U14516 ( .C1(n14231), .C2(n12358), .A(n12234), .B(n12233), .ZN(
        n12235) );
  OAI21_X1 U14517 ( .B1(n14908), .B2(n12360), .A(n12235), .ZN(P3_U3214) );
  OAI21_X1 U14518 ( .B1(n6512), .B2(n12237), .A(n12236), .ZN(n12239) );
  AOI222_X1 U14519 ( .A1(n12239), .A2(n14896), .B1(n12238), .B2(n14891), .C1(
        n12260), .C2(n14890), .ZN(n12364) );
  OAI22_X1 U14520 ( .A1(n14228), .A2(n13209), .B1(n12240), .B2(n14902), .ZN(
        n12244) );
  OAI21_X1 U14521 ( .B1(n6626), .B2(n12242), .A(n12241), .ZN(n12365) );
  NOR2_X1 U14522 ( .A1(n12365), .A2(n12305), .ZN(n12243) );
  AOI211_X1 U14523 ( .C1(n14231), .C2(n12362), .A(n12244), .B(n12243), .ZN(
        n12245) );
  OAI21_X1 U14524 ( .B1(n12364), .B2(n14908), .A(n12245), .ZN(P3_U3215) );
  XNOR2_X1 U14525 ( .A(n12246), .B(n12250), .ZN(n12248) );
  AOI222_X1 U14526 ( .A1(n12270), .A2(n14890), .B1(n14896), .B2(n12248), .C1(
        n12247), .C2(n14891), .ZN(n12369) );
  OAI21_X1 U14527 ( .B1(n12251), .B2(n12250), .A(n12249), .ZN(n12367) );
  INV_X1 U14528 ( .A(n12305), .ZN(n14828) );
  NOR2_X1 U14529 ( .A1(n12253), .A2(n12252), .ZN(n12257) );
  OAI22_X1 U14530 ( .A1(n14228), .A2(n12255), .B1(n12254), .B2(n14902), .ZN(
        n12256) );
  AOI211_X1 U14531 ( .C1(n12367), .C2(n14828), .A(n12257), .B(n12256), .ZN(
        n12258) );
  OAI21_X1 U14532 ( .B1(n12369), .B2(n14908), .A(n12258), .ZN(P3_U3216) );
  XNOR2_X1 U14533 ( .A(n12259), .B(n12266), .ZN(n12261) );
  AOI222_X1 U14534 ( .A1(n12283), .A2(n14890), .B1(n14896), .B2(n12261), .C1(
        n12260), .C2(n14891), .ZN(n12373) );
  OAI22_X1 U14535 ( .A1(n14228), .A2(n12262), .B1(n6519), .B2(n14902), .ZN(
        n12263) );
  AOI21_X1 U14536 ( .B1(n12370), .B2(n14231), .A(n12263), .ZN(n12268) );
  OAI21_X1 U14537 ( .B1(n12266), .B2(n12265), .A(n12264), .ZN(n12371) );
  NAND2_X1 U14538 ( .A1(n12371), .A2(n14828), .ZN(n12267) );
  OAI211_X1 U14539 ( .C1(n12373), .C2(n14908), .A(n12268), .B(n12267), .ZN(
        P3_U3217) );
  XNOR2_X1 U14540 ( .A(n12269), .B(n12276), .ZN(n12271) );
  AOI222_X1 U14541 ( .A1(n12297), .A2(n14890), .B1(n14896), .B2(n12271), .C1(
        n12270), .C2(n14891), .ZN(n12377) );
  OAI22_X1 U14542 ( .A1(n14228), .A2(n12273), .B1(n12272), .B2(n14902), .ZN(
        n12274) );
  AOI21_X1 U14543 ( .B1(n12374), .B2(n14231), .A(n12274), .ZN(n12279) );
  OAI21_X1 U14544 ( .B1(n12277), .B2(n12276), .A(n12275), .ZN(n12375) );
  NAND2_X1 U14545 ( .A1(n12375), .A2(n14828), .ZN(n12278) );
  OAI211_X1 U14546 ( .C1(n12377), .C2(n14908), .A(n12279), .B(n12278), .ZN(
        P3_U3218) );
  OAI211_X1 U14547 ( .C1(n12290), .C2(n12281), .A(n12280), .B(n14896), .ZN(
        n12285) );
  AOI22_X1 U14548 ( .A1(n14891), .A2(n12283), .B1(n12282), .B2(n14890), .ZN(
        n12284) );
  OAI22_X1 U14549 ( .A1(n14228), .A2(n12287), .B1(n12286), .B2(n14902), .ZN(
        n12288) );
  AOI21_X1 U14550 ( .B1(n12378), .B2(n14231), .A(n12288), .ZN(n12292) );
  XNOR2_X1 U14551 ( .A(n12289), .B(n12290), .ZN(n12379) );
  NAND2_X1 U14552 ( .A1(n12379), .A2(n14828), .ZN(n12291) );
  OAI211_X1 U14553 ( .C1(n12381), .C2(n14908), .A(n12292), .B(n12291), .ZN(
        P3_U3219) );
  XNOR2_X1 U14554 ( .A(n12293), .B(n12295), .ZN(n12385) );
  OAI211_X1 U14555 ( .C1(n12296), .C2(n12295), .A(n12294), .B(n14896), .ZN(
        n12299) );
  AOI22_X1 U14556 ( .A1(n12297), .A2(n14891), .B1(n14890), .B2(n14235), .ZN(
        n12298) );
  NAND2_X1 U14557 ( .A1(n12299), .A2(n12298), .ZN(n12382) );
  NAND2_X1 U14558 ( .A1(n12382), .A2(n14228), .ZN(n12304) );
  OAI22_X1 U14559 ( .A1(n14228), .A2(n12301), .B1(n12300), .B2(n14902), .ZN(
        n12302) );
  AOI21_X1 U14560 ( .B1(n12383), .B2(n14231), .A(n12302), .ZN(n12303) );
  OAI211_X1 U14561 ( .C1(n12305), .C2(n12385), .A(n12304), .B(n12303), .ZN(
        P3_U3220) );
  INV_X1 U14562 ( .A(n12306), .ZN(n12314) );
  NAND3_X1 U14563 ( .A1(n12309), .A2(n12308), .A3(n12307), .ZN(n12311) );
  NAND2_X1 U14564 ( .A1(n12311), .A2(n12310), .ZN(n12312) );
  OAI22_X1 U14565 ( .A1(n12315), .A2(n12314), .B1(n12313), .B2(n12312), .ZN(
        n12316) );
  INV_X1 U14566 ( .A(n12320), .ZN(P3_U3488) );
  NAND2_X1 U14567 ( .A1(n12321), .A2(n14916), .ZN(n12322) );
  OAI211_X1 U14568 ( .C1(n12386), .C2(n12324), .A(n12323), .B(n12322), .ZN(
        n12388) );
  MUX2_X1 U14569 ( .A(n12388), .B(P3_REG1_REG_28__SCAN_IN), .S(n14965), .Z(
        P3_U3487) );
  AOI22_X1 U14570 ( .A1(n12326), .A2(n14937), .B1(n14916), .B2(n12325), .ZN(
        n12327) );
  MUX2_X1 U14571 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12389), .S(n14968), .Z(
        P3_U3486) );
  AOI22_X1 U14572 ( .A1(n12330), .A2(n14937), .B1(n14916), .B2(n12329), .ZN(
        n12331) );
  NAND2_X1 U14573 ( .A1(n12332), .A2(n12331), .ZN(n12390) );
  MUX2_X1 U14574 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12390), .S(n14968), .Z(
        P3_U3485) );
  NAND2_X1 U14575 ( .A1(n12333), .A2(n14916), .ZN(n12334) );
  OAI211_X1 U14576 ( .C1(n12386), .C2(n12336), .A(n12335), .B(n12334), .ZN(
        n12391) );
  MUX2_X1 U14577 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12391), .S(n14968), .Z(
        P3_U3484) );
  NAND2_X1 U14578 ( .A1(n12337), .A2(n14916), .ZN(n12338) );
  OAI211_X1 U14579 ( .C1(n12386), .C2(n12340), .A(n12339), .B(n12338), .ZN(
        n12392) );
  MUX2_X1 U14580 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12392), .S(n14968), .Z(
        P3_U3483) );
  NAND2_X1 U14581 ( .A1(n12341), .A2(n14916), .ZN(n12342) );
  OAI211_X1 U14582 ( .C1(n12345), .C2(n12344), .A(n12343), .B(n12342), .ZN(
        n12393) );
  MUX2_X1 U14583 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12393), .S(n14968), .Z(
        P3_U3482) );
  NAND2_X1 U14584 ( .A1(n12346), .A2(n14916), .ZN(n12347) );
  OAI211_X1 U14585 ( .C1(n12386), .C2(n12349), .A(n12348), .B(n12347), .ZN(
        n12394) );
  MUX2_X1 U14586 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12394), .S(n14968), .Z(
        P3_U3481) );
  AOI21_X1 U14587 ( .B1(n14916), .B2(n12351), .A(n12350), .ZN(n12352) );
  OAI21_X1 U14588 ( .B1(n12386), .B2(n12353), .A(n12352), .ZN(n12395) );
  MUX2_X1 U14589 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n12395), .S(n14968), .Z(
        P3_U3480) );
  NAND2_X1 U14590 ( .A1(n12354), .A2(n14916), .ZN(n12355) );
  OAI211_X1 U14591 ( .C1(n12386), .C2(n12357), .A(n12356), .B(n12355), .ZN(
        n12396) );
  MUX2_X1 U14592 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12396), .S(n14968), .Z(
        P3_U3479) );
  NAND2_X1 U14593 ( .A1(n12358), .A2(n14916), .ZN(n12359) );
  OAI211_X1 U14594 ( .C1(n12386), .C2(n12361), .A(n12360), .B(n12359), .ZN(
        n12397) );
  MUX2_X1 U14595 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12397), .S(n14968), .Z(
        P3_U3478) );
  NAND2_X1 U14596 ( .A1(n12362), .A2(n14916), .ZN(n12363) );
  OAI211_X1 U14597 ( .C1(n12386), .C2(n12365), .A(n12364), .B(n12363), .ZN(
        n12398) );
  MUX2_X1 U14598 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12398), .S(n14968), .Z(
        P3_U3477) );
  AOI22_X1 U14599 ( .A1(n12367), .A2(n14946), .B1(n14916), .B2(n12366), .ZN(
        n12368) );
  NAND2_X1 U14600 ( .A1(n12369), .A2(n12368), .ZN(n12399) );
  MUX2_X1 U14601 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12399), .S(n14968), .Z(
        P3_U3476) );
  AOI22_X1 U14602 ( .A1(n12371), .A2(n14946), .B1(n14916), .B2(n12370), .ZN(
        n12372) );
  NAND2_X1 U14603 ( .A1(n12373), .A2(n12372), .ZN(n12400) );
  MUX2_X1 U14604 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12400), .S(n14968), .Z(
        P3_U3475) );
  AOI22_X1 U14605 ( .A1(n12375), .A2(n14946), .B1(n14916), .B2(n12374), .ZN(
        n12376) );
  NAND2_X1 U14606 ( .A1(n12377), .A2(n12376), .ZN(n12401) );
  MUX2_X1 U14607 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12401), .S(n14968), .Z(
        P3_U3474) );
  AOI22_X1 U14608 ( .A1(n12379), .A2(n14946), .B1(n14916), .B2(n12378), .ZN(
        n12380) );
  NAND2_X1 U14609 ( .A1(n12381), .A2(n12380), .ZN(n12402) );
  MUX2_X1 U14610 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n12402), .S(n14968), .Z(
        P3_U3473) );
  AOI21_X1 U14611 ( .B1(n12383), .B2(n14916), .A(n12382), .ZN(n12384) );
  OAI21_X1 U14612 ( .B1(n12386), .B2(n12385), .A(n12384), .ZN(n12403) );
  MUX2_X1 U14613 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12403), .S(n14968), .Z(
        P3_U3472) );
  MUX2_X1 U14614 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n12387), .S(n14968), .Z(
        P3_U3459) );
  MUX2_X1 U14615 ( .A(n12388), .B(P3_REG0_REG_28__SCAN_IN), .S(n14949), .Z(
        P3_U3455) );
  MUX2_X1 U14616 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12389), .S(n14948), .Z(
        P3_U3454) );
  MUX2_X1 U14617 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12390), .S(n14948), .Z(
        P3_U3453) );
  MUX2_X1 U14618 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12391), .S(n14948), .Z(
        P3_U3452) );
  MUX2_X1 U14619 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12392), .S(n14948), .Z(
        P3_U3451) );
  MUX2_X1 U14620 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12393), .S(n14948), .Z(
        P3_U3450) );
  MUX2_X1 U14621 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12394), .S(n14948), .Z(
        P3_U3449) );
  MUX2_X1 U14622 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n12395), .S(n14948), .Z(
        P3_U3448) );
  MUX2_X1 U14623 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12396), .S(n14948), .Z(
        P3_U3447) );
  MUX2_X1 U14624 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12397), .S(n14948), .Z(
        P3_U3446) );
  MUX2_X1 U14625 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12398), .S(n14948), .Z(
        P3_U3444) );
  MUX2_X1 U14626 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12399), .S(n14948), .Z(
        P3_U3441) );
  MUX2_X1 U14627 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12400), .S(n14948), .Z(
        P3_U3438) );
  MUX2_X1 U14628 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12401), .S(n14948), .Z(
        P3_U3435) );
  MUX2_X1 U14629 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n12402), .S(n14948), .Z(
        P3_U3432) );
  MUX2_X1 U14630 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n12403), .S(n14948), .Z(
        P3_U3429) );
  MUX2_X1 U14631 ( .A(n12405), .B(P3_D_REG_0__SCAN_IN), .S(n12404), .Z(
        P3_U3376) );
  NAND3_X1 U14632 ( .A1(n12407), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12409) );
  OAI22_X1 U14633 ( .A1(n12406), .A2(n12409), .B1(n12408), .B2(n14186), .ZN(
        n12410) );
  AOI21_X1 U14634 ( .B1(n12411), .B2(n14205), .A(n12410), .ZN(n12412) );
  INV_X1 U14635 ( .A(n12412), .ZN(P3_U3264) );
  INV_X1 U14636 ( .A(n12413), .ZN(n12415) );
  INV_X1 U14637 ( .A(n12416), .ZN(n12418) );
  OAI222_X1 U14638 ( .A1(n6473), .A2(n12419), .B1(n12423), .B2(n12418), .C1(
        n12417), .C2(n14186), .ZN(P3_U3266) );
  INV_X1 U14639 ( .A(n12420), .ZN(n12422) );
  MUX2_X1 U14640 ( .A(n12425), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI22_X1 U14641 ( .A1(n12882), .A2(n12747), .B1(n12880), .B2(n12575), .ZN(
        n12711) );
  OAI22_X1 U14642 ( .A1(n12429), .A2(n12711), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13214), .ZN(n12430) );
  AOI21_X1 U14643 ( .B1(n12716), .B2(n12558), .A(n12430), .ZN(n12431) );
  OAI22_X1 U14644 ( .A1(n12433), .A2(n12571), .B1(n12539), .B2(n12476), .ZN(
        n12434) );
  NAND2_X1 U14645 ( .A1(n12434), .A2(n12471), .ZN(n12439) );
  NOR2_X1 U14646 ( .A1(n12565), .A2(n12772), .ZN(n12437) );
  OAI22_X1 U14647 ( .A1(n12561), .A2(n12776), .B1(n12538), .B2(n12435), .ZN(
        n12436) );
  AOI211_X1 U14648 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3088), .A(n12437), 
        .B(n12436), .ZN(n12438) );
  OAI211_X1 U14649 ( .C1(n12783), .C2(n12516), .A(n12439), .B(n12438), .ZN(
        P2_U3188) );
  INV_X1 U14650 ( .A(n12440), .ZN(n12548) );
  NOR2_X1 U14651 ( .A1(n12476), .A2(n12443), .ZN(n12442) );
  AOI22_X1 U14652 ( .A1(n12548), .A2(n12533), .B1(n12442), .B2(n12441), .ZN(
        n12451) );
  OAI22_X1 U14653 ( .A1(n12465), .A2(n12777), .B1(n12443), .B2(n12773), .ZN(
        n12830) );
  AOI22_X1 U14654 ( .A1(n12444), .A2(n12830), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12445) );
  OAI21_X1 U14655 ( .B1(n12834), .B2(n12538), .A(n12445), .ZN(n12448) );
  NOR2_X1 U14656 ( .A1(n12446), .A2(n12571), .ZN(n12447) );
  AOI211_X1 U14657 ( .C1(n12956), .C2(n12569), .A(n12448), .B(n12447), .ZN(
        n12449) );
  OAI21_X1 U14658 ( .B1(n12451), .B2(n12450), .A(n12449), .ZN(P2_U3191) );
  AOI22_X1 U14659 ( .A1(n12452), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n12545), 
        .B2(n8268), .ZN(n12461) );
  AOI22_X1 U14660 ( .A1(n12492), .A2(n8273), .B1(n14695), .B2(n12569), .ZN(
        n12460) );
  INV_X1 U14661 ( .A(n12457), .ZN(n12454) );
  OAI21_X1 U14662 ( .B1(n12454), .B2(n12453), .A(n9097), .ZN(n12455) );
  NAND2_X1 U14663 ( .A1(n12533), .A2(n12455), .ZN(n12459) );
  NAND3_X1 U14664 ( .A1(n12563), .A2(n12457), .A3(n12456), .ZN(n12458) );
  NAND4_X1 U14665 ( .A1(n12461), .A2(n12460), .A3(n12459), .A4(n12458), .ZN(
        P2_U3194) );
  OAI211_X1 U14666 ( .C1(n12517), .C2(n12463), .A(n12462), .B(n12533), .ZN(
        n12469) );
  NOR2_X1 U14667 ( .A1(n12561), .A2(n12772), .ZN(n12467) );
  OAI22_X1 U14668 ( .A1(n12565), .A2(n12465), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12464), .ZN(n12466) );
  AOI211_X1 U14669 ( .C1(n12558), .C2(n12808), .A(n12467), .B(n12466), .ZN(
        n12468) );
  OAI211_X1 U14670 ( .C1(n7224), .C2(n12516), .A(n12469), .B(n12468), .ZN(
        P2_U3195) );
  NAND2_X1 U14671 ( .A1(n12471), .A2(n12470), .ZN(n12510) );
  INV_X1 U14672 ( .A(n12472), .ZN(n12474) );
  NOR2_X1 U14673 ( .A1(n12474), .A2(n12473), .ZN(n12509) );
  NAND2_X1 U14674 ( .A1(n12510), .A2(n12509), .ZN(n12508) );
  AOI21_X1 U14675 ( .B1(n12508), .B2(n12475), .A(n12571), .ZN(n12479) );
  NOR3_X1 U14676 ( .A1(n12477), .A2(n12776), .A3(n12476), .ZN(n12478) );
  OAI21_X1 U14677 ( .B1(n12479), .B2(n12478), .A(n12554), .ZN(n12485) );
  NOR2_X1 U14678 ( .A1(n12561), .A2(n12480), .ZN(n12483) );
  OAI22_X1 U14679 ( .A1(n12565), .A2(n12776), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12481), .ZN(n12482) );
  AOI211_X1 U14680 ( .C1(n12558), .C2(n12740), .A(n12483), .B(n12482), .ZN(
        n12484) );
  OAI211_X1 U14681 ( .C1(n7100), .C2(n12516), .A(n12485), .B(n12484), .ZN(
        P2_U3197) );
  OAI21_X1 U14682 ( .B1(n12488), .B2(n12487), .A(n12499), .ZN(n12489) );
  NAND2_X1 U14683 ( .A1(n12489), .A2(n12533), .ZN(n12494) );
  NAND2_X1 U14684 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14645)
         );
  INV_X1 U14685 ( .A(n14645), .ZN(n12491) );
  OAI22_X1 U14686 ( .A1(n12561), .A2(n12547), .B1(n12538), .B2(n12887), .ZN(
        n12490) );
  AOI211_X1 U14687 ( .C1(n12492), .C2(n12883), .A(n12491), .B(n12490), .ZN(
        n12493) );
  OAI211_X1 U14688 ( .C1(n12495), .C2(n12516), .A(n12494), .B(n12493), .ZN(
        P2_U3198) );
  AOI22_X1 U14689 ( .A1(n12545), .A2(n12861), .B1(n12558), .B2(n12867), .ZN(
        n12497) );
  OAI211_X1 U14690 ( .C1(n12498), .C2(n12565), .A(n12497), .B(n12496), .ZN(
        n12505) );
  INV_X1 U14691 ( .A(n12499), .ZN(n12503) );
  AOI22_X1 U14692 ( .A1(n12500), .A2(n12533), .B1(n12563), .B2(n12862), .ZN(
        n12502) );
  NOR3_X1 U14693 ( .A1(n12503), .A2(n12502), .A3(n12501), .ZN(n12504) );
  AOI211_X1 U14694 ( .C1(n12966), .C2(n12569), .A(n12505), .B(n12504), .ZN(
        n12506) );
  OAI21_X1 U14695 ( .B1(n12507), .B2(n12571), .A(n12506), .ZN(P2_U3200) );
  OAI211_X1 U14696 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n12533), .ZN(
        n12515) );
  NOR2_X1 U14697 ( .A1(n12539), .A2(n12565), .ZN(n12513) );
  INV_X1 U14698 ( .A(n12764), .ZN(n12511) );
  OAI22_X1 U14699 ( .A1(n12561), .A2(n12728), .B1(n12538), .B2(n12511), .ZN(
        n12512) );
  AOI211_X1 U14700 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3088), .A(n12513), 
        .B(n12512), .ZN(n12514) );
  OAI211_X1 U14701 ( .C1(n12766), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        P2_U3201) );
  INV_X1 U14702 ( .A(n12517), .ZN(n12528) );
  INV_X1 U14703 ( .A(n12518), .ZN(n12521) );
  AOI21_X1 U14704 ( .B1(n12521), .B2(n12520), .A(n12519), .ZN(n12522) );
  AOI21_X1 U14705 ( .B1(n12528), .B2(n12523), .A(n12522), .ZN(n12531) );
  OAI22_X1 U14706 ( .A1(n12561), .A2(n12536), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12524), .ZN(n12527) );
  OAI22_X1 U14707 ( .A1(n12565), .A2(n12525), .B1(n12538), .B2(n12821), .ZN(
        n12526) );
  AOI211_X1 U14708 ( .C1(n12951), .C2(n12569), .A(n12527), .B(n12526), .ZN(
        n12530) );
  NAND3_X1 U14709 ( .A1(n12528), .A2(n12563), .A3(n12802), .ZN(n12529) );
  OAI211_X1 U14710 ( .C1(n12531), .C2(n12571), .A(n12530), .B(n12529), .ZN(
        P2_U3205) );
  INV_X1 U14711 ( .A(n12532), .ZN(n12544) );
  AOI22_X1 U14712 ( .A1(n12534), .A2(n12533), .B1(n12563), .B2(n6968), .ZN(
        n12543) );
  INV_X1 U14713 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12535) );
  OAI22_X1 U14714 ( .A1(n12565), .A2(n12536), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12535), .ZN(n12541) );
  OAI22_X1 U14715 ( .A1(n12539), .A2(n12561), .B1(n12538), .B2(n12537), .ZN(
        n12540) );
  AOI211_X1 U14716 ( .C1(n12940), .C2(n12569), .A(n12541), .B(n12540), .ZN(
        n12542) );
  OAI21_X1 U14717 ( .B1(n12544), .B2(n12543), .A(n12542), .ZN(P2_U3207) );
  AOI22_X1 U14718 ( .A1(n12545), .A2(n12846), .B1(n12558), .B2(n12851), .ZN(
        n12546) );
  NAND2_X1 U14719 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14663)
         );
  OAI211_X1 U14720 ( .C1(n12547), .C2(n12565), .A(n12546), .B(n14663), .ZN(
        n12552) );
  AOI211_X1 U14721 ( .C1(n12550), .C2(n12549), .A(n12571), .B(n12548), .ZN(
        n12551) );
  AOI211_X1 U14722 ( .C1(n12961), .C2(n12569), .A(n12552), .B(n12551), .ZN(
        n12553) );
  INV_X1 U14723 ( .A(n12553), .ZN(P2_U3210) );
  INV_X1 U14724 ( .A(n12554), .ZN(n12557) );
  INV_X1 U14725 ( .A(n12555), .ZN(n12556) );
  AOI21_X1 U14726 ( .B1(n12564), .B2(n12557), .A(n12556), .ZN(n12572) );
  NAND2_X1 U14727 ( .A1(n12558), .A2(n12732), .ZN(n12560) );
  NAND2_X1 U14728 ( .A1(P2_U3088), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n12559)
         );
  OAI211_X1 U14729 ( .C1(n12729), .C2(n12561), .A(n12560), .B(n12559), .ZN(
        n12568) );
  NAND3_X1 U14730 ( .A1(n12564), .A2(n12563), .A3(n12562), .ZN(n12566) );
  AOI21_X1 U14731 ( .B1(n12566), .B2(n12565), .A(n12728), .ZN(n12567) );
  AOI211_X1 U14732 ( .C1(n12922), .C2(n12569), .A(n12568), .B(n12567), .ZN(
        n12570) );
  OAI21_X1 U14733 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(P2_U3212) );
  MUX2_X1 U14734 ( .A(n12573), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12588), .Z(
        P2_U3561) );
  MUX2_X1 U14735 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12574), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U14736 ( .A(n12575), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12588), .Z(
        P2_U3559) );
  MUX2_X1 U14737 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n12576), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U14738 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n12747), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U14739 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n12758), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U14740 ( .A(n12746), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12588), .Z(
        P2_U3555) );
  MUX2_X1 U14741 ( .A(n12791), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12588), .Z(
        P2_U3554) );
  MUX2_X1 U14742 ( .A(n6968), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12588), .Z(
        P2_U3553) );
  MUX2_X1 U14743 ( .A(n12817), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12588), .Z(
        P2_U3552) );
  MUX2_X1 U14744 ( .A(n12846), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12588), .Z(
        P2_U3550) );
  MUX2_X1 U14745 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n12861), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U14746 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n12881), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U14747 ( .A(n12862), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12588), .Z(
        P2_U3547) );
  MUX2_X1 U14748 ( .A(n12883), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12588), .Z(
        P2_U3546) );
  MUX2_X1 U14749 ( .A(n12577), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12588), .Z(
        P2_U3545) );
  MUX2_X1 U14750 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8326), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U14751 ( .A(n12578), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12588), .Z(
        P2_U3543) );
  MUX2_X1 U14752 ( .A(n12579), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12588), .Z(
        P2_U3542) );
  INV_X2 U14753 ( .A(P2_U3947), .ZN(n12588) );
  MUX2_X1 U14754 ( .A(n12580), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12588), .Z(
        P2_U3541) );
  MUX2_X1 U14755 ( .A(n12581), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12588), .Z(
        P2_U3540) );
  MUX2_X1 U14756 ( .A(n12582), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12588), .Z(
        P2_U3539) );
  MUX2_X1 U14757 ( .A(n12583), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12588), .Z(
        P2_U3538) );
  MUX2_X1 U14758 ( .A(n12584), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12588), .Z(
        P2_U3537) );
  MUX2_X1 U14759 ( .A(n12585), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12588), .Z(
        P2_U3536) );
  MUX2_X1 U14760 ( .A(n12586), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12588), .Z(
        P2_U3535) );
  MUX2_X1 U14761 ( .A(n12587), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12588), .Z(
        P2_U3534) );
  MUX2_X1 U14762 ( .A(n8268), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12588), .Z(
        P2_U3533) );
  MUX2_X1 U14763 ( .A(n8271), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12588), .Z(
        P2_U3532) );
  MUX2_X1 U14764 ( .A(n8273), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12588), .Z(
        P2_U3531) );
  OAI22_X1 U14765 ( .A1(n14661), .A2(n12590), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12589), .ZN(n12591) );
  AOI21_X1 U14766 ( .B1(n14535), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n12591), .ZN(
        n12600) );
  OAI211_X1 U14767 ( .C1(n12594), .C2(n12593), .A(n14652), .B(n12592), .ZN(
        n12599) );
  OAI211_X1 U14768 ( .C1(n12597), .C2(n12596), .A(n14657), .B(n12595), .ZN(
        n12598) );
  NAND3_X1 U14769 ( .A1(n12600), .A2(n12599), .A3(n12598), .ZN(P2_U3215) );
  INV_X1 U14770 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12601) );
  OAI22_X1 U14771 ( .A1(n14661), .A2(n12602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12601), .ZN(n12603) );
  AOI21_X1 U14772 ( .B1(n14535), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n12603), .ZN(
        n12612) );
  OAI211_X1 U14773 ( .C1(n12606), .C2(n12605), .A(n14652), .B(n12604), .ZN(
        n12611) );
  OAI211_X1 U14774 ( .C1(n12609), .C2(n12608), .A(n14657), .B(n12607), .ZN(
        n12610) );
  NAND3_X1 U14775 ( .A1(n12612), .A2(n12611), .A3(n12610), .ZN(P2_U3216) );
  NAND2_X1 U14776 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n12613) );
  OAI21_X1 U14777 ( .B1(n14661), .B2(n12614), .A(n12613), .ZN(n12615) );
  AOI21_X1 U14778 ( .B1(n14535), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n12615), .ZN(
        n12624) );
  OAI211_X1 U14779 ( .C1(n12618), .C2(n12617), .A(n14657), .B(n12616), .ZN(
        n12623) );
  OAI211_X1 U14780 ( .C1(n12621), .C2(n12620), .A(n14652), .B(n12619), .ZN(
        n12622) );
  NAND3_X1 U14781 ( .A1(n12624), .A2(n12623), .A3(n12622), .ZN(P2_U3220) );
  OAI211_X1 U14782 ( .C1(n12627), .C2(n12626), .A(n14657), .B(n12625), .ZN(
        n12638) );
  OAI211_X1 U14783 ( .C1(n12630), .C2(n12629), .A(n14652), .B(n12628), .ZN(
        n12637) );
  NAND2_X1 U14784 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n12633) );
  OR2_X1 U14785 ( .A1(n14661), .A2(n12631), .ZN(n12632) );
  OAI211_X1 U14786 ( .C1(n14665), .C2(n12634), .A(n12633), .B(n12632), .ZN(
        n12635) );
  INV_X1 U14787 ( .A(n12635), .ZN(n12636) );
  NAND3_X1 U14788 ( .A1(n12638), .A2(n12637), .A3(n12636), .ZN(P2_U3221) );
  OAI21_X1 U14789 ( .B1(n14661), .B2(n12640), .A(n12639), .ZN(n12641) );
  AOI21_X1 U14790 ( .B1(n14535), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n12641), .ZN(
        n12650) );
  OAI211_X1 U14791 ( .C1(n12644), .C2(n12643), .A(n14652), .B(n12642), .ZN(
        n12649) );
  OAI211_X1 U14792 ( .C1(n12647), .C2(n12646), .A(n14657), .B(n12645), .ZN(
        n12648) );
  NAND3_X1 U14793 ( .A1(n12650), .A2(n12649), .A3(n12648), .ZN(P2_U3222) );
  OAI21_X1 U14794 ( .B1(n12653), .B2(n12652), .A(n12651), .ZN(n12654) );
  NAND2_X1 U14795 ( .A1(n12654), .A2(n14657), .ZN(n12663) );
  OAI21_X1 U14796 ( .B1(n14661), .B2(n12656), .A(n12655), .ZN(n12657) );
  AOI21_X1 U14797 ( .B1(n14535), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n12657), 
        .ZN(n12662) );
  OAI211_X1 U14798 ( .C1(n12660), .C2(n12659), .A(n12658), .B(n14652), .ZN(
        n12661) );
  NAND3_X1 U14799 ( .A1(n12663), .A2(n12662), .A3(n12661), .ZN(P2_U3225) );
  AOI21_X1 U14800 ( .B1(n12670), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12664), 
        .ZN(n12665) );
  NAND2_X1 U14801 ( .A1(n12665), .A2(n14660), .ZN(n12667) );
  INV_X1 U14802 ( .A(n12665), .ZN(n12666) );
  XNOR2_X1 U14803 ( .A(n14660), .B(n12666), .ZN(n14655) );
  INV_X1 U14804 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U14805 ( .A1(n14655), .A2(n14654), .ZN(n14653) );
  NAND2_X1 U14806 ( .A1(n12667), .A2(n14653), .ZN(n12668) );
  XNOR2_X1 U14807 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12668), .ZN(n12678) );
  INV_X1 U14808 ( .A(n12678), .ZN(n12676) );
  AOI21_X1 U14809 ( .B1(n12670), .B2(P2_REG1_REG_17__SCAN_IN), .A(n12669), 
        .ZN(n12671) );
  XNOR2_X1 U14810 ( .A(n14660), .B(n12671), .ZN(n14650) );
  NOR2_X1 U14811 ( .A1(n14649), .A2(n14650), .ZN(n14648) );
  NOR2_X1 U14812 ( .A1(n12671), .A2(n14660), .ZN(n12672) );
  NOR2_X1 U14813 ( .A1(n14648), .A2(n12672), .ZN(n12674) );
  XOR2_X1 U14814 ( .A(n12674), .B(n12673), .Z(n12677) );
  OAI21_X1 U14815 ( .B1(n12677), .B2(n14633), .A(n14661), .ZN(n12675) );
  AOI21_X1 U14816 ( .B1(n12676), .B2(n14657), .A(n12675), .ZN(n12681) );
  AOI22_X1 U14817 ( .A1(n12678), .A2(n14657), .B1(n14652), .B2(n12677), .ZN(
        n12680) );
  MUX2_X1 U14818 ( .A(n12681), .B(n12680), .S(n12679), .Z(n12683) );
  NAND2_X1 U14819 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n12682)
         );
  OAI211_X1 U14820 ( .C1(n12684), .C2(n14665), .A(n12683), .B(n12682), .ZN(
        P2_U3233) );
  NAND2_X1 U14821 ( .A1(n12902), .A2(n12691), .ZN(n12690) );
  XNOR2_X1 U14822 ( .A(n12690), .B(n8217), .ZN(n12685) );
  NAND2_X1 U14823 ( .A1(n12685), .A2(n12971), .ZN(n12899) );
  OR2_X1 U14824 ( .A1(n12687), .A2(n12686), .ZN(n12900) );
  NOR2_X1 U14825 ( .A1(n12858), .A2(n12900), .ZN(n12693) );
  NOR2_X1 U14826 ( .A1(n8217), .A2(n14673), .ZN(n12688) );
  AOI211_X1 U14827 ( .C1(n14680), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12693), 
        .B(n12688), .ZN(n12689) );
  OAI21_X1 U14828 ( .B1(n12811), .B2(n12899), .A(n12689), .ZN(P2_U3234) );
  OAI211_X1 U14829 ( .C1(n12902), .C2(n12691), .A(n12971), .B(n12690), .ZN(
        n12901) );
  NOR2_X1 U14830 ( .A1(n12902), .A2(n14673), .ZN(n12692) );
  AOI211_X1 U14831 ( .C1(n14680), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12693), 
        .B(n12692), .ZN(n12694) );
  OAI21_X1 U14832 ( .B1(n12811), .B2(n12901), .A(n12694), .ZN(P2_U3235) );
  AOI21_X1 U14833 ( .B1(n12695), .B2(n12701), .A(n12774), .ZN(n12698) );
  AOI21_X1 U14834 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(n12911) );
  OAI21_X1 U14835 ( .B1(n12699), .B2(n12886), .A(n12911), .ZN(n12708) );
  OAI21_X1 U14836 ( .B1(n12702), .B2(n12701), .A(n12700), .ZN(n12912) );
  AOI22_X1 U14837 ( .A1(n12909), .A2(n12896), .B1(n14680), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n12706) );
  AOI21_X1 U14838 ( .B1(n12909), .B2(n12714), .A(n12865), .ZN(n12704) );
  AND2_X1 U14839 ( .A1(n12704), .A2(n12703), .ZN(n12908) );
  NAND2_X1 U14840 ( .A1(n12908), .A2(n14667), .ZN(n12705) );
  OAI211_X1 U14841 ( .C1(n12912), .C2(n12893), .A(n12706), .B(n12705), .ZN(
        n12707) );
  AOI21_X1 U14842 ( .B1(n12708), .B2(n12889), .A(n12707), .ZN(n12709) );
  INV_X1 U14843 ( .A(n12709), .ZN(P2_U3237) );
  XNOR2_X1 U14844 ( .A(n12710), .B(n12720), .ZN(n12713) );
  INV_X1 U14845 ( .A(n12711), .ZN(n12712) );
  AOI21_X1 U14846 ( .B1(n12713), .B2(n12879), .A(n12712), .ZN(n12919) );
  AOI21_X1 U14847 ( .B1(n12915), .B2(n12730), .A(n12865), .ZN(n12715) );
  NAND2_X1 U14848 ( .A1(n12715), .A2(n12714), .ZN(n12918) );
  AOI22_X1 U14849 ( .A1(n14680), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n12716), 
        .B2(n14669), .ZN(n12718) );
  NAND2_X1 U14850 ( .A1(n12915), .A2(n12896), .ZN(n12717) );
  OAI211_X1 U14851 ( .C1(n12918), .C2(n12811), .A(n12718), .B(n12717), .ZN(
        n12719) );
  INV_X1 U14852 ( .A(n12719), .ZN(n12723) );
  OR2_X1 U14853 ( .A1(n12721), .A2(n12720), .ZN(n12914) );
  NAND3_X1 U14854 ( .A1(n12914), .A2(n12913), .A3(n14677), .ZN(n12722) );
  OAI211_X1 U14855 ( .C1(n12919), .C2(n12858), .A(n12723), .B(n12722), .ZN(
        P2_U3238) );
  XNOR2_X1 U14856 ( .A(n12724), .B(n12725), .ZN(n12924) );
  XNOR2_X1 U14857 ( .A(n12726), .B(n12725), .ZN(n12727) );
  OAI222_X1 U14858 ( .A1(n12777), .A2(n12729), .B1(n12773), .B2(n12728), .C1(
        n12774), .C2(n12727), .ZN(n12920) );
  NAND2_X1 U14859 ( .A1(n12920), .A2(n12889), .ZN(n12737) );
  INV_X1 U14860 ( .A(n12730), .ZN(n12731) );
  AOI211_X1 U14861 ( .C1(n12922), .C2(n7103), .A(n12865), .B(n12731), .ZN(
        n12921) );
  AOI22_X1 U14862 ( .A1(n14680), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n12732), 
        .B2(n14669), .ZN(n12733) );
  OAI21_X1 U14863 ( .B1(n12734), .B2(n14673), .A(n12733), .ZN(n12735) );
  AOI21_X1 U14864 ( .B1(n12921), .B2(n14667), .A(n12735), .ZN(n12736) );
  OAI211_X1 U14865 ( .C1(n12924), .C2(n12893), .A(n12737), .B(n12736), .ZN(
        P2_U3239) );
  XOR2_X1 U14866 ( .A(n12738), .B(n12742), .Z(n12929) );
  AOI211_X1 U14867 ( .C1(n12926), .C2(n12762), .A(n12865), .B(n12739), .ZN(
        n12925) );
  AOI22_X1 U14868 ( .A1(n14680), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n12740), 
        .B2(n14669), .ZN(n12741) );
  OAI21_X1 U14869 ( .B1(n7100), .B2(n14673), .A(n12741), .ZN(n12750) );
  OR3_X1 U14870 ( .A1(n6586), .A2(n12743), .A3(n12742), .ZN(n12744) );
  NAND2_X1 U14871 ( .A1(n12745), .A2(n12744), .ZN(n12748) );
  AOI222_X1 U14872 ( .A1(n12879), .A2(n12748), .B1(n12747), .B2(n12880), .C1(
        n12746), .C2(n12882), .ZN(n12928) );
  NOR2_X1 U14873 ( .A1(n12928), .A2(n12858), .ZN(n12749) );
  AOI211_X1 U14874 ( .C1(n12925), .C2(n14667), .A(n12750), .B(n12749), .ZN(
        n12751) );
  OAI21_X1 U14875 ( .B1(n12929), .B2(n12893), .A(n12751), .ZN(P2_U3240) );
  NAND2_X1 U14876 ( .A1(n12753), .A2(n12752), .ZN(n12754) );
  AOI21_X1 U14877 ( .B1(n12757), .B2(n12756), .A(n6586), .ZN(n12760) );
  AOI22_X1 U14878 ( .A1(n12791), .A2(n12882), .B1(n12880), .B2(n12758), .ZN(
        n12759) );
  OAI21_X1 U14879 ( .B1(n12760), .B2(n12774), .A(n12759), .ZN(n12761) );
  AOI21_X1 U14880 ( .B1(n14745), .B2(n12767), .A(n12761), .ZN(n12933) );
  INV_X1 U14881 ( .A(n12762), .ZN(n12763) );
  AOI211_X1 U14882 ( .C1(n12931), .C2(n12779), .A(n12865), .B(n12763), .ZN(
        n12930) );
  AOI22_X1 U14883 ( .A1(n14680), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n12764), 
        .B2(n14669), .ZN(n12765) );
  OAI21_X1 U14884 ( .B1(n12766), .B2(n14673), .A(n12765), .ZN(n12769) );
  NOR2_X1 U14885 ( .A1(n12934), .A2(n12854), .ZN(n12768) );
  AOI211_X1 U14886 ( .C1(n12930), .C2(n14667), .A(n12769), .B(n12768), .ZN(
        n12770) );
  OAI21_X1 U14887 ( .B1(n12933), .B2(n14680), .A(n12770), .ZN(P2_U3241) );
  XNOR2_X1 U14888 ( .A(n12771), .B(n12784), .ZN(n12775) );
  OAI222_X1 U14889 ( .A1(n12777), .A2(n12776), .B1(n12775), .B2(n12774), .C1(
        n12773), .C2(n12772), .ZN(n12935) );
  AOI21_X1 U14890 ( .B1(n12778), .B2(n14669), .A(n12935), .ZN(n12788) );
  INV_X1 U14891 ( .A(n12793), .ZN(n12781) );
  INV_X1 U14892 ( .A(n12779), .ZN(n12780) );
  AOI211_X1 U14893 ( .C1(n7102), .C2(n12781), .A(n12865), .B(n12780), .ZN(
        n12936) );
  OAI22_X1 U14894 ( .A1(n12783), .A2(n14673), .B1(n12782), .B2(n12889), .ZN(
        n12786) );
  XNOR2_X1 U14895 ( .A(n6592), .B(n12784), .ZN(n12938) );
  NOR2_X1 U14896 ( .A1(n12938), .A2(n12893), .ZN(n12785) );
  AOI211_X1 U14897 ( .C1(n12936), .C2(n14667), .A(n12786), .B(n12785), .ZN(
        n12787) );
  OAI21_X1 U14898 ( .B1(n12788), .B2(n14680), .A(n12787), .ZN(P2_U3242) );
  XNOR2_X1 U14899 ( .A(n12789), .B(n6500), .ZN(n12790) );
  AOI222_X1 U14900 ( .A1(n12817), .A2(n12882), .B1(n12791), .B2(n12880), .C1(
        n12879), .C2(n12790), .ZN(n12942) );
  NOR2_X1 U14901 ( .A1(n12796), .A2(n12807), .ZN(n12792) );
  NOR3_X1 U14902 ( .A1(n12793), .A2(n12792), .A3(n12865), .ZN(n12939) );
  AOI22_X1 U14903 ( .A1(n14680), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n12794), 
        .B2(n14669), .ZN(n12795) );
  OAI21_X1 U14904 ( .B1(n12796), .B2(n14673), .A(n12795), .ZN(n12799) );
  OAI21_X1 U14905 ( .B1(n6545), .B2(n6500), .A(n12797), .ZN(n12943) );
  NOR2_X1 U14906 ( .A1(n12943), .A2(n12893), .ZN(n12798) );
  AOI211_X1 U14907 ( .C1(n12939), .C2(n14667), .A(n12799), .B(n12798), .ZN(
        n12800) );
  OAI21_X1 U14908 ( .B1(n12942), .B2(n14680), .A(n12800), .ZN(P2_U3243) );
  XNOR2_X1 U14909 ( .A(n12801), .B(n12804), .ZN(n12803) );
  AOI222_X1 U14910 ( .A1(n12879), .A2(n12803), .B1(n6968), .B2(n12880), .C1(
        n12802), .C2(n12882), .ZN(n12948) );
  XNOR2_X1 U14911 ( .A(n12805), .B(n12804), .ZN(n12949) );
  INV_X1 U14912 ( .A(n12949), .ZN(n12813) );
  AND2_X1 U14913 ( .A1(n12823), .A2(n12946), .ZN(n12806) );
  OR3_X1 U14914 ( .A1(n12807), .A2(n12806), .A3(n12865), .ZN(n12944) );
  AOI22_X1 U14915 ( .A1(n14680), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n12808), 
        .B2(n14669), .ZN(n12810) );
  NAND2_X1 U14916 ( .A1(n12946), .A2(n12896), .ZN(n12809) );
  OAI211_X1 U14917 ( .C1(n12944), .C2(n12811), .A(n12810), .B(n12809), .ZN(
        n12812) );
  AOI21_X1 U14918 ( .B1(n12813), .B2(n14677), .A(n12812), .ZN(n12814) );
  OAI21_X1 U14919 ( .B1(n12948), .B2(n14680), .A(n12814), .ZN(P2_U3244) );
  XOR2_X1 U14920 ( .A(n12818), .B(n12815), .Z(n12816) );
  AOI222_X1 U14921 ( .A1(n12846), .A2(n12882), .B1(n12817), .B2(n12880), .C1(
        n12879), .C2(n12816), .ZN(n12953) );
  XNOR2_X1 U14922 ( .A(n12819), .B(n12818), .ZN(n12954) );
  NAND2_X1 U14923 ( .A1(n14680), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U14924 ( .B1(n12886), .B2(n12821), .A(n12820), .ZN(n12822) );
  AOI21_X1 U14925 ( .B1(n12951), .B2(n12896), .A(n12822), .ZN(n12826) );
  AOI21_X1 U14926 ( .B1(n12951), .B2(n12833), .A(n12865), .ZN(n12824) );
  AND2_X1 U14927 ( .A1(n12824), .A2(n12823), .ZN(n12950) );
  NAND2_X1 U14928 ( .A1(n12950), .A2(n14667), .ZN(n12825) );
  OAI211_X1 U14929 ( .C1(n12954), .C2(n12893), .A(n12826), .B(n12825), .ZN(
        n12827) );
  INV_X1 U14930 ( .A(n12827), .ZN(n12828) );
  OAI21_X1 U14931 ( .B1(n12953), .B2(n14680), .A(n12828), .ZN(P2_U3245) );
  XOR2_X1 U14932 ( .A(n12829), .B(n12839), .Z(n12831) );
  AOI21_X1 U14933 ( .B1(n12831), .B2(n12879), .A(n12830), .ZN(n12958) );
  OR2_X1 U14934 ( .A1(n12837), .A2(n12850), .ZN(n12832) );
  AND3_X1 U14935 ( .A1(n12833), .A2(n12971), .A3(n12832), .ZN(n12955) );
  NOR2_X1 U14936 ( .A1(n12886), .A2(n12834), .ZN(n12835) );
  AOI21_X1 U14937 ( .B1(n14680), .B2(P2_REG2_REG_19__SCAN_IN), .A(n12835), 
        .ZN(n12836) );
  OAI21_X1 U14938 ( .B1(n12837), .B2(n14673), .A(n12836), .ZN(n12841) );
  XNOR2_X1 U14939 ( .A(n12838), .B(n12839), .ZN(n12959) );
  NOR2_X1 U14940 ( .A1(n12959), .A2(n12893), .ZN(n12840) );
  AOI211_X1 U14941 ( .C1(n12955), .C2(n14667), .A(n12841), .B(n12840), .ZN(
        n12842) );
  OAI21_X1 U14942 ( .B1(n12958), .B2(n14680), .A(n12842), .ZN(P2_U3246) );
  XOR2_X1 U14943 ( .A(n12843), .B(n12845), .Z(n12849) );
  AOI21_X1 U14944 ( .B1(n12845), .B2(n12844), .A(n6553), .ZN(n12964) );
  AOI22_X1 U14945 ( .A1(n12846), .A2(n12880), .B1(n12882), .B2(n12881), .ZN(
        n12847) );
  OAI21_X1 U14946 ( .B1(n12964), .B2(n6485), .A(n12847), .ZN(n12848) );
  AOI21_X1 U14947 ( .B1(n12849), .B2(n12879), .A(n12848), .ZN(n12963) );
  AOI211_X1 U14948 ( .C1(n12961), .C2(n6497), .A(n12865), .B(n12850), .ZN(
        n12960) );
  AOI22_X1 U14949 ( .A1(n14680), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n12851), 
        .B2(n14669), .ZN(n12852) );
  OAI21_X1 U14950 ( .B1(n12853), .B2(n14673), .A(n12852), .ZN(n12856) );
  NOR2_X1 U14951 ( .A1(n12964), .A2(n12854), .ZN(n12855) );
  AOI211_X1 U14952 ( .C1(n12960), .C2(n14667), .A(n12856), .B(n12855), .ZN(
        n12857) );
  OAI21_X1 U14953 ( .B1(n12963), .B2(n12858), .A(n12857), .ZN(P2_U3247) );
  XOR2_X1 U14954 ( .A(n12859), .B(n12863), .Z(n12860) );
  AOI222_X1 U14955 ( .A1(n12862), .A2(n12882), .B1(n12861), .B2(n12880), .C1(
        n12879), .C2(n12860), .ZN(n12968) );
  XNOR2_X1 U14956 ( .A(n12864), .B(n12863), .ZN(n12969) );
  INV_X1 U14957 ( .A(n12969), .ZN(n12872) );
  AOI21_X1 U14958 ( .B1(n12966), .B2(n12874), .A(n12865), .ZN(n12866) );
  AND2_X1 U14959 ( .A1(n12866), .A2(n6497), .ZN(n12965) );
  NAND2_X1 U14960 ( .A1(n12965), .A2(n14667), .ZN(n12869) );
  AOI22_X1 U14961 ( .A1(n14680), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12867), 
        .B2(n14669), .ZN(n12868) );
  OAI211_X1 U14962 ( .C1(n12870), .C2(n14673), .A(n12869), .B(n12868), .ZN(
        n12871) );
  AOI21_X1 U14963 ( .B1(n12872), .B2(n14677), .A(n12871), .ZN(n12873) );
  OAI21_X1 U14964 ( .B1(n12968), .B2(n14680), .A(n12873), .ZN(P2_U3248) );
  INV_X1 U14965 ( .A(n12874), .ZN(n12875) );
  AOI21_X1 U14966 ( .B1(n12970), .B2(n12876), .A(n12875), .ZN(n12972) );
  XNOR2_X1 U14967 ( .A(n12877), .B(n12891), .ZN(n12878) );
  AOI222_X1 U14968 ( .A1(n12883), .A2(n12882), .B1(n12881), .B2(n12880), .C1(
        n12879), .C2(n12878), .ZN(n12974) );
  INV_X1 U14969 ( .A(n12974), .ZN(n12884) );
  AOI21_X1 U14970 ( .B1(n12885), .B2(n12972), .A(n12884), .ZN(n12898) );
  INV_X1 U14971 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12888) );
  OAI22_X1 U14972 ( .A1(n12889), .A2(n12888), .B1(n12887), .B2(n12886), .ZN(
        n12895) );
  OAI21_X1 U14973 ( .B1(n12892), .B2(n12891), .A(n12890), .ZN(n12975) );
  NOR2_X1 U14974 ( .A1(n12975), .A2(n12893), .ZN(n12894) );
  AOI211_X1 U14975 ( .C1(n12896), .C2(n12970), .A(n12895), .B(n12894), .ZN(
        n12897) );
  OAI21_X1 U14976 ( .B1(n12898), .B2(n14680), .A(n12897), .ZN(P2_U3249) );
  OAI211_X1 U14977 ( .C1(n8217), .C2(n14756), .A(n12899), .B(n12900), .ZN(
        n12977) );
  MUX2_X1 U14978 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n12977), .S(n14779), .Z(
        P2_U3530) );
  OAI211_X1 U14979 ( .C1(n12902), .C2(n14756), .A(n12901), .B(n12900), .ZN(
        n12978) );
  MUX2_X1 U14980 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n12978), .S(n14779), .Z(
        P2_U3529) );
  AOI21_X1 U14981 ( .B1(n14738), .B2(n12904), .A(n12903), .ZN(n12905) );
  AOI21_X1 U14982 ( .B1(n14738), .B2(n12909), .A(n12908), .ZN(n12910) );
  OAI211_X1 U14983 ( .C1(n14720), .C2(n12912), .A(n12911), .B(n12910), .ZN(
        n12979) );
  MUX2_X1 U14984 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n12979), .S(n14779), .Z(
        P2_U3527) );
  NAND3_X1 U14985 ( .A1(n12914), .A2(n12913), .A3(n14274), .ZN(n12917) );
  NAND2_X1 U14986 ( .A1(n12915), .A2(n14738), .ZN(n12916) );
  NAND4_X1 U14987 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12980) );
  MUX2_X1 U14988 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n12980), .S(n14779), .Z(
        P2_U3526) );
  AOI211_X1 U14989 ( .C1(n14738), .C2(n12922), .A(n12921), .B(n12920), .ZN(
        n12923) );
  OAI21_X1 U14990 ( .B1(n14720), .B2(n12924), .A(n12923), .ZN(n12981) );
  MUX2_X1 U14991 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n12981), .S(n14779), .Z(
        P2_U3525) );
  AOI21_X1 U14992 ( .B1(n14738), .B2(n12926), .A(n12925), .ZN(n12927) );
  OAI211_X1 U14993 ( .C1(n14720), .C2(n12929), .A(n12928), .B(n12927), .ZN(
        n12982) );
  MUX2_X1 U14994 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n12982), .S(n14779), .Z(
        P2_U3524) );
  AOI21_X1 U14995 ( .B1(n14738), .B2(n12931), .A(n12930), .ZN(n12932) );
  OAI211_X1 U14996 ( .C1(n14740), .C2(n12934), .A(n12933), .B(n12932), .ZN(
        n12983) );
  MUX2_X1 U14997 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n12983), .S(n14779), .Z(
        P2_U3523) );
  AOI211_X1 U14998 ( .C1(n14738), .C2(n7102), .A(n12936), .B(n12935), .ZN(
        n12937) );
  OAI21_X1 U14999 ( .B1(n14720), .B2(n12938), .A(n12937), .ZN(n12984) );
  MUX2_X1 U15000 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n12984), .S(n14779), .Z(
        P2_U3522) );
  AOI21_X1 U15001 ( .B1(n14738), .B2(n12940), .A(n12939), .ZN(n12941) );
  OAI211_X1 U15002 ( .C1(n14720), .C2(n12943), .A(n12942), .B(n12941), .ZN(
        n12985) );
  MUX2_X1 U15003 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n12985), .S(n14779), .Z(
        P2_U3521) );
  INV_X1 U15004 ( .A(n12944), .ZN(n12945) );
  AOI21_X1 U15005 ( .B1(n14738), .B2(n12946), .A(n12945), .ZN(n12947) );
  OAI211_X1 U15006 ( .C1(n14720), .C2(n12949), .A(n12948), .B(n12947), .ZN(
        n12986) );
  MUX2_X1 U15007 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n12986), .S(n14779), .Z(
        P2_U3520) );
  AOI21_X1 U15008 ( .B1(n14738), .B2(n12951), .A(n12950), .ZN(n12952) );
  OAI211_X1 U15009 ( .C1(n14720), .C2(n12954), .A(n12953), .B(n12952), .ZN(
        n12987) );
  MUX2_X1 U15010 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n12987), .S(n14779), .Z(
        P2_U3519) );
  AOI21_X1 U15011 ( .B1(n14738), .B2(n12956), .A(n12955), .ZN(n12957) );
  OAI211_X1 U15012 ( .C1(n14720), .C2(n12959), .A(n12958), .B(n12957), .ZN(
        n12988) );
  MUX2_X1 U15013 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n12988), .S(n14779), .Z(
        P2_U3518) );
  AOI21_X1 U15014 ( .B1(n14738), .B2(n12961), .A(n12960), .ZN(n12962) );
  OAI211_X1 U15015 ( .C1(n12964), .C2(n14740), .A(n12963), .B(n12962), .ZN(
        n12989) );
  MUX2_X1 U15016 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n12989), .S(n14779), .Z(
        P2_U3517) );
  AOI21_X1 U15017 ( .B1(n14738), .B2(n12966), .A(n12965), .ZN(n12967) );
  OAI211_X1 U15018 ( .C1(n14720), .C2(n12969), .A(n12968), .B(n12967), .ZN(
        n12990) );
  MUX2_X1 U15019 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n12990), .S(n14779), .Z(
        P2_U3516) );
  AOI22_X1 U15020 ( .A1(n12972), .A2(n12971), .B1(n14738), .B2(n12970), .ZN(
        n12973) );
  OAI211_X1 U15021 ( .C1(n14720), .C2(n12975), .A(n12974), .B(n12973), .ZN(
        n12991) );
  MUX2_X1 U15022 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n12991), .S(n14779), .Z(
        P2_U3515) );
  MUX2_X1 U15023 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n12976), .S(n14779), .Z(
        P2_U3510) );
  MUX2_X1 U15024 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n12977), .S(n14764), .Z(
        P2_U3498) );
  MUX2_X1 U15025 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n12978), .S(n14764), .Z(
        P2_U3497) );
  MUX2_X1 U15026 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n12979), .S(n14764), .Z(
        P2_U3495) );
  MUX2_X1 U15027 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n12980), .S(n14764), .Z(
        P2_U3494) );
  MUX2_X1 U15028 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n12981), .S(n14764), .Z(
        P2_U3493) );
  MUX2_X1 U15029 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n12982), .S(n14764), .Z(
        P2_U3492) );
  MUX2_X1 U15030 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n12983), .S(n14764), .Z(
        P2_U3491) );
  MUX2_X1 U15031 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n12984), .S(n14764), .Z(
        P2_U3490) );
  MUX2_X1 U15032 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n12985), .S(n14764), .Z(
        P2_U3489) );
  MUX2_X1 U15033 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n12986), .S(n14764), .Z(
        P2_U3488) );
  MUX2_X1 U15034 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n12987), .S(n14764), .Z(
        P2_U3487) );
  MUX2_X1 U15035 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n12988), .S(n14764), .Z(
        P2_U3486) );
  MUX2_X1 U15036 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n12989), .S(n14764), .Z(
        P2_U3484) );
  MUX2_X1 U15037 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n12990), .S(n14764), .Z(
        P2_U3481) );
  MUX2_X1 U15038 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n12991), .S(n14764), .Z(
        P2_U3478) );
  INV_X1 U15039 ( .A(n12992), .ZN(n14159) );
  NOR4_X1 U15040 ( .A1(n7569), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7929), .A4(
        P2_U3088), .ZN(n12993) );
  AOI21_X1 U15041 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n12998), .A(n12993), 
        .ZN(n12994) );
  OAI21_X1 U15042 ( .B1(n14159), .B2(n13012), .A(n12994), .ZN(P2_U3296) );
  INV_X1 U15043 ( .A(n13563), .ZN(n14161) );
  OAI222_X1 U15044 ( .A1(P2_U3088), .A2(n12996), .B1(n13012), .B2(n14161), 
        .C1(n12995), .C2(n13010), .ZN(P2_U3298) );
  AOI21_X1 U15045 ( .B1(n12998), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n12997), 
        .ZN(n12999) );
  OAI21_X1 U15046 ( .B1(n13000), .B2(n13012), .A(n12999), .ZN(P2_U3299) );
  INV_X1 U15047 ( .A(n13001), .ZN(n14164) );
  OAI222_X1 U15048 ( .A1(P2_U3088), .A2(n13003), .B1(n13012), .B2(n14164), 
        .C1(n13002), .C2(n13010), .ZN(P2_U3300) );
  INV_X1 U15049 ( .A(n13004), .ZN(n13007) );
  INV_X1 U15050 ( .A(n13005), .ZN(n14169) );
  OAI222_X1 U15051 ( .A1(P2_U3088), .A2(n13007), .B1(n13012), .B2(n14169), 
        .C1(n13006), .C2(n13010), .ZN(P2_U3301) );
  INV_X1 U15052 ( .A(n13009), .ZN(n14171) );
  OAI222_X1 U15053 ( .A1(n13013), .A2(P2_U3088), .B1(n13012), .B2(n14171), 
        .C1(n13011), .C2(n13010), .ZN(P2_U3302) );
  INV_X1 U15054 ( .A(n13014), .ZN(n13015) );
  MUX2_X1 U15055 ( .A(n13015), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15056 ( .A(n13016), .ZN(n13019) );
  INV_X1 U15057 ( .A(n13017), .ZN(n13018) );
  AOI22_X2 U15058 ( .A1(n13021), .A2(n13020), .B1(n13019), .B2(n13018), .ZN(
        n14289) );
  OAI22_X1 U15059 ( .A1(n14315), .A2(n13064), .B1(n14016), .B2(n13063), .ZN(
        n13023) );
  XNOR2_X1 U15060 ( .A(n13023), .B(n13022), .ZN(n13025) );
  OAI22_X1 U15061 ( .A1(n14315), .A2(n13063), .B1(n14016), .B2(n13062), .ZN(
        n13024) );
  NOR2_X1 U15062 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  AOI21_X1 U15063 ( .B1(n13025), .B2(n13024), .A(n13026), .ZN(n14290) );
  NAND2_X1 U15064 ( .A1(n14289), .A2(n14290), .ZN(n14288) );
  INV_X1 U15065 ( .A(n13026), .ZN(n13027) );
  OAI22_X1 U15066 ( .A1(n7119), .A2(n13064), .B1(n14001), .B2(n13063), .ZN(
        n13028) );
  XNOR2_X1 U15067 ( .A(n13028), .B(n13022), .ZN(n13029) );
  OAI22_X1 U15068 ( .A1(n7119), .A2(n13063), .B1(n14001), .B2(n13062), .ZN(
        n13417) );
  OAI22_X1 U15069 ( .A1(n14008), .A2(n13064), .B1(n14014), .B2(n13063), .ZN(
        n13030) );
  XNOR2_X1 U15070 ( .A(n13030), .B(n13022), .ZN(n13034) );
  OR2_X1 U15071 ( .A1(n14008), .A2(n13063), .ZN(n13032) );
  NAND2_X1 U15072 ( .A1(n13655), .A2(n13313), .ZN(n13031) );
  NAND2_X1 U15073 ( .A1(n13032), .A2(n13031), .ZN(n13033) );
  NOR2_X1 U15074 ( .A1(n13034), .A2(n13033), .ZN(n13035) );
  AOI21_X1 U15075 ( .B1(n13034), .B2(n13033), .A(n13035), .ZN(n13348) );
  INV_X1 U15076 ( .A(n13035), .ZN(n13036) );
  NAND2_X1 U15077 ( .A1(n13346), .A2(n13036), .ZN(n13358) );
  NAND2_X1 U15078 ( .A1(n14126), .A2(n13311), .ZN(n13038) );
  NAND2_X1 U15079 ( .A1(n13966), .A2(n9725), .ZN(n13037) );
  NAND2_X1 U15080 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  XNOR2_X1 U15081 ( .A(n13039), .B(n13022), .ZN(n13042) );
  NAND2_X1 U15082 ( .A1(n14126), .A2(n9725), .ZN(n13041) );
  NAND2_X1 U15083 ( .A1(n13966), .A2(n13313), .ZN(n13040) );
  NAND2_X1 U15084 ( .A1(n13041), .A2(n13040), .ZN(n13043) );
  NAND2_X1 U15085 ( .A1(n13042), .A2(n13043), .ZN(n13359) );
  NAND2_X1 U15086 ( .A1(n13358), .A2(n13359), .ZN(n13357) );
  INV_X1 U15087 ( .A(n13042), .ZN(n13045) );
  INV_X1 U15088 ( .A(n13043), .ZN(n13044) );
  NAND2_X1 U15089 ( .A1(n13045), .A2(n13044), .ZN(n13361) );
  NAND2_X1 U15090 ( .A1(n13357), .A2(n13361), .ZN(n13395) );
  NAND2_X1 U15091 ( .A1(n13972), .A2(n13311), .ZN(n13047) );
  NAND2_X1 U15092 ( .A1(n13654), .A2(n9725), .ZN(n13046) );
  NAND2_X1 U15093 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  XNOR2_X1 U15094 ( .A(n13048), .B(n13022), .ZN(n13049) );
  AOI22_X1 U15095 ( .A1(n13972), .A2(n9725), .B1(n13313), .B2(n13654), .ZN(
        n13050) );
  XNOR2_X1 U15096 ( .A(n13049), .B(n13050), .ZN(n13396) );
  INV_X1 U15097 ( .A(n13049), .ZN(n13051) );
  NAND2_X1 U15098 ( .A1(n13051), .A2(n13050), .ZN(n13052) );
  AND2_X1 U15099 ( .A1(n13965), .A2(n13313), .ZN(n13053) );
  AOI21_X1 U15100 ( .B1(n14116), .B2(n9725), .A(n13053), .ZN(n13058) );
  NAND2_X1 U15101 ( .A1(n14116), .A2(n13311), .ZN(n13055) );
  NAND2_X1 U15102 ( .A1(n13965), .A2(n9725), .ZN(n13054) );
  NAND2_X1 U15103 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  XNOR2_X1 U15104 ( .A(n13056), .B(n13022), .ZN(n13060) );
  XOR2_X1 U15105 ( .A(n13058), .B(n13060), .Z(n13301) );
  INV_X1 U15106 ( .A(n13301), .ZN(n13057) );
  INV_X1 U15107 ( .A(n13058), .ZN(n13059) );
  NAND2_X1 U15108 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  OAI22_X1 U15109 ( .A1(n14108), .A2(n13063), .B1(n13531), .B2(n13062), .ZN(
        n13066) );
  OAI22_X1 U15110 ( .A1(n14108), .A2(n13064), .B1(n13531), .B2(n13063), .ZN(
        n13065) );
  XNOR2_X1 U15111 ( .A(n13065), .B(n13022), .ZN(n13067) );
  XOR2_X1 U15112 ( .A(n13066), .B(n13067), .Z(n13377) );
  NAND2_X1 U15113 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  AOI22_X1 U15114 ( .A1(n13923), .A2(n13311), .B1(n9725), .B2(n13652), .ZN(
        n13069) );
  XNOR2_X1 U15115 ( .A(n13069), .B(n13022), .ZN(n13071) );
  AOI22_X1 U15116 ( .A1(n13923), .A2(n9725), .B1(n13313), .B2(n13652), .ZN(
        n13070) );
  XNOR2_X1 U15117 ( .A(n13071), .B(n13070), .ZN(n13329) );
  NAND2_X1 U15118 ( .A1(n13071), .A2(n13070), .ZN(n13072) );
  NAND2_X1 U15119 ( .A1(n13326), .A2(n13072), .ZN(n13384) );
  NAND2_X1 U15120 ( .A1(n14094), .A2(n13311), .ZN(n13074) );
  NAND2_X1 U15121 ( .A1(n13651), .A2(n9725), .ZN(n13073) );
  NAND2_X1 U15122 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  XNOR2_X1 U15123 ( .A(n13075), .B(n13022), .ZN(n13076) );
  AOI22_X1 U15124 ( .A1(n14094), .A2(n9725), .B1(n13313), .B2(n13651), .ZN(
        n13077) );
  XNOR2_X1 U15125 ( .A(n13076), .B(n13077), .ZN(n13385) );
  INV_X1 U15126 ( .A(n13076), .ZN(n13078) );
  NAND2_X1 U15127 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  NAND2_X1 U15128 ( .A1(n14087), .A2(n13311), .ZN(n13081) );
  NAND2_X1 U15129 ( .A1(n13876), .A2(n9725), .ZN(n13080) );
  NAND2_X1 U15130 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  XNOR2_X1 U15131 ( .A(n13082), .B(n13022), .ZN(n13083) );
  AOI22_X1 U15132 ( .A1(n14087), .A2(n9725), .B1(n13313), .B2(n13876), .ZN(
        n13084) );
  XNOR2_X1 U15133 ( .A(n13083), .B(n13084), .ZN(n13118) );
  INV_X1 U15134 ( .A(n13083), .ZN(n13085) );
  NAND2_X1 U15135 ( .A1(n14083), .A2(n13311), .ZN(n13087) );
  NAND2_X1 U15136 ( .A1(n13858), .A2(n9725), .ZN(n13086) );
  NAND2_X1 U15137 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  XNOR2_X1 U15138 ( .A(n13088), .B(n13022), .ZN(n13089) );
  AOI22_X1 U15139 ( .A1(n14083), .A2(n9725), .B1(n13313), .B2(n13858), .ZN(
        n13090) );
  XNOR2_X1 U15140 ( .A(n13089), .B(n13090), .ZN(n13369) );
  INV_X1 U15141 ( .A(n13089), .ZN(n13091) );
  NAND2_X1 U15142 ( .A1(n13091), .A2(n13090), .ZN(n13092) );
  NAND2_X1 U15143 ( .A1(n14074), .A2(n13311), .ZN(n13094) );
  NAND2_X1 U15144 ( .A1(n13875), .A2(n9725), .ZN(n13093) );
  NAND2_X1 U15145 ( .A1(n13094), .A2(n13093), .ZN(n13095) );
  XNOR2_X1 U15146 ( .A(n13095), .B(n13022), .ZN(n13096) );
  AOI22_X1 U15147 ( .A1(n14074), .A2(n9725), .B1(n13313), .B2(n13875), .ZN(
        n13097) );
  XNOR2_X1 U15148 ( .A(n13096), .B(n13097), .ZN(n13337) );
  INV_X1 U15149 ( .A(n13096), .ZN(n13098) );
  NAND2_X1 U15150 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND2_X1 U15151 ( .A1(n13839), .A2(n13311), .ZN(n13101) );
  NAND2_X1 U15152 ( .A1(n13859), .A2(n9725), .ZN(n13100) );
  NAND2_X1 U15153 ( .A1(n13101), .A2(n13100), .ZN(n13102) );
  XNOR2_X1 U15154 ( .A(n13102), .B(n13022), .ZN(n13105) );
  AOI22_X1 U15155 ( .A1(n13839), .A2(n9725), .B1(n13313), .B2(n13859), .ZN(
        n13103) );
  XNOR2_X1 U15156 ( .A(n13105), .B(n13103), .ZN(n13406) );
  INV_X1 U15157 ( .A(n13103), .ZN(n13104) );
  AOI22_X1 U15158 ( .A1(n14063), .A2(n9725), .B1(n13313), .B2(n13835), .ZN(
        n13306) );
  NAND2_X1 U15159 ( .A1(n14063), .A2(n13311), .ZN(n13107) );
  NAND2_X1 U15160 ( .A1(n13835), .A2(n9725), .ZN(n13106) );
  NAND2_X1 U15161 ( .A1(n13107), .A2(n13106), .ZN(n13108) );
  XNOR2_X1 U15162 ( .A(n13108), .B(n13022), .ZN(n13308) );
  XOR2_X1 U15163 ( .A(n13306), .B(n13308), .Z(n13309) );
  XNOR2_X1 U15164 ( .A(n13310), .B(n13309), .ZN(n13109) );
  NAND2_X1 U15165 ( .A1(n13109), .A2(n14366), .ZN(n13116) );
  NAND2_X1 U15166 ( .A1(n13859), .A2(n14416), .ZN(n13111) );
  NAND2_X1 U15167 ( .A1(n13798), .A2(n14413), .ZN(n13110) );
  NAND2_X1 U15168 ( .A1(n13111), .A2(n13110), .ZN(n13819) );
  INV_X1 U15169 ( .A(n13825), .ZN(n13113) );
  OAI22_X1 U15170 ( .A1(n14376), .A2(n13113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13112), .ZN(n13114) );
  AOI21_X1 U15171 ( .B1(n13819), .B2(n14373), .A(n13114), .ZN(n13115) );
  OAI211_X1 U15172 ( .C1(n13827), .C2(n13393), .A(n13116), .B(n13115), .ZN(
        P1_U3214) );
  XOR2_X1 U15173 ( .A(n13118), .B(n13117), .Z(n13124) );
  AND2_X1 U15174 ( .A1(n13858), .A2(n14413), .ZN(n13119) );
  AOI21_X1 U15175 ( .B1(n13651), .B2(n14416), .A(n13119), .ZN(n13900) );
  NOR2_X1 U15176 ( .A1(n13900), .A2(n13332), .ZN(n13122) );
  INV_X1 U15177 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13120) );
  OAI22_X1 U15178 ( .A1(n13893), .A2(n14376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13120), .ZN(n13121) );
  AOI211_X1 U15179 ( .C1(n14087), .C2(n14300), .A(n13122), .B(n13121), .ZN(
        n13123) );
  OAI21_X1 U15180 ( .B1(n13124), .B2(n13425), .A(n13123), .ZN(P1_U3216) );
  AOI22_X1 U15181 ( .A1(n13251), .A2(keyinput117), .B1(keyinput96), .B2(n13126), .ZN(n13125) );
  OAI221_X1 U15182 ( .B1(n13251), .B2(keyinput117), .C1(n13126), .C2(
        keyinput96), .A(n13125), .ZN(n13135) );
  AOI22_X1 U15183 ( .A1(n13128), .A2(keyinput110), .B1(n10072), .B2(keyinput75), .ZN(n13127) );
  OAI221_X1 U15184 ( .B1(n13128), .B2(keyinput110), .C1(n10072), .C2(
        keyinput75), .A(n13127), .ZN(n13134) );
  AOI22_X1 U15185 ( .A1(n13130), .A2(keyinput89), .B1(n14771), .B2(keyinput79), 
        .ZN(n13129) );
  OAI221_X1 U15186 ( .B1(n13130), .B2(keyinput89), .C1(n14771), .C2(keyinput79), .A(n13129), .ZN(n13133) );
  INV_X1 U15187 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n13245) );
  INV_X1 U15188 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U15189 ( .A1(n13245), .A2(keyinput111), .B1(keyinput124), .B2(
        n14489), .ZN(n13131) );
  OAI221_X1 U15190 ( .B1(n13245), .B2(keyinput111), .C1(n14489), .C2(
        keyinput124), .A(n13131), .ZN(n13132) );
  NOR4_X1 U15191 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n13154) );
  AOI22_X1 U15192 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput87), .B1(
        P3_IR_REG_26__SCAN_IN), .B2(keyinput114), .ZN(n13136) );
  OAI221_X1 U15193 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput87), .C1(
        P3_IR_REG_26__SCAN_IN), .C2(keyinput114), .A(n13136), .ZN(n13143) );
  AOI22_X1 U15194 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput66), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput121), .ZN(n13137) );
  OAI221_X1 U15195 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput66), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput121), .A(n13137), .ZN(n13142)
         );
  AOI22_X1 U15196 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(keyinput64), .B1(
        P2_REG2_REG_20__SCAN_IN), .B2(keyinput103), .ZN(n13138) );
  OAI221_X1 U15197 ( .B1(P3_IR_REG_20__SCAN_IN), .B2(keyinput64), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput103), .A(n13138), .ZN(n13141) );
  AOI22_X1 U15198 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput104), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput122), .ZN(n13139) );
  OAI221_X1 U15199 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput104), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput122), .A(n13139), .ZN(n13140) );
  NOR4_X1 U15200 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13153) );
  AOI22_X1 U15201 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput102), .B1(SI_29_), .B2(keyinput127), .ZN(n13144) );
  OAI221_X1 U15202 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput102), .C1(
        SI_29_), .C2(keyinput127), .A(n13144), .ZN(n13151) );
  AOI22_X1 U15203 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(keyinput78), .B1(
        P2_REG0_REG_27__SCAN_IN), .B2(keyinput72), .ZN(n13145) );
  OAI221_X1 U15204 ( .B1(P3_IR_REG_24__SCAN_IN), .B2(keyinput78), .C1(
        P2_REG0_REG_27__SCAN_IN), .C2(keyinput72), .A(n13145), .ZN(n13150) );
  AOI22_X1 U15205 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput77), .B1(
        P2_REG0_REG_22__SCAN_IN), .B2(keyinput101), .ZN(n13146) );
  OAI221_X1 U15206 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput77), .C1(
        P2_REG0_REG_22__SCAN_IN), .C2(keyinput101), .A(n13146), .ZN(n13149) );
  AOI22_X1 U15207 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(keyinput93), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput74), .ZN(n13147) );
  OAI221_X1 U15208 ( .B1(P3_IR_REG_17__SCAN_IN), .B2(keyinput93), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput74), .A(n13147), .ZN(n13148) );
  NOR4_X1 U15209 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n13148), .ZN(
        n13152) );
  AND3_X1 U15210 ( .A1(n13154), .A2(n13153), .A3(n13152), .ZN(n13207) );
  AOI22_X1 U15211 ( .A1(P3_REG0_REG_30__SCAN_IN), .A2(keyinput80), .B1(
        P2_REG2_REG_9__SCAN_IN), .B2(keyinput115), .ZN(n13155) );
  OAI221_X1 U15212 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(keyinput80), .C1(
        P2_REG2_REG_9__SCAN_IN), .C2(keyinput115), .A(n13155), .ZN(n13162) );
  AOI22_X1 U15213 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(keyinput91), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput82), .ZN(n13156) );
  OAI221_X1 U15214 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(keyinput91), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput82), .A(n13156), .ZN(n13161) );
  AOI22_X1 U15215 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput105), .B1(
        P2_ADDR_REG_19__SCAN_IN), .B2(keyinput83), .ZN(n13157) );
  OAI221_X1 U15216 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput105), .C1(
        P2_ADDR_REG_19__SCAN_IN), .C2(keyinput83), .A(n13157), .ZN(n13160) );
  AOI22_X1 U15217 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput118), .B1(
        P3_REG2_REG_1__SCAN_IN), .B2(keyinput92), .ZN(n13158) );
  OAI221_X1 U15218 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput118), .C1(
        P3_REG2_REG_1__SCAN_IN), .C2(keyinput92), .A(n13158), .ZN(n13159) );
  NOR4_X1 U15219 ( .A1(n13162), .A2(n13161), .A3(n13160), .A4(n13159), .ZN(
        n13187) );
  AOI22_X1 U15220 ( .A1(n13164), .A2(keyinput67), .B1(n13209), .B2(keyinput120), .ZN(n13163) );
  OAI221_X1 U15221 ( .B1(n13164), .B2(keyinput67), .C1(n13209), .C2(
        keyinput120), .A(n13163), .ZN(n13170) );
  XNOR2_X1 U15222 ( .A(n14562), .B(keyinput84), .ZN(n13169) );
  XNOR2_X1 U15223 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput112), .ZN(n13167)
         );
  XNOR2_X1 U15224 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput81), .ZN(n13166) );
  XNOR2_X1 U15225 ( .A(keyinput119), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n13165)
         );
  NAND3_X1 U15226 ( .A1(n13167), .A2(n13166), .A3(n13165), .ZN(n13168) );
  NOR3_X1 U15227 ( .A1(n13170), .A2(n13169), .A3(n13168), .ZN(n13186) );
  INV_X1 U15228 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U15229 ( .A1(keyinput98), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n13172), 
        .B2(keyinput95), .ZN(n13171) );
  OAI221_X1 U15230 ( .B1(keyinput98), .B2(P2_REG1_REG_12__SCAN_IN), .C1(n13172), .C2(keyinput95), .A(n13171), .ZN(n13178) );
  XNOR2_X1 U15231 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput107), .ZN(n13176) );
  XNOR2_X1 U15232 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput70), .ZN(n13175) );
  XNOR2_X1 U15233 ( .A(P3_IR_REG_2__SCAN_IN), .B(keyinput108), .ZN(n13174) );
  XNOR2_X1 U15234 ( .A(keyinput68), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n13173) );
  NAND4_X1 U15235 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13177) );
  NOR2_X1 U15236 ( .A1(n13178), .A2(n13177), .ZN(n13185) );
  AOI22_X1 U15237 ( .A1(n10009), .A2(keyinput106), .B1(keyinput99), .B2(n13246), .ZN(n13179) );
  OAI221_X1 U15238 ( .B1(n10009), .B2(keyinput106), .C1(n13246), .C2(
        keyinput99), .A(n13179), .ZN(n13183) );
  INV_X1 U15239 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U15240 ( .A1(n14437), .A2(keyinput123), .B1(n13181), .B2(keyinput86), .ZN(n13180) );
  OAI221_X1 U15241 ( .B1(n14437), .B2(keyinput123), .C1(n13181), .C2(
        keyinput86), .A(n13180), .ZN(n13182) );
  NOR2_X1 U15242 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  AND4_X1 U15243 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13206) );
  AOI22_X1 U15244 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(keyinput88), .B1(
        P3_REG2_REG_23__SCAN_IN), .B2(keyinput126), .ZN(n13188) );
  OAI221_X1 U15245 ( .B1(P1_REG0_REG_8__SCAN_IN), .B2(keyinput88), .C1(
        P3_REG2_REG_23__SCAN_IN), .C2(keyinput126), .A(n13188), .ZN(n13195) );
  AOI22_X1 U15246 ( .A1(P3_REG0_REG_12__SCAN_IN), .A2(keyinput71), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput97), .ZN(n13189) );
  OAI221_X1 U15247 ( .B1(P3_REG0_REG_12__SCAN_IN), .B2(keyinput71), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput97), .A(n13189), .ZN(n13194) );
  AOI22_X1 U15248 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(keyinput73), .B1(
        P3_IR_REG_27__SCAN_IN), .B2(keyinput65), .ZN(n13190) );
  OAI221_X1 U15249 ( .B1(P1_REG0_REG_23__SCAN_IN), .B2(keyinput73), .C1(
        P3_IR_REG_27__SCAN_IN), .C2(keyinput65), .A(n13190), .ZN(n13193) );
  AOI22_X1 U15250 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput76), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput94), .ZN(n13191) );
  OAI221_X1 U15251 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput76), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput94), .A(n13191), .ZN(n13192) );
  NOR4_X1 U15252 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13205) );
  AOI22_X1 U15253 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput113), .B1(
        P3_REG2_REG_4__SCAN_IN), .B2(keyinput125), .ZN(n13196) );
  OAI221_X1 U15254 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput113), .C1(
        P3_REG2_REG_4__SCAN_IN), .C2(keyinput125), .A(n13196), .ZN(n13203) );
  AOI22_X1 U15255 ( .A1(P1_D_REG_22__SCAN_IN), .A2(keyinput109), .B1(SI_9_), 
        .B2(keyinput116), .ZN(n13197) );
  OAI221_X1 U15256 ( .B1(P1_D_REG_22__SCAN_IN), .B2(keyinput109), .C1(SI_9_), 
        .C2(keyinput116), .A(n13197), .ZN(n13202) );
  AOI22_X1 U15257 ( .A1(P1_REG0_REG_31__SCAN_IN), .A2(keyinput90), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput69), .ZN(n13198) );
  OAI221_X1 U15258 ( .B1(P1_REG0_REG_31__SCAN_IN), .B2(keyinput90), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput69), .A(n13198), .ZN(n13201) );
  AOI22_X1 U15259 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(keyinput85), .B1(
        P2_D_REG_6__SCAN_IN), .B2(keyinput100), .ZN(n13199) );
  OAI221_X1 U15260 ( .B1(P1_REG1_REG_21__SCAN_IN), .B2(keyinput85), .C1(
        P2_D_REG_6__SCAN_IN), .C2(keyinput100), .A(n13199), .ZN(n13200) );
  NOR4_X1 U15261 ( .A1(n13203), .A2(n13202), .A3(n13201), .A4(n13200), .ZN(
        n13204) );
  NAND4_X1 U15262 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        n13296) );
  AOI22_X1 U15263 ( .A1(n13210), .A2(keyinput51), .B1(keyinput56), .B2(n13209), 
        .ZN(n13208) );
  OAI221_X1 U15264 ( .B1(n13210), .B2(keyinput51), .C1(n13209), .C2(keyinput56), .A(n13208), .ZN(n13219) );
  INV_X1 U15265 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U15266 ( .A1(n14436), .A2(keyinput45), .B1(keyinput55), .B2(n13212), 
        .ZN(n13211) );
  OAI221_X1 U15267 ( .B1(n14436), .B2(keyinput45), .C1(n13212), .C2(keyinput55), .A(n13211), .ZN(n13218) );
  AOI22_X1 U15268 ( .A1(n13214), .A2(keyinput33), .B1(keyinput59), .B2(n14437), 
        .ZN(n13213) );
  OAI221_X1 U15269 ( .B1(n13214), .B2(keyinput33), .C1(n14437), .C2(keyinput59), .A(n13213), .ZN(n13217) );
  AOI22_X1 U15270 ( .A1(n8870), .A2(keyinput4), .B1(n14281), .B2(keyinput34), 
        .ZN(n13215) );
  OAI221_X1 U15271 ( .B1(n8870), .B2(keyinput4), .C1(n14281), .C2(keyinput34), 
        .A(n13215), .ZN(n13216) );
  NOR4_X1 U15272 ( .A1(n13219), .A2(n13218), .A3(n13217), .A4(n13216), .ZN(
        n13295) );
  AOI22_X1 U15273 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput3), .B1(
        P2_REG0_REG_22__SCAN_IN), .B2(keyinput37), .ZN(n13220) );
  OAI221_X1 U15274 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput3), .C1(
        P2_REG0_REG_22__SCAN_IN), .C2(keyinput37), .A(n13220), .ZN(n13228) );
  AOI22_X1 U15275 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(keyinput60), .B1(
        P3_IR_REG_27__SCAN_IN), .B2(keyinput1), .ZN(n13221) );
  OAI221_X1 U15276 ( .B1(P1_REG0_REG_7__SCAN_IN), .B2(keyinput60), .C1(
        P3_IR_REG_27__SCAN_IN), .C2(keyinput1), .A(n13221), .ZN(n13227) );
  AOI22_X1 U15277 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput20), .B1(n13223), 
        .B2(keyinput49), .ZN(n13222) );
  OAI221_X1 U15278 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput20), .C1(n13223), 
        .C2(keyinput49), .A(n13222), .ZN(n13226) );
  AOI22_X1 U15279 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(keyinput11), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput5), .ZN(n13224) );
  OAI221_X1 U15280 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(keyinput11), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput5), .A(n13224), .ZN(n13225) );
  NOR4_X1 U15281 ( .A1(n13228), .A2(n13227), .A3(n13226), .A4(n13225), .ZN(
        n13294) );
  OAI22_X1 U15282 ( .A1(P3_REG0_REG_12__SCAN_IN), .A2(keyinput7), .B1(
        keyinput23), .B2(P1_D_REG_8__SCAN_IN), .ZN(n13229) );
  AOI221_X1 U15283 ( .B1(P3_REG0_REG_12__SCAN_IN), .B2(keyinput7), .C1(
        P1_D_REG_8__SCAN_IN), .C2(keyinput23), .A(n13229), .ZN(n13236) );
  OAI22_X1 U15284 ( .A1(SI_29_), .A2(keyinput63), .B1(keyinput50), .B2(
        P3_IR_REG_26__SCAN_IN), .ZN(n13230) );
  AOI221_X1 U15285 ( .B1(SI_29_), .B2(keyinput63), .C1(P3_IR_REG_26__SCAN_IN), 
        .C2(keyinput50), .A(n13230), .ZN(n13235) );
  OAI22_X1 U15286 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput19), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput17), .ZN(n13231) );
  AOI221_X1 U15287 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput19), .C1(
        keyinput17), .C2(P1_REG2_REG_1__SCAN_IN), .A(n13231), .ZN(n13234) );
  OAI22_X1 U15288 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput30), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput54), .ZN(n13232) );
  AOI221_X1 U15289 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput30), .C1(
        keyinput54), .C2(P1_IR_REG_23__SCAN_IN), .A(n13232), .ZN(n13233) );
  NAND4_X1 U15290 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13243) );
  AOI22_X1 U15291 ( .A1(n12782), .A2(keyinput12), .B1(keyinput42), .B2(n10009), 
        .ZN(n13237) );
  OAI221_X1 U15292 ( .B1(n12782), .B2(keyinput12), .C1(n10009), .C2(keyinput42), .A(n13237), .ZN(n13242) );
  INV_X1 U15293 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13240) );
  INV_X1 U15294 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U15295 ( .A1(n13240), .A2(keyinput8), .B1(keyinput2), .B2(n13239), 
        .ZN(n13238) );
  OAI221_X1 U15296 ( .B1(n13240), .B2(keyinput8), .C1(n13239), .C2(keyinput2), 
        .A(n13238), .ZN(n13241) );
  NOR3_X1 U15297 ( .A1(n13243), .A2(n13242), .A3(n13241), .ZN(n13292) );
  AOI22_X1 U15298 ( .A1(n13246), .A2(keyinput35), .B1(n13245), .B2(keyinput47), 
        .ZN(n13244) );
  OAI221_X1 U15299 ( .B1(n13246), .B2(keyinput35), .C1(n13245), .C2(keyinput47), .A(n13244), .ZN(n13262) );
  XNOR2_X1 U15300 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput32), .ZN(n13250)
         );
  XNOR2_X1 U15301 ( .A(P1_REG1_REG_22__SCAN_IN), .B(keyinput38), .ZN(n13249)
         );
  XNOR2_X1 U15302 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput40), .ZN(n13248) );
  XNOR2_X1 U15303 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput29), .ZN(n13247) );
  AND4_X1 U15304 ( .A1(n13250), .A2(n13249), .A3(n13248), .A4(n13247), .ZN(
        n13255) );
  XNOR2_X1 U15305 ( .A(keyinput53), .B(n13251), .ZN(n13253) );
  XNOR2_X1 U15306 ( .A(keyinput15), .B(n14771), .ZN(n13252) );
  NOR2_X1 U15307 ( .A1(n13253), .A2(n13252), .ZN(n13254) );
  NAND2_X1 U15308 ( .A1(n13255), .A2(n13254), .ZN(n13261) );
  XNOR2_X1 U15309 ( .A(P3_IR_REG_2__SCAN_IN), .B(keyinput44), .ZN(n13259) );
  XNOR2_X1 U15310 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput0), .ZN(n13258) );
  XNOR2_X1 U15311 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput14), .ZN(n13257) );
  XNOR2_X1 U15312 ( .A(keyinput22), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n13256)
         );
  NAND4_X1 U15313 ( .A1(n13259), .A2(n13258), .A3(n13257), .A4(n13256), .ZN(
        n13260) );
  NOR3_X1 U15314 ( .A1(n13262), .A2(n13261), .A3(n13260), .ZN(n13291) );
  OAI22_X1 U15315 ( .A1(P3_REG2_REG_1__SCAN_IN), .A2(keyinput28), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput58), .ZN(n13263) );
  AOI221_X1 U15316 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(keyinput28), .C1(
        keyinput58), .C2(P1_IR_REG_0__SCAN_IN), .A(n13263), .ZN(n13270) );
  OAI22_X1 U15317 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(keyinput27), .B1(
        P2_REG1_REG_31__SCAN_IN), .B2(keyinput41), .ZN(n13264) );
  AOI221_X1 U15318 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(keyinput27), .C1(
        keyinput41), .C2(P2_REG1_REG_31__SCAN_IN), .A(n13264), .ZN(n13269) );
  OAI22_X1 U15319 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput6), .B1(
        P3_REG2_REG_4__SCAN_IN), .B2(keyinput61), .ZN(n13265) );
  AOI221_X1 U15320 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput6), .C1(keyinput61), 
        .C2(P3_REG2_REG_4__SCAN_IN), .A(n13265), .ZN(n13268) );
  OAI22_X1 U15321 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput36), .B1(keyinput62), 
        .B2(P3_REG2_REG_23__SCAN_IN), .ZN(n13266) );
  AOI221_X1 U15322 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput36), .C1(
        P3_REG2_REG_23__SCAN_IN), .C2(keyinput62), .A(n13266), .ZN(n13267) );
  NAND4_X1 U15323 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        n13280) );
  OAI22_X1 U15324 ( .A1(P2_D_REG_28__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput48), .ZN(n13271) );
  AOI221_X1 U15325 ( .B1(P2_D_REG_28__SCAN_IN), .B2(keyinput10), .C1(
        keyinput48), .C2(P2_REG3_REG_20__SCAN_IN), .A(n13271), .ZN(n13278) );
  OAI22_X1 U15326 ( .A1(P3_REG0_REG_30__SCAN_IN), .A2(keyinput16), .B1(
        keyinput24), .B2(P1_REG0_REG_8__SCAN_IN), .ZN(n13272) );
  AOI221_X1 U15327 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(keyinput16), .C1(
        P1_REG0_REG_8__SCAN_IN), .C2(keyinput24), .A(n13272), .ZN(n13277) );
  OAI22_X1 U15328 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(keyinput39), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(keyinput46), .ZN(n13273) );
  AOI221_X1 U15329 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(keyinput39), .C1(
        keyinput46), .C2(P3_DATAO_REG_29__SCAN_IN), .A(n13273), .ZN(n13276) );
  OAI22_X1 U15330 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput43), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput18), .ZN(n13274) );
  AOI221_X1 U15331 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput43), .C1(
        keyinput18), .C2(P1_REG3_REG_23__SCAN_IN), .A(n13274), .ZN(n13275) );
  NAND4_X1 U15332 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13279) );
  NOR2_X1 U15333 ( .A1(n13280), .A2(n13279), .ZN(n13290) );
  OAI22_X1 U15334 ( .A1(SI_9_), .A2(keyinput52), .B1(keyinput26), .B2(
        P1_REG0_REG_31__SCAN_IN), .ZN(n13281) );
  AOI221_X1 U15335 ( .B1(SI_9_), .B2(keyinput52), .C1(P1_REG0_REG_31__SCAN_IN), 
        .C2(keyinput26), .A(n13281), .ZN(n13288) );
  OAI22_X1 U15336 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput13), .B1(keyinput9), 
        .B2(P1_REG0_REG_23__SCAN_IN), .ZN(n13282) );
  AOI221_X1 U15337 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput13), .C1(
        P1_REG0_REG_23__SCAN_IN), .C2(keyinput9), .A(n13282), .ZN(n13287) );
  OAI22_X1 U15338 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(keyinput57), .B1(
        keyinput31), .B2(P2_ADDR_REG_17__SCAN_IN), .ZN(n13283) );
  AOI221_X1 U15339 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(keyinput57), .C1(
        P2_ADDR_REG_17__SCAN_IN), .C2(keyinput31), .A(n13283), .ZN(n13286) );
  OAI22_X1 U15340 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(keyinput25), .B1(
        keyinput21), .B2(P1_REG1_REG_21__SCAN_IN), .ZN(n13284) );
  AOI221_X1 U15341 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput21), .A(n13284), .ZN(n13285) );
  AND4_X1 U15342 ( .A1(n13288), .A2(n13287), .A3(n13286), .A4(n13285), .ZN(
        n13289) );
  AND4_X1 U15343 ( .A1(n13292), .A2(n13291), .A3(n13290), .A4(n13289), .ZN(
        n13293) );
  NAND4_X1 U15344 ( .A1(n13296), .A2(n13295), .A3(n13294), .A4(n13293), .ZN(
        n13305) );
  OAI22_X1 U15345 ( .A1(n13531), .A2(n14013), .B1(n13982), .B2(n14015), .ZN(
        n14115) );
  NAND2_X1 U15346 ( .A1(n14115), .A2(n14373), .ZN(n13297) );
  NAND2_X1 U15347 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13778)
         );
  OAI211_X1 U15348 ( .C1(n14376), .C2(n13954), .A(n13297), .B(n13778), .ZN(
        n13303) );
  INV_X1 U15349 ( .A(n13298), .ZN(n13299) );
  AOI211_X1 U15350 ( .C1(n13301), .C2(n13300), .A(n13425), .B(n13299), .ZN(
        n13302) );
  AOI211_X1 U15351 ( .C1(n14300), .C2(n14116), .A(n13303), .B(n13302), .ZN(
        n13304) );
  XOR2_X1 U15352 ( .A(n13305), .B(n13304), .Z(P1_U3219) );
  INV_X1 U15353 ( .A(n13306), .ZN(n13307) );
  AOI22_X1 U15354 ( .A1(n14058), .A2(n13311), .B1(n9725), .B2(n13798), .ZN(
        n13312) );
  XNOR2_X1 U15355 ( .A(n13312), .B(n13022), .ZN(n13315) );
  AOI22_X1 U15356 ( .A1(n14058), .A2(n9725), .B1(n13313), .B2(n13798), .ZN(
        n13314) );
  XNOR2_X1 U15357 ( .A(n13315), .B(n13314), .ZN(n13316) );
  XNOR2_X1 U15358 ( .A(n13317), .B(n13316), .ZN(n13325) );
  INV_X1 U15359 ( .A(n13318), .ZN(n13320) );
  OAI22_X1 U15360 ( .A1(n14376), .A2(n13320), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13319), .ZN(n13323) );
  INV_X1 U15361 ( .A(n13650), .ZN(n13607) );
  OAI22_X1 U15362 ( .A1(n13607), .A2(n13400), .B1(n13321), .B2(n13399), .ZN(
        n13322) );
  AOI211_X1 U15363 ( .C1(n14058), .C2(n14300), .A(n13323), .B(n13322), .ZN(
        n13324) );
  OAI21_X1 U15364 ( .B1(n13325), .B2(n13425), .A(n13324), .ZN(P1_U3220) );
  INV_X1 U15365 ( .A(n13326), .ZN(n13327) );
  AOI21_X1 U15366 ( .B1(n13329), .B2(n13328), .A(n13327), .ZN(n13335) );
  AND2_X1 U15367 ( .A1(n13653), .A2(n14416), .ZN(n13330) );
  AOI21_X1 U15368 ( .B1(n13651), .B2(n14413), .A(n13330), .ZN(n14099) );
  AOI22_X1 U15369 ( .A1(n13926), .A2(n13403), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13331) );
  OAI21_X1 U15370 ( .B1(n14099), .B2(n13332), .A(n13331), .ZN(n13333) );
  AOI21_X1 U15371 ( .B1(n13923), .B2(n14300), .A(n13333), .ZN(n13334) );
  OAI21_X1 U15372 ( .B1(n13335), .B2(n13425), .A(n13334), .ZN(P1_U3223) );
  XOR2_X1 U15373 ( .A(n13337), .B(n13336), .Z(n13345) );
  INV_X1 U15374 ( .A(n13338), .ZN(n13862) );
  OAI22_X1 U15375 ( .A1(n14376), .A2(n13862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13339), .ZN(n13343) );
  OAI22_X1 U15376 ( .A1(n13341), .A2(n13400), .B1(n13340), .B2(n13399), .ZN(
        n13342) );
  AOI211_X1 U15377 ( .C1(n14074), .C2(n14300), .A(n13343), .B(n13342), .ZN(
        n13344) );
  OAI21_X1 U15378 ( .B1(n13345), .B2(n13425), .A(n13344), .ZN(P1_U3225) );
  OAI21_X1 U15379 ( .B1(n13348), .B2(n13347), .A(n13346), .ZN(n13355) );
  INV_X1 U15380 ( .A(n14005), .ZN(n13350) );
  OAI21_X1 U15381 ( .B1(n14376), .B2(n13350), .A(n13349), .ZN(n13351) );
  INV_X1 U15382 ( .A(n13351), .ZN(n13353) );
  INV_X1 U15383 ( .A(n14001), .ZN(n13656) );
  AOI22_X1 U15384 ( .A1(n13656), .A2(n13419), .B1(n13420), .B2(n13966), .ZN(
        n13352) );
  OAI211_X1 U15385 ( .C1(n14008), .C2(n13393), .A(n13353), .B(n13352), .ZN(
        n13354) );
  AOI21_X1 U15386 ( .B1(n13355), .B2(n14366), .A(n13354), .ZN(n13356) );
  INV_X1 U15387 ( .A(n13356), .ZN(P1_U3226) );
  INV_X1 U15388 ( .A(n13357), .ZN(n13362) );
  AOI21_X1 U15389 ( .B1(n13359), .B2(n13361), .A(n13358), .ZN(n13360) );
  AOI21_X1 U15390 ( .B1(n13362), .B2(n13361), .A(n13360), .ZN(n13367) );
  AOI22_X1 U15391 ( .A1(n13655), .A2(n13419), .B1(n13420), .B2(n13654), .ZN(
        n13363) );
  NAND2_X1 U15392 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13734)
         );
  OAI211_X1 U15393 ( .C1(n14376), .C2(n13364), .A(n13363), .B(n13734), .ZN(
        n13365) );
  AOI21_X1 U15394 ( .B1(n14126), .B2(n14300), .A(n13365), .ZN(n13366) );
  OAI21_X1 U15395 ( .B1(n13367), .B2(n13425), .A(n13366), .ZN(P1_U3228) );
  XOR2_X1 U15396 ( .A(n13369), .B(n13368), .Z(n13375) );
  NAND2_X1 U15397 ( .A1(n13876), .A2(n13419), .ZN(n13371) );
  AOI22_X1 U15398 ( .A1(n13403), .A2(n13882), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13370) );
  OAI211_X1 U15399 ( .C1(n13372), .C2(n13400), .A(n13371), .B(n13370), .ZN(
        n13373) );
  AOI21_X1 U15400 ( .B1(n14083), .B2(n14300), .A(n13373), .ZN(n13374) );
  OAI21_X1 U15401 ( .B1(n13375), .B2(n13425), .A(n13374), .ZN(P1_U3229) );
  OAI211_X1 U15402 ( .C1(n13378), .C2(n13377), .A(n13376), .B(n14366), .ZN(
        n13382) );
  OAI22_X1 U15403 ( .A1(n13387), .A2(n14013), .B1(n13401), .B2(n14015), .ZN(
        n13941) );
  OAI22_X1 U15404 ( .A1(n13942), .A2(n14376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13379), .ZN(n13380) );
  AOI21_X1 U15405 ( .B1(n13941), .B2(n14373), .A(n13380), .ZN(n13381) );
  OAI211_X1 U15406 ( .C1(n14108), .C2(n13393), .A(n13382), .B(n13381), .ZN(
        P1_U3233) );
  OAI21_X1 U15407 ( .B1(n13385), .B2(n13384), .A(n13383), .ZN(n13386) );
  NAND2_X1 U15408 ( .A1(n13386), .A2(n14366), .ZN(n13392) );
  OAI22_X1 U15409 ( .A1(n13388), .A2(n14013), .B1(n13387), .B2(n14015), .ZN(
        n14093) );
  INV_X1 U15410 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13389) );
  OAI22_X1 U15411 ( .A1(n13911), .A2(n14376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13389), .ZN(n13390) );
  AOI21_X1 U15412 ( .B1(n14093), .B2(n14373), .A(n13390), .ZN(n13391) );
  OAI211_X1 U15413 ( .C1(n13393), .C2(n13915), .A(n13392), .B(n13391), .ZN(
        P1_U3235) );
  INV_X1 U15414 ( .A(n14364), .ZN(n13413) );
  NAND2_X1 U15415 ( .A1(n13972), .A2(n14499), .ZN(n14122) );
  OAI21_X1 U15416 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(n13397) );
  NAND2_X1 U15417 ( .A1(n13397), .A2(n14366), .ZN(n13405) );
  INV_X1 U15418 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n13398) );
  NOR2_X1 U15419 ( .A1(n13398), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13745) );
  OAI22_X1 U15420 ( .A1(n13401), .A2(n13400), .B1(n14002), .B2(n13399), .ZN(
        n13402) );
  AOI211_X1 U15421 ( .C1(n13403), .C2(n13971), .A(n13745), .B(n13402), .ZN(
        n13404) );
  OAI211_X1 U15422 ( .C1(n13413), .C2(n14122), .A(n13405), .B(n13404), .ZN(
        P1_U3238) );
  XNOR2_X1 U15423 ( .A(n13407), .B(n13406), .ZN(n13415) );
  NAND2_X1 U15424 ( .A1(n13839), .A2(n14499), .ZN(n14070) );
  INV_X1 U15425 ( .A(n13842), .ZN(n13409) );
  OAI22_X1 U15426 ( .A1(n14376), .A2(n13409), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13408), .ZN(n13410) );
  INV_X1 U15427 ( .A(n13410), .ZN(n13412) );
  AOI22_X1 U15428 ( .A1(n13420), .A2(n13835), .B1(n13419), .B2(n13875), .ZN(
        n13411) );
  OAI211_X1 U15429 ( .C1(n14070), .C2(n13413), .A(n13412), .B(n13411), .ZN(
        n13414) );
  AOI21_X1 U15430 ( .B1(n13415), .B2(n14366), .A(n13414), .ZN(n13416) );
  INV_X1 U15431 ( .A(n13416), .ZN(P1_U3240) );
  XNOR2_X1 U15432 ( .A(n13418), .B(n13417), .ZN(n13426) );
  INV_X1 U15433 ( .A(n14019), .ZN(n13422) );
  AOI22_X1 U15434 ( .A1(n13420), .A2(n13655), .B1(n13657), .B2(n13419), .ZN(
        n13421) );
  NAND2_X1 U15435 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14389)
         );
  OAI211_X1 U15436 ( .C1(n13422), .C2(n14376), .A(n13421), .B(n14389), .ZN(
        n13423) );
  AOI21_X1 U15437 ( .B1(n14307), .B2(n14300), .A(n13423), .ZN(n13424) );
  OAI21_X1 U15438 ( .B1(n13426), .B2(n13425), .A(n13424), .ZN(P1_U3241) );
  NAND2_X1 U15439 ( .A1(n13428), .A2(n13427), .ZN(n13429) );
  NAND2_X1 U15440 ( .A1(n13429), .A2(n13605), .ZN(n13585) );
  AOI21_X1 U15441 ( .B1(n9226), .B2(n13600), .A(n13432), .ZN(n13443) );
  NAND3_X1 U15442 ( .A1(n13437), .A2(n13436), .A3(n13435), .ZN(n13442) );
  INV_X1 U15443 ( .A(n13438), .ZN(n13440) );
  NAND3_X1 U15444 ( .A1(n13440), .A2(n6477), .A3(n13439), .ZN(n13441) );
  OAI211_X1 U15445 ( .C1(n13444), .C2(n13443), .A(n13442), .B(n13441), .ZN(
        n13445) );
  NAND2_X1 U15446 ( .A1(n13445), .A2(n13610), .ZN(n13449) );
  MUX2_X1 U15447 ( .A(n13447), .B(n13446), .S(n6477), .Z(n13448) );
  NAND3_X1 U15448 ( .A1(n13449), .A2(n13616), .A3(n13448), .ZN(n13453) );
  NAND2_X1 U15449 ( .A1(n14363), .A2(n13600), .ZN(n13451) );
  NAND2_X1 U15450 ( .A1(n6747), .A2(n6477), .ZN(n13450) );
  MUX2_X1 U15451 ( .A(n13451), .B(n13450), .S(n14415), .Z(n13452) );
  NAND2_X1 U15452 ( .A1(n13453), .A2(n13452), .ZN(n13457) );
  MUX2_X1 U15453 ( .A(n13454), .B(n14461), .S(n6477), .Z(n13456) );
  MUX2_X1 U15454 ( .A(n13608), .B(n13666), .S(n6477), .Z(n13455) );
  OAI21_X1 U15455 ( .B1(n13457), .B2(n13456), .A(n13455), .ZN(n13459) );
  NAND2_X1 U15456 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  NAND2_X1 U15457 ( .A1(n13459), .A2(n13458), .ZN(n13461) );
  MUX2_X1 U15458 ( .A(n14414), .B(n14468), .S(n13600), .Z(n13462) );
  MUX2_X1 U15459 ( .A(n14414), .B(n14468), .S(n6477), .Z(n13460) );
  INV_X1 U15460 ( .A(n13462), .ZN(n13463) );
  MUX2_X1 U15461 ( .A(n13665), .B(n13464), .S(n6477), .Z(n13467) );
  MUX2_X1 U15462 ( .A(n13665), .B(n13464), .S(n13600), .Z(n13465) );
  MUX2_X1 U15463 ( .A(n13664), .B(n14484), .S(n13600), .Z(n13470) );
  MUX2_X1 U15464 ( .A(n13664), .B(n14484), .S(n6477), .Z(n13468) );
  INV_X1 U15465 ( .A(n13470), .ZN(n13471) );
  MUX2_X1 U15466 ( .A(n13663), .B(n13472), .S(n6477), .Z(n13476) );
  MUX2_X1 U15467 ( .A(n13472), .B(n13663), .S(n6477), .Z(n13473) );
  NAND2_X1 U15468 ( .A1(n13474), .A2(n13473), .ZN(n13479) );
  INV_X1 U15469 ( .A(n13475), .ZN(n13477) );
  NAND2_X1 U15470 ( .A1(n13477), .A2(n7268), .ZN(n13478) );
  MUX2_X1 U15471 ( .A(n13662), .B(n14498), .S(n13600), .Z(n13481) );
  MUX2_X1 U15472 ( .A(n13662), .B(n14498), .S(n6477), .Z(n13480) );
  MUX2_X1 U15473 ( .A(n13661), .B(n13482), .S(n6477), .Z(n13484) );
  MUX2_X1 U15474 ( .A(n13661), .B(n13482), .S(n13600), .Z(n13483) );
  INV_X1 U15475 ( .A(n13484), .ZN(n13485) );
  MUX2_X1 U15476 ( .A(n13660), .B(n14301), .S(n13600), .Z(n13488) );
  MUX2_X1 U15477 ( .A(n13660), .B(n14301), .S(n6477), .Z(n13486) );
  INV_X1 U15478 ( .A(n13488), .ZN(n13489) );
  MUX2_X1 U15479 ( .A(n13659), .B(n13490), .S(n6477), .Z(n13494) );
  MUX2_X1 U15480 ( .A(n13659), .B(n13490), .S(n13600), .Z(n13491) );
  NAND2_X1 U15481 ( .A1(n13492), .A2(n13491), .ZN(n13498) );
  INV_X1 U15482 ( .A(n13493), .ZN(n13496) );
  INV_X1 U15483 ( .A(n13494), .ZN(n13495) );
  NAND2_X1 U15484 ( .A1(n13496), .A2(n13495), .ZN(n13497) );
  MUX2_X1 U15485 ( .A(n13658), .B(n13499), .S(n13600), .Z(n13502) );
  MUX2_X1 U15486 ( .A(n13658), .B(n13499), .S(n6477), .Z(n13500) );
  INV_X1 U15487 ( .A(n13502), .ZN(n13503) );
  NAND2_X1 U15488 ( .A1(n13509), .A2(n13505), .ZN(n13507) );
  OAI21_X1 U15489 ( .B1(n14315), .B2(n13657), .A(n13508), .ZN(n13506) );
  MUX2_X1 U15490 ( .A(n13507), .B(n13506), .S(n6477), .Z(n13511) );
  MUX2_X1 U15491 ( .A(n13509), .B(n13508), .S(n13600), .Z(n13510) );
  MUX2_X1 U15492 ( .A(n14014), .B(n14008), .S(n13600), .Z(n13515) );
  MUX2_X1 U15493 ( .A(n13655), .B(n14132), .S(n6477), .Z(n13514) );
  NAND2_X1 U15494 ( .A1(n13515), .A2(n13514), .ZN(n13512) );
  NAND4_X1 U15495 ( .A1(n13513), .A2(n13967), .A3(n13512), .A4(n13977), .ZN(
        n13526) );
  MUX2_X1 U15496 ( .A(n13966), .B(n14126), .S(n6477), .Z(n13519) );
  INV_X1 U15497 ( .A(n13514), .ZN(n13517) );
  INV_X1 U15498 ( .A(n13515), .ZN(n13516) );
  NAND3_X1 U15499 ( .A1(n13977), .A2(n13517), .A3(n13516), .ZN(n13518) );
  OAI21_X1 U15500 ( .B1(n13520), .B2(n13519), .A(n13518), .ZN(n13521) );
  NAND2_X1 U15501 ( .A1(n13967), .A2(n13521), .ZN(n13525) );
  NAND2_X1 U15502 ( .A1(n13972), .A2(n13600), .ZN(n13523) );
  OR2_X1 U15503 ( .A1(n13972), .A2(n13600), .ZN(n13522) );
  MUX2_X1 U15504 ( .A(n13523), .B(n13522), .S(n13654), .Z(n13524) );
  NAND2_X1 U15505 ( .A1(n13526), .A2(n7522), .ZN(n13530) );
  NAND2_X1 U15506 ( .A1(n14116), .A2(n6477), .ZN(n13528) );
  OR2_X1 U15507 ( .A1(n14116), .A2(n6477), .ZN(n13527) );
  MUX2_X1 U15508 ( .A(n13528), .B(n13527), .S(n13965), .Z(n13529) );
  NAND2_X1 U15509 ( .A1(n13530), .A2(n13529), .ZN(n13534) );
  MUX2_X1 U15510 ( .A(n13531), .B(n14108), .S(n13600), .Z(n13533) );
  MUX2_X1 U15511 ( .A(n13653), .B(n13946), .S(n6477), .Z(n13532) );
  OAI21_X1 U15512 ( .B1(n13534), .B2(n13533), .A(n13532), .ZN(n13536) );
  NAND2_X1 U15513 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  MUX2_X1 U15514 ( .A(n13652), .B(n13923), .S(n6477), .Z(n13538) );
  MUX2_X1 U15515 ( .A(n13652), .B(n13923), .S(n13600), .Z(n13537) );
  MUX2_X1 U15516 ( .A(n13651), .B(n14094), .S(n13600), .Z(n13541) );
  MUX2_X1 U15517 ( .A(n13651), .B(n14094), .S(n6477), .Z(n13539) );
  INV_X1 U15518 ( .A(n13541), .ZN(n13542) );
  MUX2_X1 U15519 ( .A(n13876), .B(n14087), .S(n6477), .Z(n13545) );
  MUX2_X1 U15520 ( .A(n13876), .B(n14087), .S(n13600), .Z(n13543) );
  MUX2_X1 U15521 ( .A(n13858), .B(n14083), .S(n13600), .Z(n13548) );
  MUX2_X1 U15522 ( .A(n13858), .B(n14083), .S(n6477), .Z(n13546) );
  INV_X1 U15523 ( .A(n13548), .ZN(n13549) );
  MUX2_X1 U15524 ( .A(n13875), .B(n14074), .S(n6477), .Z(n13552) );
  MUX2_X1 U15525 ( .A(n13875), .B(n14074), .S(n13600), .Z(n13550) );
  NAND2_X1 U15526 ( .A1(n13551), .A2(n13550), .ZN(n13555) );
  INV_X1 U15527 ( .A(n13552), .ZN(n13553) );
  NAND2_X1 U15528 ( .A1(n6574), .A2(n13553), .ZN(n13554) );
  MUX2_X1 U15529 ( .A(n13859), .B(n13839), .S(n13600), .Z(n13557) );
  MUX2_X1 U15530 ( .A(n13859), .B(n13839), .S(n6477), .Z(n13556) );
  INV_X1 U15531 ( .A(n13557), .ZN(n13558) );
  MUX2_X1 U15532 ( .A(n13835), .B(n14063), .S(n6477), .Z(n13560) );
  MUX2_X1 U15533 ( .A(n14063), .B(n13835), .S(n6477), .Z(n13559) );
  MUX2_X1 U15534 ( .A(n13798), .B(n14058), .S(n13600), .Z(n13562) );
  MUX2_X1 U15535 ( .A(n13798), .B(n14058), .S(n6477), .Z(n13561) );
  NAND2_X1 U15536 ( .A1(n13563), .A2(n13595), .ZN(n13565) );
  OR2_X1 U15537 ( .A1(n13574), .A2(n14160), .ZN(n13564) );
  MUX2_X1 U15538 ( .A(n13650), .B(n14049), .S(n6477), .Z(n13567) );
  NAND2_X1 U15539 ( .A1(n13566), .A2(n13567), .ZN(n13571) );
  MUX2_X1 U15540 ( .A(n14049), .B(n13650), .S(n6477), .Z(n13570) );
  INV_X1 U15541 ( .A(n13566), .ZN(n13569) );
  INV_X1 U15542 ( .A(n13567), .ZN(n13568) );
  NAND2_X1 U15543 ( .A1(n13572), .A2(n13595), .ZN(n13576) );
  OR2_X1 U15544 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  INV_X1 U15545 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U15546 ( .A1(n9739), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U15547 ( .A1(n8606), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n13577) );
  OAI211_X1 U15548 ( .C1(n9795), .C2(n13788), .A(n13578), .B(n13577), .ZN(
        n13804) );
  INV_X1 U15549 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n13583) );
  NAND2_X1 U15550 ( .A1(n13579), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n13582) );
  NAND2_X1 U15551 ( .A1(n13580), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13581) );
  OAI211_X1 U15552 ( .C1(n13584), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13782) );
  INV_X1 U15553 ( .A(n13782), .ZN(n13601) );
  OAI21_X1 U15554 ( .B1(n13601), .B2(n13600), .A(n13585), .ZN(n13586) );
  AOI22_X1 U15555 ( .A1(n13791), .A2(n13600), .B1(n13804), .B2(n13586), .ZN(
        n13592) );
  OAI21_X1 U15556 ( .B1(n13782), .B2(n13587), .A(n13804), .ZN(n13588) );
  INV_X1 U15557 ( .A(n13588), .ZN(n13589) );
  MUX2_X1 U15558 ( .A(n13589), .B(n13791), .S(n6477), .Z(n13590) );
  INV_X1 U15559 ( .A(n13592), .ZN(n13593) );
  XNOR2_X1 U15560 ( .A(n14041), .B(n13782), .ZN(n13634) );
  NAND2_X1 U15561 ( .A1(n13597), .A2(n13596), .ZN(n13599) );
  NAND2_X1 U15562 ( .A1(n13599), .A2(n13598), .ZN(n13606) );
  NOR2_X1 U15563 ( .A1(n13782), .A2(n13600), .ZN(n13603) );
  NOR2_X1 U15564 ( .A1(n13601), .A2(n6477), .ZN(n13602) );
  MUX2_X1 U15565 ( .A(n13603), .B(n13602), .S(n14041), .Z(n13637) );
  NAND2_X1 U15566 ( .A1(n13605), .A2(n13604), .ZN(n13636) );
  NAND2_X1 U15567 ( .A1(n13606), .A2(n13636), .ZN(n13643) );
  XOR2_X1 U15568 ( .A(n13804), .B(n13791), .Z(n13633) );
  XNOR2_X1 U15569 ( .A(n14049), .B(n13607), .ZN(n13795) );
  XNOR2_X1 U15570 ( .A(n13666), .B(n13608), .ZN(n14425) );
  NAND4_X1 U15571 ( .A1(n13610), .A2(n14029), .A3(n13609), .A4(n14425), .ZN(
        n13612) );
  NOR3_X1 U15572 ( .A1(n13612), .A2(n14396), .A3(n13611), .ZN(n13615) );
  NAND4_X1 U15573 ( .A1(n13616), .A2(n13615), .A3(n13614), .A4(n13613), .ZN(
        n13618) );
  NOR2_X1 U15574 ( .A1(n13618), .A2(n13617), .ZN(n13621) );
  NAND4_X1 U15575 ( .A1(n13622), .A2(n13621), .A3(n13620), .A4(n13619), .ZN(
        n13623) );
  NOR2_X1 U15576 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  AND4_X1 U15577 ( .A1(n13977), .A2(n14024), .A3(n13625), .A4(n7255), .ZN(
        n13627) );
  NAND4_X1 U15578 ( .A1(n13950), .A2(n13627), .A3(n13967), .A4(n13626), .ZN(
        n13628) );
  OR4_X1 U15579 ( .A1(n13907), .A2(n13939), .A3(n13921), .A4(n13628), .ZN(
        n13629) );
  NOR4_X1 U15580 ( .A1(n13852), .A2(n13871), .A3(n13890), .A4(n13629), .ZN(
        n13630) );
  NAND4_X1 U15581 ( .A1(n13631), .A2(n13822), .A3(n13838), .A4(n13630), .ZN(
        n13632) );
  XNOR2_X1 U15582 ( .A(n13635), .B(n13928), .ZN(n13641) );
  INV_X1 U15583 ( .A(n13636), .ZN(n13640) );
  INV_X1 U15584 ( .A(n13637), .ZN(n13638) );
  NOR2_X1 U15585 ( .A1(n13638), .A2(n13643), .ZN(n13639) );
  AOI211_X1 U15586 ( .C1(n13641), .C2(n13640), .A(n13639), .B(n13645), .ZN(
        n13642) );
  OAI21_X1 U15587 ( .B1(n13644), .B2(n13643), .A(n13642), .ZN(n13648) );
  NOR3_X1 U15588 ( .A1(n14136), .A2(n14163), .A3(n14015), .ZN(n13647) );
  OAI21_X1 U15589 ( .B1(n13645), .B2(n8661), .A(P1_B_REG_SCAN_IN), .ZN(n13646)
         );
  OAI22_X1 U15590 ( .A1(n13649), .A2(n13648), .B1(n13647), .B2(n13646), .ZN(
        P1_U3242) );
  MUX2_X1 U15591 ( .A(n13782), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13668), .Z(
        P1_U3591) );
  MUX2_X1 U15592 ( .A(n13804), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13668), .Z(
        P1_U3590) );
  MUX2_X1 U15593 ( .A(n13650), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13668), .Z(
        P1_U3589) );
  MUX2_X1 U15594 ( .A(n13798), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13668), .Z(
        P1_U3588) );
  MUX2_X1 U15595 ( .A(n13835), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13668), .Z(
        P1_U3587) );
  MUX2_X1 U15596 ( .A(n13859), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13668), .Z(
        P1_U3586) );
  MUX2_X1 U15597 ( .A(n13875), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13668), .Z(
        P1_U3585) );
  MUX2_X1 U15598 ( .A(n13858), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13668), .Z(
        P1_U3584) );
  MUX2_X1 U15599 ( .A(n13876), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13668), .Z(
        P1_U3583) );
  MUX2_X1 U15600 ( .A(n13651), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13668), .Z(
        P1_U3582) );
  MUX2_X1 U15601 ( .A(n13652), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13668), .Z(
        P1_U3581) );
  MUX2_X1 U15602 ( .A(n13653), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13668), .Z(
        P1_U3580) );
  MUX2_X1 U15603 ( .A(n13965), .B(P1_DATAO_REG_19__SCAN_IN), .S(n13668), .Z(
        P1_U3579) );
  MUX2_X1 U15604 ( .A(n13654), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13668), .Z(
        P1_U3578) );
  MUX2_X1 U15605 ( .A(n13966), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13668), .Z(
        P1_U3577) );
  MUX2_X1 U15606 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13655), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15607 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13656), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15608 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13657), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15609 ( .A(n13658), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13668), .Z(
        P1_U3573) );
  MUX2_X1 U15610 ( .A(n13659), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13668), .Z(
        P1_U3572) );
  MUX2_X1 U15611 ( .A(n13660), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13668), .Z(
        P1_U3571) );
  MUX2_X1 U15612 ( .A(n13661), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13668), .Z(
        P1_U3570) );
  MUX2_X1 U15613 ( .A(n13662), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13668), .Z(
        P1_U3569) );
  MUX2_X1 U15614 ( .A(n13663), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13668), .Z(
        P1_U3568) );
  MUX2_X1 U15615 ( .A(n13664), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13668), .Z(
        P1_U3567) );
  MUX2_X1 U15616 ( .A(n13665), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13668), .Z(
        P1_U3566) );
  MUX2_X1 U15617 ( .A(n14414), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13668), .Z(
        P1_U3565) );
  MUX2_X1 U15618 ( .A(n13666), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13668), .Z(
        P1_U3564) );
  MUX2_X1 U15619 ( .A(n14415), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13668), .Z(
        P1_U3563) );
  MUX2_X1 U15620 ( .A(n13667), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13668), .Z(
        P1_U3562) );
  MUX2_X1 U15621 ( .A(n9226), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13668), .Z(
        P1_U3561) );
  NAND2_X1 U15622 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13672) );
  INV_X1 U15623 ( .A(n13669), .ZN(n13671) );
  AOI211_X1 U15624 ( .C1(n13672), .C2(n13671), .A(n13670), .B(n13737), .ZN(
        n13673) );
  INV_X1 U15625 ( .A(n13673), .ZN(n13682) );
  INV_X1 U15626 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13674) );
  OAI22_X1 U15627 ( .A1(n14391), .A2(n8418), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13674), .ZN(n13675) );
  AOI21_X1 U15628 ( .B1(n13676), .B2(n14383), .A(n13675), .ZN(n13681) );
  OAI211_X1 U15629 ( .C1(n13679), .C2(n13678), .A(n14387), .B(n13677), .ZN(
        n13680) );
  NAND3_X1 U15630 ( .A1(n13682), .A2(n13681), .A3(n13680), .ZN(P1_U3244) );
  OAI21_X1 U15631 ( .B1(n13685), .B2(n13684), .A(n13683), .ZN(n13686) );
  NAND2_X1 U15632 ( .A1(n13686), .A2(n14386), .ZN(n13699) );
  INV_X1 U15633 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13688) );
  OAI21_X1 U15634 ( .B1(n14391), .B2(n13688), .A(n13687), .ZN(n13689) );
  AOI21_X1 U15635 ( .B1(n13690), .B2(n14383), .A(n13689), .ZN(n13698) );
  MUX2_X1 U15636 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9818), .S(n13691), .Z(
        n13692) );
  NAND3_X1 U15637 ( .A1(n13694), .A2(n13693), .A3(n13692), .ZN(n13695) );
  NAND3_X1 U15638 ( .A1(n14387), .A2(n13696), .A3(n13695), .ZN(n13697) );
  NAND3_X1 U15639 ( .A1(n13699), .A2(n13698), .A3(n13697), .ZN(P1_U3248) );
  OAI21_X1 U15640 ( .B1(n13702), .B2(n13701), .A(n13700), .ZN(n13703) );
  NAND2_X1 U15641 ( .A1(n13703), .A2(n14386), .ZN(n13713) );
  AOI21_X1 U15642 ( .B1(n13746), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n13704), .ZN(
        n13712) );
  MUX2_X1 U15643 ( .A(n9199), .B(P1_REG2_REG_8__SCAN_IN), .S(n13709), .Z(
        n13705) );
  NAND3_X1 U15644 ( .A1(n13707), .A2(n13706), .A3(n13705), .ZN(n13708) );
  NAND3_X1 U15645 ( .A1(n14387), .A2(n13722), .A3(n13708), .ZN(n13711) );
  NAND2_X1 U15646 ( .A1(n14383), .A2(n13709), .ZN(n13710) );
  NAND4_X1 U15647 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        P1_U3251) );
  OAI21_X1 U15648 ( .B1(n13716), .B2(n13715), .A(n13714), .ZN(n13717) );
  NAND2_X1 U15649 ( .A1(n13717), .A2(n14386), .ZN(n13729) );
  INV_X1 U15650 ( .A(n13718), .ZN(n13719) );
  AOI21_X1 U15651 ( .B1(n13746), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n13719), .ZN(
        n13728) );
  MUX2_X1 U15652 ( .A(n9202), .B(P1_REG2_REG_9__SCAN_IN), .S(n13725), .Z(
        n13720) );
  NAND3_X1 U15653 ( .A1(n13722), .A2(n13721), .A3(n13720), .ZN(n13723) );
  NAND3_X1 U15654 ( .A1(n14387), .A2(n13724), .A3(n13723), .ZN(n13727) );
  NAND2_X1 U15655 ( .A1(n14383), .A2(n13725), .ZN(n13726) );
  NAND4_X1 U15656 ( .A1(n13729), .A2(n13728), .A3(n13727), .A4(n13726), .ZN(
        P1_U3252) );
  NAND2_X1 U15657 ( .A1(n13731), .A2(n13730), .ZN(n13733) );
  XNOR2_X1 U15658 ( .A(n13748), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U15659 ( .A1(n13732), .A2(n13733), .ZN(n13747) );
  OAI211_X1 U15660 ( .C1(n13733), .C2(n13732), .A(n14387), .B(n13747), .ZN(
        n13743) );
  OAI21_X1 U15661 ( .B1(n14391), .B2(n8450), .A(n13734), .ZN(n13741) );
  XNOR2_X1 U15662 ( .A(n13752), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13738) );
  AOI211_X1 U15663 ( .C1(n13739), .C2(n13738), .A(n13751), .B(n13737), .ZN(
        n13740) );
  AOI211_X1 U15664 ( .C1(n14383), .C2(n13752), .A(n13741), .B(n13740), .ZN(
        n13742) );
  NAND2_X1 U15665 ( .A1(n13743), .A2(n13742), .ZN(P1_U3260) );
  NOR2_X1 U15666 ( .A1(n13772), .A2(n13760), .ZN(n13744) );
  AOI211_X1 U15667 ( .C1(n13746), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n13745), 
        .B(n13744), .ZN(n13759) );
  INV_X1 U15668 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13749) );
  OAI21_X1 U15669 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13766) );
  XNOR2_X1 U15670 ( .A(n13760), .B(n13766), .ZN(n13750) );
  NAND2_X1 U15671 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13750), .ZN(n13769) );
  OAI211_X1 U15672 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13750), .A(n14387), 
        .B(n13769), .ZN(n13758) );
  INV_X1 U15673 ( .A(n13753), .ZN(n13756) );
  INV_X1 U15674 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13754) );
  NOR2_X1 U15675 ( .A1(n13754), .A2(n13753), .ZN(n13762) );
  INV_X1 U15676 ( .A(n13762), .ZN(n13755) );
  OAI211_X1 U15677 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13756), .A(n14386), 
        .B(n13755), .ZN(n13757) );
  NAND3_X1 U15678 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(P1_U3261) );
  NOR2_X1 U15679 ( .A1(n13761), .A2(n13760), .ZN(n13763) );
  NOR2_X1 U15680 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  NAND2_X1 U15681 ( .A1(n13767), .A2(n13766), .ZN(n13768) );
  NAND2_X1 U15682 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  XOR2_X1 U15683 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13770), .Z(n13774) );
  AOI22_X1 U15684 ( .A1(n13771), .A2(n14386), .B1(n14387), .B2(n13774), .ZN(
        n13777) );
  INV_X1 U15685 ( .A(n13775), .ZN(n13776) );
  MUX2_X1 U15686 ( .A(n13777), .B(n13776), .S(n13928), .Z(n13779) );
  OAI211_X1 U15687 ( .C1(n7560), .C2(n14391), .A(n13779), .B(n13778), .ZN(
        P1_U3262) );
  OR2_X2 U15688 ( .A1(n13808), .A2(n14049), .ZN(n13810) );
  INV_X1 U15689 ( .A(P1_B_REG_SCAN_IN), .ZN(n13780) );
  NOR2_X1 U15690 ( .A1(n14163), .A2(n13780), .ZN(n13781) );
  NOR2_X1 U15691 ( .A1(n14013), .A2(n13781), .ZN(n13803) );
  NAND2_X1 U15692 ( .A1(n13782), .A2(n13803), .ZN(n14042) );
  NOR2_X1 U15693 ( .A1(n14042), .A2(n6479), .ZN(n13789) );
  NOR2_X1 U15694 ( .A1(n14041), .A2(n14422), .ZN(n13783) );
  AOI211_X1 U15695 ( .C1(n6479), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13789), .B(
        n13783), .ZN(n13784) );
  OAI21_X1 U15696 ( .B1(n14022), .B2(n14040), .A(n13784), .ZN(P1_U3263) );
  INV_X1 U15697 ( .A(n13791), .ZN(n14044) );
  INV_X1 U15698 ( .A(n13810), .ZN(n13787) );
  INV_X1 U15699 ( .A(n13785), .ZN(n13786) );
  OAI211_X1 U15700 ( .C1(n14044), .C2(n13787), .A(n13786), .B(n14429), .ZN(
        n14043) );
  NOR2_X1 U15701 ( .A1(n14419), .A2(n13788), .ZN(n13790) );
  AOI211_X1 U15702 ( .C1(n13791), .C2(n14033), .A(n13790), .B(n13789), .ZN(
        n13792) );
  OAI21_X1 U15703 ( .B1(n14043), .B2(n14022), .A(n13792), .ZN(P1_U3264) );
  XNOR2_X1 U15704 ( .A(n13796), .B(n13801), .ZN(n13797) );
  NAND2_X1 U15705 ( .A1(n13797), .A2(n14411), .ZN(n14053) );
  NAND2_X1 U15706 ( .A1(n13798), .A2(n14416), .ZN(n14047) );
  AND2_X1 U15707 ( .A1(n14053), .A2(n14047), .ZN(n13815) );
  NAND2_X1 U15708 ( .A1(n14058), .A2(n13798), .ZN(n13799) );
  NAND2_X1 U15709 ( .A1(n13800), .A2(n13799), .ZN(n13802) );
  XNOR2_X1 U15710 ( .A(n13802), .B(n13801), .ZN(n14045) );
  NAND2_X1 U15711 ( .A1(n14045), .A2(n14433), .ZN(n13814) );
  NAND2_X1 U15712 ( .A1(n13804), .A2(n13803), .ZN(n14046) );
  AOI22_X1 U15713 ( .A1(n6479), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n13805), 
        .B2(n14400), .ZN(n13806) );
  OAI21_X1 U15714 ( .B1(n14046), .B2(n13807), .A(n13806), .ZN(n13812) );
  NAND2_X1 U15715 ( .A1(n13808), .A2(n14049), .ZN(n13809) );
  NAND3_X1 U15716 ( .A1(n13810), .A2(n14429), .A3(n13809), .ZN(n14051) );
  NOR2_X1 U15717 ( .A1(n14051), .A2(n14022), .ZN(n13811) );
  AOI211_X1 U15718 ( .C1(n14033), .C2(n14049), .A(n13812), .B(n13811), .ZN(
        n13813) );
  OAI211_X1 U15719 ( .C1(n6479), .C2(n13815), .A(n13814), .B(n13813), .ZN(
        P1_U3356) );
  NAND2_X1 U15720 ( .A1(n13816), .A2(n13822), .ZN(n13817) );
  INV_X1 U15721 ( .A(n13819), .ZN(n13823) );
  NAND2_X1 U15722 ( .A1(n14067), .A2(n14419), .ZN(n13830) );
  AOI211_X1 U15723 ( .C1(n14063), .C2(n13840), .A(n14076), .B(n6527), .ZN(
        n14062) );
  AOI22_X1 U15724 ( .A1(n6479), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13825), 
        .B2(n14400), .ZN(n13826) );
  OAI21_X1 U15725 ( .B1(n13827), .B2(n14422), .A(n13826), .ZN(n13828) );
  AOI21_X1 U15726 ( .B1(n14062), .B2(n14432), .A(n13828), .ZN(n13829) );
  OAI211_X1 U15727 ( .C1(n14065), .C2(n13886), .A(n13830), .B(n13829), .ZN(
        P1_U3266) );
  NAND3_X1 U15728 ( .A1(n13849), .A2(n13832), .A3(n13831), .ZN(n13833) );
  NAND2_X1 U15729 ( .A1(n13834), .A2(n13833), .ZN(n13836) );
  AOI222_X1 U15730 ( .A1(n14411), .A2(n13836), .B1(n13835), .B2(n14413), .C1(
        n13875), .C2(n14416), .ZN(n14071) );
  XNOR2_X1 U15731 ( .A(n13837), .B(n13838), .ZN(n14068) );
  NAND2_X1 U15732 ( .A1(n14068), .A2(n14433), .ZN(n13848) );
  INV_X1 U15733 ( .A(n13857), .ZN(n13841) );
  INV_X1 U15734 ( .A(n13839), .ZN(n13844) );
  OAI211_X1 U15735 ( .C1(n13841), .C2(n13844), .A(n14429), .B(n13840), .ZN(
        n14069) );
  INV_X1 U15736 ( .A(n14069), .ZN(n13846) );
  AOI22_X1 U15737 ( .A1(n6479), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13842), 
        .B2(n14400), .ZN(n13843) );
  OAI21_X1 U15738 ( .B1(n13844), .B2(n14422), .A(n13843), .ZN(n13845) );
  AOI21_X1 U15739 ( .B1(n13846), .B2(n14432), .A(n13845), .ZN(n13847) );
  OAI211_X1 U15740 ( .C1(n6479), .C2(n14071), .A(n13848), .B(n13847), .ZN(
        P1_U3267) );
  INV_X1 U15741 ( .A(n13849), .ZN(n13850) );
  AOI21_X1 U15742 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(n14081) );
  AOI21_X1 U15743 ( .B1(n13854), .B2(n13853), .A(n6563), .ZN(n14079) );
  OR2_X1 U15744 ( .A1(n13880), .A2(n13855), .ZN(n13856) );
  NAND2_X1 U15745 ( .A1(n13857), .A2(n13856), .ZN(n14077) );
  NAND2_X1 U15746 ( .A1(n14432), .A2(n14429), .ZN(n13892) );
  NAND2_X1 U15747 ( .A1(n13858), .A2(n14416), .ZN(n13861) );
  NAND2_X1 U15748 ( .A1(n13859), .A2(n14413), .ZN(n13860) );
  NAND2_X1 U15749 ( .A1(n13861), .A2(n13860), .ZN(n14073) );
  NOR2_X1 U15750 ( .A1(n14421), .A2(n13862), .ZN(n13863) );
  OAI21_X1 U15751 ( .B1(n14073), .B2(n13863), .A(n14419), .ZN(n13865) );
  NAND2_X1 U15752 ( .A1(n6479), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U15753 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  AOI21_X1 U15754 ( .B1(n14074), .B2(n14033), .A(n13866), .ZN(n13867) );
  OAI21_X1 U15755 ( .B1(n14077), .B2(n13892), .A(n13867), .ZN(n13868) );
  AOI21_X1 U15756 ( .B1(n14079), .B2(n14433), .A(n13868), .ZN(n13869) );
  OAI21_X1 U15757 ( .B1(n14081), .B2(n13962), .A(n13869), .ZN(P1_U3268) );
  OAI21_X1 U15758 ( .B1(n13872), .B2(n13871), .A(n13870), .ZN(n13885) );
  OAI211_X1 U15759 ( .C1(n13874), .C2(n7373), .A(n13873), .B(n14411), .ZN(
        n13878) );
  AOI22_X1 U15760 ( .A1(n13876), .A2(n14416), .B1(n14413), .B2(n13875), .ZN(
        n13877) );
  NAND2_X1 U15761 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  AOI21_X1 U15762 ( .B1(n13885), .B2(n14507), .A(n13879), .ZN(n14085) );
  AOI211_X1 U15763 ( .C1(n14083), .C2(n13881), .A(n14076), .B(n13880), .ZN(
        n14082) );
  AOI22_X1 U15764 ( .A1(n6479), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13882), 
        .B2(n14400), .ZN(n13883) );
  OAI21_X1 U15765 ( .B1(n13884), .B2(n14422), .A(n13883), .ZN(n13888) );
  INV_X1 U15766 ( .A(n13885), .ZN(n14086) );
  NOR2_X1 U15767 ( .A1(n14086), .A2(n13886), .ZN(n13887) );
  AOI211_X1 U15768 ( .C1(n14082), .C2(n14432), .A(n13888), .B(n13887), .ZN(
        n13889) );
  OAI21_X1 U15769 ( .B1(n6479), .B2(n14085), .A(n13889), .ZN(P1_U3269) );
  XNOR2_X1 U15770 ( .A(n13891), .B(n13890), .ZN(n14091) );
  INV_X1 U15771 ( .A(n13892), .ZN(n14034) );
  XNOR2_X1 U15772 ( .A(n13896), .B(n13909), .ZN(n14088) );
  INV_X1 U15773 ( .A(n13893), .ZN(n13894) );
  AOI22_X1 U15774 ( .A1(n13894), .A2(n14400), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n6479), .ZN(n13895) );
  OAI21_X1 U15775 ( .B1(n13896), .B2(n14422), .A(n13895), .ZN(n13904) );
  OAI21_X1 U15776 ( .B1(n13899), .B2(n13898), .A(n13897), .ZN(n13902) );
  INV_X1 U15777 ( .A(n13900), .ZN(n13901) );
  AOI21_X1 U15778 ( .B1(n13902), .B2(n14411), .A(n13901), .ZN(n14090) );
  NOR2_X1 U15779 ( .A1(n14090), .A2(n6479), .ZN(n13903) );
  AOI211_X1 U15780 ( .C1(n14034), .C2(n14088), .A(n13904), .B(n13903), .ZN(
        n13905) );
  OAI21_X1 U15781 ( .B1(n14091), .B2(n14025), .A(n13905), .ZN(P1_U3270) );
  XOR2_X1 U15782 ( .A(n13907), .B(n13906), .Z(n14098) );
  XNOR2_X1 U15783 ( .A(n13908), .B(n13907), .ZN(n14095) );
  INV_X1 U15784 ( .A(n13962), .ZN(n14031) );
  INV_X1 U15785 ( .A(n13909), .ZN(n13910) );
  AOI211_X1 U15786 ( .C1(n14094), .C2(n13924), .A(n14076), .B(n13910), .ZN(
        n14092) );
  NAND2_X1 U15787 ( .A1(n14092), .A2(n14432), .ZN(n13914) );
  OAI22_X1 U15788 ( .A1(n13911), .A2(n14421), .B1(n13245), .B2(n14419), .ZN(
        n13912) );
  AOI21_X1 U15789 ( .B1(n14093), .B2(n14419), .A(n13912), .ZN(n13913) );
  OAI211_X1 U15790 ( .C1(n14422), .C2(n13915), .A(n13914), .B(n13913), .ZN(
        n13916) );
  AOI21_X1 U15791 ( .B1(n14095), .B2(n14031), .A(n13916), .ZN(n13917) );
  OAI21_X1 U15792 ( .B1(n14098), .B2(n14025), .A(n13917), .ZN(P1_U3271) );
  XNOR2_X1 U15793 ( .A(n13918), .B(n13919), .ZN(n14104) );
  INV_X1 U15794 ( .A(n14104), .ZN(n13932) );
  AOI22_X1 U15795 ( .A1(n13923), .A2(n14033), .B1(n6479), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n13931) );
  XNOR2_X1 U15796 ( .A(n13920), .B(n13921), .ZN(n13922) );
  AND2_X1 U15797 ( .A1(n13922), .A2(n14411), .ZN(n14103) );
  AOI21_X1 U15798 ( .B1(n13940), .B2(n13923), .A(n14076), .ZN(n13925) );
  NAND2_X1 U15799 ( .A1(n13925), .A2(n13924), .ZN(n14100) );
  NAND2_X1 U15800 ( .A1(n13926), .A2(n14400), .ZN(n13927) );
  OAI211_X1 U15801 ( .C1(n14100), .C2(n13928), .A(n14099), .B(n13927), .ZN(
        n13929) );
  OAI21_X1 U15802 ( .B1(n14103), .B2(n13929), .A(n14419), .ZN(n13930) );
  OAI211_X1 U15803 ( .C1(n13932), .C2(n14025), .A(n13931), .B(n13930), .ZN(
        P1_U3272) );
  INV_X1 U15804 ( .A(n13933), .ZN(n13935) );
  OAI21_X1 U15805 ( .B1(n13935), .B2(n13939), .A(n13934), .ZN(n14112) );
  INV_X1 U15806 ( .A(n13936), .ZN(n13937) );
  AOI21_X1 U15807 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(n14110) );
  OAI211_X1 U15808 ( .C1(n14108), .C2(n13953), .A(n14429), .B(n13940), .ZN(
        n14107) );
  INV_X1 U15809 ( .A(n13941), .ZN(n14106) );
  INV_X1 U15810 ( .A(n13942), .ZN(n13943) );
  AOI22_X1 U15811 ( .A1(n6479), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n13943), 
        .B2(n14400), .ZN(n13944) );
  OAI21_X1 U15812 ( .B1(n14106), .B2(n6479), .A(n13944), .ZN(n13945) );
  AOI21_X1 U15813 ( .B1(n13946), .B2(n14033), .A(n13945), .ZN(n13947) );
  OAI21_X1 U15814 ( .B1(n14107), .B2(n14022), .A(n13947), .ZN(n13948) );
  AOI21_X1 U15815 ( .B1(n14110), .B2(n14031), .A(n13948), .ZN(n13949) );
  OAI21_X1 U15816 ( .B1(n14112), .B2(n14025), .A(n13949), .ZN(P1_U3273) );
  XNOR2_X1 U15817 ( .A(n13951), .B(n13950), .ZN(n14119) );
  XNOR2_X1 U15818 ( .A(n13952), .B(n11112), .ZN(n14113) );
  NAND2_X1 U15819 ( .A1(n14113), .A2(n14433), .ZN(n13961) );
  AOI211_X1 U15820 ( .C1(n14116), .C2(n13969), .A(n14076), .B(n13953), .ZN(
        n14114) );
  INV_X1 U15821 ( .A(n14116), .ZN(n13958) );
  INV_X1 U15822 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n13955) );
  OAI22_X1 U15823 ( .A1(n14419), .A2(n13955), .B1(n13954), .B2(n14421), .ZN(
        n13956) );
  AOI21_X1 U15824 ( .B1(n14115), .B2(n14419), .A(n13956), .ZN(n13957) );
  OAI21_X1 U15825 ( .B1(n13958), .B2(n14422), .A(n13957), .ZN(n13959) );
  AOI21_X1 U15826 ( .B1(n14114), .B2(n14432), .A(n13959), .ZN(n13960) );
  OAI211_X1 U15827 ( .C1(n14119), .C2(n13962), .A(n13961), .B(n13960), .ZN(
        P1_U3274) );
  XOR2_X1 U15828 ( .A(n13963), .B(n13967), .Z(n13964) );
  AOI222_X1 U15829 ( .A1(n13966), .A2(n14416), .B1(n13965), .B2(n14413), .C1(
        n14411), .C2(n13964), .ZN(n14123) );
  XNOR2_X1 U15830 ( .A(n13968), .B(n13967), .ZN(n14120) );
  AOI21_X1 U15831 ( .B1(n13972), .B2(n13986), .A(n14076), .ZN(n13970) );
  NAND2_X1 U15832 ( .A1(n13970), .A2(n13969), .ZN(n14121) );
  AOI22_X1 U15833 ( .A1(n6479), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13971), 
        .B2(n14400), .ZN(n13974) );
  NAND2_X1 U15834 ( .A1(n13972), .A2(n14033), .ZN(n13973) );
  OAI211_X1 U15835 ( .C1(n14121), .C2(n14022), .A(n13974), .B(n13973), .ZN(
        n13975) );
  AOI21_X1 U15836 ( .B1(n14120), .B2(n14433), .A(n13975), .ZN(n13976) );
  OAI21_X1 U15837 ( .B1(n6479), .B2(n14123), .A(n13976), .ZN(P1_U3275) );
  XNOR2_X1 U15838 ( .A(n13978), .B(n13977), .ZN(n14129) );
  NOR2_X1 U15839 ( .A1(n13979), .A2(n14422), .ZN(n13993) );
  AOI21_X1 U15840 ( .B1(n13981), .B2(n13980), .A(n14501), .ZN(n13985) );
  OAI22_X1 U15841 ( .A1(n13982), .A2(n14013), .B1(n14014), .B2(n14015), .ZN(
        n13983) );
  AOI21_X1 U15842 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n14128) );
  INV_X1 U15843 ( .A(n14003), .ZN(n13988) );
  INV_X1 U15844 ( .A(n13986), .ZN(n13987) );
  AOI211_X1 U15845 ( .C1(n14126), .C2(n13988), .A(n14076), .B(n13987), .ZN(
        n14125) );
  AOI22_X1 U15846 ( .A1(n14125), .A2(n13990), .B1(n14400), .B2(n13989), .ZN(
        n13991) );
  AOI21_X1 U15847 ( .B1(n14128), .B2(n13991), .A(n6479), .ZN(n13992) );
  AOI211_X1 U15848 ( .C1(n6479), .C2(P1_REG2_REG_17__SCAN_IN), .A(n13993), .B(
        n13992), .ZN(n13994) );
  OAI21_X1 U15849 ( .B1(n14129), .B2(n14025), .A(n13994), .ZN(P1_U3276) );
  XNOR2_X1 U15850 ( .A(n13995), .B(n13999), .ZN(n14134) );
  INV_X1 U15851 ( .A(n13996), .ZN(n13997) );
  AOI21_X1 U15852 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14000) );
  OAI222_X1 U15853 ( .A1(n14013), .A2(n14002), .B1(n14015), .B2(n14001), .C1(
        n14501), .C2(n14000), .ZN(n14130) );
  OAI21_X1 U15854 ( .B1(n6617), .B2(n14008), .A(n14429), .ZN(n14004) );
  NOR2_X1 U15855 ( .A1(n14004), .A2(n14003), .ZN(n14131) );
  NAND2_X1 U15856 ( .A1(n14131), .A2(n14432), .ZN(n14007) );
  AOI22_X1 U15857 ( .A1(n6479), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14005), 
        .B2(n14400), .ZN(n14006) );
  OAI211_X1 U15858 ( .C1(n14008), .C2(n14422), .A(n14007), .B(n14006), .ZN(
        n14009) );
  AOI21_X1 U15859 ( .B1(n14130), .B2(n14419), .A(n14009), .ZN(n14010) );
  OAI21_X1 U15860 ( .B1(n14134), .B2(n14025), .A(n14010), .ZN(P1_U3277) );
  XOR2_X1 U15861 ( .A(n14024), .B(n14011), .Z(n14312) );
  XNOR2_X1 U15862 ( .A(n14012), .B(n7119), .ZN(n14018) );
  OAI22_X1 U15863 ( .A1(n14016), .A2(n14015), .B1(n14014), .B2(n14013), .ZN(
        n14017) );
  AOI21_X1 U15864 ( .B1(n14018), .B2(n14429), .A(n14017), .ZN(n14309) );
  AOI22_X1 U15865 ( .A1(n6479), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14019), 
        .B2(n14400), .ZN(n14021) );
  NAND2_X1 U15866 ( .A1(n14307), .A2(n14033), .ZN(n14020) );
  OAI211_X1 U15867 ( .C1(n14309), .C2(n14022), .A(n14021), .B(n14020), .ZN(
        n14027) );
  AOI21_X1 U15868 ( .B1(n14024), .B2(n14023), .A(n6622), .ZN(n14310) );
  NOR2_X1 U15869 ( .A1(n14310), .A2(n14025), .ZN(n14026) );
  AOI211_X1 U15870 ( .C1(n14031), .C2(n14312), .A(n14027), .B(n14026), .ZN(
        n14028) );
  INV_X1 U15871 ( .A(n14028), .ZN(P1_U3278) );
  INV_X1 U15872 ( .A(n14029), .ZN(n14030) );
  OAI21_X1 U15873 ( .B1(n14433), .B2(n14031), .A(n14030), .ZN(n14039) );
  AOI22_X1 U15874 ( .A1(n6479), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14400), .ZN(n14038) );
  OAI21_X1 U15875 ( .B1(n14034), .B2(n14033), .A(n14032), .ZN(n14037) );
  NAND2_X1 U15876 ( .A1(n14035), .A2(n14419), .ZN(n14036) );
  NAND4_X1 U15877 ( .A1(n14039), .A2(n14038), .A3(n14037), .A4(n14036), .ZN(
        P1_U3293) );
  MUX2_X1 U15878 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14139), .S(n14534), .Z(
        P1_U3559) );
  OAI211_X1 U15879 ( .C1(n14044), .C2(n14512), .A(n14043), .B(n14042), .ZN(
        n14140) );
  MUX2_X1 U15880 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14140), .S(n14534), .Z(
        P1_U3558) );
  NAND2_X1 U15881 ( .A1(n14045), .A2(n14515), .ZN(n14055) );
  NAND2_X1 U15882 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  AOI21_X1 U15883 ( .B1(n14049), .B2(n14499), .A(n14048), .ZN(n14050) );
  AND2_X1 U15884 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U15885 ( .A1(n14055), .A2(n14054), .ZN(n14141) );
  MUX2_X1 U15886 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14141), .S(n14534), .Z(
        P1_U3557) );
  NAND2_X1 U15887 ( .A1(n14056), .A2(n14515), .ZN(n14061) );
  AOI21_X1 U15888 ( .B1(n14499), .B2(n14058), .A(n14057), .ZN(n14059) );
  MUX2_X1 U15889 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14142), .S(n14534), .Z(
        P1_U3556) );
  AOI21_X1 U15890 ( .B1(n14499), .B2(n14063), .A(n14062), .ZN(n14064) );
  OAI21_X1 U15891 ( .B1(n14065), .B2(n14503), .A(n14064), .ZN(n14066) );
  MUX2_X1 U15892 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14143), .S(n14534), .Z(
        P1_U3555) );
  NAND2_X1 U15893 ( .A1(n14068), .A2(n14515), .ZN(n14072) );
  NAND4_X1 U15894 ( .A1(n14072), .A2(n14071), .A3(n14070), .A4(n14069), .ZN(
        n14144) );
  MUX2_X1 U15895 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14144), .S(n14534), .Z(
        P1_U3554) );
  AOI21_X1 U15896 ( .B1(n14074), .B2(n14499), .A(n14073), .ZN(n14075) );
  OAI21_X1 U15897 ( .B1(n14077), .B2(n14076), .A(n14075), .ZN(n14078) );
  AOI21_X1 U15898 ( .B1(n14079), .B2(n14515), .A(n14078), .ZN(n14080) );
  OAI21_X1 U15899 ( .B1(n14501), .B2(n14081), .A(n14080), .ZN(n14145) );
  MUX2_X1 U15900 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14145), .S(n14534), .Z(
        P1_U3553) );
  AOI21_X1 U15901 ( .B1(n14499), .B2(n14083), .A(n14082), .ZN(n14084) );
  OAI211_X1 U15902 ( .C1(n14086), .C2(n14503), .A(n14085), .B(n14084), .ZN(
        n14146) );
  MUX2_X1 U15903 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14146), .S(n14534), .Z(
        P1_U3552) );
  AOI22_X1 U15904 ( .A1(n14088), .A2(n14429), .B1(n14499), .B2(n14087), .ZN(
        n14089) );
  OAI211_X1 U15905 ( .C1(n14091), .C2(n14316), .A(n14090), .B(n14089), .ZN(
        n14147) );
  MUX2_X1 U15906 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14147), .S(n14534), .Z(
        P1_U3551) );
  AOI211_X1 U15907 ( .C1(n14499), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        n14097) );
  NAND2_X1 U15908 ( .A1(n14095), .A2(n14411), .ZN(n14096) );
  OAI211_X1 U15909 ( .C1(n14098), .C2(n14316), .A(n14097), .B(n14096), .ZN(
        n14148) );
  MUX2_X1 U15910 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14148), .S(n14534), .Z(
        P1_U3550) );
  OAI211_X1 U15911 ( .C1(n14101), .C2(n14512), .A(n14100), .B(n14099), .ZN(
        n14102) );
  AOI211_X1 U15912 ( .C1(n14104), .C2(n14515), .A(n14103), .B(n14102), .ZN(
        n14105) );
  INV_X1 U15913 ( .A(n14105), .ZN(n14149) );
  MUX2_X1 U15914 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14149), .S(n14534), .Z(
        P1_U3549) );
  OAI211_X1 U15915 ( .C1(n14108), .C2(n14512), .A(n14107), .B(n14106), .ZN(
        n14109) );
  AOI21_X1 U15916 ( .B1(n14110), .B2(n14411), .A(n14109), .ZN(n14111) );
  OAI21_X1 U15917 ( .B1(n14112), .B2(n14316), .A(n14111), .ZN(n14150) );
  MUX2_X1 U15918 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14150), .S(n14534), .Z(
        P1_U3548) );
  NAND2_X1 U15919 ( .A1(n14113), .A2(n14515), .ZN(n14118) );
  AOI211_X1 U15920 ( .C1(n14499), .C2(n14116), .A(n14115), .B(n14114), .ZN(
        n14117) );
  OAI211_X1 U15921 ( .C1(n14501), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        n14151) );
  MUX2_X1 U15922 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14151), .S(n14534), .Z(
        P1_U3547) );
  NAND2_X1 U15923 ( .A1(n14120), .A2(n14515), .ZN(n14124) );
  NAND4_X1 U15924 ( .A1(n14124), .A2(n14123), .A3(n14122), .A4(n14121), .ZN(
        n14152) );
  MUX2_X1 U15925 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14152), .S(n14534), .Z(
        P1_U3546) );
  AOI21_X1 U15926 ( .B1(n14499), .B2(n14126), .A(n14125), .ZN(n14127) );
  OAI211_X1 U15927 ( .C1(n14129), .C2(n14316), .A(n14128), .B(n14127), .ZN(
        n14153) );
  MUX2_X1 U15928 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14153), .S(n14534), .Z(
        P1_U3545) );
  AOI211_X1 U15929 ( .C1(n14499), .C2(n14132), .A(n14131), .B(n14130), .ZN(
        n14133) );
  OAI21_X1 U15930 ( .B1(n14134), .B2(n14316), .A(n14133), .ZN(n14154) );
  MUX2_X1 U15931 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14154), .S(n14534), .Z(
        P1_U3544) );
  NOR2_X1 U15932 ( .A1(n14136), .A2(n14135), .ZN(n14138) );
  MUX2_X1 U15933 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14139), .S(n14519), .Z(
        P1_U3527) );
  MUX2_X1 U15934 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14140), .S(n14519), .Z(
        P1_U3526) );
  MUX2_X1 U15935 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14141), .S(n14519), .Z(
        P1_U3525) );
  MUX2_X1 U15936 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14142), .S(n14519), .Z(
        P1_U3524) );
  MUX2_X1 U15937 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14143), .S(n14519), .Z(
        P1_U3523) );
  MUX2_X1 U15938 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14144), .S(n14519), .Z(
        P1_U3522) );
  MUX2_X1 U15939 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14145), .S(n14519), .Z(
        P1_U3521) );
  MUX2_X1 U15940 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14146), .S(n14519), .Z(
        P1_U3520) );
  MUX2_X1 U15941 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14147), .S(n14519), .Z(
        P1_U3519) );
  MUX2_X1 U15942 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14148), .S(n14519), .Z(
        P1_U3518) );
  MUX2_X1 U15943 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14149), .S(n14519), .Z(
        P1_U3517) );
  MUX2_X1 U15944 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14150), .S(n14519), .Z(
        P1_U3516) );
  MUX2_X1 U15945 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14151), .S(n14519), .Z(
        P1_U3515) );
  MUX2_X1 U15946 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14152), .S(n14519), .Z(
        P1_U3513) );
  MUX2_X1 U15947 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14153), .S(n14519), .Z(
        P1_U3510) );
  MUX2_X1 U15948 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14154), .S(n14519), .Z(
        P1_U3507) );
  NOR4_X1 U15949 ( .A1(n6746), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14155), .A4(
        P1_U3086), .ZN(n14156) );
  AOI21_X1 U15950 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14157), .A(n14156), 
        .ZN(n14158) );
  OAI21_X1 U15951 ( .B1(n14159), .B2(n14165), .A(n14158), .ZN(P1_U3324) );
  OAI222_X1 U15952 ( .A1(n14165), .A2(n14161), .B1(n8564), .B2(P1_U3086), .C1(
        n14160), .C2(n14166), .ZN(P1_U3326) );
  OAI222_X1 U15953 ( .A1(n14165), .A2(n14164), .B1(n14163), .B2(P1_U3086), 
        .C1(n14162), .C2(n14166), .ZN(P1_U3328) );
  OAI222_X1 U15954 ( .A1(n14165), .A2(n14169), .B1(n14168), .B2(P1_U3086), 
        .C1(n7241), .C2(n14166), .ZN(P1_U3329) );
  OAI222_X1 U15955 ( .A1(n14166), .A2(n14172), .B1(n14165), .B2(n14171), .C1(
        P1_U3086), .C2(n14170), .ZN(P1_U3330) );
  MUX2_X1 U15956 ( .A(n14173), .B(n8661), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U15957 ( .A(n14174), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15958 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14666) );
  XNOR2_X1 U15959 ( .A(n14666), .B(n14175), .ZN(SUB_1596_U62) );
  AOI21_X1 U15960 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14176) );
  OAI21_X1 U15961 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14176), 
        .ZN(U28) );
  AOI21_X1 U15962 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14177) );
  OAI21_X1 U15963 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14177), 
        .ZN(U29) );
  AOI21_X1 U15964 ( .B1(n14180), .B2(n14179), .A(n14178), .ZN(n14181) );
  XOR2_X1 U15965 ( .A(n14181), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  INV_X1 U15966 ( .A(n14182), .ZN(n14183) );
  INV_X1 U15967 ( .A(n14186), .ZN(n14204) );
  AOI22_X1 U15968 ( .A1(n14183), .A2(n14205), .B1(SI_9_), .B2(n14204), .ZN(
        n14184) );
  OAI21_X1 U15969 ( .B1(P3_U3151), .B2(n14185), .A(n14184), .ZN(P3_U3286) );
  INV_X1 U15970 ( .A(SI_13_), .ZN(n14187) );
  OAI22_X1 U15971 ( .A1(n14188), .A2(n12423), .B1(n14187), .B2(n14186), .ZN(
        n14189) );
  INV_X1 U15972 ( .A(n14189), .ZN(n14190) );
  OAI21_X1 U15973 ( .B1(P3_U3151), .B2(n14191), .A(n14190), .ZN(P3_U3282) );
  XOR2_X1 U15974 ( .A(n14193), .B(n14192), .Z(SUB_1596_U57) );
  AOI22_X1 U15975 ( .A1(n14194), .A2(n14205), .B1(SI_14_), .B2(n14204), .ZN(
        n14195) );
  OAI21_X1 U15976 ( .B1(n6473), .B2(n14196), .A(n14195), .ZN(P3_U3281) );
  AOI22_X1 U15977 ( .A1(n14197), .A2(n14205), .B1(SI_15_), .B2(n14204), .ZN(
        n14198) );
  OAI21_X1 U15978 ( .B1(P3_U3151), .B2(n14199), .A(n14198), .ZN(P3_U3280) );
  AOI22_X1 U15979 ( .A1(n14200), .A2(n14205), .B1(SI_16_), .B2(n14204), .ZN(
        n14201) );
  OAI21_X1 U15980 ( .B1(n6473), .B2(n14202), .A(n14201), .ZN(P3_U3279) );
  XNOR2_X1 U15981 ( .A(n14203), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  AOI22_X1 U15982 ( .A1(n14206), .A2(n14205), .B1(SI_18_), .B2(n14204), .ZN(
        n14207) );
  OAI21_X1 U15983 ( .B1(n6473), .B2(n14208), .A(n14207), .ZN(P3_U3277) );
  XOR2_X1 U15984 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14209), .Z(SUB_1596_U54) );
  AOI21_X1 U15985 ( .B1(n14212), .B2(n14211), .A(n14210), .ZN(n14213) );
  XOR2_X1 U15986 ( .A(n14213), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  OAI211_X1 U15987 ( .C1(n14216), .C2(n14512), .A(n14215), .B(n14214), .ZN(
        n14217) );
  AOI21_X1 U15988 ( .B1(n14218), .B2(n14515), .A(n14217), .ZN(n14221) );
  INV_X1 U15989 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14219) );
  AOI22_X1 U15990 ( .A1(n14519), .A2(n14221), .B1(n14219), .B2(n14517), .ZN(
        P1_U3495) );
  AOI22_X1 U15991 ( .A1(n14534), .A2(n14221), .B1(n14220), .B2(n14532), .ZN(
        P1_U3540) );
  XOR2_X1 U15992 ( .A(n14222), .B(n14223), .Z(SUB_1596_U63) );
  AOI21_X1 U15993 ( .B1(n14247), .B2(n14228), .A(n14226), .ZN(n14233) );
  NOR2_X1 U15994 ( .A1(n14228), .A2(n14227), .ZN(n14229) );
  AOI21_X1 U15995 ( .B1(n14245), .B2(n14231), .A(n14229), .ZN(n14230) );
  NAND2_X1 U15996 ( .A1(n14233), .A2(n14230), .ZN(P3_U3202) );
  AOI22_X1 U15997 ( .A1(n14248), .A2(n14231), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14908), .ZN(n14232) );
  NAND2_X1 U15998 ( .A1(n14233), .A2(n14232), .ZN(P3_U3203) );
  XNOR2_X1 U15999 ( .A(n14234), .B(n10926), .ZN(n14236) );
  AOI222_X1 U16000 ( .A1(n14237), .A2(n14890), .B1(n14896), .B2(n14236), .C1(
        n14235), .C2(n14891), .ZN(n14253) );
  INV_X1 U16001 ( .A(n14238), .ZN(n14239) );
  AOI22_X1 U16002 ( .A1(n14908), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n14884), 
        .B2(n14239), .ZN(n14244) );
  OAI21_X1 U16003 ( .B1(n14241), .B2(n10926), .A(n14240), .ZN(n14256) );
  NOR2_X1 U16004 ( .A1(n14242), .A2(n14886), .ZN(n14255) );
  AOI22_X1 U16005 ( .A1(n14256), .A2(n14828), .B1(n14255), .B2(n14861), .ZN(
        n14243) );
  OAI211_X1 U16006 ( .C1(n14908), .C2(n14253), .A(n14244), .B(n14243), .ZN(
        P3_U3222) );
  AOI21_X1 U16007 ( .B1(n14245), .B2(n14916), .A(n14247), .ZN(n14258) );
  INV_X1 U16008 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U16009 ( .A1(n14968), .A2(n14258), .B1(n14246), .B2(n14965), .ZN(
        P3_U3490) );
  AOI21_X1 U16010 ( .B1(n14248), .B2(n14916), .A(n14247), .ZN(n14259) );
  INV_X1 U16011 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U16012 ( .A1(n14968), .A2(n14259), .B1(n14249), .B2(n14965), .ZN(
        P3_U3489) );
  AOI211_X1 U16013 ( .C1(n14252), .C2(n14946), .A(n14251), .B(n14250), .ZN(
        n14261) );
  AOI22_X1 U16014 ( .A1(n14968), .A2(n14261), .B1(n10220), .B2(n14965), .ZN(
        P3_U3471) );
  INV_X1 U16015 ( .A(n14253), .ZN(n14254) );
  AOI211_X1 U16016 ( .C1(n14946), .C2(n14256), .A(n14255), .B(n14254), .ZN(
        n14262) );
  INV_X1 U16017 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14257) );
  AOI22_X1 U16018 ( .A1(n14968), .A2(n14262), .B1(n14257), .B2(n14965), .ZN(
        P3_U3470) );
  AOI22_X1 U16019 ( .A1(n14949), .A2(n11457), .B1(n14258), .B2(n14948), .ZN(
        P3_U3458) );
  AOI22_X1 U16020 ( .A1(n14949), .A2(n14260), .B1(n14259), .B2(n14948), .ZN(
        P3_U3457) );
  AOI22_X1 U16021 ( .A1(n14949), .A2(n10927), .B1(n14261), .B2(n14948), .ZN(
        P3_U3426) );
  AOI22_X1 U16022 ( .A1(n14949), .A2(n10826), .B1(n14262), .B2(n14948), .ZN(
        P3_U3423) );
  OAI21_X1 U16023 ( .B1(n14264), .B2(n14756), .A(n14263), .ZN(n14266) );
  AOI211_X1 U16024 ( .C1(n14267), .C2(n14274), .A(n14266), .B(n14265), .ZN(
        n14283) );
  INV_X1 U16025 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U16026 ( .A1(n14779), .A2(n14283), .B1(n14268), .B2(n14777), .ZN(
        P2_U3513) );
  OAI21_X1 U16027 ( .B1(n14270), .B2(n14756), .A(n14269), .ZN(n14272) );
  AOI211_X1 U16028 ( .C1(n14274), .C2(n14273), .A(n14272), .B(n14271), .ZN(
        n14285) );
  AOI22_X1 U16029 ( .A1(n14779), .A2(n14285), .B1(n10439), .B2(n14777), .ZN(
        P2_U3512) );
  INV_X1 U16030 ( .A(n14740), .ZN(n14761) );
  OAI21_X1 U16031 ( .B1(n14276), .B2(n14756), .A(n14275), .ZN(n14277) );
  AOI21_X1 U16032 ( .B1(n14278), .B2(n14761), .A(n14277), .ZN(n14279) );
  AOI22_X1 U16033 ( .A1(n14779), .A2(n14287), .B1(n14281), .B2(n14777), .ZN(
        P2_U3511) );
  INV_X1 U16034 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U16035 ( .A1(n14764), .A2(n14283), .B1(n14282), .B2(n14762), .ZN(
        P2_U3472) );
  INV_X1 U16036 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U16037 ( .A1(n14764), .A2(n14285), .B1(n14284), .B2(n14762), .ZN(
        P2_U3469) );
  INV_X1 U16038 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U16039 ( .A1(n14764), .A2(n14287), .B1(n14286), .B2(n14762), .ZN(
        P2_U3466) );
  OAI21_X1 U16040 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14292) );
  AOI222_X1 U16041 ( .A1(n14293), .A2(n14373), .B1(n14292), .B2(n14366), .C1(
        n14291), .C2(n14300), .ZN(n14295) );
  OAI211_X1 U16042 ( .C1(n14376), .C2(n14296), .A(n14295), .B(n14294), .ZN(
        P1_U3215) );
  OAI21_X1 U16043 ( .B1(n14299), .B2(n14298), .A(n14297), .ZN(n14302) );
  AOI222_X1 U16044 ( .A1(n14303), .A2(n14373), .B1(n14302), .B2(n14366), .C1(
        n14301), .C2(n14300), .ZN(n14305) );
  OAI211_X1 U16045 ( .C1(n14376), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        P1_U3236) );
  NAND2_X1 U16046 ( .A1(n14307), .A2(n14499), .ZN(n14308) );
  OAI211_X1 U16047 ( .C1(n14310), .C2(n14316), .A(n14309), .B(n14308), .ZN(
        n14311) );
  AOI21_X1 U16048 ( .B1(n14411), .B2(n14312), .A(n14311), .ZN(n14335) );
  AOI22_X1 U16049 ( .A1(n14534), .A2(n14335), .B1(n14381), .B2(n14532), .ZN(
        P1_U3543) );
  OAI211_X1 U16050 ( .C1(n14315), .C2(n14512), .A(n14314), .B(n14313), .ZN(
        n14320) );
  NOR3_X1 U16051 ( .A1(n14318), .A2(n14317), .A3(n14316), .ZN(n14319) );
  AOI211_X1 U16052 ( .C1(n14321), .C2(n14411), .A(n14320), .B(n14319), .ZN(
        n14337) );
  AOI22_X1 U16053 ( .A1(n14534), .A2(n14337), .B1(n9942), .B2(n14532), .ZN(
        P1_U3542) );
  NOR2_X1 U16054 ( .A1(n14322), .A2(n14501), .ZN(n14327) );
  OAI211_X1 U16055 ( .C1(n14325), .C2(n14512), .A(n14324), .B(n14323), .ZN(
        n14326) );
  AOI211_X1 U16056 ( .C1(n14328), .C2(n14515), .A(n14327), .B(n14326), .ZN(
        n14339) );
  AOI22_X1 U16057 ( .A1(n14534), .A2(n14339), .B1(n9867), .B2(n14532), .ZN(
        P1_U3541) );
  OAI211_X1 U16058 ( .C1(n14331), .C2(n14512), .A(n14330), .B(n14329), .ZN(
        n14332) );
  AOI21_X1 U16059 ( .B1(n14333), .B2(n14515), .A(n14332), .ZN(n14341) );
  AOI22_X1 U16060 ( .A1(n14534), .A2(n14341), .B1(n9420), .B2(n14532), .ZN(
        P1_U3539) );
  INV_X1 U16061 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U16062 ( .A1(n14519), .A2(n14335), .B1(n14334), .B2(n14517), .ZN(
        P1_U3504) );
  INV_X1 U16063 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U16064 ( .A1(n14519), .A2(n14337), .B1(n14336), .B2(n14517), .ZN(
        P1_U3501) );
  INV_X1 U16065 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16066 ( .A1(n14519), .A2(n14339), .B1(n14338), .B2(n14517), .ZN(
        P1_U3498) );
  INV_X1 U16067 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U16068 ( .A1(n14519), .A2(n14341), .B1(n14340), .B2(n14517), .ZN(
        P1_U3492) );
  NOR2_X1 U16069 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  XOR2_X1 U16070 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14344), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16071 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n14348) );
  XOR2_X1 U16072 ( .A(n14348), .B(n14590), .Z(SUB_1596_U68) );
  AOI21_X1 U16073 ( .B1(n14350), .B2(n14349), .A(n6625), .ZN(n14351) );
  XOR2_X1 U16074 ( .A(n14351), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16075 ( .B1(n14354), .B2(n14353), .A(n14352), .ZN(n14355) );
  XOR2_X1 U16076 ( .A(n14355), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16077 ( .B1(n14358), .B2(n14357), .A(n14356), .ZN(n14359) );
  XOR2_X1 U16078 ( .A(n14359), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  INV_X1 U16079 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14647) );
  NOR2_X1 U16080 ( .A1(n14361), .A2(n14360), .ZN(n14362) );
  XNOR2_X1 U16081 ( .A(n14647), .B(n14362), .ZN(SUB_1596_U64) );
  NAND2_X1 U16082 ( .A1(n14363), .A2(n14499), .ZN(n14454) );
  INV_X1 U16083 ( .A(n14454), .ZN(n14365) );
  AOI22_X1 U16084 ( .A1(n14365), .A2(n14364), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14375) );
  OAI211_X1 U16085 ( .C1(n14369), .C2(n14368), .A(n14367), .B(n14366), .ZN(
        n14370) );
  INV_X1 U16086 ( .A(n14370), .ZN(n14371) );
  AOI21_X1 U16087 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n14374) );
  OAI211_X1 U16088 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14376), .A(n14375), .B(
        n14374), .ZN(P1_U3218) );
  AOI21_X1 U16089 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14378), .A(n14377), 
        .ZN(n14379) );
  INV_X1 U16090 ( .A(n14379), .ZN(n14388) );
  OAI21_X1 U16091 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14385) );
  AOI222_X1 U16092 ( .A1(n14388), .A2(n14387), .B1(n14386), .B2(n14385), .C1(
        n14384), .C2(n14383), .ZN(n14390) );
  OAI211_X1 U16093 ( .C1(n14392), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        P1_U3258) );
  XNOR2_X1 U16094 ( .A(n14393), .B(n14394), .ZN(n14479) );
  XNOR2_X1 U16095 ( .A(n14395), .B(n14396), .ZN(n14397) );
  NOR2_X1 U16096 ( .A1(n14397), .A2(n14501), .ZN(n14399) );
  AOI211_X1 U16097 ( .C1(n14479), .C2(n14507), .A(n14399), .B(n14398), .ZN(
        n14476) );
  AOI22_X1 U16098 ( .A1(n6479), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n14401), .B2(
        n14400), .ZN(n14402) );
  OAI21_X1 U16099 ( .B1(n14422), .B2(n14475), .A(n14402), .ZN(n14403) );
  INV_X1 U16100 ( .A(n14403), .ZN(n14409) );
  OAI211_X1 U16101 ( .C1(n14475), .C2(n14405), .A(n14404), .B(n14429), .ZN(
        n14474) );
  INV_X1 U16102 ( .A(n14474), .ZN(n14406) );
  AOI22_X1 U16103 ( .A1(n14479), .A2(n14407), .B1(n14432), .B2(n14406), .ZN(
        n14408) );
  OAI211_X1 U16104 ( .C1(n6479), .C2(n14476), .A(n14409), .B(n14408), .ZN(
        P1_U3287) );
  XNOR2_X1 U16105 ( .A(n14410), .B(n14425), .ZN(n14412) );
  NAND2_X1 U16106 ( .A1(n14412), .A2(n14411), .ZN(n14418) );
  AOI22_X1 U16107 ( .A1(n14416), .A2(n14415), .B1(n14414), .B2(n14413), .ZN(
        n14417) );
  NAND2_X1 U16108 ( .A1(n14418), .A2(n14417), .ZN(n14463) );
  MUX2_X1 U16109 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14463), .S(n14419), .Z(
        n14424) );
  OAI22_X1 U16110 ( .A1(n14422), .A2(n14461), .B1(n14421), .B2(n14420), .ZN(
        n14423) );
  NOR2_X1 U16111 ( .A1(n14424), .A2(n14423), .ZN(n14435) );
  XNOR2_X1 U16112 ( .A(n14426), .B(n14425), .ZN(n14464) );
  INV_X1 U16113 ( .A(n14427), .ZN(n14430) );
  OAI211_X1 U16114 ( .C1(n14430), .C2(n14461), .A(n14429), .B(n14428), .ZN(
        n14460) );
  INV_X1 U16115 ( .A(n14460), .ZN(n14431) );
  AOI22_X1 U16116 ( .A1(n14464), .A2(n14433), .B1(n14432), .B2(n14431), .ZN(
        n14434) );
  NAND2_X1 U16117 ( .A1(n14435), .A2(n14434), .ZN(P1_U3289) );
  AND2_X1 U16118 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14439), .ZN(P1_U3294) );
  AND2_X1 U16119 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14439), .ZN(P1_U3295) );
  AND2_X1 U16120 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14439), .ZN(P1_U3296) );
  AND2_X1 U16121 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14439), .ZN(P1_U3297) );
  AND2_X1 U16122 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14439), .ZN(P1_U3298) );
  AND2_X1 U16123 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14439), .ZN(P1_U3299) );
  AND2_X1 U16124 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14439), .ZN(P1_U3300) );
  AND2_X1 U16125 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14439), .ZN(P1_U3301) );
  AND2_X1 U16126 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14439), .ZN(P1_U3302) );
  INV_X1 U16127 ( .A(n14439), .ZN(n14438) );
  NOR2_X1 U16128 ( .A1(n14438), .A2(n14436), .ZN(P1_U3303) );
  AND2_X1 U16129 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14439), .ZN(P1_U3304) );
  AND2_X1 U16130 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14439), .ZN(P1_U3305) );
  AND2_X1 U16131 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14439), .ZN(P1_U3306) );
  AND2_X1 U16132 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14439), .ZN(P1_U3307) );
  AND2_X1 U16133 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14439), .ZN(P1_U3308) );
  AND2_X1 U16134 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14439), .ZN(P1_U3309) );
  AND2_X1 U16135 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14439), .ZN(P1_U3310) );
  AND2_X1 U16136 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14439), .ZN(P1_U3311) );
  NOR2_X1 U16137 ( .A1(n14438), .A2(n14437), .ZN(P1_U3312) );
  AND2_X1 U16138 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14439), .ZN(P1_U3313) );
  AND2_X1 U16139 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14439), .ZN(P1_U3314) );
  AND2_X1 U16140 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14439), .ZN(P1_U3315) );
  AND2_X1 U16141 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14439), .ZN(P1_U3316) );
  AND2_X1 U16142 ( .A1(n14439), .A2(P1_D_REG_8__SCAN_IN), .ZN(P1_U3317) );
  AND2_X1 U16143 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14439), .ZN(P1_U3318) );
  AND2_X1 U16144 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14439), .ZN(P1_U3319) );
  AND2_X1 U16145 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14439), .ZN(P1_U3320) );
  AND2_X1 U16146 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14439), .ZN(P1_U3321) );
  AND2_X1 U16147 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14439), .ZN(P1_U3322) );
  AND2_X1 U16148 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14439), .ZN(P1_U3323) );
  INV_X1 U16149 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U16150 ( .A1(n14519), .A2(n14441), .B1(n14440), .B2(n14517), .ZN(
        P1_U3459) );
  INV_X1 U16151 ( .A(n14503), .ZN(n14480) );
  OAI21_X1 U16152 ( .B1(n9158), .B2(n14512), .A(n14442), .ZN(n14444) );
  AOI211_X1 U16153 ( .C1(n14480), .C2(n14445), .A(n14444), .B(n14443), .ZN(
        n14521) );
  INV_X1 U16154 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U16155 ( .A1(n14519), .A2(n14521), .B1(n14446), .B2(n14517), .ZN(
        P1_U3462) );
  OAI21_X1 U16156 ( .B1(n14448), .B2(n14512), .A(n14447), .ZN(n14450) );
  AOI211_X1 U16157 ( .C1(n14480), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14522) );
  INV_X1 U16158 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U16159 ( .A1(n14519), .A2(n14522), .B1(n14452), .B2(n14517), .ZN(
        P1_U3465) );
  NAND2_X1 U16160 ( .A1(n14453), .A2(n14480), .ZN(n14456) );
  NAND3_X1 U16161 ( .A1(n14456), .A2(n14455), .A3(n14454), .ZN(n14457) );
  NOR2_X1 U16162 ( .A1(n14458), .A2(n14457), .ZN(n14523) );
  INV_X1 U16163 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16164 ( .A1(n14519), .A2(n14523), .B1(n14459), .B2(n14517), .ZN(
        P1_U3468) );
  OAI21_X1 U16165 ( .B1(n14461), .B2(n14512), .A(n14460), .ZN(n14462) );
  AOI211_X1 U16166 ( .C1(n14464), .C2(n14515), .A(n14463), .B(n14462), .ZN(
        n14524) );
  INV_X1 U16167 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U16168 ( .A1(n14519), .A2(n14524), .B1(n14465), .B2(n14517), .ZN(
        P1_U3471) );
  INV_X1 U16169 ( .A(n14470), .ZN(n14472) );
  AOI211_X1 U16170 ( .C1(n14499), .C2(n14468), .A(n14467), .B(n14466), .ZN(
        n14469) );
  OAI21_X1 U16171 ( .B1(n14503), .B2(n14470), .A(n14469), .ZN(n14471) );
  AOI21_X1 U16172 ( .B1(n14507), .B2(n14472), .A(n14471), .ZN(n14526) );
  INV_X1 U16173 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U16174 ( .A1(n14519), .A2(n14526), .B1(n14473), .B2(n14517), .ZN(
        P1_U3474) );
  OAI21_X1 U16175 ( .B1(n14475), .B2(n14512), .A(n14474), .ZN(n14478) );
  INV_X1 U16176 ( .A(n14476), .ZN(n14477) );
  AOI211_X1 U16177 ( .C1(n14480), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14528) );
  INV_X1 U16178 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U16179 ( .A1(n14519), .A2(n14528), .B1(n14481), .B2(n14517), .ZN(
        P1_U3477) );
  INV_X1 U16180 ( .A(n14486), .ZN(n14488) );
  AOI211_X1 U16181 ( .C1(n14499), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14485) );
  OAI21_X1 U16182 ( .B1(n14486), .B2(n14503), .A(n14485), .ZN(n14487) );
  AOI21_X1 U16183 ( .B1(n14507), .B2(n14488), .A(n14487), .ZN(n14529) );
  AOI22_X1 U16184 ( .A1(n14519), .A2(n14529), .B1(n14489), .B2(n14517), .ZN(
        P1_U3480) );
  OAI211_X1 U16185 ( .C1(n14492), .C2(n14512), .A(n14491), .B(n14490), .ZN(
        n14493) );
  AOI21_X1 U16186 ( .B1(n14494), .B2(n14515), .A(n14493), .ZN(n14530) );
  INV_X1 U16187 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14495) );
  AOI22_X1 U16188 ( .A1(n14519), .A2(n14530), .B1(n14495), .B2(n14517), .ZN(
        P1_U3483) );
  AOI211_X1 U16189 ( .C1(n14499), .C2(n14498), .A(n14497), .B(n14496), .ZN(
        n14500) );
  OAI21_X1 U16190 ( .B1(n14502), .B2(n14501), .A(n14500), .ZN(n14506) );
  NOR2_X1 U16191 ( .A1(n14504), .A2(n14503), .ZN(n14505) );
  AOI211_X1 U16192 ( .C1(n14508), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14531) );
  INV_X1 U16193 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U16194 ( .A1(n14519), .A2(n14531), .B1(n14509), .B2(n14517), .ZN(
        P1_U3486) );
  OAI211_X1 U16195 ( .C1(n14513), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14514) );
  AOI21_X1 U16196 ( .B1(n14516), .B2(n14515), .A(n14514), .ZN(n14533) );
  INV_X1 U16197 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U16198 ( .A1(n14519), .A2(n14533), .B1(n14518), .B2(n14517), .ZN(
        P1_U3489) );
  INV_X1 U16199 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14520) );
  AOI22_X1 U16200 ( .A1(n14534), .A2(n14521), .B1(n14520), .B2(n14532), .ZN(
        P1_U3529) );
  AOI22_X1 U16201 ( .A1(n14534), .A2(n14522), .B1(n8850), .B2(n14532), .ZN(
        P1_U3530) );
  AOI22_X1 U16202 ( .A1(n14534), .A2(n14523), .B1(n8851), .B2(n14532), .ZN(
        P1_U3531) );
  AOI22_X1 U16203 ( .A1(n14534), .A2(n14524), .B1(n8870), .B2(n14532), .ZN(
        P1_U3532) );
  INV_X1 U16204 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U16205 ( .A1(n14534), .A2(n14526), .B1(n14525), .B2(n14532), .ZN(
        P1_U3533) );
  INV_X1 U16206 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14527) );
  AOI22_X1 U16207 ( .A1(n14534), .A2(n14528), .B1(n14527), .B2(n14532), .ZN(
        P1_U3534) );
  AOI22_X1 U16208 ( .A1(n14534), .A2(n14529), .B1(n8970), .B2(n14532), .ZN(
        P1_U3535) );
  AOI22_X1 U16209 ( .A1(n14534), .A2(n14530), .B1(n9195), .B2(n14532), .ZN(
        P1_U3536) );
  AOI22_X1 U16210 ( .A1(n14534), .A2(n14531), .B1(n9196), .B2(n14532), .ZN(
        P1_U3537) );
  AOI22_X1 U16211 ( .A1(n14534), .A2(n14533), .B1(n9193), .B2(n14532), .ZN(
        P1_U3538) );
  NOR2_X1 U16212 ( .A1(n14535), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI211_X1 U16213 ( .C1(n14538), .C2(n14537), .A(n14657), .B(n14536), .ZN(
        n14544) );
  OAI21_X1 U16214 ( .B1(n14541), .B2(n14540), .A(n14539), .ZN(n14542) );
  OR2_X1 U16215 ( .A1(n14633), .A2(n14542), .ZN(n14543) );
  OAI211_X1 U16216 ( .C1(n14661), .C2(n14545), .A(n14544), .B(n14543), .ZN(
        n14546) );
  INV_X1 U16217 ( .A(n14546), .ZN(n14548) );
  NAND2_X1 U16218 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14547) );
  OAI211_X1 U16219 ( .C1(n14665), .C2(n14980), .A(n14548), .B(n14547), .ZN(
        P2_U3217) );
  OAI211_X1 U16220 ( .C1(n14551), .C2(n14550), .A(n14657), .B(n14549), .ZN(
        n14552) );
  INV_X1 U16221 ( .A(n14552), .ZN(n14559) );
  OAI21_X1 U16222 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n14557) );
  OAI22_X1 U16223 ( .A1(n14633), .A2(n14557), .B1(n14556), .B2(n14661), .ZN(
        n14558) );
  NOR2_X1 U16224 ( .A1(n14559), .A2(n14558), .ZN(n14561) );
  OAI211_X1 U16225 ( .C1(n14665), .C2(n14562), .A(n14561), .B(n14560), .ZN(
        P2_U3218) );
  INV_X1 U16226 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n14972) );
  OAI211_X1 U16227 ( .C1(n14565), .C2(n14564), .A(n14657), .B(n14563), .ZN(
        n14566) );
  INV_X1 U16228 ( .A(n14566), .ZN(n14573) );
  OAI21_X1 U16229 ( .B1(n14569), .B2(n14568), .A(n14567), .ZN(n14571) );
  OAI22_X1 U16230 ( .A1(n14633), .A2(n14571), .B1(n14570), .B2(n14661), .ZN(
        n14572) );
  NOR2_X1 U16231 ( .A1(n14573), .A2(n14572), .ZN(n14575) );
  NAND2_X1 U16232 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14574) );
  OAI211_X1 U16233 ( .C1(n14665), .C2(n14972), .A(n14575), .B(n14574), .ZN(
        P2_U3219) );
  OAI21_X1 U16234 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14579) );
  NAND2_X1 U16235 ( .A1(n14579), .A2(n14657), .ZN(n14585) );
  OAI21_X1 U16236 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n14583) );
  NAND2_X1 U16237 ( .A1(n14583), .A2(n14652), .ZN(n14584) );
  OAI211_X1 U16238 ( .C1(n14661), .C2(n14586), .A(n14585), .B(n14584), .ZN(
        n14587) );
  INV_X1 U16239 ( .A(n14587), .ZN(n14589) );
  OAI211_X1 U16240 ( .C1(n14590), .C2(n14665), .A(n14589), .B(n14588), .ZN(
        P2_U3226) );
  AOI21_X1 U16241 ( .B1(n14592), .B2(n14591), .A(n14637), .ZN(n14594) );
  NAND2_X1 U16242 ( .A1(n14594), .A2(n14593), .ZN(n14600) );
  AOI21_X1 U16243 ( .B1(n14596), .B2(n14595), .A(n14633), .ZN(n14598) );
  NAND2_X1 U16244 ( .A1(n14598), .A2(n14597), .ZN(n14599) );
  OAI211_X1 U16245 ( .C1(n14661), .C2(n14601), .A(n14600), .B(n14599), .ZN(
        n14602) );
  INV_X1 U16246 ( .A(n14602), .ZN(n14604) );
  NAND2_X1 U16247 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14603)
         );
  OAI211_X1 U16248 ( .C1(n14605), .C2(n14665), .A(n14604), .B(n14603), .ZN(
        P2_U3227) );
  INV_X1 U16249 ( .A(n14606), .ZN(n14616) );
  OAI21_X1 U16250 ( .B1(n14607), .B2(P2_REG2_REG_14__SCAN_IN), .A(n14657), 
        .ZN(n14608) );
  INV_X1 U16251 ( .A(n14608), .ZN(n14615) );
  OAI21_X1 U16252 ( .B1(n14610), .B2(n14609), .A(n14652), .ZN(n14613) );
  OAI22_X1 U16253 ( .A1(n14613), .A2(n14612), .B1(n14611), .B2(n14661), .ZN(
        n14614) );
  AOI21_X1 U16254 ( .B1(n14616), .B2(n14615), .A(n14614), .ZN(n14618) );
  OAI211_X1 U16255 ( .C1(n14619), .C2(n14665), .A(n14618), .B(n14617), .ZN(
        P2_U3228) );
  INV_X1 U16256 ( .A(n14661), .ZN(n14644) );
  AOI211_X1 U16257 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14637), .ZN(
        n14628) );
  INV_X1 U16258 ( .A(n14623), .ZN(n14626) );
  INV_X1 U16259 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14625) );
  AOI211_X1 U16260 ( .C1(n14626), .C2(n14625), .A(n14633), .B(n14624), .ZN(
        n14627) );
  AOI211_X1 U16261 ( .C1(n14644), .C2(n14629), .A(n14628), .B(n14627), .ZN(
        n14631) );
  NAND2_X1 U16262 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14630)
         );
  OAI211_X1 U16263 ( .C1(n14632), .C2(n14665), .A(n14631), .B(n14630), .ZN(
        P2_U3229) );
  AOI211_X1 U16264 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14642) );
  AOI211_X1 U16265 ( .C1(n14640), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14641) );
  AOI211_X1 U16266 ( .C1(n14644), .C2(n14643), .A(n14642), .B(n14641), .ZN(
        n14646) );
  OAI211_X1 U16267 ( .C1(n14647), .C2(n14665), .A(n14646), .B(n14645), .ZN(
        P2_U3230) );
  AOI21_X1 U16268 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(n14651) );
  NAND2_X1 U16269 ( .A1(n14652), .A2(n14651), .ZN(n14659) );
  OAI21_X1 U16270 ( .B1(n14655), .B2(n14654), .A(n14653), .ZN(n14656) );
  NAND2_X1 U16271 ( .A1(n14657), .A2(n14656), .ZN(n14658) );
  OAI211_X1 U16272 ( .C1(n14661), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        n14662) );
  INV_X1 U16273 ( .A(n14662), .ZN(n14664) );
  OAI211_X1 U16274 ( .C1(n14666), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        P2_U3232) );
  NAND2_X1 U16275 ( .A1(n14668), .A2(n14667), .ZN(n14672) );
  AOI22_X1 U16276 ( .A1(n14680), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14670), 
        .B2(n14669), .ZN(n14671) );
  OAI211_X1 U16277 ( .C1(n14674), .C2(n14673), .A(n14672), .B(n14671), .ZN(
        n14675) );
  AOI21_X1 U16278 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14678) );
  OAI21_X1 U16279 ( .B1(n14680), .B2(n14679), .A(n14678), .ZN(P2_U3258) );
  INV_X1 U16280 ( .A(n14685), .ZN(n14687) );
  AND2_X1 U16281 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14682), .ZN(P2_U3266) );
  AND2_X1 U16282 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14682), .ZN(P2_U3267) );
  AND2_X1 U16283 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14682), .ZN(P2_U3268) );
  AND2_X1 U16284 ( .A1(n14682), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3269) );
  AND2_X1 U16285 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14682), .ZN(P2_U3270) );
  AND2_X1 U16286 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14682), .ZN(P2_U3271) );
  AND2_X1 U16287 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14682), .ZN(P2_U3272) );
  AND2_X1 U16288 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14682), .ZN(P2_U3273) );
  AND2_X1 U16289 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14682), .ZN(P2_U3274) );
  AND2_X1 U16290 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14682), .ZN(P2_U3275) );
  AND2_X1 U16291 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14682), .ZN(P2_U3276) );
  AND2_X1 U16292 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14682), .ZN(P2_U3277) );
  AND2_X1 U16293 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14682), .ZN(P2_U3278) );
  AND2_X1 U16294 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14682), .ZN(P2_U3279) );
  AND2_X1 U16295 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14682), .ZN(P2_U3280) );
  AND2_X1 U16296 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14682), .ZN(P2_U3281) );
  AND2_X1 U16297 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14682), .ZN(P2_U3282) );
  AND2_X1 U16298 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14682), .ZN(P2_U3283) );
  AND2_X1 U16299 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14682), .ZN(P2_U3284) );
  AND2_X1 U16300 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14682), .ZN(P2_U3285) );
  AND2_X1 U16301 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14682), .ZN(P2_U3286) );
  AND2_X1 U16302 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14682), .ZN(P2_U3287) );
  AND2_X1 U16303 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14682), .ZN(P2_U3288) );
  AND2_X1 U16304 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14682), .ZN(P2_U3289) );
  AND2_X1 U16305 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14682), .ZN(P2_U3290) );
  AND2_X1 U16306 ( .A1(n14682), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3291) );
  AND2_X1 U16307 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14682), .ZN(P2_U3292) );
  AND2_X1 U16308 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14682), .ZN(P2_U3293) );
  AND2_X1 U16309 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14682), .ZN(P2_U3294) );
  AND2_X1 U16310 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14682), .ZN(P2_U3295) );
  AOI22_X1 U16311 ( .A1(n14685), .A2(n14684), .B1(n14683), .B2(n14687), .ZN(
        P2_U3416) );
  AOI21_X1 U16312 ( .B1(n14688), .B2(n14687), .A(n14686), .ZN(P2_U3417) );
  OAI211_X1 U16313 ( .C1(n14691), .C2(n14740), .A(n14690), .B(n14689), .ZN(
        n14692) );
  INV_X1 U16314 ( .A(n14692), .ZN(n14766) );
  INV_X1 U16315 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U16316 ( .A1(n14764), .A2(n14766), .B1(n14693), .B2(n14762), .ZN(
        P2_U3430) );
  AOI21_X1 U16317 ( .B1(n14738), .B2(n14695), .A(n14694), .ZN(n14696) );
  OAI211_X1 U16318 ( .C1(n14698), .C2(n14740), .A(n14697), .B(n14696), .ZN(
        n14699) );
  INV_X1 U16319 ( .A(n14699), .ZN(n14767) );
  INV_X1 U16320 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14700) );
  AOI22_X1 U16321 ( .A1(n14764), .A2(n14767), .B1(n14700), .B2(n14762), .ZN(
        P2_U3433) );
  INV_X1 U16322 ( .A(n14705), .ZN(n14707) );
  INV_X1 U16323 ( .A(n14701), .ZN(n14702) );
  AOI211_X1 U16324 ( .C1(n14738), .C2(n8267), .A(n14703), .B(n14702), .ZN(
        n14704) );
  OAI21_X1 U16325 ( .B1(n14705), .B2(n14740), .A(n14704), .ZN(n14706) );
  AOI21_X1 U16326 ( .B1(n14745), .B2(n14707), .A(n14706), .ZN(n14768) );
  INV_X1 U16327 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14708) );
  AOI22_X1 U16328 ( .A1(n14764), .A2(n14768), .B1(n14708), .B2(n14762), .ZN(
        P2_U3436) );
  OAI21_X1 U16329 ( .B1(n14710), .B2(n14756), .A(n14709), .ZN(n14711) );
  NOR2_X1 U16330 ( .A1(n14712), .A2(n14711), .ZN(n14715) );
  OR2_X1 U16331 ( .A1(n14713), .A2(n14720), .ZN(n14714) );
  AND2_X1 U16332 ( .A1(n14715), .A2(n14714), .ZN(n14769) );
  INV_X1 U16333 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16334 ( .A1(n14764), .A2(n14769), .B1(n14716), .B2(n14762), .ZN(
        P2_U3439) );
  AND2_X1 U16335 ( .A1(n14738), .A2(n14717), .ZN(n14718) );
  NOR2_X1 U16336 ( .A1(n14719), .A2(n14718), .ZN(n14723) );
  OR2_X1 U16337 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  INV_X1 U16338 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U16339 ( .A1(n14764), .A2(n14770), .B1(n14725), .B2(n14762), .ZN(
        P2_U3442) );
  INV_X1 U16340 ( .A(n14729), .ZN(n14733) );
  AOI21_X1 U16341 ( .B1(n14738), .B2(n14727), .A(n14726), .ZN(n14728) );
  OAI21_X1 U16342 ( .B1(n14729), .B2(n14740), .A(n14728), .ZN(n14732) );
  INV_X1 U16343 ( .A(n14730), .ZN(n14731) );
  AOI211_X1 U16344 ( .C1(n14745), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        n14772) );
  INV_X1 U16345 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16346 ( .A1(n14764), .A2(n14772), .B1(n14734), .B2(n14762), .ZN(
        P2_U3445) );
  INV_X1 U16347 ( .A(n14735), .ZN(n14743) );
  AOI21_X1 U16348 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14739) );
  OAI21_X1 U16349 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14742) );
  AOI211_X1 U16350 ( .C1(n14745), .C2(n14744), .A(n14743), .B(n14742), .ZN(
        n14774) );
  INV_X1 U16351 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U16352 ( .A1(n14764), .A2(n14774), .B1(n14746), .B2(n14762), .ZN(
        P2_U3448) );
  INV_X1 U16353 ( .A(n14747), .ZN(n14752) );
  OAI21_X1 U16354 ( .B1(n14749), .B2(n14756), .A(n14748), .ZN(n14751) );
  AOI211_X1 U16355 ( .C1(n14761), .C2(n14752), .A(n14751), .B(n14750), .ZN(
        n14776) );
  INV_X1 U16356 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U16357 ( .A1(n14764), .A2(n14776), .B1(n14753), .B2(n14762), .ZN(
        P2_U3454) );
  INV_X1 U16358 ( .A(n14754), .ZN(n14760) );
  OAI21_X1 U16359 ( .B1(n14757), .B2(n14756), .A(n14755), .ZN(n14759) );
  AOI211_X1 U16360 ( .C1(n14761), .C2(n14760), .A(n14759), .B(n14758), .ZN(
        n14778) );
  INV_X1 U16361 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U16362 ( .A1(n14764), .A2(n14778), .B1(n14763), .B2(n14762), .ZN(
        P2_U3460) );
  AOI22_X1 U16363 ( .A1(n14779), .A2(n14766), .B1(n14765), .B2(n14777), .ZN(
        P2_U3499) );
  AOI22_X1 U16364 ( .A1(n14779), .A2(n14767), .B1(n8915), .B2(n14777), .ZN(
        P2_U3500) );
  AOI22_X1 U16365 ( .A1(n14779), .A2(n14768), .B1(n8914), .B2(n14777), .ZN(
        P2_U3501) );
  AOI22_X1 U16366 ( .A1(n14779), .A2(n14769), .B1(n8918), .B2(n14777), .ZN(
        P2_U3502) );
  AOI22_X1 U16367 ( .A1(n14779), .A2(n14770), .B1(n8920), .B2(n14777), .ZN(
        P2_U3503) );
  AOI22_X1 U16368 ( .A1(n14779), .A2(n14772), .B1(n14771), .B2(n14777), .ZN(
        P2_U3504) );
  AOI22_X1 U16369 ( .A1(n14779), .A2(n14774), .B1(n14773), .B2(n14777), .ZN(
        P2_U3505) );
  AOI22_X1 U16370 ( .A1(n14779), .A2(n14776), .B1(n14775), .B2(n14777), .ZN(
        P2_U3507) );
  AOI22_X1 U16371 ( .A1(n14779), .A2(n14778), .B1(n8988), .B2(n14777), .ZN(
        P2_U3509) );
  NOR2_X1 U16372 ( .A1(P3_U3897), .A2(n14780), .ZN(P3_U3150) );
  OAI21_X1 U16373 ( .B1(n14783), .B2(n14782), .A(n14781), .ZN(n14800) );
  OAI21_X1 U16374 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(n14787) );
  AND2_X1 U16375 ( .A1(n14788), .A2(n14787), .ZN(n14799) );
  AND3_X1 U16376 ( .A1(n14791), .A2(n14790), .A3(n14789), .ZN(n14793) );
  OAI21_X1 U16377 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(n14795) );
  OAI21_X1 U16378 ( .B1(n14797), .B2(n14796), .A(n14795), .ZN(n14798) );
  AOI211_X1 U16379 ( .C1(n14801), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14803) );
  OAI211_X1 U16380 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        P3_U3188) );
  XNOR2_X1 U16381 ( .A(n14806), .B(n10920), .ZN(n14808) );
  AOI222_X1 U16382 ( .A1(n14809), .A2(n14890), .B1(n14896), .B2(n14808), .C1(
        n14807), .C2(n14891), .ZN(n14943) );
  AOI22_X1 U16383 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n14908), .B1(n14884), 
        .B2(n14810), .ZN(n14817) );
  INV_X1 U16384 ( .A(n14811), .ZN(n14812) );
  AOI21_X1 U16385 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n14947) );
  NOR2_X1 U16386 ( .A1(n14815), .A2(n14886), .ZN(n14945) );
  AOI22_X1 U16387 ( .A1(n14947), .A2(n14828), .B1(n14945), .B2(n14861), .ZN(
        n14816) );
  OAI211_X1 U16388 ( .C1(n14908), .C2(n14943), .A(n14817), .B(n14816), .ZN(
        P3_U3223) );
  AOI21_X1 U16389 ( .B1(n6621), .B2(n14826), .A(n14873), .ZN(n14822) );
  OAI22_X1 U16390 ( .A1(n14819), .A2(n14869), .B1(n14818), .B2(n14867), .ZN(
        n14820) );
  AOI21_X1 U16391 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14939) );
  INV_X1 U16392 ( .A(n14823), .ZN(n14824) );
  AOI22_X1 U16393 ( .A1(n14908), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n14884), 
        .B2(n14824), .ZN(n14830) );
  XNOR2_X1 U16394 ( .A(n14825), .B(n14826), .ZN(n14942) );
  NOR2_X1 U16395 ( .A1(n14827), .A2(n14886), .ZN(n14941) );
  AOI22_X1 U16396 ( .A1(n14942), .A2(n14828), .B1(n14941), .B2(n14861), .ZN(
        n14829) );
  OAI211_X1 U16397 ( .C1(n14908), .C2(n14939), .A(n14830), .B(n14829), .ZN(
        P3_U3224) );
  XNOR2_X1 U16398 ( .A(n14836), .B(n14831), .ZN(n14840) );
  INV_X1 U16399 ( .A(n14840), .ZN(n14930) );
  OAI22_X1 U16400 ( .A1(n14833), .A2(n14869), .B1(n14832), .B2(n14867), .ZN(
        n14834) );
  INV_X1 U16401 ( .A(n14834), .ZN(n14839) );
  OAI211_X1 U16402 ( .C1(n14837), .C2(n14836), .A(n14835), .B(n14896), .ZN(
        n14838) );
  OAI211_X1 U16403 ( .C1(n14840), .C2(n14900), .A(n14839), .B(n14838), .ZN(
        n14928) );
  AOI21_X1 U16404 ( .B1(n14881), .B2(n14930), .A(n14928), .ZN(n14846) );
  NOR2_X1 U16405 ( .A1(n14841), .A2(n14886), .ZN(n14929) );
  INV_X1 U16406 ( .A(n14842), .ZN(n14843) );
  AOI22_X1 U16407 ( .A1(n14861), .A2(n14929), .B1(n14884), .B2(n14843), .ZN(
        n14844) );
  OAI221_X1 U16408 ( .B1(n14908), .B2(n14846), .C1(n14228), .C2(n14845), .A(
        n14844), .ZN(P3_U3227) );
  NAND3_X1 U16409 ( .A1(n14848), .A2(n14852), .A3(n14847), .ZN(n14849) );
  NAND2_X1 U16410 ( .A1(n14850), .A2(n14849), .ZN(n14923) );
  XNOR2_X1 U16411 ( .A(n14852), .B(n14851), .ZN(n14857) );
  AOI22_X1 U16412 ( .A1(n14854), .A2(n14891), .B1(n14890), .B2(n14853), .ZN(
        n14856) );
  NAND2_X1 U16413 ( .A1(n14923), .A2(n14878), .ZN(n14855) );
  OAI211_X1 U16414 ( .C1(n14857), .C2(n14873), .A(n14856), .B(n14855), .ZN(
        n14921) );
  AOI21_X1 U16415 ( .B1(n14881), .B2(n14923), .A(n14921), .ZN(n14864) );
  NOR2_X1 U16416 ( .A1(n14858), .A2(n14886), .ZN(n14922) );
  INV_X1 U16417 ( .A(n14859), .ZN(n14860) );
  AOI22_X1 U16418 ( .A1(n14861), .A2(n14922), .B1(n14884), .B2(n14860), .ZN(
        n14862) );
  OAI221_X1 U16419 ( .B1(n14908), .B2(n14864), .C1(n14228), .C2(n14863), .A(
        n14862), .ZN(P3_U3229) );
  OAI21_X1 U16420 ( .B1(n14866), .B2(n7410), .A(n14865), .ZN(n14915) );
  OAI22_X1 U16421 ( .A1(n14870), .A2(n14869), .B1(n14868), .B2(n14867), .ZN(
        n14877) );
  NAND3_X1 U16422 ( .A1(n7410), .A2(n14871), .A3(n14893), .ZN(n14874) );
  AOI21_X1 U16423 ( .B1(n14875), .B2(n14874), .A(n14873), .ZN(n14876) );
  AOI211_X1 U16424 ( .C1(n14878), .C2(n14915), .A(n14877), .B(n14876), .ZN(
        n14879) );
  INV_X1 U16425 ( .A(n14879), .ZN(n14913) );
  NOR2_X1 U16426 ( .A1(n14880), .A2(n14886), .ZN(n14914) );
  AOI22_X1 U16427 ( .A1(n14915), .A2(n14881), .B1(n14914), .B2(n14901), .ZN(
        n14882) );
  INV_X1 U16428 ( .A(n14882), .ZN(n14883) );
  AOI211_X1 U16429 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n14884), .A(n14913), .B(
        n14883), .ZN(n14885) );
  AOI22_X1 U16430 ( .A1(n14908), .A2(n9043), .B1(n14885), .B2(n14228), .ZN(
        P3_U3231) );
  NOR2_X1 U16431 ( .A1(n14887), .A2(n14886), .ZN(n14911) );
  XNOR2_X1 U16432 ( .A(n14888), .B(n14894), .ZN(n14909) );
  AOI22_X1 U16433 ( .A1(n14892), .A2(n14891), .B1(n14890), .B2(n14889), .ZN(
        n14899) );
  OAI21_X1 U16434 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14897) );
  NAND2_X1 U16435 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  OAI211_X1 U16436 ( .C1(n14909), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        n14910) );
  AOI21_X1 U16437 ( .B1(n14911), .B2(n14901), .A(n14910), .ZN(n14907) );
  OAI22_X1 U16438 ( .A1(n14909), .A2(n14904), .B1(n14903), .B2(n14902), .ZN(
        n14905) );
  INV_X1 U16439 ( .A(n14905), .ZN(n14906) );
  OAI221_X1 U16440 ( .B1(n14908), .B2(n14907), .C1(n14228), .C2(n9385), .A(
        n14906), .ZN(P3_U3232) );
  INV_X1 U16441 ( .A(n14909), .ZN(n14912) );
  AOI211_X1 U16442 ( .C1(n14937), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14950) );
  AOI22_X1 U16443 ( .A1(n14949), .A2(n9386), .B1(n14950), .B2(n14948), .ZN(
        P3_U3393) );
  AOI211_X1 U16444 ( .C1(n14937), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        n14952) );
  AOI22_X1 U16445 ( .A1(n14949), .A2(n8908), .B1(n14952), .B2(n14948), .ZN(
        P3_U3396) );
  AOI22_X1 U16446 ( .A1(n14918), .A2(n14937), .B1(n14917), .B2(n14916), .ZN(
        n14919) );
  AND2_X1 U16447 ( .A1(n14920), .A2(n14919), .ZN(n14954) );
  AOI22_X1 U16448 ( .A1(n14949), .A2(n9517), .B1(n14954), .B2(n14948), .ZN(
        P3_U3399) );
  AOI211_X1 U16449 ( .C1(n14937), .C2(n14923), .A(n14922), .B(n14921), .ZN(
        n14956) );
  AOI22_X1 U16450 ( .A1(n14949), .A2(n9606), .B1(n14956), .B2(n14948), .ZN(
        P3_U3402) );
  INV_X1 U16451 ( .A(n14924), .ZN(n14925) );
  AOI211_X1 U16452 ( .C1(n14927), .C2(n14937), .A(n14926), .B(n14925), .ZN(
        n14957) );
  AOI22_X1 U16453 ( .A1(n14949), .A2(n10009), .B1(n14957), .B2(n14948), .ZN(
        P3_U3405) );
  INV_X1 U16454 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14931) );
  AOI211_X1 U16455 ( .C1(n14930), .C2(n14937), .A(n14929), .B(n14928), .ZN(
        n14959) );
  AOI22_X1 U16456 ( .A1(n14949), .A2(n14931), .B1(n14959), .B2(n14948), .ZN(
        P3_U3408) );
  AOI211_X1 U16457 ( .C1(n14937), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        n14960) );
  AOI22_X1 U16458 ( .A1(n14949), .A2(n10069), .B1(n14960), .B2(n14948), .ZN(
        P3_U3411) );
  AOI211_X1 U16459 ( .C1(n14938), .C2(n14937), .A(n14936), .B(n14935), .ZN(
        n14962) );
  AOI22_X1 U16460 ( .A1(n14949), .A2(n10162), .B1(n14962), .B2(n14948), .ZN(
        P3_U3414) );
  INV_X1 U16461 ( .A(n14939), .ZN(n14940) );
  AOI211_X1 U16462 ( .C1(n14942), .C2(n14946), .A(n14941), .B(n14940), .ZN(
        n14964) );
  AOI22_X1 U16463 ( .A1(n14949), .A2(n10371), .B1(n14964), .B2(n14948), .ZN(
        P3_U3417) );
  INV_X1 U16464 ( .A(n14943), .ZN(n14944) );
  AOI211_X1 U16465 ( .C1(n14947), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14967) );
  AOI22_X1 U16466 ( .A1(n14949), .A2(n10615), .B1(n14967), .B2(n14948), .ZN(
        P3_U3420) );
  AOI22_X1 U16467 ( .A1(n14968), .A2(n14950), .B1(n9027), .B2(n14965), .ZN(
        P3_U3460) );
  INV_X1 U16468 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U16469 ( .A1(n14968), .A2(n14952), .B1(n14951), .B2(n14965), .ZN(
        P3_U3461) );
  INV_X1 U16470 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U16471 ( .A1(n14968), .A2(n14954), .B1(n14953), .B2(n14965), .ZN(
        P3_U3462) );
  AOI22_X1 U16472 ( .A1(n14968), .A2(n14956), .B1(n14955), .B2(n14965), .ZN(
        P3_U3463) );
  AOI22_X1 U16473 ( .A1(n14968), .A2(n14957), .B1(n9281), .B2(n14965), .ZN(
        P3_U3464) );
  AOI22_X1 U16474 ( .A1(n14968), .A2(n14959), .B1(n14958), .B2(n14965), .ZN(
        P3_U3465) );
  AOI22_X1 U16475 ( .A1(n14968), .A2(n14960), .B1(n9682), .B2(n14965), .ZN(
        P3_U3466) );
  AOI22_X1 U16476 ( .A1(n14968), .A2(n14962), .B1(n14961), .B2(n14965), .ZN(
        P3_U3467) );
  INV_X1 U16477 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16478 ( .A1(n14968), .A2(n14964), .B1(n14963), .B2(n14965), .ZN(
        P3_U3468) );
  AOI22_X1 U16479 ( .A1(n14968), .A2(n14967), .B1(n14966), .B2(n14965), .ZN(
        P3_U3469) );
  XOR2_X1 U16480 ( .A(n14970), .B(n14969), .Z(SUB_1596_U59) );
  XOR2_X1 U16481 ( .A(n14972), .B(n14971), .Z(SUB_1596_U58) );
  AOI21_X1 U16482 ( .B1(n14974), .B2(n14973), .A(n14983), .ZN(SUB_1596_U53) );
  XOR2_X1 U16483 ( .A(n14975), .B(n14976), .Z(SUB_1596_U56) );
  OAI21_X1 U16484 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14981) );
  XOR2_X1 U16485 ( .A(n14981), .B(n14980), .Z(SUB_1596_U60) );
  XOR2_X1 U16486 ( .A(n14983), .B(n14982), .Z(SUB_1596_U5) );
  BUF_X2 U7232 ( .A(n8604), .Z(n11208) );
  CLKBUF_X2 U7243 ( .A(n8800), .Z(n6476) );
  CLKBUF_X1 U7257 ( .A(n9074), .Z(n9262) );
  CLKBUF_X1 U7285 ( .A(n8616), .Z(n8617) );
  INV_X1 U7449 ( .A(n9262), .ZN(n11743) );
  CLKBUF_X1 U10860 ( .A(n9072), .Z(n6485) );
  CLKBUF_X1 U11665 ( .A(n7657), .Z(n6832) );
endmodule

