

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181;

  AOI21_X1 U4790 ( .B1(n4671), .B2(n4669), .A(n4668), .ZN(n4667) );
  CLKBUF_X2 U4791 ( .A(n9234), .Z(n4292) );
  XNOR2_X1 U4792 ( .A(n5511), .B(n5510), .ZN(n7450) );
  OAI21_X1 U4793 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(n5480) );
  NAND2_X1 U4794 ( .A1(n4713), .A2(n4715), .ZN(n5467) );
  NAND2_X2 U4795 ( .A1(n5915), .A2(n5914), .ZN(n6992) );
  INV_X2 U4796 ( .A(n5158), .ZN(n7914) );
  OR2_X1 U4797 ( .A1(n5906), .A2(n5905), .ZN(n5917) );
  BUF_X1 U4798 ( .A(n5128), .Z(n5685) );
  AND2_X1 U4799 ( .A1(n5759), .A2(n8220), .ZN(n5820) );
  AND2_X1 U4800 ( .A1(n6181), .A2(n6180), .ZN(n4390) );
  AND2_X2 U4801 ( .A1(n8220), .A2(n7630), .ZN(n5837) );
  BUF_X1 U4803 ( .A(n5773), .Z(n5774) );
  INV_X4 U4804 ( .A(n10141), .ZN(n9677) );
  INV_X1 U4805 ( .A(n7840), .ZN(n7776) );
  NAND2_X1 U4806 ( .A1(n8144), .A2(n7965), .ZN(n8127) );
  OR2_X1 U4807 ( .A1(n9919), .A2(n7487), .ZN(n8008) );
  NAND2_X1 U4808 ( .A1(n5087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4522) );
  INV_X1 U4809 ( .A(n6231), .ZN(n6846) );
  OR2_X1 U4810 ( .A1(n7275), .A2(n7186), .ZN(n7675) );
  NAND2_X1 U4811 ( .A1(n5002), .A2(n4286), .ZN(n5128) );
  MUX2_X1 U4812 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4926), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4927) );
  INV_X1 U4813 ( .A(n8523), .ZN(n8504) );
  OR2_X1 U4814 ( .A1(n8376), .A2(n9910), .ZN(n8011) );
  AND3_X1 U4815 ( .A1(n5114), .A2(n5113), .A3(n5112), .ZN(n7099) );
  NAND2_X1 U4816 ( .A1(n4764), .A2(n4762), .ZN(n6009) );
  NAND2_X1 U4817 ( .A1(n7644), .A2(n9713), .ZN(n7775) );
  OAI21_X1 U4818 ( .B1(n6158), .B2(n6157), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6159) );
  NAND2_X1 U4819 ( .A1(n5270), .A2(n5269), .ZN(n5279) );
  OAI222_X1 U4820 ( .A1(n8646), .A2(n8505), .B1(n8633), .B2(n8504), .C1(n8650), 
        .C2(n8503), .ZN(n8671) );
  AND2_X1 U4821 ( .A1(n7109), .A2(n8128), .ZN(n9862) );
  NAND2_X1 U4822 ( .A1(n5304), .A2(n5303), .ZN(n7496) );
  NAND2_X1 U4823 ( .A1(n8072), .A2(n8073), .ZN(n8582) );
  INV_X1 U4824 ( .A(n5845), .ZN(n6210) );
  XNOR2_X1 U4825 ( .A(n6159), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6181) );
  XNOR2_X1 U4826 ( .A(n5279), .B(n5278), .ZN(n6543) );
  NAND4_X1 U4828 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n8980)
         );
  XNOR2_X1 U4829 ( .A(n6111), .B(n6110), .ZN(n7840) );
  INV_X1 U4830 ( .A(n5819), .ZN(n6139) );
  AND3_X2 U4831 ( .A1(n5979), .A2(n4835), .A3(n4761), .ZN(n4500) );
  AND3_X2 U4832 ( .A1(n5979), .A2(n4460), .A3(n4761), .ZN(n6108) );
  BUF_X2 U4833 ( .A(n5150), .Z(n4284) );
  AOI21_X2 U4834 ( .B1(n8060), .B2(n4376), .A(n4375), .ZN(n4374) );
  NAND2_X2 U4835 ( .A1(n9521), .A2(n9522), .ZN(n7284) );
  INV_X1 U4836 ( .A(n5819), .ZN(n4285) );
  AOI21_X2 U4837 ( .B1(n8500), .B2(n8107), .A(n8106), .ZN(n8489) );
  NAND2_X1 U4838 ( .A1(n4927), .A2(n5087), .ZN(n4286) );
  NAND2_X1 U4839 ( .A1(n4927), .A2(n5087), .ZN(n4287) );
  NAND2_X1 U4840 ( .A1(n4927), .A2(n5087), .ZN(n5675) );
  AOI21_X2 U4841 ( .B1(n9802), .B2(n5012), .A(n6883), .ZN(n6888) );
  INV_X1 U4842 ( .A(n6433), .ZN(n4288) );
  INV_X2 U4843 ( .A(n6433), .ZN(n6448) );
  OR2_X2 U4844 ( .A1(n9322), .A2(n9405), .ZN(n9302) );
  NOR2_X2 U4845 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7076) );
  OAI222_X1 U4846 ( .A1(P1_U3086), .A2(n7840), .B1(n9478), .B2(n7388), .C1(
        n7387), .C2(n8222), .ZN(P1_U3334) );
  NAND2_X2 U4847 ( .A1(n6109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6111) );
  XNOR2_X2 U4848 ( .A(n4522), .B(n4924), .ZN(n5002) );
  OAI21_X2 U4849 ( .B1(n9169), .B2(n9175), .A(n7733), .ZN(n9151) );
  AOI21_X2 U4850 ( .B1(n9191), .B2(n6075), .A(n6074), .ZN(n9174) );
  NAND2_X2 U4851 ( .A1(n5282), .A2(n5281), .ZN(n9919) );
  NOR2_X2 U4853 ( .A1(n9793), .A2(n9794), .ZN(n9792) );
  XNOR2_X2 U4854 ( .A(n5491), .B(n5481), .ZN(n7343) );
  AOI22_X2 U4855 ( .A1(n9335), .A2(n9334), .B1(n8969), .B2(n9415), .ZN(n9321)
         );
  OAI22_X2 U4856 ( .A1(n6009), .A2(n6008), .B1(n6132), .B2(n8958), .ZN(n9335)
         );
  NOR2_X2 U4857 ( .A1(n5013), .A2(n9816), .ZN(n5015) );
  NAND3_X1 U4858 ( .A1(n4834), .A2(n8848), .A3(n6396), .ZN(n8847) );
  NAND2_X1 U4859 ( .A1(n9439), .A2(n8962), .ZN(n7734) );
  INV_X1 U4860 ( .A(n7257), .ZN(n9905) );
  AND3_X1 U4861 ( .A1(n5197), .A2(n5196), .A3(n5195), .ZN(n8204) );
  INV_X1 U4862 ( .A(n6943), .ZN(n9703) );
  AND3_X1 U4863 ( .A1(n5173), .A2(n5172), .A3(n5171), .ZN(n8215) );
  INV_X1 U4864 ( .A(n5149), .ZN(n9871) );
  AND2_X1 U4865 ( .A1(n4595), .A2(n4594), .ZN(n8726) );
  BUF_X2 U4866 ( .A(n5177), .Z(n5438) );
  INV_X2 U4867 ( .A(n6249), .ZN(n5834) );
  INV_X4 U4868 ( .A(n5685), .ZN(n4289) );
  BUF_X2 U4869 ( .A(n5179), .Z(n4290) );
  CLKBUF_X2 U4870 ( .A(n6235), .Z(n7053) );
  AND4_X2 U4872 ( .A1(n5746), .A2(n5744), .A3(n5745), .A4(n5743), .ZN(n5979)
         );
  INV_X2 U4873 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI21_X1 U4874 ( .B1(n4487), .B2(n4490), .A(n4380), .ZN(n4482) );
  AOI21_X1 U4875 ( .B1(n8832), .B2(n6478), .A(n6477), .ZN(n6479) );
  AND2_X1 U4876 ( .A1(n4495), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U4877 ( .A1(n4812), .A2(n4810), .ZN(n8879) );
  AND2_X1 U4878 ( .A1(n9146), .A2(n9142), .ZN(n6153) );
  NAND2_X1 U4879 ( .A1(n4461), .A2(n7749), .ZN(n7759) );
  OAI21_X1 U4880 ( .B1(n8345), .B2(n4632), .A(n4631), .ZN(n8194) );
  AND2_X1 U4881 ( .A1(n9356), .A2(n9750), .ZN(n4428) );
  AOI21_X1 U4882 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n7894) );
  NAND2_X1 U4883 ( .A1(n8847), .A2(n8848), .ZN(n6406) );
  OR2_X2 U4884 ( .A1(n9109), .A2(n7758), .ZN(n7901) );
  NAND2_X1 U4885 ( .A1(n6205), .A2(n6204), .ZN(n9109) );
  NAND2_X1 U4886 ( .A1(n7925), .A2(n7920), .ZN(n8105) );
  NAND2_X1 U4887 ( .A1(n6209), .A2(n6208), .ZN(n9115) );
  XNOR2_X1 U4888 ( .A(n6189), .B(n6188), .ZN(n6192) );
  NAND2_X1 U4889 ( .A1(n5621), .A2(n5620), .ZN(n6189) );
  AOI21_X2 U4890 ( .B1(n7607), .B2(n6210), .A(n4371), .ZN(n9439) );
  AND2_X1 U4891 ( .A1(n4674), .A2(n4672), .ZN(n4671) );
  OR2_X1 U4892 ( .A1(n4819), .A2(n4445), .ZN(n4443) );
  NAND2_X1 U4893 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  OR2_X1 U4894 ( .A1(n8612), .A2(n8611), .ZN(n8704) );
  NAND2_X1 U4895 ( .A1(n5776), .A2(n5775), .ZN(n9380) );
  OR2_X1 U4896 ( .A1(n6346), .A2(n6345), .ZN(n4818) );
  INV_X1 U4897 ( .A(n9275), .ZN(n7634) );
  NAND2_X1 U4898 ( .A1(n5501), .A2(n5500), .ZN(n8772) );
  OR2_X1 U4899 ( .A1(n9453), .A2(n8967), .ZN(n7633) );
  AOI21_X2 U4900 ( .B1(n7450), .B2(n6210), .A(n4364), .ZN(n9453) );
  NAND2_X2 U4901 ( .A1(n6037), .A2(n6036), .ZN(n9265) );
  AOI22_X1 U4902 ( .A1(n8235), .A2(n8234), .B1(n8153), .B2(n8152), .ZN(n8356)
         );
  NAND2_X1 U4903 ( .A1(n5483), .A2(n5482), .ZN(n8778) );
  OR2_X1 U4904 ( .A1(n6035), .A2(n9296), .ZN(n9258) );
  OAI21_X1 U4905 ( .B1(n7286), .B2(n4802), .A(n4801), .ZN(n4800) );
  NAND2_X1 U4906 ( .A1(n5794), .A2(n5793), .ZN(n9399) );
  AND2_X1 U4907 ( .A1(n4441), .A2(n6314), .ZN(n4440) );
  NAND2_X1 U4908 ( .A1(n6086), .A2(n6085), .ZN(n8963) );
  AOI21_X1 U4909 ( .B1(n4831), .B2(n4829), .A(n4828), .ZN(n4827) );
  AOI22_X1 U4910 ( .A1(n7358), .A2(n7357), .B1(n7356), .B2(n7355), .ZN(n7360)
         );
  NOR2_X1 U4911 ( .A1(n5966), .A2(n8972), .ZN(n4293) );
  NAND2_X1 U4912 ( .A1(n6073), .A2(n6072), .ZN(n8964) );
  AND2_X1 U4913 ( .A1(n6126), .A2(n7671), .ZN(n7848) );
  NAND2_X1 U4914 ( .A1(n5766), .A2(n5765), .ZN(n8966) );
  NAND2_X1 U4915 ( .A1(n5987), .A2(n5986), .ZN(n9430) );
  NAND2_X1 U4916 ( .A1(n4720), .A2(n4718), .ZN(n5399) );
  AOI21_X1 U4917 ( .B1(n9249), .B2(n6139), .A(n6053), .ZN(n9234) );
  INV_X4 U4918 ( .A(n8184), .ZN(n4291) );
  OR2_X1 U4919 ( .A1(n6503), .A2(n9943), .ZN(n6731) );
  MUX2_X1 U4920 ( .A(n7977), .B(n7976), .S(n8128), .Z(n7978) );
  NAND4_X2 U4921 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n7143)
         );
  OR2_X1 U4922 ( .A1(n7101), .A2(n7099), .ZN(n7970) );
  OR2_X1 U4923 ( .A1(n7098), .A2(n8726), .ZN(n6894) );
  NAND4_X2 U4924 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n7101)
         );
  BUF_X1 U4925 ( .A(n6225), .Z(n8983) );
  NAND4_X2 U4926 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n9861)
         );
  INV_X1 U4927 ( .A(n6446), .ZN(n6409) );
  NAND2_X1 U4928 ( .A1(n5816), .A2(n4886), .ZN(n7043) );
  CLKBUF_X3 U4929 ( .A(n5175), .Z(n7134) );
  NAND2_X1 U4930 ( .A1(n5094), .A2(n5095), .ZN(n5175) );
  NAND2_X1 U4931 ( .A1(n5094), .A2(n8819), .ZN(n5177) );
  NAND4_X1 U4932 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n8982)
         );
  CLKBUF_X1 U4933 ( .A(n5179), .Z(n7137) );
  NAND2_X1 U4934 ( .A1(n5096), .A2(n8819), .ZN(n5179) );
  CLKBUF_X3 U4935 ( .A(n5820), .Z(n7751) );
  INV_X1 U4936 ( .A(n6032), .ZN(n7752) );
  OAI211_X1 U4937 ( .C1(n5845), .C2(n6522), .A(n4687), .B(n4686), .ZN(n6235)
         );
  INV_X1 U4938 ( .A(n5821), .ZN(n6032) );
  AND2_X1 U4939 ( .A1(n4884), .A2(n4737), .ZN(n4735) );
  NAND2_X2 U4940 ( .A1(n6138), .A2(n6217), .ZN(n6548) );
  NAND2_X1 U4941 ( .A1(n4635), .A2(n4333), .ZN(n5087) );
  XNOR2_X1 U4942 ( .A(n4740), .B(n5772), .ZN(n6217) );
  OR2_X1 U4943 ( .A1(n5771), .A2(n9473), .ZN(n4740) );
  MUX2_X1 U4944 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5768), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5770) );
  NOR2_X2 U4945 ( .A1(n5767), .A2(n5754), .ZN(n5756) );
  INV_X4 U4946 ( .A(n5774), .ZN(n6514) );
  CLKBUF_X2 U4947 ( .A(n5003), .Z(n9771) );
  XNOR2_X1 U4948 ( .A(n6114), .B(n6113), .ZN(n7296) );
  INV_X1 U4949 ( .A(n5773), .ZN(n5325) );
  OAI21_X1 U4950 ( .B1(n5138), .B2(n5107), .A(n5106), .ZN(n5131) );
  NOR2_X1 U4951 ( .A1(n4949), .A2(n4953), .ZN(n5003) );
  NAND2_X1 U4952 ( .A1(n4500), .A2(n4760), .ZN(n5767) );
  NOR2_X1 U4953 ( .A1(n4759), .A2(n5830), .ZN(n4758) );
  NAND2_X1 U4954 ( .A1(n4865), .A2(n5083), .ZN(n4864) );
  NAND2_X2 U4955 ( .A1(n5105), .A2(n5104), .ZN(n5138) );
  NAND2_X1 U4956 ( .A1(n5004), .A2(n4948), .ZN(n4955) );
  AND2_X2 U4957 ( .A1(n4423), .A2(n4422), .ZN(n5004) );
  AND3_X1 U4958 ( .A1(n4895), .A2(n4894), .A3(n4893), .ZN(n4898) );
  AND3_X1 U4959 ( .A1(n10058), .A2(n6107), .A3(n6174), .ZN(n5750) );
  NOR2_X1 U4960 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5744) );
  INV_X1 U4961 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10058) );
  INV_X1 U4962 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5982) );
  INV_X1 U4963 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6107) );
  NOR2_X1 U4964 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5740) );
  INV_X1 U4965 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6174) );
  AND2_X1 U4966 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7077) );
  NOR2_X2 U4967 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5826) );
  INV_X1 U4968 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5772) );
  INV_X4 U4969 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X2 U4970 ( .A1(n5594), .A2(n5575), .ZN(n8517) );
  NAND2_X2 U4971 ( .A1(n7909), .A2(n7900), .ZN(n6229) );
  NOR2_X2 U4972 ( .A1(n5862), .A2(n6777), .ZN(n5881) );
  OR2_X2 U4973 ( .A1(n8748), .A2(n8504), .ZN(n8101) );
  NOR2_X2 U4974 ( .A1(n9177), .A2(n9192), .ZN(n9176) );
  INV_X2 U4975 ( .A(n8100), .ZN(n8512) );
  AND2_X2 U4976 ( .A1(n8090), .A2(n8101), .ZN(n8100) );
  OAI21_X1 U4977 ( .B1(n8113), .B2(n8105), .A(n8114), .ZN(n8119) );
  OAI211_X2 U4978 ( .C1(n8111), .C2(n8501), .A(n8110), .B(n8109), .ZN(n8114)
         );
  NOR2_X2 U4979 ( .A1(n5917), .A2(n5916), .ZN(n5933) );
  NAND2_X2 U4980 ( .A1(n5580), .A2(n5579), .ZN(n8523) );
  NOR2_X4 U4981 ( .A1(n9265), .A2(n9279), .ZN(n9264) );
  NAND2_X1 U4982 ( .A1(n9109), .A2(n7758), .ZN(n7893) );
  OR2_X1 U4983 ( .A1(n5715), .A2(n8368), .ZN(n7925) );
  NOR2_X1 U4984 ( .A1(n4550), .A2(n4864), .ZN(n4547) );
  INV_X1 U4985 ( .A(n5138), .ZN(n5773) );
  NAND2_X1 U4986 ( .A1(n5566), .A2(n5565), .ZN(n5582) );
  INV_X1 U4987 ( .A(n8400), .ZN(n4580) );
  NAND2_X1 U4988 ( .A1(n4498), .A2(n4492), .ZN(n4491) );
  INV_X1 U4989 ( .A(n7835), .ZN(n4497) );
  INV_X1 U4990 ( .A(n7768), .ZN(n4492) );
  AND2_X1 U4991 ( .A1(n9157), .A2(n4745), .ZN(n4741) );
  NAND2_X1 U4992 ( .A1(n9177), .A2(n8963), .ZN(n4745) );
  AND2_X1 U4993 ( .A1(n4507), .A2(n7716), .ZN(n4506) );
  OR2_X1 U4994 ( .A1(n4508), .A2(n7713), .ZN(n4501) );
  INV_X1 U4995 ( .A(n7708), .ZN(n4509) );
  AND2_X1 U4996 ( .A1(n7283), .A2(n8468), .ZN(n5712) );
  NAND2_X1 U4997 ( .A1(n5366), .A2(n4324), .ZN(n4720) );
  NAND2_X1 U4998 ( .A1(n5380), .A2(SI_14_), .ZN(n4722) );
  INV_X1 U4999 ( .A(n8163), .ZN(n4601) );
  AND2_X1 U5000 ( .A1(n8125), .A2(n7920), .ZN(n8112) );
  NAND2_X1 U5001 ( .A1(n6695), .A2(n4645), .ZN(n6679) );
  AOI21_X1 U5002 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6568), .A(n7378), .ZN(
        n5017) );
  NOR2_X1 U5003 ( .A1(n8444), .A2(n4421), .ZN(n5023) );
  AND2_X1 U5004 ( .A1(n8443), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U5005 ( .A1(n5657), .A2(n4880), .ZN(n5656) );
  NAND2_X1 U5006 ( .A1(n8648), .A2(n5654), .ZN(n8629) );
  NAND2_X1 U5007 ( .A1(n4906), .A2(n4634), .ZN(n4636) );
  NOR3_X1 U5008 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4906) );
  INV_X1 U5009 ( .A(n4455), .ZN(n4454) );
  NOR2_X1 U5010 ( .A1(n9159), .A2(n6474), .ZN(n6213) );
  INV_X1 U5011 ( .A(n4778), .ZN(n4777) );
  INV_X1 U5012 ( .A(n9422), .ZN(n4766) );
  AOI21_X1 U5013 ( .B1(n4769), .B2(n4293), .A(n4354), .ZN(n4767) );
  NAND2_X1 U5014 ( .A1(n6548), .A2(n4300), .ZN(n4687) );
  NAND2_X1 U5015 ( .A1(n6117), .A2(n7042), .ZN(n7041) );
  NAND2_X2 U5016 ( .A1(n7776), .A2(n7296), .ZN(n6231) );
  NOR2_X1 U5017 ( .A1(n4836), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4835) );
  NAND2_X1 U5018 ( .A1(n4837), .A2(n5772), .ZN(n4836) );
  INV_X1 U5019 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4837) );
  NAND2_X1 U5020 ( .A1(n5604), .A2(n5603), .ZN(n5617) );
  AND2_X1 U5021 ( .A1(n5546), .A2(n5532), .ZN(n5544) );
  AOI21_X1 U5022 ( .B1(n5434), .B2(n4716), .A(n4304), .ZN(n4715) );
  NAND2_X1 U5023 ( .A1(n5350), .A2(n5349), .ZN(n5366) );
  INV_X1 U5024 ( .A(n5256), .ZN(n4710) );
  NOR2_X1 U5025 ( .A1(n5278), .A2(n4712), .ZN(n4711) );
  OAI21_X1 U5026 ( .B1(n6514), .B2(n4417), .A(n4416), .ZN(n5252) );
  NAND2_X1 U5027 ( .A1(n6514), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4416) );
  AND2_X1 U5028 ( .A1(n4617), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U5029 ( .A1(n8185), .A2(n8246), .ZN(n8267) );
  AND2_X1 U5030 ( .A1(n4609), .A2(n4607), .ZN(n4296) );
  INV_X1 U5031 ( .A(n7243), .ZN(n4607) );
  INV_X1 U5032 ( .A(n4864), .ZN(n4545) );
  INV_X1 U5033 ( .A(n5438), .ZN(n5625) );
  NAND3_X1 U5034 ( .A1(n4574), .A2(n4346), .A3(n4575), .ZN(n4573) );
  NOR2_X1 U5035 ( .A1(n8409), .A2(n4373), .ZN(n5021) );
  XNOR2_X1 U5036 ( .A(n5671), .B(n8105), .ZN(n4543) );
  AOI22_X1 U5037 ( .A1(n8513), .A2(n5668), .B1(n5667), .B2(n8504), .ZN(n8502)
         );
  OAI21_X1 U5038 ( .B1(n8616), .B2(n8618), .A(n7930), .ZN(n8612) );
  INV_X1 U5039 ( .A(n5155), .ZN(n5206) );
  AOI21_X1 U5040 ( .B1(n8567), .B2(n8078), .A(n8080), .ZN(n8555) );
  OR2_X1 U5041 ( .A1(n7568), .A2(n7563), .ZN(n8031) );
  NAND2_X1 U5042 ( .A1(n5774), .A2(n5128), .ZN(n5158) );
  XNOR2_X1 U5043 ( .A(n4919), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7965) );
  INV_X1 U5044 ( .A(n4550), .ZN(n4548) );
  INV_X1 U5045 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4900) );
  AND2_X1 U5046 ( .A1(n4938), .A2(n4937), .ZN(n5368) );
  XNOR2_X1 U5047 ( .A(n6177), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U5048 ( .A1(n8879), .A2(n8880), .ZN(n6481) );
  NAND2_X1 U5049 ( .A1(n4489), .A2(n4493), .ZN(n4488) );
  INV_X1 U5050 ( .A(n7902), .ZN(n4494) );
  INV_X1 U5051 ( .A(n4285), .ZN(n6081) );
  NAND2_X1 U5052 ( .A1(n6213), .A2(n6212), .ZN(n9132) );
  NAND2_X1 U5053 ( .A1(n4725), .A2(n6211), .ZN(n7742) );
  INV_X1 U5054 ( .A(n6213), .ZN(n9131) );
  AND2_X1 U5055 ( .A1(n7801), .A2(n4321), .ZN(n4743) );
  INV_X1 U5056 ( .A(n6465), .ZN(n6460) );
  NAND2_X1 U5057 ( .A1(n9240), .A2(n4794), .ZN(n4790) );
  AOI21_X1 U5058 ( .B1(n6536), .B2(n6538), .A(n6540), .ZN(n6842) );
  NAND2_X1 U5059 ( .A1(n6077), .A2(n6076), .ZN(n9177) );
  AND2_X1 U5060 ( .A1(n6496), .A2(n6226), .ZN(n7907) );
  XNOR2_X1 U5061 ( .A(n6202), .B(n6201), .ZN(n8813) );
  OAI21_X1 U5062 ( .B1(n6207), .B2(n6206), .A(n6198), .ZN(n6202) );
  OR2_X1 U5063 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5754) );
  NAND2_X1 U5064 ( .A1(n5300), .A2(n5301), .ZN(n5312) );
  NAND2_X1 U5065 ( .A1(n5160), .A2(n5159), .ZN(n5169) );
  NAND2_X1 U5066 ( .A1(n4323), .A2(n4385), .ZN(n4384) );
  INV_X1 U5067 ( .A(n8469), .ZN(n4385) );
  NAND2_X1 U5068 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  OAI211_X1 U5069 ( .C1(n7767), .C2(n7766), .A(n7893), .B(n7765), .ZN(n7903)
         );
  INV_X1 U5070 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U5071 ( .A1(n4690), .A2(n9665), .ZN(n4689) );
  OAI22_X1 U5072 ( .A1(n9127), .A2(n9721), .B1(n9124), .B2(n9123), .ZN(n9125)
         );
  NAND2_X1 U5073 ( .A1(n7653), .A2(n7650), .ZN(n7649) );
  INV_X1 U5074 ( .A(n4472), .ZN(n4471) );
  OAI21_X1 U5075 ( .B1(n4473), .B2(n4314), .A(n4476), .ZN(n4472) );
  NAND2_X1 U5076 ( .A1(n7663), .A2(n7897), .ZN(n4476) );
  OR2_X1 U5077 ( .A1(n4360), .A2(n7897), .ZN(n4473) );
  OR2_X1 U5078 ( .A1(n4314), .A2(n7897), .ZN(n4474) );
  MUX2_X1 U5079 ( .A(n7704), .B(n7813), .S(n7760), .Z(n7705) );
  NOR2_X1 U5080 ( .A1(n7806), .A2(n7760), .ZN(n4513) );
  NOR2_X1 U5081 ( .A1(n4514), .A2(n7717), .ZN(n4505) );
  NAND2_X1 U5082 ( .A1(n7814), .A2(n7760), .ZN(n4514) );
  MUX2_X1 U5083 ( .A(n7720), .B(n7719), .S(n7760), .Z(n7721) );
  INV_X1 U5084 ( .A(n8570), .ZN(n4563) );
  NAND2_X1 U5085 ( .A1(n6894), .A2(n7970), .ZN(n7966) );
  INV_X1 U5086 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4887) );
  INV_X1 U5087 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4888) );
  AND2_X1 U5088 ( .A1(n9380), .A2(n8966), .ZN(n4798) );
  NOR2_X1 U5089 ( .A1(n5380), .A2(SI_14_), .ZN(n4721) );
  INV_X1 U5090 ( .A(n7564), .ZN(n4615) );
  NAND2_X1 U5091 ( .A1(n4311), .A2(n7489), .ZN(n4619) );
  INV_X1 U5092 ( .A(n7490), .ZN(n4620) );
  NOR2_X1 U5093 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  NAND2_X1 U5094 ( .A1(n4643), .A2(n6679), .ZN(n6696) );
  NAND2_X1 U5095 ( .A1(n4957), .A2(n6695), .ZN(n6673) );
  NAND2_X1 U5096 ( .A1(n5008), .A2(n6678), .ZN(n6682) );
  INV_X1 U5097 ( .A(n6724), .ZN(n4592) );
  OR2_X1 U5098 ( .A1(n6728), .A2(n4359), .ZN(n4382) );
  AND2_X1 U5099 ( .A1(n6879), .A2(n4983), .ZN(n4985) );
  OAI21_X1 U5100 ( .B1(n4538), .B2(n4536), .A(n5643), .ZN(n4535) );
  AND2_X1 U5101 ( .A1(n4299), .A2(n4883), .ZN(n4538) );
  OAI21_X1 U5102 ( .B1(n7933), .B2(n4527), .A(n5637), .ZN(n4526) );
  INV_X1 U5103 ( .A(n5636), .ZN(n4527) );
  OR2_X1 U5104 ( .A1(n5693), .A2(n5711), .ZN(n5724) );
  AND2_X1 U5105 ( .A1(n8748), .A2(n8504), .ZN(n7927) );
  NOR2_X1 U5106 ( .A1(n8095), .A2(n4849), .ZN(n4848) );
  AND2_X1 U5107 ( .A1(n4850), .A2(n5508), .ZN(n4849) );
  OR2_X1 U5108 ( .A1(n8760), .A2(n8246), .ZN(n8094) );
  INV_X1 U5109 ( .A(n8557), .ZN(n4555) );
  INV_X1 U5110 ( .A(n8556), .ZN(n4552) );
  NAND2_X1 U5111 ( .A1(n4558), .A2(n4563), .ZN(n4557) );
  OAI21_X1 U5112 ( .B1(n4561), .B2(n5661), .A(n8569), .ZN(n4558) );
  NAND2_X1 U5113 ( .A1(n4560), .A2(n4563), .ZN(n4559) );
  OR2_X1 U5114 ( .A1(n8702), .A2(n8165), .ZN(n8053) );
  NOR2_X1 U5115 ( .A1(n8652), .A2(n4516), .ZN(n4515) );
  INV_X1 U5116 ( .A(n5652), .ZN(n4516) );
  OR2_X1 U5117 ( .A1(n8805), .A2(n8634), .ZN(n8048) );
  INV_X1 U5118 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5119 ( .A1(n4917), .A2(n4336), .ZN(n4381) );
  INV_X1 U5120 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4921) );
  OAI22_X1 U5121 ( .A1(n5004), .A2(n4658), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        P2_IR_REG_2__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U5122 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4658) );
  NAND2_X1 U5123 ( .A1(n6298), .A2(n6297), .ZN(n4832) );
  INV_X1 U5124 ( .A(n4833), .ZN(n4828) );
  AOI21_X1 U5125 ( .B1(n6310), .B2(n6311), .A(n4320), .ZN(n4833) );
  INV_X1 U5126 ( .A(n6297), .ZN(n4829) );
  NAND2_X1 U5127 ( .A1(n6290), .A2(n6289), .ZN(n7031) );
  INV_X1 U5128 ( .A(n4823), .ZN(n4822) );
  XNOR2_X1 U5129 ( .A(n6266), .B(n6446), .ZN(n6270) );
  INV_X1 U5130 ( .A(n7748), .ZN(n7749) );
  NAND2_X1 U5131 ( .A1(n4463), .A2(n4462), .ZN(n4461) );
  MUX2_X1 U5132 ( .A(n7885), .B(n7747), .S(n7760), .Z(n7748) );
  INV_X1 U5133 ( .A(n7630), .ZN(n5759) );
  AND2_X1 U5134 ( .A1(n5760), .A2(n7630), .ZN(n5821) );
  NAND2_X1 U5135 ( .A1(n7628), .A2(n6210), .ZN(n4725) );
  NAND2_X1 U5136 ( .A1(n4789), .A2(n4341), .ZN(n4787) );
  NAND2_X1 U5137 ( .A1(n9453), .A2(n4292), .ZN(n4793) );
  NOR2_X1 U5138 ( .A1(n4798), .A2(n4795), .ZN(n4794) );
  INV_X1 U5139 ( .A(n6054), .ZN(n4795) );
  NOR2_X1 U5140 ( .A1(n4798), .A2(n4793), .ZN(n4792) );
  INV_X1 U5141 ( .A(n4779), .ZN(n4776) );
  INV_X1 U5142 ( .A(n4664), .ZN(n4663) );
  OAI21_X1 U5143 ( .B1(n9341), .B2(n4665), .A(n7698), .ZN(n4664) );
  INV_X1 U5144 ( .A(n7868), .ZN(n4665) );
  NOR2_X1 U5145 ( .A1(n7460), .A2(n4431), .ZN(n4430) );
  INV_X1 U5146 ( .A(n4432), .ZN(n4431) );
  INV_X1 U5147 ( .A(n6131), .ZN(n4682) );
  NAND2_X1 U5148 ( .A1(n9642), .A2(n6347), .ZN(n4771) );
  OR2_X1 U5149 ( .A1(n7294), .A2(n7338), .ZN(n4877) );
  INV_X1 U5150 ( .A(n7685), .ZN(n4684) );
  NAND2_X1 U5151 ( .A1(n7297), .A2(n6131), .ZN(n4685) );
  OAI21_X1 U5152 ( .B1(n6192), .B2(n6191), .A(n6190), .ZN(n6207) );
  OR2_X1 U5153 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NAND2_X1 U5154 ( .A1(n4695), .A2(n5546), .ZN(n4694) );
  NAND2_X1 U5155 ( .A1(n4697), .A2(n4699), .ZN(n4695) );
  AND2_X1 U5156 ( .A1(n5565), .A2(n5551), .ZN(n5563) );
  AND2_X1 U5157 ( .A1(n4839), .A2(n6110), .ZN(n4838) );
  NAND2_X1 U5158 ( .A1(n4739), .A2(SI_20_), .ZN(n4738) );
  OAI21_X1 U5159 ( .B1(n5312), .B2(n4728), .A(n4726), .ZN(n5350) );
  INV_X1 U5160 ( .A(n4727), .ZN(n4726) );
  OAI21_X1 U5161 ( .B1(n4733), .B2(n4728), .A(n5343), .ZN(n4727) );
  INV_X1 U5162 ( .A(n4729), .ZN(n4728) );
  AND2_X1 U5163 ( .A1(n5365), .A2(n5348), .ZN(n5349) );
  NOR2_X1 U5164 ( .A1(n5323), .A2(n4734), .ZN(n4733) );
  INV_X1 U5165 ( .A(n5311), .ZN(n4734) );
  OR2_X1 U5166 ( .A1(n5953), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U5167 ( .A1(n5826), .A2(n5741), .ZN(n5829) );
  NAND2_X1 U5168 ( .A1(n7077), .A2(n5103), .ZN(n5104) );
  INV_X1 U5169 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5170 ( .A1(n4604), .A2(n4602), .ZN(n7323) );
  NOR2_X1 U5171 ( .A1(n4605), .A2(n4603), .ZN(n4602) );
  INV_X1 U5172 ( .A(n7258), .ZN(n4603) );
  INV_X1 U5173 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6699) );
  OAI21_X1 U5174 ( .B1(n8156), .B2(n4601), .A(n8333), .ZN(n4600) );
  NOR2_X1 U5175 ( .A1(n4601), .A2(n4598), .ZN(n4597) );
  INV_X1 U5176 ( .A(n8355), .ZN(n4598) );
  NAND2_X1 U5177 ( .A1(n4618), .A2(n4311), .ZN(n4617) );
  INV_X1 U5178 ( .A(n7561), .ZN(n4618) );
  NOR2_X1 U5179 ( .A1(n8183), .A2(n8328), .ZN(n4626) );
  INV_X1 U5180 ( .A(n4623), .ZN(n4622) );
  INV_X1 U5181 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6676) );
  AND3_X1 U5182 ( .A1(n5507), .A2(n5506), .A3(n5505), .ZN(n8180) );
  AND3_X1 U5183 ( .A1(n5490), .A2(n5489), .A3(n5488), .ZN(n8315) );
  OR2_X1 U5184 ( .A1(n5175), .A2(n6822), .ZN(n5118) );
  NAND2_X1 U5185 ( .A1(n4573), .A2(n4572), .ZN(n6645) );
  AND2_X1 U5186 ( .A1(n4951), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4572) );
  AOI21_X1 U5187 ( .B1(n6731), .B2(n6729), .A(n6730), .ZN(n6728) );
  NAND2_X1 U5188 ( .A1(n4591), .A2(n4592), .ZN(n4590) );
  NAND2_X1 U5189 ( .A1(n4971), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6725) );
  XNOR2_X1 U5190 ( .A(n4382), .B(n5249), .ZN(n9803) );
  NOR2_X1 U5191 ( .A1(n5011), .A2(n5249), .ZN(n6885) );
  INV_X1 U5192 ( .A(n4382), .ZN(n5011) );
  NAND2_X1 U5193 ( .A1(n9803), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U5194 ( .A1(n4565), .A2(n4564), .ZN(n9814) );
  NAND2_X1 U5195 ( .A1(n4985), .A2(n9816), .ZN(n4564) );
  OR2_X1 U5196 ( .A1(n4985), .A2(n9816), .ZN(n4565) );
  NOR2_X1 U5197 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  INV_X1 U5198 ( .A(n5015), .ZN(n4647) );
  NOR2_X1 U5199 ( .A1(n7368), .A2(n4577), .ZN(n4988) );
  NOR2_X1 U5200 ( .A1(n7384), .A2(n7404), .ZN(n4577) );
  XNOR2_X1 U5201 ( .A(n4388), .B(n8425), .ZN(n8427) );
  NAND2_X1 U5202 ( .A1(n4579), .A2(n4578), .ZN(n4388) );
  NAND2_X1 U5203 ( .A1(n8408), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U5204 ( .A1(n8427), .A2(n8656), .ZN(n8426) );
  NAND2_X1 U5205 ( .A1(n5022), .A2(n4642), .ZN(n4637) );
  OR2_X1 U5206 ( .A1(n8418), .A2(n4639), .ZN(n4638) );
  NAND2_X1 U5207 ( .A1(n4642), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4639) );
  OR2_X1 U5208 ( .A1(n5574), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U5209 ( .A1(n5536), .A2(n5535), .ZN(n5556) );
  INV_X1 U5210 ( .A(n5537), .ZN(n5536) );
  OR2_X1 U5211 ( .A1(n5519), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5537) );
  OR2_X1 U5212 ( .A1(n5502), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5519) );
  OR2_X1 U5213 ( .A1(n5471), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5486) );
  AOI21_X1 U5214 ( .B1(n8637), .B2(n5660), .A(n4875), .ZN(n8589) );
  OR2_X1 U5215 ( .A1(n5371), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5388) );
  OR2_X1 U5216 ( .A1(n7345), .A2(n7943), .ZN(n7347) );
  OR2_X1 U5217 ( .A1(n5262), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5285) );
  INV_X1 U5218 ( .A(n7222), .ZN(n4539) );
  OR2_X1 U5219 ( .A1(n5221), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U5220 ( .A1(n7098), .A2(n4593), .ZN(n6898) );
  INV_X1 U5221 ( .A(n8726), .ZN(n4593) );
  AND3_X1 U5222 ( .A1(n6749), .A2(n5674), .A3(n9928), .ZN(n7401) );
  NAND2_X1 U5223 ( .A1(n5624), .A2(n5623), .ZN(n5715) );
  OR2_X1 U5224 ( .A1(n8672), .A2(n8514), .ZN(n5669) );
  XNOR2_X1 U5225 ( .A(n8495), .B(n8505), .ZN(n8491) );
  NAND2_X1 U5226 ( .A1(n8521), .A2(n4517), .ZN(n8513) );
  OR2_X1 U5227 ( .A1(n8754), .A2(n8535), .ZN(n4517) );
  AND2_X1 U5228 ( .A1(n4519), .A2(n4518), .ZN(n8522) );
  NAND2_X1 U5229 ( .A1(n8760), .A2(n8549), .ZN(n4518) );
  NAND2_X1 U5230 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  NAND2_X1 U5231 ( .A1(n8533), .A2(n8246), .ZN(n4520) );
  AOI21_X1 U5232 ( .B1(n4848), .B2(n4846), .A(n4845), .ZN(n4844) );
  INV_X1 U5233 ( .A(n4850), .ZN(n4846) );
  INV_X1 U5234 ( .A(n8094), .ZN(n4845) );
  INV_X1 U5235 ( .A(n4848), .ZN(n4847) );
  AND2_X1 U5236 ( .A1(n4851), .A2(n5662), .ZN(n4850) );
  OR2_X1 U5237 ( .A1(n8766), .A2(n8560), .ZN(n5664) );
  OR2_X1 U5238 ( .A1(n8092), .A2(n8540), .ZN(n8547) );
  OR2_X1 U5239 ( .A1(n8555), .A2(n5508), .ZN(n4852) );
  AOI21_X1 U5240 ( .B1(n8704), .B2(n4859), .A(n4353), .ZN(n8567) );
  AND2_X1 U5241 ( .A1(n4860), .A2(n8072), .ZN(n4859) );
  NAND2_X1 U5242 ( .A1(n8589), .A2(n5661), .ZN(n4562) );
  NAND2_X1 U5243 ( .A1(n4562), .A2(n4560), .ZN(n8581) );
  AOI21_X1 U5244 ( .B1(n8596), .B2(n4861), .A(n7960), .ZN(n4860) );
  INV_X1 U5245 ( .A(n8053), .ZN(n4861) );
  OAI21_X1 U5246 ( .B1(n8628), .B2(n5412), .A(n8061), .ZN(n8616) );
  INV_X1 U5247 ( .A(n9862), .ZN(n8633) );
  AND4_X1 U5248 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n8647)
         );
  NAND2_X1 U5249 ( .A1(n5684), .A2(n8128), .ZN(n8646) );
  NAND2_X1 U5250 ( .A1(n4529), .A2(n4528), .ZN(n7574) );
  AOI21_X1 U5251 ( .B1(n4530), .B2(n7555), .A(n4343), .ZN(n4528) );
  NAND2_X1 U5252 ( .A1(n5647), .A2(n7558), .ZN(n7441) );
  INV_X1 U5253 ( .A(n8646), .ZN(n9860) );
  NOR2_X1 U5254 ( .A1(n6751), .A2(n6535), .ZN(n6764) );
  INV_X1 U5255 ( .A(n8650), .ZN(n9866) );
  INV_X1 U5256 ( .A(n7603), .ZN(n5694) );
  INV_X1 U5257 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5258 ( .A1(n8814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U5259 ( .A(n5093), .B(n5092), .ZN(n5095) );
  OR2_X1 U5260 ( .A1(n5091), .A2(n5090), .ZN(n5093) );
  NOR2_X1 U5261 ( .A1(n4302), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5262 ( .A1(n4900), .A2(n4868), .ZN(n4867) );
  INV_X1 U5263 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5083) );
  OR2_X1 U5264 ( .A1(n4972), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4975) );
  OR2_X1 U5265 ( .A1(n4955), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4961) );
  INV_X1 U5266 ( .A(n5004), .ZN(n4574) );
  NAND2_X1 U5267 ( .A1(n4571), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5268 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4422), .ZN(n4571) );
  NAND2_X1 U5269 ( .A1(n4297), .A2(n4319), .ZN(n4455) );
  AND2_X1 U5270 ( .A1(n9686), .A2(n6449), .ZN(n6237) );
  NOR2_X1 U5271 ( .A1(n4453), .A2(n4452), .ZN(n4451) );
  INV_X1 U5272 ( .A(n4820), .ZN(n4452) );
  NOR3_X1 U5273 ( .A1(n4822), .A2(n4307), .A3(n4454), .ZN(n4453) );
  AOI21_X1 U5274 ( .B1(n4823), .B2(n4821), .A(n6383), .ZN(n4820) );
  INV_X1 U5275 ( .A(n7284), .ZN(n4807) );
  OAI21_X1 U5276 ( .B1(n7286), .B2(n7285), .A(n6325), .ZN(n4809) );
  CLKBUF_X1 U5277 ( .A(n6280), .Z(n6805) );
  NAND2_X1 U5278 ( .A1(n6270), .A2(n6271), .ZN(n6277) );
  AND2_X1 U5279 ( .A1(n8917), .A2(n4322), .ZN(n4823) );
  NAND2_X1 U5280 ( .A1(n6393), .A2(n6392), .ZN(n4834) );
  XNOR2_X1 U5281 ( .A(n6230), .B(n6446), .ZN(n6242) );
  AND2_X1 U5282 ( .A1(n6235), .A2(n6448), .ZN(n6236) );
  NAND2_X1 U5283 ( .A1(n5759), .A2(n5760), .ZN(n5819) );
  AOI21_X1 U5284 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9587), .A(n9582), .ZN(
        n9592) );
  AOI21_X1 U5285 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9062), .A(n9591), .ZN(
        n9063) );
  INV_X1 U5286 ( .A(n8961), .ZN(n9127) );
  INV_X1 U5287 ( .A(n4793), .ZN(n4791) );
  INV_X1 U5288 ( .A(n4792), .ZN(n4788) );
  OAI22_X1 U5289 ( .A1(n9255), .A2(n6046), .B1(n8968), .B2(n9265), .ZN(n9240)
         );
  AOI21_X1 U5290 ( .B1(n6035), .B2(n8871), .A(n9273), .ZN(n9255) );
  AND2_X1 U5291 ( .A1(n4295), .A2(n4310), .ZN(n4779) );
  NAND2_X1 U5292 ( .A1(n4295), .A2(n4344), .ZN(n4778) );
  AND2_X1 U5293 ( .A1(n9405), .A2(n9295), .ZN(n4782) );
  AND2_X1 U5294 ( .A1(n7874), .A2(n7638), .ZN(n9310) );
  NAND2_X1 U5295 ( .A1(n9342), .A2(n9341), .ZN(n4662) );
  AND2_X1 U5296 ( .A1(n7690), .A2(n7868), .ZN(n9341) );
  NAND2_X1 U5297 ( .A1(n7430), .A2(n6133), .ZN(n9342) );
  NOR2_X1 U5298 ( .A1(n7460), .A2(n9344), .ZN(n6008) );
  NAND2_X1 U5299 ( .A1(n5970), .A2(n5969), .ZN(n6339) );
  NAND2_X1 U5300 ( .A1(n5958), .A2(n5957), .ZN(n7275) );
  AND2_X1 U5301 ( .A1(n7675), .A2(n7860), .ZN(n7270) );
  NAND2_X1 U5302 ( .A1(n7269), .A2(n7270), .ZN(n7297) );
  OR2_X1 U5303 ( .A1(n6992), .A2(n8975), .ZN(n5923) );
  INV_X1 U5304 ( .A(n7785), .ZN(n4691) );
  NAND2_X1 U5305 ( .A1(n4751), .A2(n4753), .ZN(n6987) );
  AOI21_X1 U5306 ( .B1(n6966), .B2(n4754), .A(n4340), .ZN(n4753) );
  NAND2_X1 U5307 ( .A1(n7011), .A2(n4477), .ZN(n7010) );
  NAND2_X1 U5308 ( .A1(n9662), .A2(n6119), .ZN(n6120) );
  NAND2_X1 U5309 ( .A1(n6095), .A2(n6094), .ZN(n6474) );
  AND2_X1 U5310 ( .A1(n6163), .A2(n6180), .ZN(n6536) );
  AND2_X1 U5311 ( .A1(n4760), .A2(n5752), .ZN(n4499) );
  XNOR2_X1 U5312 ( .A(n5617), .B(n5616), .ZN(n7631) );
  XNOR2_X1 U5313 ( .A(n5602), .B(n5601), .ZN(n7607) );
  XNOR2_X1 U5314 ( .A(n5582), .B(n5581), .ZN(n7602) );
  XNOR2_X1 U5315 ( .A(n5545), .B(n5544), .ZN(n7527) );
  NAND2_X1 U5316 ( .A1(n4714), .A2(n5435), .ZN(n5451) );
  OR2_X1 U5317 ( .A1(n5433), .A2(n5434), .ZN(n4714) );
  INV_X1 U5318 ( .A(n5399), .ZN(n5398) );
  NOR2_X1 U5319 ( .A1(n4732), .A2(n5330), .ZN(n4729) );
  NAND2_X1 U5320 ( .A1(n5312), .A2(n4733), .ZN(n4730) );
  NAND2_X1 U5321 ( .A1(n4705), .A2(n4703), .ZN(n5300) );
  INV_X1 U5322 ( .A(n4704), .ZN(n4703) );
  AND2_X1 U5323 ( .A1(n5311), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U5324 ( .A1(n5251), .A2(n5250), .ZN(n5257) );
  NAND2_X1 U5325 ( .A1(n5257), .A2(n5256), .ZN(n5270) );
  NAND2_X1 U5326 ( .A1(n5169), .A2(n5168), .ZN(n5185) );
  NAND2_X1 U5327 ( .A1(n5370), .A2(n5369), .ZN(n8240) );
  NAND2_X1 U5328 ( .A1(n4628), .A2(n8328), .ZN(n4627) );
  AND4_X1 U5329 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n7556)
         );
  INV_X1 U5330 ( .A(n8375), .ZN(n7487) );
  INV_X1 U5331 ( .A(n8655), .ZN(n8153) );
  NAND2_X1 U5332 ( .A1(n4608), .A2(n4609), .ZN(n7242) );
  OR2_X1 U5333 ( .A1(n7241), .A2(n7240), .ZN(n4608) );
  INV_X1 U5334 ( .A(n8514), .ZN(n8348) );
  XNOR2_X1 U5335 ( .A(n4916), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8144) );
  OAI21_X1 U5336 ( .B1(n7959), .B2(n7958), .A(n7957), .ZN(n8140) );
  INV_X1 U5337 ( .A(n8315), .ZN(n8584) );
  XNOR2_X1 U5338 ( .A(n4981), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6882) );
  XNOR2_X1 U5339 ( .A(n4988), .B(n7476), .ZN(n7464) );
  NOR2_X1 U5340 ( .A1(n7464), .A2(n5315), .ZN(n7463) );
  OR2_X1 U5341 ( .A1(n8382), .A2(n4992), .ZN(n4581) );
  INV_X1 U5342 ( .A(n5020), .ZN(n4652) );
  INV_X1 U5343 ( .A(n4579), .ZN(n8399) );
  OR2_X1 U5344 ( .A1(n8418), .A2(n8713), .ZN(n4641) );
  XNOR2_X1 U5345 ( .A(n5021), .B(n5383), .ZN(n8418) );
  NAND2_X1 U5346 ( .A1(n4409), .A2(n4315), .ZN(n4569) );
  AND2_X1 U5347 ( .A1(n5077), .A2(n8461), .ZN(n5078) );
  INV_X1 U5348 ( .A(n4567), .ZN(n8453) );
  NAND2_X1 U5349 ( .A1(n4569), .A2(n4568), .ZN(n4567) );
  INV_X1 U5350 ( .A(n5000), .ZN(n4568) );
  NOR2_X1 U5351 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  AND2_X1 U5352 ( .A1(n5027), .A2(n5675), .ZN(n9821) );
  NAND2_X1 U5353 ( .A1(n4542), .A2(n4540), .ZN(n4840) );
  NOR2_X1 U5354 ( .A1(n4318), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5355 ( .A1(n4543), .A2(n9866), .ZN(n4542) );
  INV_X1 U5356 ( .A(n5686), .ZN(n4541) );
  NAND2_X1 U5357 ( .A1(n5457), .A2(n5456), .ZN(n8695) );
  OR2_X1 U5358 ( .A1(n6570), .A2(n5158), .ZN(n5304) );
  AND2_X1 U5359 ( .A1(n7283), .A2(n5673), .ZN(n9873) );
  AND2_X1 U5360 ( .A1(n6820), .A2(n8607), .ZN(n9881) );
  INV_X1 U5361 ( .A(n8731), .ZN(n8667) );
  INV_X1 U5362 ( .A(n5715), .ZN(n8482) );
  NAND2_X1 U5363 ( .A1(n5334), .A2(n5333), .ZN(n7568) );
  OR2_X1 U5364 ( .A1(n9936), .A2(n9928), .ZN(n8740) );
  XNOR2_X1 U5365 ( .A(n5086), .B(n4868), .ZN(n8468) );
  INV_X1 U5366 ( .A(n4998), .ZN(n4866) );
  NAND2_X1 U5367 ( .A1(n4450), .A2(n4455), .ZN(n8861) );
  NAND2_X1 U5368 ( .A1(n8898), .A2(n4307), .ZN(n4450) );
  NAND2_X1 U5369 ( .A1(n6025), .A2(n6024), .ZN(n9325) );
  NAND2_X1 U5370 ( .A1(n4459), .A2(n8911), .ZN(n4458) );
  NAND2_X1 U5371 ( .A1(n8851), .A2(n4369), .ZN(n4459) );
  NAND2_X1 U5372 ( .A1(n6461), .A2(n9326), .ZN(n8943) );
  AND2_X1 U5373 ( .A1(n6483), .A2(n6482), .ZN(n6429) );
  OAI21_X1 U5374 ( .B1(n9442), .B2(n9528), .A(n6490), .ZN(n6491) );
  NAND2_X1 U5375 ( .A1(n4484), .A2(n7484), .ZN(n4481) );
  NAND2_X1 U5376 ( .A1(n7484), .A2(n7905), .ZN(n4380) );
  INV_X1 U5377 ( .A(n4487), .ZN(n4483) );
  OAI21_X1 U5378 ( .B1(n4480), .B2(n4485), .A(n7910), .ZN(n4479) );
  OR2_X1 U5379 ( .A1(n4486), .A2(n7911), .ZN(n4480) );
  NAND2_X1 U5380 ( .A1(n7903), .A2(n4482), .ZN(n4478) );
  OR2_X1 U5381 ( .A1(n9178), .A2(n6081), .ZN(n6086) );
  AND2_X1 U5382 ( .A1(n4744), .A2(n4321), .ZN(n6103) );
  NAND2_X1 U5383 ( .A1(n6460), .A2(n7907), .ZN(n9326) );
  INV_X1 U5384 ( .A(n6474), .ZN(n9145) );
  NAND2_X1 U5385 ( .A1(n5932), .A2(n5931), .ZN(n7158) );
  NOR2_X1 U5386 ( .A1(n4413), .A2(n9357), .ZN(n4412) );
  NOR2_X1 U5387 ( .A1(n4428), .A2(n4688), .ZN(n4427) );
  INV_X1 U5388 ( .A(n9177), .ZN(n9442) );
  NAND2_X1 U5389 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5792) );
  MUX2_X1 U5390 ( .A(n8003), .B(n8002), .S(n8127), .Z(n8014) );
  AND2_X1 U5391 ( .A1(n7843), .A2(n7760), .ZN(n4470) );
  NOR2_X1 U5392 ( .A1(n4468), .A2(n4467), .ZN(n4466) );
  NAND2_X1 U5393 ( .A1(n7651), .A2(n9713), .ZN(n4467) );
  NOR2_X1 U5394 ( .A1(n7646), .A2(n7645), .ZN(n4468) );
  INV_X1 U5395 ( .A(n6125), .ZN(n7662) );
  NAND2_X1 U5396 ( .A1(n4469), .A2(n4464), .ZN(n7653) );
  OAI21_X1 U5397 ( .B1(n4466), .B2(n4465), .A(n7897), .ZN(n4464) );
  NAND2_X1 U5398 ( .A1(n7842), .A2(n4470), .ZN(n4469) );
  INV_X1 U5399 ( .A(n7647), .ZN(n4465) );
  OAI21_X1 U5400 ( .B1(n7659), .B2(n4474), .A(n4471), .ZN(n7664) );
  NAND2_X1 U5401 ( .A1(n7646), .A2(n9713), .ZN(n7842) );
  INV_X1 U5402 ( .A(n8076), .ZN(n4405) );
  INV_X1 U5403 ( .A(n6117), .ZN(n7772) );
  INV_X1 U5404 ( .A(n4511), .ZN(n4510) );
  AOI21_X1 U5405 ( .B1(n7708), .B2(n7710), .A(n4512), .ZN(n4511) );
  AOI211_X1 U5406 ( .C1(n7730), .C2(n7729), .A(n7823), .B(n7728), .ZN(n7731)
         );
  OR2_X1 U5407 ( .A1(n4591), .A2(n4878), .ZN(n4584) );
  INV_X1 U5408 ( .A(n4583), .ZN(n4582) );
  INV_X1 U5409 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4892) );
  AOI21_X1 U5410 ( .B1(n7740), .B2(n7897), .A(n4347), .ZN(n4463) );
  AND2_X1 U5411 ( .A1(n7744), .A2(n7760), .ZN(n7745) );
  NAND2_X1 U5412 ( .A1(n4725), .A2(n4723), .ZN(n7827) );
  NOR2_X1 U5413 ( .A1(n7741), .A2(n4724), .ZN(n4723) );
  INV_X1 U5414 ( .A(n6211), .ZN(n4724) );
  OR2_X1 U5415 ( .A1(n9265), .A2(n7769), .ZN(n7712) );
  NAND2_X1 U5416 ( .A1(n6980), .A2(n7783), .ZN(n6125) );
  NAND2_X1 U5417 ( .A1(n5746), .A2(n5744), .ZN(n4759) );
  AOI21_X1 U5418 ( .B1(n4700), .B2(n5528), .A(n4698), .ZN(n4697) );
  INV_X1 U5419 ( .A(n5544), .ZN(n4698) );
  INV_X1 U5420 ( .A(n5492), .ZN(n5493) );
  NOR2_X1 U5421 ( .A1(n5450), .A2(n4717), .ZN(n4716) );
  INV_X1 U5422 ( .A(n5435), .ZN(n4717) );
  INV_X1 U5423 ( .A(n5414), .ZN(n5416) );
  NAND2_X1 U5424 ( .A1(n4720), .A2(n4326), .ZN(n5397) );
  INV_X1 U5425 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5102) );
  AND2_X1 U5426 ( .A1(n4630), .A2(n8324), .ZN(n4629) );
  INV_X1 U5427 ( .A(n8183), .ZN(n4630) );
  NAND2_X1 U5428 ( .A1(n5691), .A2(n5690), .ZN(n7095) );
  OAI21_X1 U5429 ( .B1(n4629), .B2(n8560), .A(n4624), .ZN(n4623) );
  NAND2_X1 U5430 ( .A1(n4625), .A2(n8183), .ZN(n4624) );
  INV_X1 U5431 ( .A(n8324), .ZN(n4625) );
  OR2_X1 U5432 ( .A1(n7488), .A2(n7487), .ZN(n7489) );
  NOR2_X1 U5433 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4897) );
  INV_X1 U5434 ( .A(n4867), .ZN(n4865) );
  NAND2_X1 U5435 ( .A1(n7926), .A2(n8127), .ZN(n8117) );
  INV_X1 U5436 ( .A(n8445), .ZN(n4642) );
  NAND2_X1 U5437 ( .A1(n5426), .A2(n8294), .ZN(n5439) );
  INV_X1 U5438 ( .A(n5427), .ZN(n5426) );
  OR2_X1 U5439 ( .A1(n5305), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5316) );
  OR2_X1 U5440 ( .A1(n8377), .A2(n9905), .ZN(n8010) );
  OR2_X1 U5441 ( .A1(n8778), .A2(n8315), .ZN(n8071) );
  AOI21_X1 U5442 ( .B1(n7944), .B2(n4531), .A(n4350), .ZN(n4530) );
  INV_X1 U5443 ( .A(n7558), .ZN(n4531) );
  XNOR2_X1 U5444 ( .A(n8380), .B(n5149), .ZN(n9858) );
  AND2_X1 U5445 ( .A1(n7966), .A2(n7969), .ZN(n9859) );
  NAND2_X1 U5446 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  INV_X1 U5447 ( .A(n5712), .ZN(n7096) );
  NOR2_X1 U5448 ( .A1(n5720), .A2(n5719), .ZN(n6747) );
  INV_X1 U5449 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n4935) );
  OR2_X1 U5450 ( .A1(n4941), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4939) );
  NOR2_X1 U5451 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4890) );
  NOR2_X1 U5452 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4889) );
  AND3_X1 U5453 ( .A1(n4973), .A2(n4888), .A3(n4887), .ZN(n4891) );
  INV_X1 U5454 ( .A(n6379), .ZN(n4821) );
  NAND2_X1 U5455 ( .A1(n7332), .A2(n4803), .ZN(n4802) );
  AOI21_X1 U5456 ( .B1(n7332), .B2(n7333), .A(n4804), .ZN(n4801) );
  INV_X1 U5457 ( .A(n6335), .ZN(n4804) );
  NOR2_X1 U5458 ( .A1(n6349), .A2(n6351), .ZN(n4442) );
  NAND2_X1 U5459 ( .A1(n9103), .A2(n7840), .ZN(n4498) );
  INV_X1 U5460 ( .A(n4498), .ZN(n4493) );
  AOI21_X1 U5461 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9542), .A(n9538), .ZN(
        n9553) );
  OR2_X1 U5462 ( .A1(n6474), .A2(n9127), .ZN(n7828) );
  INV_X1 U5463 ( .A(n8963), .ZN(n7724) );
  OR2_X1 U5464 ( .A1(n6135), .A2(n9194), .ZN(n7812) );
  NOR2_X1 U5465 ( .A1(n9211), .A2(n4436), .ZN(n4435) );
  INV_X1 U5466 ( .A(n4437), .ZN(n4436) );
  OR2_X1 U5467 ( .A1(n9211), .A2(n9235), .ZN(n7809) );
  NOR2_X1 U5468 ( .A1(n9380), .A2(n9248), .ZN(n4437) );
  INV_X1 U5469 ( .A(n4676), .ZN(n4669) );
  INV_X1 U5470 ( .A(n7715), .ZN(n4668) );
  NAND2_X1 U5471 ( .A1(n7712), .A2(n9256), .ZN(n7813) );
  NOR2_X1 U5472 ( .A1(n7813), .A2(n4677), .ZN(n4676) );
  INV_X1 U5473 ( .A(n9294), .ZN(n4677) );
  OR2_X1 U5474 ( .A1(n9415), .A2(n6020), .ZN(n7690) );
  NOR2_X1 U5475 ( .A1(n6339), .A2(n9430), .ZN(n4432) );
  INV_X1 U5476 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5988) );
  INV_X1 U5477 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5905) );
  NOR2_X1 U5478 ( .A1(n4755), .A2(n7658), .ZN(n4752) );
  INV_X1 U5479 ( .A(n6966), .ZN(n4755) );
  INV_X1 U5480 ( .A(n5899), .ZN(n4754) );
  INV_X1 U5481 ( .A(n7645), .ZN(n7644) );
  NOR2_X1 U5482 ( .A1(n9154), .A2(n6136), .ZN(n6137) );
  NOR2_X1 U5483 ( .A1(n6137), .A2(n7801), .ZN(n9121) );
  INV_X1 U5484 ( .A(n8981), .ZN(n9720) );
  AND2_X1 U5485 ( .A1(n5603), .A2(n5589), .ZN(n5601) );
  AND2_X1 U5486 ( .A1(n5583), .A2(n5571), .ZN(n5581) );
  INV_X1 U5487 ( .A(n5528), .ZN(n4699) );
  INV_X1 U5488 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U5489 ( .A1(n5420), .A2(n5419), .ZN(n5435) );
  INV_X1 U5490 ( .A(SI_17_), .ZN(n5419) );
  INV_X1 U5491 ( .A(n4721), .ZN(n4718) );
  NAND2_X1 U5492 ( .A1(n5277), .A2(n4708), .ZN(n4707) );
  INV_X1 U5493 ( .A(n5293), .ZN(n4708) );
  NOR2_X1 U5494 ( .A1(n4710), .A2(n4707), .ZN(n4706) );
  OR2_X1 U5495 ( .A1(n5900), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5927) );
  NOR2_X1 U5496 ( .A1(n5877), .A2(n5876), .ZN(n5980) );
  OAI21_X1 U5497 ( .B1(n5325), .B2(n5156), .A(n4692), .ZN(n5164) );
  OAI21_X1 U5498 ( .B1(n5138), .B2(n5137), .A(n5136), .ZN(n5139) );
  NAND2_X1 U5499 ( .A1(n5138), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U5500 ( .A1(n8182), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U5501 ( .A1(n8182), .A2(n8324), .ZN(n4621) );
  OR2_X1 U5502 ( .A1(n4620), .A2(n4619), .ZN(n4616) );
  NAND2_X1 U5503 ( .A1(n5387), .A2(n5386), .ZN(n5406) );
  INV_X1 U5504 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5386) );
  INV_X1 U5505 ( .A(n5388), .ZN(n5387) );
  OR2_X1 U5506 ( .A1(n5406), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5427) );
  AND2_X1 U5507 ( .A1(n8267), .A2(n8187), .ZN(n8301) );
  INV_X1 U5508 ( .A(n4613), .ZN(n4612) );
  AOI21_X1 U5509 ( .B1(n4349), .B2(n4617), .A(n4301), .ZN(n4613) );
  NAND2_X1 U5510 ( .A1(n7490), .A2(n7489), .ZN(n7562) );
  NOR2_X1 U5511 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  NOR2_X1 U5512 ( .A1(n8158), .A2(n8605), .ZN(n8162) );
  NAND2_X1 U5513 ( .A1(n8277), .A2(n8156), .ZN(n8291) );
  NAND2_X1 U5514 ( .A1(n4611), .A2(n4610), .ZN(n4609) );
  INV_X1 U5515 ( .A(n7239), .ZN(n4611) );
  NOR2_X1 U5516 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  INV_X1 U5517 ( .A(n7956), .ZN(n7957) );
  OAI21_X1 U5518 ( .B1(n7955), .B2(n7965), .A(n8135), .ZN(n7956) );
  NAND2_X1 U5519 ( .A1(n5219), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U5520 ( .A1(n4379), .A2(n4378), .ZN(n9774) );
  NAND2_X1 U5521 ( .A1(n9771), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4378) );
  OR2_X1 U5522 ( .A1(n9771), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U5523 ( .A1(n9774), .A2(n9773), .ZN(n9772) );
  OAI21_X1 U5524 ( .B1(n5003), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4389), .ZN(
        n9781) );
  NAND2_X1 U5525 ( .A1(n4383), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U5526 ( .A1(n4959), .A2(n6673), .ZN(n6702) );
  NAND2_X1 U5527 ( .A1(n4970), .A2(n6723), .ZN(n6501) );
  NAND2_X1 U5528 ( .A1(n5010), .A2(n6527), .ZN(n6729) );
  OAI21_X1 U5529 ( .B1(n9792), .B2(n4982), .A(n6874), .ZN(n6879) );
  NAND2_X1 U5530 ( .A1(n7571), .A2(n4914), .ZN(n5721) );
  NOR2_X1 U5531 ( .A1(n5694), .A2(n5687), .ZN(n4914) );
  NOR2_X1 U5532 ( .A1(n5018), .A2(n7471), .ZN(n7416) );
  INV_X1 U5533 ( .A(n4653), .ZN(n8388) );
  NOR2_X1 U5534 ( .A1(n7420), .A2(n4990), .ZN(n4410) );
  NAND2_X1 U5535 ( .A1(n4654), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4651) );
  INV_X1 U5536 ( .A(n8410), .ZN(n4654) );
  OR2_X1 U5537 ( .A1(n8389), .A2(n10050), .ZN(n4653) );
  AND2_X1 U5538 ( .A1(n8443), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4411) );
  NOR2_X1 U5539 ( .A1(n9846), .A2(n9847), .ZN(n9845) );
  NAND2_X1 U5540 ( .A1(n4657), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4656) );
  AND2_X1 U5541 ( .A1(n5614), .A2(n5613), .ZN(n8505) );
  NAND2_X1 U5542 ( .A1(n5555), .A2(n5554), .ZN(n5574) );
  INV_X1 U5543 ( .A(n5486), .ZN(n5485) );
  NAND2_X1 U5544 ( .A1(n5458), .A2(n8253), .ZN(n5471) );
  INV_X1 U5545 ( .A(n5459), .ZN(n5458) );
  NAND2_X1 U5546 ( .A1(n8704), .A2(n8053), .ZN(n8597) );
  INV_X1 U5547 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5355) );
  INV_X1 U5548 ( .A(n5357), .ZN(n5356) );
  OR2_X1 U5549 ( .A1(n5316), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U5550 ( .A1(n5335), .A2(n7412), .ZN(n5357) );
  INV_X1 U5551 ( .A(n5336), .ZN(n5335) );
  NAND2_X1 U5552 ( .A1(n4855), .A2(n4853), .ZN(n7444) );
  AOI21_X1 U5553 ( .B1(n7943), .B2(n4856), .A(n4854), .ZN(n4853) );
  AND2_X1 U5554 ( .A1(n8008), .A2(n8020), .ZN(n4856) );
  INV_X1 U5555 ( .A(n4535), .ZN(n4534) );
  NAND2_X1 U5556 ( .A1(n5284), .A2(n5283), .ZN(n5305) );
  INV_X1 U5557 ( .A(n5285), .ZN(n5284) );
  NAND2_X1 U5558 ( .A1(n4533), .A2(n4537), .ZN(n7348) );
  NAND2_X1 U5559 ( .A1(n4539), .A2(n4538), .ZN(n4533) );
  INV_X1 U5560 ( .A(n5243), .ZN(n5242) );
  AND2_X1 U5561 ( .A1(n8010), .A2(n7311), .ZN(n8004) );
  AND3_X1 U5562 ( .A1(n5238), .A2(n5237), .A3(n5236), .ZN(n7246) );
  AOI21_X1 U5563 ( .B1(n4525), .B2(n4527), .A(n4337), .ZN(n4524) );
  INV_X1 U5564 ( .A(n4526), .ZN(n4525) );
  INV_X1 U5565 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U5566 ( .A1(n7084), .A2(n5636), .ZN(n7144) );
  NAND2_X1 U5567 ( .A1(n5635), .A2(n7933), .ZN(n7084) );
  NAND2_X1 U5568 ( .A1(n9857), .A2(n7974), .ZN(n7004) );
  INV_X1 U5569 ( .A(n8468), .ZN(n5673) );
  OR2_X1 U5570 ( .A1(n6813), .A2(n6812), .ZN(n5720) );
  INV_X1 U5571 ( .A(n8491), .ZN(n4395) );
  NAND2_X1 U5572 ( .A1(n8492), .A2(n9860), .ZN(n4393) );
  NOR2_X1 U5573 ( .A1(n8106), .A2(n7928), .ZN(n8499) );
  NAND2_X1 U5574 ( .A1(n4843), .A2(n4842), .ZN(n8511) );
  AOI21_X1 U5575 ( .B1(n4351), .B2(n4844), .A(n8088), .ZN(n4842) );
  NAND2_X1 U5576 ( .A1(n8522), .A2(n8528), .ZN(n8521) );
  AND2_X1 U5577 ( .A1(n5518), .A2(n5517), .ZN(n5663) );
  AOI21_X1 U5578 ( .B1(n4554), .B2(n4559), .A(n4552), .ZN(n4551) );
  AND2_X1 U5579 ( .A1(n4557), .A2(n4555), .ZN(n4554) );
  NAND2_X1 U5580 ( .A1(n4556), .A2(n4557), .ZN(n8568) );
  OR2_X1 U5581 ( .A1(n8589), .A2(n4559), .ZN(n4556) );
  AND2_X1 U5582 ( .A1(n8071), .A2(n8078), .ZN(n8570) );
  AND2_X1 U5583 ( .A1(n8597), .A2(n8596), .ZN(n8697) );
  OAI21_X1 U5584 ( .B1(n8645), .B2(n5394), .A(n8059), .ZN(n8628) );
  AND4_X1 U5585 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n8635)
         );
  NAND2_X1 U5586 ( .A1(n8629), .A2(n8630), .ZN(n8637) );
  AND4_X1 U5587 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n8634)
         );
  INV_X1 U5588 ( .A(n8215), .ZN(n9886) );
  OR2_X1 U5589 ( .A1(n8127), .A2(n7096), .ZN(n6749) );
  OR2_X1 U5590 ( .A1(n7401), .A2(n9926), .ZN(n9933) );
  XNOR2_X1 U5591 ( .A(n4920), .B(n4921), .ZN(n7090) );
  AND2_X1 U5592 ( .A1(n5721), .A2(n6562), .ZN(n6761) );
  AND2_X1 U5593 ( .A1(n4635), .A2(n4357), .ZN(n5091) );
  INV_X1 U5594 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U5595 ( .A(n4905), .B(n4904), .ZN(n5695) );
  INV_X1 U5596 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U5597 ( .A1(n4912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5598 ( .A1(n4902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U5599 ( .A1(n4910), .A2(n4903), .ZN(n4912) );
  INV_X1 U5600 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4903) );
  AND2_X1 U5601 ( .A1(n4944), .A2(n4893), .ZN(n4946) );
  AND2_X1 U5602 ( .A1(n4961), .A2(n4956), .ZN(n5157) );
  MUX2_X1 U5603 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4954), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n4956) );
  INV_X1 U5604 ( .A(n8840), .ZN(n4817) );
  AND2_X1 U5605 ( .A1(n8913), .A2(n6405), .ZN(n8849) );
  OAI21_X1 U5606 ( .B1(n7031), .B2(n4830), .A(n4827), .ZN(n4441) );
  INV_X1 U5607 ( .A(n4831), .ZN(n4830) );
  AND2_X1 U5608 ( .A1(n6310), .A2(n4832), .ZN(n4831) );
  NAND2_X1 U5609 ( .A1(n5737), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6048) );
  AOI21_X1 U5610 ( .B1(n4813), .B2(n4815), .A(n4811), .ZN(n4810) );
  INV_X1 U5611 ( .A(n6418), .ZN(n4811) );
  XNOR2_X1 U5612 ( .A(n6426), .B(n6427), .ZN(n8880) );
  INV_X1 U5613 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6013) );
  OR2_X1 U5614 ( .A1(n6014), .A2(n6013), .ZN(n6027) );
  INV_X1 U5615 ( .A(n4814), .ZN(n4813) );
  OAI21_X1 U5616 ( .B1(n8849), .B2(n4815), .A(n8912), .ZN(n4814) );
  INV_X1 U5617 ( .A(n8913), .ZN(n4815) );
  NAND2_X1 U5618 ( .A1(n6273), .A2(n6272), .ZN(n4825) );
  OR2_X1 U5619 ( .A1(n5796), .A2(n5783), .ZN(n5785) );
  NAND2_X1 U5620 ( .A1(n5736), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6039) );
  INV_X1 U5621 ( .A(n5785), .ZN(n5736) );
  NAND2_X1 U5622 ( .A1(n5733), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5972) );
  INV_X1 U5623 ( .A(n5960), .ZN(n5733) );
  INV_X1 U5624 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5971) );
  OR2_X1 U5625 ( .A1(n5972), .A2(n5971), .ZN(n5989) );
  INV_X1 U5626 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5944) );
  OR2_X1 U5627 ( .A1(n5945), .A2(n5944), .ZN(n5960) );
  XNOR2_X1 U5628 ( .A(n6248), .B(n6446), .ZN(n6251) );
  NAND2_X1 U5629 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  NAND2_X1 U5630 ( .A1(n5735), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6029) );
  INV_X1 U5631 ( .A(n6027), .ZN(n5735) );
  OR2_X1 U5632 ( .A1(n6029), .A2(n8936), .ZN(n5796) );
  INV_X1 U5633 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U5634 ( .A1(n6281), .A2(n6805), .ZN(n6773) );
  OR2_X1 U5635 ( .A1(n5989), .A2(n5988), .ZN(n6002) );
  NAND2_X1 U5636 ( .A1(n5734), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6014) );
  INV_X1 U5637 ( .A(n6002), .ZN(n5734) );
  NAND2_X1 U5638 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  NOR2_X1 U5639 ( .A1(n7904), .A2(n4325), .ZN(n4486) );
  INV_X1 U5640 ( .A(n6115), .ZN(n7909) );
  INV_X1 U5641 ( .A(n5837), .ZN(n5852) );
  INV_X1 U5642 ( .A(n7751), .ZN(n6099) );
  INV_X1 U5643 ( .A(n6032), .ZN(n6140) );
  AND3_X1 U5644 ( .A1(n5807), .A2(n5806), .A3(n5805), .ZN(n5810) );
  AOI21_X1 U5645 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6610), .A(n9492), .ZN(
        n9507) );
  AOI21_X1 U5646 ( .B1(n9489), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9484), .ZN(
        n9569) );
  NOR2_X1 U5647 ( .A1(n9065), .A2(n9611), .ZN(n9068) );
  AND2_X1 U5648 ( .A1(n9134), .A2(n6090), .ZN(n9163) );
  OAI21_X1 U5649 ( .B1(n9240), .B2(n4787), .A(n4785), .ZN(n4796) );
  INV_X1 U5650 ( .A(n4786), .ZN(n4785) );
  OAI21_X1 U5651 ( .B1(n4787), .B2(n4794), .A(n4797), .ZN(n4786) );
  AND2_X1 U5652 ( .A1(n7812), .A2(n7729), .ZN(n9190) );
  NAND2_X1 U5653 ( .A1(n9264), .A2(n4433), .ZN(n9192) );
  AND2_X1 U5654 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  AND2_X1 U5655 ( .A1(n6079), .A2(n6068), .ZN(n9195) );
  NOR2_X1 U5656 ( .A1(n4792), .A2(n9218), .ZN(n4789) );
  INV_X1 U5657 ( .A(n9202), .ZN(n9208) );
  NAND2_X1 U5658 ( .A1(n9264), .A2(n4435), .ZN(n9209) );
  OR2_X1 U5659 ( .A1(n6048), .A2(n6047), .ZN(n6050) );
  NAND2_X1 U5660 ( .A1(n5738), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6058) );
  INV_X1 U5661 ( .A(n6050), .ZN(n5738) );
  NAND2_X1 U5662 ( .A1(n9264), .A2(n9453), .ZN(n9245) );
  INV_X1 U5663 ( .A(n4675), .ZN(n4674) );
  OAI21_X1 U5664 ( .B1(n7813), .B2(n7878), .A(n7815), .ZN(n4675) );
  NAND2_X1 U5665 ( .A1(n9293), .A2(n4676), .ZN(n4673) );
  INV_X1 U5666 ( .A(n4672), .ZN(n4508) );
  NAND2_X1 U5667 ( .A1(n4776), .A2(n4778), .ZN(n4775) );
  NAND2_X1 U5668 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  NOR2_X1 U5669 ( .A1(n9399), .A2(n9302), .ZN(n9287) );
  AOI21_X1 U5670 ( .B1(n4663), .B2(n4665), .A(n4661), .ZN(n4660) );
  INV_X1 U5671 ( .A(n7697), .ZN(n4661) );
  AND2_X1 U5672 ( .A1(n7305), .A2(n4303), .ZN(n9336) );
  NAND2_X1 U5673 ( .A1(n7305), .A2(n4430), .ZN(n9337) );
  INV_X1 U5674 ( .A(n4681), .ZN(n4679) );
  AOI21_X1 U5675 ( .B1(n4683), .B2(n4682), .A(n7691), .ZN(n4681) );
  INV_X1 U5676 ( .A(n7791), .ZN(n7432) );
  INV_X1 U5677 ( .A(n4765), .ZN(n4764) );
  NOR2_X1 U5678 ( .A1(n4766), .A2(n4770), .ZN(n4763) );
  NAND2_X1 U5679 ( .A1(n7305), .A2(n4772), .ZN(n9426) );
  NAND2_X1 U5680 ( .A1(n4768), .A2(n4767), .ZN(n9421) );
  NAND2_X1 U5681 ( .A1(n7268), .A2(n4769), .ZN(n4768) );
  AOI21_X1 U5682 ( .B1(n4691), .B2(n4750), .A(n4339), .ZN(n4749) );
  INV_X1 U5683 ( .A(n5923), .ZN(n4750) );
  AND2_X1 U5684 ( .A1(n7017), .A2(n9727), .ZN(n7125) );
  NOR2_X1 U5685 ( .A1(n6909), .A2(n6852), .ZN(n7019) );
  INV_X1 U5686 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5892) );
  OR2_X1 U5687 ( .A1(n5893), .A2(n5892), .ZN(n5906) );
  AOI21_X1 U5688 ( .B1(n6907), .B2(n6906), .A(n6123), .ZN(n6961) );
  AND2_X1 U5689 ( .A1(n6146), .A2(n8995), .ZN(n9343) );
  OR2_X1 U5690 ( .A1(n9709), .A2(n6267), .ZN(n9710) );
  INV_X1 U5691 ( .A(n8982), .ZN(n6941) );
  AND2_X1 U5692 ( .A1(n7041), .A2(n6118), .ZN(n9662) );
  NAND2_X1 U5693 ( .A1(n7041), .A2(n4678), .ZN(n7047) );
  OR2_X1 U5694 ( .A1(n6117), .A2(n7042), .ZN(n4678) );
  NOR2_X1 U5695 ( .A1(n7053), .A2(n9686), .ZN(n9671) );
  AND2_X1 U5696 ( .A1(n7742), .A2(n9416), .ZN(n4688) );
  AND2_X1 U5697 ( .A1(n9133), .A2(n9132), .ZN(n9357) );
  INV_X1 U5698 ( .A(n9740), .ZN(n9711) );
  INV_X1 U5699 ( .A(n5844), .ZN(n6023) );
  INV_X1 U5700 ( .A(n6548), .ZN(n6022) );
  NAND2_X1 U5701 ( .A1(n4685), .A2(n4683), .ZN(n9424) );
  NAND2_X1 U5702 ( .A1(n4685), .A2(n7685), .ZN(n9423) );
  OR2_X1 U5703 ( .A1(n5872), .A2(n5871), .ZN(n6952) );
  NOR2_X1 U5704 ( .A1(n6183), .A2(n6841), .ZN(n6185) );
  INV_X1 U5705 ( .A(n9750), .ZN(n9683) );
  NOR2_X1 U5706 ( .A1(n6161), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U5707 ( .A1(n6174), .A2(n6156), .ZN(n6157) );
  INV_X1 U5708 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U5709 ( .A1(n6158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6175) );
  AND2_X1 U5710 ( .A1(n4870), .A2(n6113), .ZN(n4839) );
  INV_X1 U5711 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4460) );
  INV_X1 U5712 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6113) );
  XNOR2_X1 U5713 ( .A(n5480), .B(n5468), .ZN(n7281) );
  INV_X1 U5714 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U5715 ( .A1(n5366), .A2(n5365), .ZN(n5381) );
  AND2_X1 U5716 ( .A1(n5967), .A2(n5956), .ZN(n9060) );
  NAND2_X1 U5717 ( .A1(n5312), .A2(n5311), .ZN(n5324) );
  OAI21_X1 U5718 ( .B1(n5257), .B2(n4702), .A(n4701), .ZN(n5295) );
  INV_X1 U5719 ( .A(n4711), .ZN(n4702) );
  AOI21_X1 U5720 ( .B1(n4711), .B2(n4710), .A(n4709), .ZN(n4701) );
  AND2_X1 U5721 ( .A1(n5269), .A2(n5255), .ZN(n5256) );
  AND2_X1 U5722 ( .A1(n5250), .A2(n5232), .ZN(n5233) );
  AND2_X1 U5723 ( .A1(n5228), .A2(n5213), .ZN(n5214) );
  NAND2_X1 U5724 ( .A1(n5185), .A2(n5184), .ZN(n5193) );
  NAND2_X1 U5725 ( .A1(n5138), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5108) );
  AND2_X1 U5726 ( .A1(n4604), .A2(n4606), .ZN(n7259) );
  OR2_X1 U5727 ( .A1(n8343), .A2(n8504), .ZN(n4631) );
  AND2_X1 U5728 ( .A1(n8343), .A2(n8504), .ZN(n4632) );
  AND2_X1 U5729 ( .A1(n5543), .A2(n5542), .ZN(n8246) );
  INV_X1 U5730 ( .A(n4600), .ZN(n4599) );
  AND2_X1 U5731 ( .A1(n7140), .A2(n5630), .ZN(n8368) );
  XOR2_X1 U5732 ( .A(n4291), .B(n8491), .Z(n8227) );
  AND2_X1 U5733 ( .A1(n5272), .A2(n5271), .ZN(n9910) );
  AND3_X1 U5734 ( .A1(n5477), .A2(n5476), .A3(n5475), .ZN(n8590) );
  AND2_X1 U5735 ( .A1(n4616), .A2(n4614), .ZN(n7587) );
  NAND2_X1 U5736 ( .A1(n4616), .A2(n4617), .ZN(n7565) );
  AND2_X1 U5737 ( .A1(n5525), .A2(n5524), .ZN(n8328) );
  AND2_X1 U5738 ( .A1(n7110), .A2(n7109), .ZN(n8358) );
  AND2_X1 U5739 ( .A1(n6758), .A2(n6757), .ZN(n8352) );
  NAND2_X1 U5740 ( .A1(n6762), .A2(n8607), .ZN(n8350) );
  INV_X1 U5741 ( .A(n8352), .ZN(n8354) );
  OR2_X1 U5742 ( .A1(n7091), .A2(n7479), .ZN(n8362) );
  AND2_X1 U5743 ( .A1(n7140), .A2(n7139), .ZN(n8474) );
  INV_X1 U5744 ( .A(n8505), .ZN(n8369) );
  NAND2_X1 U5745 ( .A1(n5600), .A2(n5599), .ZN(n8514) );
  INV_X1 U5746 ( .A(n8246), .ZN(n8549) );
  INV_X1 U5747 ( .A(n8180), .ZN(n8573) );
  INV_X1 U5748 ( .A(n8634), .ZN(n8370) );
  OR2_X1 U5749 ( .A1(n5175), .A2(n6642), .ZN(n5100) );
  OR2_X1 U5750 ( .A1(n4284), .A2(n5115), .ZN(n5119) );
  OR2_X1 U5751 ( .A1(n5721), .A2(n6754), .ZN(n8381) );
  NAND2_X1 U5752 ( .A1(n4573), .A2(n4951), .ZN(n6643) );
  NAND2_X1 U5753 ( .A1(n4589), .A2(n4590), .ZN(n6727) );
  INV_X1 U5754 ( .A(n4565), .ZN(n4986) );
  NOR2_X1 U5755 ( .A1(n4989), .A2(n7463), .ZN(n7411) );
  NOR2_X1 U5756 ( .A1(n8426), .A2(n4994), .ZN(n8436) );
  INV_X1 U5757 ( .A(n4388), .ZN(n4993) );
  INV_X1 U5758 ( .A(n5022), .ZN(n4640) );
  NAND2_X1 U5759 ( .A1(n5607), .A2(n5606), .ZN(n8495) );
  NAND2_X1 U5760 ( .A1(n5591), .A2(n5590), .ZN(n8672) );
  AND2_X1 U5761 ( .A1(n5534), .A2(n5533), .ZN(n8533) );
  NAND2_X1 U5762 ( .A1(n5437), .A2(n5436), .ZN(n8702) );
  NOR2_X1 U5763 ( .A1(n8040), .A2(n8037), .ZN(n4862) );
  OR2_X1 U5764 ( .A1(n9928), .A2(n9873), .ZN(n8532) );
  NAND2_X1 U5765 ( .A1(n7347), .A2(n8008), .ZN(n7398) );
  NAND2_X1 U5766 ( .A1(n4539), .A2(n4883), .ZN(n7314) );
  OAI211_X1 U5767 ( .C1(n5206), .C2(n4417), .A(n5260), .B(n5259), .ZN(n7257)
         );
  INV_X1 U5768 ( .A(n5638), .ZN(n9895) );
  INV_X1 U5769 ( .A(n9877), .ZN(n8607) );
  NAND2_X1 U5770 ( .A1(n9878), .A2(n6895), .ZN(n8661) );
  NAND2_X1 U5771 ( .A1(n5685), .A2(n8827), .ZN(n4594) );
  NAND2_X1 U5772 ( .A1(n5127), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4595) );
  INV_X1 U5773 ( .A(n9928), .ZN(n9920) );
  AND2_X1 U5774 ( .A1(n6761), .A2(n6760), .ZN(n9877) );
  NAND2_X1 U5775 ( .A1(n7917), .A2(n7916), .ZN(n8727) );
  NAND2_X1 U5776 ( .A1(n7913), .A2(n7912), .ZN(n8731) );
  INV_X1 U5777 ( .A(n8495), .ZN(n8741) );
  AOI21_X1 U5778 ( .B1(n4394), .B2(n9866), .A(n4391), .ZN(n8735) );
  NAND2_X1 U5779 ( .A1(n4393), .A2(n4392), .ZN(n4391) );
  XNOR2_X1 U5780 ( .A(n8490), .B(n4395), .ZN(n4394) );
  NAND2_X1 U5781 ( .A1(n8514), .A2(n9862), .ZN(n4392) );
  NAND2_X1 U5782 ( .A1(n5573), .A2(n5572), .ZN(n8748) );
  NAND2_X1 U5783 ( .A1(n5553), .A2(n5552), .ZN(n8754) );
  NAND2_X1 U5784 ( .A1(n4841), .A2(n4844), .ZN(n8529) );
  OR2_X1 U5785 ( .A1(n8555), .A2(n4847), .ZN(n4841) );
  INV_X1 U5786 ( .A(n8533), .ZN(n8760) );
  AND2_X1 U5787 ( .A1(n4852), .A2(n4850), .ZN(n8541) );
  INV_X1 U5788 ( .A(n5663), .ZN(n8766) );
  NAND2_X1 U5789 ( .A1(n4852), .A2(n5662), .ZN(n8546) );
  AND2_X1 U5790 ( .A1(n4562), .A2(n4313), .ZN(n8583) );
  OR2_X1 U5791 ( .A1(n8704), .A2(n5661), .ZN(n4857) );
  NAND2_X1 U5792 ( .A1(n5425), .A2(n5424), .ZN(n8793) );
  NAND2_X1 U5793 ( .A1(n5405), .A2(n5404), .ZN(n8799) );
  NAND2_X1 U5794 ( .A1(n5385), .A2(n5384), .ZN(n8805) );
  NAND2_X1 U5795 ( .A1(n5653), .A2(n5652), .ZN(n8651) );
  NAND2_X1 U5796 ( .A1(n5354), .A2(n5353), .ZN(n7589) );
  NOR2_X1 U5797 ( .A1(n9936), .A2(n9911), .ZN(n8807) );
  NAND2_X1 U5798 ( .A1(n7441), .A2(n7944), .ZN(n7514) );
  INV_X1 U5799 ( .A(n8740), .ZN(n8806) );
  AND2_X1 U5800 ( .A1(n7090), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6562) );
  INV_X1 U5801 ( .A(n5095), .ZN(n8819) );
  AND2_X1 U5802 ( .A1(n4909), .A2(n4925), .ZN(n7603) );
  INV_X1 U5803 ( .A(n5695), .ZN(n7571) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7452) );
  INV_X1 U5805 ( .A(n8144), .ZN(n7451) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7344) );
  XNOR2_X1 U5807 ( .A(n5084), .B(n5083), .ZN(n7283) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7253) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7162) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10035) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6893) );
  INV_X1 U5812 ( .A(n5403), .ZN(n8443) );
  INV_X1 U5813 ( .A(n5368), .ZN(n8408) );
  AND2_X1 U5814 ( .A1(n6514), .A2(P2_U3151), .ZN(n8823) );
  INV_X1 U5815 ( .A(n6882), .ZN(n6544) );
  NAND2_X1 U5816 ( .A1(n4977), .A2(n4980), .ZN(n6531) );
  INV_X1 U5817 ( .A(n5207), .ZN(n6527) );
  INV_X1 U5818 ( .A(n5157), .ZN(n6695) );
  AND2_X1 U5819 ( .A1(n6178), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6496) );
  NAND2_X1 U5820 ( .A1(n4818), .A2(n4816), .ZN(n8839) );
  XNOR2_X1 U5821 ( .A(n6260), .B(n6261), .ZN(n6714) );
  AOI21_X1 U5822 ( .B1(n4451), .B2(n4309), .A(n4448), .ZN(n4447) );
  INV_X1 U5823 ( .A(n8870), .ZN(n4448) );
  OAI21_X1 U5824 ( .B1(n8898), .B2(n4309), .A(n4451), .ZN(n8869) );
  NAND2_X1 U5825 ( .A1(n4806), .A2(n4808), .ZN(n4805) );
  INV_X1 U5826 ( .A(n4809), .ZN(n4808) );
  NAND2_X1 U5827 ( .A1(n4807), .A2(n4803), .ZN(n4806) );
  NAND2_X1 U5828 ( .A1(n4826), .A2(n6263), .ZN(n6804) );
  NAND2_X1 U5829 ( .A1(n4825), .A2(n6277), .ZN(n6807) );
  NAND2_X1 U5830 ( .A1(n4824), .A2(n4823), .ZN(n8916) );
  AND2_X1 U5831 ( .A1(n4824), .A2(n4322), .ZN(n8915) );
  NAND2_X1 U5832 ( .A1(n8861), .A2(n6379), .ZN(n4824) );
  AOI21_X1 U5833 ( .B1(n7286), .B2(n7284), .A(n7285), .ZN(n7334) );
  NAND2_X1 U5834 ( .A1(n8898), .A2(n8902), .ZN(n8935) );
  INV_X1 U5835 ( .A(n8943), .ZN(n9528) );
  AND3_X1 U5836 ( .A1(n5815), .A2(n5814), .A3(n5813), .ZN(n4886) );
  NAND2_X1 U5837 ( .A1(n9011), .A2(n9012), .ZN(n9010) );
  AOI21_X1 U5838 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9075), .A(n9073), .ZN(
        n9084) );
  OR2_X1 U5839 ( .A1(n9622), .A2(n9621), .ZN(n9631) );
  OR2_X1 U5840 ( .A1(n9145), .A2(n9127), .ZN(n4873) );
  AND2_X1 U5841 ( .A1(n4742), .A2(n4745), .ZN(n9158) );
  NAND2_X1 U5842 ( .A1(n4790), .A2(n4788), .ZN(n9222) );
  AOI21_X1 U5843 ( .B1(n9240), .B2(n6054), .A(n4791), .ZN(n9220) );
  NAND2_X1 U5844 ( .A1(n4774), .A2(n4778), .ZN(n9286) );
  NAND2_X1 U5845 ( .A1(n4773), .A2(n4779), .ZN(n4774) );
  NAND2_X1 U5846 ( .A1(n4780), .A2(n4783), .ZN(n9301) );
  NAND2_X1 U5847 ( .A1(n4773), .A2(n4310), .ZN(n4780) );
  NAND2_X1 U5848 ( .A1(n4662), .A2(n7868), .ZN(n9316) );
  AOI21_X1 U5849 ( .B1(n7266), .B2(n7267), .A(n4293), .ZN(n7304) );
  NAND2_X1 U5850 ( .A1(n7118), .A2(n4691), .ZN(n7117) );
  NAND2_X1 U5851 ( .A1(n6989), .A2(n5923), .ZN(n7118) );
  NAND2_X1 U5852 ( .A1(n6967), .A2(n6966), .ZN(n6965) );
  NAND2_X1 U5853 ( .A1(n7010), .A2(n5899), .ZN(n6967) );
  NAND2_X1 U5854 ( .A1(n6972), .A2(n6848), .ZN(n10150) );
  OR2_X1 U5855 ( .A1(n9677), .A2(n9103), .ZN(n9655) );
  NOR2_X1 U5856 ( .A1(n6223), .A2(n6222), .ZN(n9537) );
  NAND2_X1 U5857 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  NAND2_X1 U5858 ( .A1(n9109), .A2(n9416), .ZN(n6221) );
  INV_X1 U5859 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4399) );
  INV_X1 U5860 ( .A(n9265), .ZN(n9457) );
  INV_X1 U5861 ( .A(n9325), .ZN(n9466) );
  INV_X1 U5862 ( .A(n9430), .ZN(n9642) );
  INV_X1 U5863 ( .A(n9651), .ZN(n7025) );
  NAND2_X1 U5864 ( .A1(n9753), .A2(n9416), .ZN(n9469) );
  INV_X1 U5865 ( .A(n9678), .ZN(n9679) );
  INV_X1 U5866 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5757) );
  OR2_X1 U5867 ( .A1(n5756), .A2(n9473), .ZN(n5758) );
  NAND2_X1 U5868 ( .A1(n5755), .A2(n9474), .ZN(n7630) );
  MUX2_X1 U5869 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5753), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5755) );
  NAND2_X1 U5870 ( .A1(n5767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5768) );
  CLKBUF_X1 U5871 ( .A(n6217), .Z(n8994) );
  XNOR2_X1 U5872 ( .A(n6155), .B(n6154), .ZN(n7601) );
  INV_X1 U5873 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7486) );
  XNOR2_X1 U5874 ( .A(n5527), .B(n5526), .ZN(n7483) );
  INV_X1 U5875 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7387) );
  INV_X1 U5876 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10016) );
  INV_X1 U5877 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7254) );
  INV_X1 U5878 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7165) );
  INV_X1 U5879 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10111) );
  XNOR2_X1 U5880 ( .A(n5968), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U5881 ( .A1(n4730), .A2(n4729), .ZN(n5344) );
  OR2_X1 U5882 ( .A1(n5300), .A2(n5301), .ZN(n5302) );
  INV_X1 U5883 ( .A(n5169), .ZN(n5166) );
  OR2_X1 U5884 ( .A1(n8146), .A2(n8145), .ZN(n4387) );
  INV_X1 U5885 ( .A(n4581), .ZN(n8401) );
  INV_X1 U5886 ( .A(n4641), .ZN(n8417) );
  INV_X1 U5887 ( .A(n4569), .ZN(n5001) );
  NAND2_X1 U5888 ( .A1(n4567), .A2(n8452), .ZN(n4566) );
  NAND2_X1 U5889 ( .A1(n4840), .A2(n9878), .ZN(n8486) );
  OAI22_X1 U5890 ( .A1(n8482), .A2(n8670), .B1(n9954), .B2(n10127), .ZN(n5716)
         );
  NOR2_X1 U5891 ( .A1(n5728), .A2(n5730), .ZN(n5731) );
  NOR2_X1 U5892 ( .A1(n9934), .A2(n5729), .ZN(n5730) );
  NOR2_X1 U5893 ( .A1(n8482), .A2(n8740), .ZN(n5728) );
  AND2_X1 U5894 ( .A1(n6458), .A2(n9531), .ZN(n6478) );
  NAND2_X1 U5895 ( .A1(n4457), .A2(n4456), .ZN(P1_U3229) );
  AOI21_X1 U5896 ( .B1(n8943), .B2(n9211), .A(n8914), .ZN(n4456) );
  NAND2_X1 U5897 ( .A1(n4458), .A2(n9531), .ZN(n4457) );
  NOR2_X1 U5898 ( .A1(n6484), .A2(n6483), .ZN(n6494) );
  INV_X1 U5899 ( .A(n4479), .ZN(n4420) );
  NAND2_X1 U5900 ( .A1(n4482), .A2(n4483), .ZN(n4418) );
  OR2_X1 U5901 ( .A1(n4481), .A2(n7903), .ZN(n4419) );
  MUX2_X1 U5902 ( .A(n9105), .B(n9104), .S(n9103), .Z(n9107) );
  NAND2_X1 U5903 ( .A1(n4426), .A2(n4425), .ZN(P1_U3551) );
  NAND2_X1 U5904 ( .A1(n9768), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4425) );
  OAI21_X1 U5905 ( .B1(n6186), .B2(n9768), .A(n4396), .ZN(n6187) );
  NAND2_X1 U5906 ( .A1(n9768), .A2(n6098), .ZN(n4396) );
  NOR2_X1 U5907 ( .A1(n4368), .A2(n4398), .ZN(n4397) );
  INV_X2 U5908 ( .A(n5206), .ZN(n7915) );
  NOR2_X1 U5909 ( .A1(n4627), .A2(n8302), .ZN(n4294) );
  OR2_X1 U5910 ( .A1(n9405), .A2(n9295), .ZN(n4295) );
  XNOR2_X1 U5911 ( .A(n6175), .B(n6174), .ZN(n6115) );
  NAND2_X1 U5912 ( .A1(n4500), .A2(n4499), .ZN(n5769) );
  INV_X1 U5913 ( .A(n7285), .ZN(n4803) );
  INV_X1 U5914 ( .A(n5661), .ZN(n8596) );
  XNOR2_X1 U5915 ( .A(n4978), .B(P2_IR_REG_7__SCAN_IN), .ZN(n5249) );
  INV_X1 U5916 ( .A(n5249), .ZN(n4587) );
  NAND2_X1 U5917 ( .A1(n6374), .A2(n6373), .ZN(n4297) );
  AND4_X1 U5918 ( .A1(n4544), .A2(n4899), .A3(n4896), .A4(n4898), .ZN(n4298)
         );
  NAND2_X1 U5919 ( .A1(n4621), .A2(n8183), .ZN(n8300) );
  OR2_X1 U5920 ( .A1(n5642), .A2(n7938), .ZN(n4299) );
  AND2_X1 U5921 ( .A1(n5774), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U5922 ( .A1(n4866), .A2(n4900), .ZN(n5085) );
  AND2_X1 U5923 ( .A1(n7588), .A2(n8372), .ZN(n4301) );
  OR2_X1 U5924 ( .A1(n4636), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4302) );
  AND2_X1 U5925 ( .A1(n4430), .A2(n4429), .ZN(n4303) );
  AND2_X1 U5926 ( .A1(n5449), .A2(SI_18_), .ZN(n4304) );
  INV_X1 U5927 ( .A(n6339), .ZN(n4772) );
  NOR2_X1 U5928 ( .A1(n7610), .A2(n7611), .ZN(n4305) );
  NAND2_X1 U5929 ( .A1(n7097), .A2(n7096), .ZN(n7100) );
  INV_X1 U5930 ( .A(n7100), .ZN(n8184) );
  AND2_X1 U5931 ( .A1(n4592), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U5932 ( .A1(n5096), .A2(n5095), .ZN(n5150) );
  INV_X1 U5933 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4973) );
  OAI21_X1 U5934 ( .B1(n6406), .B2(n4815), .A(n4813), .ZN(n8911) );
  AND2_X1 U5935 ( .A1(n4297), .A2(n8902), .ZN(n4307) );
  INV_X1 U5936 ( .A(n5666), .ZN(n8097) );
  OR2_X1 U5937 ( .A1(n8754), .A2(n5631), .ZN(n5666) );
  NAND2_X1 U5938 ( .A1(n5470), .A2(n5469), .ZN(n8784) );
  AND2_X1 U5939 ( .A1(n7660), .A2(n7760), .ZN(n4308) );
  OR2_X1 U5940 ( .A1(n4822), .A2(n4454), .ZN(n4309) );
  NAND2_X1 U5941 ( .A1(n5804), .A2(n5803), .ZN(n9405) );
  OR2_X1 U5942 ( .A1(n9325), .A2(n9346), .ZN(n4310) );
  NAND2_X1 U5943 ( .A1(n7560), .A2(n7559), .ZN(n4311) );
  AND2_X1 U5944 ( .A1(n9292), .A2(n7878), .ZN(n4312) );
  XNOR2_X1 U5945 ( .A(n5089), .B(n5088), .ZN(n5096) );
  OR2_X1 U5946 ( .A1(n9861), .A2(n8215), .ZN(n7991) );
  NAND2_X1 U5947 ( .A1(n8695), .A2(n8604), .ZN(n4313) );
  NAND2_X1 U5948 ( .A1(n4912), .A2(n4913), .ZN(n5687) );
  AND2_X1 U5949 ( .A1(n4308), .A2(n7662), .ZN(n4314) );
  OR2_X1 U5950 ( .A1(n5423), .A2(n4997), .ZN(n4315) );
  INV_X1 U5951 ( .A(n8023), .ZN(n4854) );
  AND2_X1 U5952 ( .A1(n4790), .A2(n4789), .ZN(n4316) );
  AND2_X1 U5953 ( .A1(n4674), .A2(n4673), .ZN(n4317) );
  NAND2_X1 U5954 ( .A1(n5943), .A2(n5942), .ZN(n7233) );
  AND2_X1 U5955 ( .A1(n8480), .A2(n7401), .ZN(n4318) );
  AND2_X1 U5956 ( .A1(n8933), .A2(n8932), .ZN(n4319) );
  AND2_X1 U5957 ( .A1(n7198), .A2(n6312), .ZN(n4320) );
  NAND2_X1 U5958 ( .A1(n4917), .A2(n4633), .ZN(n4925) );
  OR2_X1 U5959 ( .A1(n9162), .A2(n8962), .ZN(n4321) );
  NAND2_X1 U5960 ( .A1(n7633), .A2(n7715), .ZN(n9241) );
  NAND2_X1 U5961 ( .A1(n8848), .A2(n4834), .ZN(n8924) );
  OR2_X1 U5962 ( .A1(n8858), .A2(n8859), .ZN(n4322) );
  NAND2_X1 U5963 ( .A1(n6000), .A2(n5999), .ZN(n7460) );
  OR2_X1 U5964 ( .A1(n8465), .A2(n9826), .ZN(n4323) );
  OR2_X1 U5965 ( .A1(n8784), .A2(n8590), .ZN(n8072) );
  NOR2_X1 U5966 ( .A1(n9422), .A2(n4684), .ZN(n4683) );
  AND2_X1 U5967 ( .A1(n7853), .A2(n7665), .ZN(n7785) );
  AND2_X1 U5968 ( .A1(n5365), .A2(n4722), .ZN(n4324) );
  INV_X1 U5969 ( .A(n9211), .ZN(n9448) );
  NAND2_X1 U5970 ( .A1(n6056), .A2(n6055), .ZN(n9211) );
  AND2_X1 U5971 ( .A1(n7898), .A2(n7897), .ZN(n4325) );
  NOR2_X1 U5972 ( .A1(n4721), .A2(n4719), .ZN(n4326) );
  NOR2_X1 U5973 ( .A1(n5650), .A2(n7575), .ZN(n4327) );
  AND2_X1 U5974 ( .A1(n7256), .A2(n8378), .ZN(n4328) );
  INV_X1 U5975 ( .A(n4878), .ZN(n4588) );
  NAND2_X1 U5976 ( .A1(n9264), .A2(n4437), .ZN(n4438) );
  AND2_X1 U5977 ( .A1(n4306), .A2(n4587), .ZN(n4329) );
  AOI21_X1 U5978 ( .B1(n7659), .B2(n7658), .A(n4308), .ZN(n4475) );
  NOR2_X1 U5979 ( .A1(n6522), .A2(n6514), .ZN(n4330) );
  NAND2_X1 U5980 ( .A1(n7313), .A2(n5641), .ZN(n4331) );
  OR2_X1 U5981 ( .A1(n4816), .A2(n4445), .ZN(n4332) );
  AND2_X1 U5982 ( .A1(n4923), .A2(n4869), .ZN(n4333) );
  INV_X1 U5983 ( .A(n4490), .ZN(n4489) );
  NAND2_X1 U5984 ( .A1(n4497), .A2(n4491), .ZN(n4490) );
  AND2_X1 U5985 ( .A1(n4653), .A2(n4652), .ZN(n4334) );
  AND2_X1 U5986 ( .A1(n4641), .A2(n4640), .ZN(n4335) );
  AND2_X1 U5987 ( .A1(n4901), .A2(n4634), .ZN(n4336) );
  NOR2_X1 U5988 ( .A1(n8379), .A2(n5638), .ZN(n4337) );
  AND2_X1 U5989 ( .A1(n6127), .A2(n6963), .ZN(n7658) );
  INV_X1 U5990 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4422) );
  INV_X1 U5991 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4634) );
  INV_X1 U5992 ( .A(n4770), .ZN(n4769) );
  OAI21_X1 U5993 ( .B1(n4293), .B2(n7267), .A(n7298), .ZN(n4770) );
  INV_X1 U5994 ( .A(n4732), .ZN(n4731) );
  NOR2_X1 U5995 ( .A1(n5322), .A2(SI_11_), .ZN(n4732) );
  NAND2_X1 U5996 ( .A1(n4446), .A2(n4445), .ZN(n4338) );
  AND2_X1 U5997 ( .A1(n8048), .A2(n8059), .ZN(n8652) );
  NOR2_X1 U5998 ( .A1(n7158), .A2(n8974), .ZN(n4339) );
  NOR2_X1 U5999 ( .A1(n7178), .A2(n8976), .ZN(n4340) );
  NAND2_X1 U6000 ( .A1(n9448), .A2(n9235), .ZN(n4341) );
  AND2_X1 U6001 ( .A1(n6348), .A2(n4817), .ZN(n4342) );
  AND2_X1 U6002 ( .A1(n5648), .A2(n7563), .ZN(n4343) );
  INV_X1 U6003 ( .A(n4784), .ZN(n4783) );
  NOR2_X1 U6004 ( .A1(n9466), .A2(n8937), .ZN(n4784) );
  OR2_X1 U6005 ( .A1(n4782), .A2(n4784), .ZN(n4344) );
  AND2_X1 U6006 ( .A1(n7640), .A2(n7685), .ZN(n7790) );
  AND2_X1 U6007 ( .A1(n4549), .A2(n4547), .ZN(n4917) );
  OR2_X1 U6008 ( .A1(n4998), .A2(n4867), .ZN(n4345) );
  OR2_X1 U6009 ( .A1(n6822), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4346) );
  INV_X1 U6010 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6154) );
  OR2_X1 U6011 ( .A1(n9122), .A2(n7745), .ZN(n4347) );
  INV_X1 U6012 ( .A(n6351), .ZN(n4445) );
  INV_X1 U6013 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U6014 ( .A1(n5127), .A2(n9771), .ZN(n4348) );
  AND2_X1 U6015 ( .A1(n4619), .A2(n4615), .ZN(n4349) );
  NAND2_X1 U6016 ( .A1(n4885), .A2(n7513), .ZN(n4350) );
  AND2_X1 U6017 ( .A1(n4847), .A2(n5666), .ZN(n4351) );
  NAND2_X1 U6018 ( .A1(n7332), .A2(n4803), .ZN(n4352) );
  NAND2_X1 U6019 ( .A1(n4858), .A2(n8073), .ZN(n4353) );
  AND2_X1 U6020 ( .A1(n4772), .A2(n5978), .ZN(n4354) );
  INV_X1 U6021 ( .A(n5277), .ZN(n4709) );
  INV_X1 U6022 ( .A(n4561), .ZN(n4560) );
  NAND2_X1 U6023 ( .A1(n8582), .A2(n4313), .ZN(n4561) );
  AND2_X1 U6024 ( .A1(n8480), .A2(n9926), .ZN(n4355) );
  AND2_X1 U6025 ( .A1(n4844), .A2(n5666), .ZN(n4356) );
  AND3_X1 U6026 ( .A1(n4923), .A2(n4869), .A3(n4924), .ZN(n4357) );
  AND3_X1 U6027 ( .A1(n4825), .A2(n6277), .A3(n6263), .ZN(n4358) );
  AND2_X1 U6028 ( .A1(n9922), .A2(n8374), .ZN(n8007) );
  AND2_X1 U6029 ( .A1(n6531), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4359) );
  AND2_X1 U6030 ( .A1(n5663), .A2(n8560), .ZN(n8092) );
  INV_X1 U6031 ( .A(n8092), .ZN(n4851) );
  AND2_X1 U6032 ( .A1(n7658), .A2(n7662), .ZN(n4360) );
  AND2_X1 U6033 ( .A1(n4689), .A2(n9126), .ZN(n4361) );
  INV_X1 U6034 ( .A(n7713), .ZN(n4512) );
  AND2_X1 U6035 ( .A1(n4590), .A2(n4588), .ZN(n4362) );
  INV_X1 U6036 ( .A(n4537), .ZN(n4536) );
  NAND2_X1 U6037 ( .A1(n4299), .A2(n4331), .ZN(n4537) );
  OR2_X1 U6038 ( .A1(n4513), .A2(n4505), .ZN(n4363) );
  INV_X1 U6039 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6110) );
  INV_X1 U6040 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U6041 ( .A1(n6115), .A2(n9103), .ZN(n7760) );
  INV_X1 U6042 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U6043 ( .A1(n6066), .A2(n6065), .ZN(n9194) );
  INV_X1 U6044 ( .A(n9194), .ZN(n4434) );
  NAND2_X1 U6045 ( .A1(n5979), .A2(n4761), .ZN(n5997) );
  XNOR2_X1 U6046 ( .A(n6192), .B(SI_29_), .ZN(n7628) );
  NOR2_X1 U6047 ( .A1(n5844), .A2(n7453), .ZN(n4364) );
  NAND2_X1 U6048 ( .A1(n8291), .A2(n8163), .ZN(n8332) );
  AND2_X1 U6049 ( .A1(n4857), .A2(n4860), .ZN(n4365) );
  INV_X1 U6050 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U6051 ( .A1(n7305), .A2(n4432), .ZN(n4366) );
  OR2_X1 U6052 ( .A1(n4947), .A2(n4946), .ZN(n6568) );
  INV_X1 U6053 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4893) );
  INV_X1 U6054 ( .A(n5631), .ZN(n8535) );
  AND2_X1 U6055 ( .A1(n4805), .A2(n7332), .ZN(n4367) );
  NOR2_X1 U6056 ( .A1(n9145), .A2(n9469), .ZN(n4368) );
  AND2_X1 U6057 ( .A1(n6417), .A2(n8913), .ZN(n4369) );
  NAND2_X1 U6058 ( .A1(n8291), .A2(n8290), .ZN(n4370) );
  INV_X1 U6059 ( .A(n5478), .ZN(n4739) );
  INV_X1 U6060 ( .A(n5526), .ZN(n4700) );
  AND2_X1 U6061 ( .A1(n5528), .A2(n5516), .ZN(n5526) );
  NAND2_X1 U6062 ( .A1(n6012), .A2(n6011), .ZN(n9415) );
  INV_X1 U6063 ( .A(n9415), .ZN(n4429) );
  NOR2_X1 U6064 ( .A1(n5844), .A2(n7626), .ZN(n4371) );
  OAI21_X1 U6065 ( .B1(n9708), .B2(n5861), .A(n5860), .ZN(n6905) );
  NAND2_X1 U6066 ( .A1(n5689), .A2(n7603), .ZN(n5693) );
  NAND2_X1 U6067 ( .A1(n4549), .A2(n4548), .ZN(n4998) );
  NAND2_X1 U6068 ( .A1(n4863), .A2(n8036), .ZN(n7582) );
  INV_X1 U6069 ( .A(SI_15_), .ZN(n4719) );
  NAND2_X1 U6070 ( .A1(n4381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4920) );
  AND2_X1 U6071 ( .A1(n4608), .A2(n4296), .ZN(n4372) );
  AND2_X1 U6072 ( .A1(n8408), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4373) );
  INV_X1 U6073 ( .A(n4606), .ZN(n4605) );
  AOI21_X1 U6074 ( .B1(n4296), .B2(n7240), .A(n4328), .ZN(n4606) );
  AND2_X1 U6075 ( .A1(n6462), .A2(n6453), .ZN(n9531) );
  AND2_X2 U6076 ( .A1(n6185), .A2(n6464), .ZN(n9770) );
  INV_X1 U6077 ( .A(n9665), .ZN(n9719) );
  OR2_X1 U6078 ( .A1(n7768), .A2(n7899), .ZN(n9665) );
  INV_X1 U6079 ( .A(n7900), .ZN(n9103) );
  AND2_X1 U6080 ( .A1(n5722), .A2(n5672), .ZN(n8650) );
  NAND2_X1 U6081 ( .A1(n4377), .A2(n6672), .ZN(n6670) );
  INV_X1 U6082 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5107) );
  MUX2_X1 U6083 ( .A(n8029), .B(n8028), .S(n8127), .Z(n8035) );
  NAND2_X1 U6084 ( .A1(n4414), .A2(n8077), .ZN(n4406) );
  INV_X1 U6085 ( .A(n4374), .ZN(n4415) );
  NAND2_X1 U6086 ( .A1(n8058), .A2(n8128), .ZN(n4375) );
  NOR2_X1 U6087 ( .A1(n8114), .A2(n8113), .ZN(n8121) );
  MUX2_X1 U6088 ( .A(n8000), .B(n7999), .S(n8128), .Z(n8006) );
  NAND4_X1 U6089 ( .A1(n5004), .A2(n4891), .A3(n4889), .A4(n4890), .ZN(n4929)
         );
  OAI21_X1 U6090 ( .B1(n7980), .B2(n9865), .A(n7979), .ZN(n7982) );
  OR2_X1 U6091 ( .A1(n8118), .A2(n8117), .ZN(n8131) );
  NAND2_X1 U6092 ( .A1(n8024), .A2(n8023), .ZN(n8027) );
  NAND2_X1 U6093 ( .A1(n8018), .A2(n8019), .ZN(n8024) );
  AND2_X1 U6094 ( .A1(n8061), .A2(n8048), .ZN(n4376) );
  NAND2_X1 U6095 ( .A1(n8047), .A2(n8652), .ZN(n8060) );
  NAND2_X1 U6096 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  OAI21_X1 U6097 ( .B1(n8089), .B2(n8088), .A(n8100), .ZN(n8091) );
  NAND2_X1 U6098 ( .A1(n6662), .A2(n6661), .ZN(n6660) );
  XNOR2_X1 U6099 ( .A(n6243), .B(n6242), .ZN(n6662) );
  INV_X1 U6100 ( .A(n4800), .ZN(n4799) );
  INV_X1 U6101 ( .A(n6349), .ZN(n4816) );
  NAND2_X1 U6102 ( .A1(n4730), .A2(n4731), .ZN(n5331) );
  NAND2_X1 U6103 ( .A1(n4744), .A2(n4743), .ZN(n9128) );
  NOR2_X1 U6104 ( .A1(n9274), .A2(n7634), .ZN(n9273) );
  NAND2_X1 U6105 ( .A1(n9435), .A2(n9770), .ZN(n4426) );
  NAND2_X1 U6106 ( .A1(n6346), .A2(n6345), .ZN(n6348) );
  OAI21_X1 U6107 ( .B1(n4767), .B2(n4766), .A(n4771), .ZN(n4765) );
  OAI211_X1 U6108 ( .C1(n4781), .C2(n4777), .A(n6033), .B(n4775), .ZN(n6034)
         );
  INV_X1 U6109 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U6110 ( .A1(n4638), .A2(n4637), .ZN(n8444) );
  NAND2_X1 U6111 ( .A1(n4570), .A2(n6673), .ZN(n4377) );
  NAND2_X1 U6112 ( .A1(n8988), .A2(n6584), .ZN(n9011) );
  NOR2_X1 U6113 ( .A1(n8383), .A2(n8384), .ZN(n8382) );
  XNOR2_X1 U6114 ( .A(n4991), .B(n5352), .ZN(n8383) );
  NAND2_X1 U6115 ( .A1(n4362), .A2(n4589), .ZN(n4979) );
  NAND4_X1 U6116 ( .A1(n4420), .A2(n4419), .A3(n4418), .A4(n4478), .ZN(
        P1_U3242) );
  NAND2_X1 U6117 ( .A1(n5418), .A2(n5417), .ZN(n5433) );
  NAND2_X1 U6118 ( .A1(n5495), .A2(n5494), .ZN(n5511) );
  NAND2_X1 U6119 ( .A1(n5584), .A2(n5583), .ZN(n5602) );
  INV_X1 U6120 ( .A(n7834), .ZN(n4496) );
  AOI21_X1 U6121 ( .B1(n4506), .B2(n4510), .A(n4363), .ZN(n4503) );
  NAND2_X1 U6122 ( .A1(n4504), .A2(n4503), .ZN(n7723) );
  NAND2_X1 U6123 ( .A1(n7739), .A2(n7760), .ZN(n4462) );
  AOI21_X1 U6124 ( .B1(n7707), .B2(n7706), .A(n7705), .ZN(n7708) );
  INV_X1 U6125 ( .A(n5693), .ZN(n5691) );
  AOI21_X1 U6126 ( .B1(n4620), .B2(n4614), .A(n4612), .ZN(n7591) );
  NAND2_X1 U6127 ( .A1(n8270), .A2(n8191), .ZN(n8345) );
  NAND2_X1 U6128 ( .A1(n8194), .A2(n8193), .ZN(n8226) );
  NOR2_X1 U6129 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  OAI21_X1 U6130 ( .B1(n8171), .B2(n8170), .A(n4881), .ZN(n8310) );
  OAI21_X1 U6131 ( .B1(n8182), .B2(n4626), .A(n4622), .ZN(n8188) );
  OAI22_X1 U6132 ( .A1(n7611), .A2(n7610), .B1(n7101), .B2(n7102), .ZN(n7618)
         );
  NAND2_X1 U6133 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(n4950), .ZN(n4576) );
  INV_X1 U6134 ( .A(n6696), .ZN(n4383) );
  AOI21_X1 U6135 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6626), .A(n7414), .ZN(
        n5019) );
  XNOR2_X1 U6136 ( .A(n5023), .B(n5423), .ZN(n9838) );
  NOR2_X1 U6137 ( .A1(n9837), .A2(n5024), .ZN(n5026) );
  NAND2_X1 U6138 ( .A1(n5026), .A2(n5025), .ZN(n4408) );
  INV_X1 U6139 ( .A(n4955), .ZN(n4953) );
  AOI21_X1 U6140 ( .B1(n4386), .B2(n9821), .A(n4384), .ZN(n8470) );
  XNOR2_X1 U6141 ( .A(n8457), .B(n8458), .ZN(n4386) );
  OAI21_X1 U6142 ( .B1(n8148), .B2(n8147), .A(n4387), .ZN(P2_U3296) );
  NAND2_X1 U6143 ( .A1(n4406), .A2(n4405), .ZN(n4404) );
  NAND2_X1 U6144 ( .A1(n4402), .A2(n4401), .ZN(n8093) );
  NAND2_X1 U6145 ( .A1(n5257), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U6146 ( .A1(n4742), .A2(n4741), .ZN(n4744) );
  NAND2_X1 U6147 ( .A1(n9128), .A2(n4873), .ZN(n9130) );
  INV_X1 U6148 ( .A(n4427), .ZN(n4413) );
  NAND2_X1 U6149 ( .A1(n4361), .A2(n4412), .ZN(n9435) );
  OAI21_X1 U6150 ( .B1(n4592), .B2(n4878), .A(n4587), .ZN(n4583) );
  NAND2_X1 U6151 ( .A1(n4584), .A2(n4582), .ZN(n4586) );
  XNOR2_X1 U6152 ( .A(n4566), .B(n8459), .ZN(n8471) );
  NAND2_X1 U6153 ( .A1(n5003), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U6154 ( .A1(n9780), .A2(n9781), .ZN(n9779) );
  NAND2_X1 U6155 ( .A1(n5024), .A2(n4657), .ZN(n4655) );
  NOR2_X1 U6156 ( .A1(n7409), .A2(n4410), .ZN(n4991) );
  NOR2_X1 U6157 ( .A1(n8434), .A2(n4411), .ZN(n4997) );
  NOR2_X1 U6158 ( .A1(n5023), .A2(n5423), .ZN(n5024) );
  NAND2_X1 U6159 ( .A1(n4496), .A2(n7900), .ZN(n4495) );
  NAND2_X1 U6160 ( .A1(n5480), .A2(n4738), .ZN(n4736) );
  AOI21_X1 U6161 ( .B1(n5527), .B2(n4697), .A(n4694), .ZN(n4693) );
  NAND2_X2 U6162 ( .A1(n4390), .A2(n6179), .ZN(n6226) );
  NAND2_X2 U6163 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  INV_X1 U6164 ( .A(n8534), .ZN(n4521) );
  NAND2_X1 U6165 ( .A1(n4553), .A2(n4551), .ZN(n8559) );
  OAI22_X1 U6166 ( .A1(n4711), .A2(n4707), .B1(n5293), .B2(n5294), .ZN(n4704)
         );
  NAND2_X1 U6167 ( .A1(n7182), .A2(n7856), .ZN(n6130) );
  OR2_X1 U6168 ( .A1(n6637), .A2(n6921), .ZN(n6639) );
  NAND2_X1 U6169 ( .A1(n6639), .A2(n5006), .ZN(n9780) );
  NAND2_X1 U6170 ( .A1(n5164), .A2(SI_3_), .ZN(n5184) );
  OAI21_X1 U6171 ( .B1(n9293), .B2(n4670), .A(n4667), .ZN(n9231) );
  NAND2_X2 U6172 ( .A1(n5904), .A2(n5903), .ZN(n7178) );
  NAND2_X1 U6173 ( .A1(n4400), .A2(n4397), .ZN(P1_U3518) );
  NOR2_X1 U6174 ( .A1(n9753), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U6175 ( .A1(n6186), .A2(n9753), .ZN(n4400) );
  NOR2_X1 U6176 ( .A1(n5015), .A2(n5014), .ZN(n9811) );
  NAND2_X1 U6177 ( .A1(n6129), .A2(n7858), .ZN(n7120) );
  XNOR2_X1 U6178 ( .A(n5019), .B(n5352), .ZN(n8389) );
  AOI21_X1 U6179 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6544), .A(n6888), .ZN(
        n5013) );
  NAND2_X1 U6180 ( .A1(n4826), .A2(n4358), .ZN(n6280) );
  NAND2_X1 U6181 ( .A1(n4439), .A2(n6279), .ZN(n6774) );
  NAND2_X1 U6182 ( .A1(n8949), .A2(n8948), .ZN(n8947) );
  NAND2_X1 U6183 ( .A1(n4449), .A2(n4447), .ZN(n8868) );
  NAND2_X4 U6184 ( .A1(n6846), .A2(n6226), .ZN(n6433) );
  MUX2_X2 U6185 ( .A(n7973), .B(n7972), .S(n8128), .Z(n7980) );
  NAND2_X1 U6186 ( .A1(n8133), .A2(n8132), .ZN(n8138) );
  INV_X1 U6187 ( .A(n4929), .ZN(n4549) );
  OR3_X1 U6188 ( .A1(n8772), .A2(n8127), .A3(n8180), .ZN(n4401) );
  NOR2_X1 U6189 ( .A1(n8556), .A2(n8081), .ZN(n4403) );
  INV_X1 U6190 ( .A(n4635), .ZN(n4908) );
  AOI21_X1 U6191 ( .B1(n4408), .B2(n4407), .A(n9852), .ZN(n5080) );
  INV_X1 U6192 ( .A(n8456), .ZN(n4407) );
  NAND2_X1 U6193 ( .A1(n5020), .A2(n4654), .ZN(n4650) );
  INV_X1 U6194 ( .A(n9845), .ZN(n4409) );
  NAND2_X1 U6195 ( .A1(n4586), .A2(n4585), .ZN(n4982) );
  NOR2_X1 U6196 ( .A1(n7370), .A2(n7369), .ZN(n7368) );
  NOR2_X1 U6197 ( .A1(n9121), .A2(n9120), .ZN(n4424) );
  XNOR2_X1 U6198 ( .A(n4424), .B(n9129), .ZN(n4690) );
  NAND3_X1 U6199 ( .A1(n8070), .A2(n8069), .A3(n8068), .ZN(n4414) );
  NAND2_X1 U6200 ( .A1(n4415), .A2(n8049), .ZN(n8052) );
  NAND2_X1 U6201 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  INV_X1 U6202 ( .A(n4485), .ZN(n4484) );
  NOR3_X1 U6203 ( .A1(n5080), .A2(n5079), .A3(n5078), .ZN(n5081) );
  NAND2_X1 U6204 ( .A1(n4736), .A2(n4735), .ZN(n5495) );
  INV_X1 U6205 ( .A(n9241), .ZN(n4672) );
  NAND2_X1 U6206 ( .A1(n9185), .A2(n7812), .ZN(n9169) );
  NOR2_X2 U6207 ( .A1(n5742), .A2(n5829), .ZN(n4761) );
  NAND4_X1 U6208 ( .A1(n5740), .A2(n5842), .A3(n5875), .A4(n5982), .ZN(n5742)
         );
  INV_X1 U6209 ( .A(n4438), .ZN(n9225) );
  NAND2_X1 U6210 ( .A1(n6774), .A2(n6775), .ZN(n6282) );
  NAND2_X1 U6211 ( .A1(n6280), .A2(n6277), .ZN(n4439) );
  NOR2_X2 U6212 ( .A1(n6315), .A2(n4440), .ZN(n9521) );
  NOR2_X2 U6213 ( .A1(n4441), .A2(n6314), .ZN(n6315) );
  NAND2_X1 U6214 ( .A1(n4819), .A2(n4442), .ZN(n4444) );
  NAND3_X1 U6215 ( .A1(n4444), .A2(n4443), .A3(n4332), .ZN(n8949) );
  NAND2_X1 U6216 ( .A1(n4819), .A2(n4816), .ZN(n4446) );
  NAND2_X1 U6217 ( .A1(n8898), .A2(n4451), .ZN(n4449) );
  NAND4_X1 U6218 ( .A1(n5979), .A2(n4761), .A3(n4460), .A4(n4870), .ZN(n6112)
         );
  INV_X1 U6219 ( .A(n7658), .ZN(n4477) );
  NOR2_X2 U6220 ( .A1(n7904), .A2(n4494), .ZN(n4485) );
  NAND2_X2 U6221 ( .A1(n6548), .A2(n5774), .ZN(n5844) );
  NAND2_X2 U6222 ( .A1(n5769), .A2(n5770), .ZN(n6138) );
  OAI211_X1 U6223 ( .C1(n4509), .C2(n4508), .A(n4502), .B(n4501), .ZN(n4507)
         );
  NAND3_X1 U6224 ( .A1(n7708), .A2(n7710), .A3(n4672), .ZN(n4502) );
  NAND2_X1 U6225 ( .A1(n7709), .A2(n4506), .ZN(n4504) );
  XNOR2_X2 U6226 ( .A(n7053), .B(n6225), .ZN(n6117) );
  NAND2_X1 U6227 ( .A1(n5653), .A2(n4515), .ZN(n8648) );
  OAI211_X1 U6228 ( .C1(n5158), .C2(n6515), .A(n4348), .B(n5148), .ZN(n5149)
         );
  NAND2_X1 U6229 ( .A1(n5635), .A2(n4525), .ZN(n4523) );
  NAND2_X1 U6230 ( .A1(n4524), .A2(n4523), .ZN(n7211) );
  NAND2_X1 U6231 ( .A1(n5647), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U6232 ( .A1(n4532), .A2(n4534), .ZN(n5645) );
  NAND2_X1 U6233 ( .A1(n7222), .A2(n4537), .ZN(n4532) );
  AND2_X1 U6234 ( .A1(n4897), .A2(n4901), .ZN(n4544) );
  NAND3_X1 U6235 ( .A1(n4549), .A2(n4545), .A3(n4298), .ZN(n4915) );
  AND2_X1 U6236 ( .A1(n4896), .A2(n4897), .ZN(n4546) );
  NAND3_X1 U6237 ( .A1(n4546), .A2(n4898), .A3(n4899), .ZN(n4550) );
  NAND2_X1 U6238 ( .A1(n8589), .A2(n4554), .ZN(n4553) );
  NAND3_X1 U6239 ( .A1(n4959), .A2(n6673), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6671) );
  NAND2_X1 U6240 ( .A1(n4959), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U6241 ( .A1(n4574), .A2(n4575), .ZN(n6523) );
  NAND2_X1 U6242 ( .A1(n4971), .A2(n4329), .ZN(n4585) );
  INV_X1 U6243 ( .A(n6723), .ZN(n4591) );
  NAND2_X1 U6244 ( .A1(n4971), .A2(n4306), .ZN(n4589) );
  NAND2_X1 U6245 ( .A1(n8356), .A2(n8355), .ZN(n8277) );
  NAND2_X1 U6246 ( .A1(n4596), .A2(n4599), .ZN(n8167) );
  NAND2_X1 U6247 ( .A1(n8356), .A2(n4597), .ZN(n4596) );
  NAND2_X1 U6248 ( .A1(n7241), .A2(n4296), .ZN(n4604) );
  INV_X1 U6249 ( .A(n8379), .ZN(n4610) );
  NAND2_X1 U6250 ( .A1(n8300), .A2(n4628), .ZN(n8243) );
  NAND2_X1 U6251 ( .A1(n8226), .A2(n8225), .ZN(n8228) );
  NOR2_X2 U6252 ( .A1(n4915), .A2(n4636), .ZN(n4635) );
  OAI21_X1 U6253 ( .B1(n4979), .B2(n4587), .A(n6877), .ZN(n9794) );
  NAND2_X1 U6254 ( .A1(n6670), .A2(n4966), .ZN(n4969) );
  NAND2_X1 U6255 ( .A1(n4968), .A2(n5207), .ZN(n4970) );
  NAND2_X1 U6256 ( .A1(n4644), .A2(n5157), .ZN(n4643) );
  INV_X1 U6257 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U6258 ( .A1(n9779), .A2(n5007), .ZN(n4645) );
  INV_X1 U6259 ( .A(n9811), .ZN(n4646) );
  AOI21_X1 U6260 ( .B1(n4646), .B2(n4647), .A(n4648), .ZN(n7378) );
  OAI21_X1 U6261 ( .B1(n5015), .B2(P2_REG1_REG_9__SCAN_IN), .A(n4649), .ZN(
        n4648) );
  INV_X1 U6262 ( .A(n7379), .ZN(n4649) );
  NOR2_X1 U6263 ( .A1(n9809), .A2(n5015), .ZN(n7380) );
  AND2_X1 U6264 ( .A1(n9811), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9809) );
  OAI21_X1 U6265 ( .B1(n8389), .B2(n4651), .A(n4650), .ZN(n8409) );
  OAI21_X1 U6266 ( .B1(n9838), .B2(n4656), .A(n4655), .ZN(n8456) );
  NOR2_X1 U6267 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
  INV_X1 U6268 ( .A(n5025), .ZN(n4657) );
  NAND2_X1 U6269 ( .A1(n9342), .A2(n4663), .ZN(n4659) );
  NAND2_X1 U6270 ( .A1(n4659), .A2(n4660), .ZN(n9309) );
  NAND3_X1 U6271 ( .A1(n5979), .A2(n4761), .A3(n4760), .ZN(n4666) );
  INV_X1 U6272 ( .A(n4671), .ZN(n4670) );
  XNOR2_X1 U6273 ( .A(n6117), .B(n7040), .ZN(n9694) );
  INV_X1 U6274 ( .A(n7297), .ZN(n4680) );
  AOI21_X2 U6275 ( .B1(n4680), .B2(n4683), .A(n4679), .ZN(n7431) );
  OR2_X1 U6276 ( .A1(n6548), .A2(n6599), .ZN(n4686) );
  NAND2_X2 U6277 ( .A1(n6548), .A2(n6514), .ZN(n5845) );
  OR2_X2 U6278 ( .A1(n7120), .A2(n4691), .ZN(n7182) );
  NAND2_X1 U6279 ( .A1(n5325), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4692) );
  INV_X1 U6280 ( .A(n4693), .ZN(n5564) );
  AOI21_X1 U6281 ( .B1(n5527), .B2(n5526), .A(n4699), .ZN(n4696) );
  INV_X1 U6282 ( .A(n4696), .ZN(n5545) );
  INV_X1 U6283 ( .A(n5269), .ZN(n4712) );
  NAND2_X1 U6284 ( .A1(n5433), .A2(n4716), .ZN(n4713) );
  NAND2_X1 U6285 ( .A1(n4736), .A2(n4737), .ZN(n5491) );
  NAND2_X1 U6286 ( .A1(n5478), .A2(n5479), .ZN(n4737) );
  NAND2_X1 U6287 ( .A1(n9174), .A2(n6087), .ZN(n4742) );
  OAI21_X1 U6288 ( .B1(n6989), .B2(n7785), .A(n4749), .ZN(n7181) );
  INV_X1 U6289 ( .A(n4746), .ZN(n5952) );
  AOI21_X1 U6290 ( .B1(n6989), .B2(n4749), .A(n4747), .ZN(n4746) );
  NAND2_X1 U6291 ( .A1(n4748), .A2(n4877), .ZN(n4747) );
  NAND2_X1 U6292 ( .A1(n4749), .A2(n7785), .ZN(n4748) );
  NAND2_X1 U6293 ( .A1(n7011), .A2(n4752), .ZN(n4751) );
  NOR2_X1 U6294 ( .A1(n4756), .A2(n5742), .ZN(n4757) );
  NAND3_X1 U6295 ( .A1(n5743), .A2(n5745), .A3(n6154), .ZN(n4756) );
  INV_X1 U6296 ( .A(n5751), .ZN(n4760) );
  NAND3_X1 U6297 ( .A1(n4760), .A2(n4758), .A3(n4757), .ZN(n6161) );
  NAND2_X1 U6298 ( .A1(n7266), .A2(n4763), .ZN(n4762) );
  INV_X1 U6299 ( .A(n6009), .ZN(n7429) );
  INV_X1 U6300 ( .A(n9321), .ZN(n4781) );
  CLKBUF_X1 U6301 ( .A(n4781), .Z(n4773) );
  INV_X1 U6302 ( .A(n4796), .ZN(n9191) );
  NAND2_X1 U6303 ( .A1(n9211), .A2(n8965), .ZN(n4797) );
  OAI21_X2 U6304 ( .B1(n7284), .B2(n4352), .A(n4799), .ZN(n7390) );
  NAND2_X1 U6305 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
  NAND2_X1 U6306 ( .A1(n6406), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6307 ( .A1(n6406), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U6308 ( .A1(n4342), .A2(n4818), .ZN(n4819) );
  INV_X1 U6309 ( .A(n4819), .ZN(n8838) );
  NAND2_X1 U6310 ( .A1(n6713), .A2(n6714), .ZN(n4826) );
  OAI21_X1 U6311 ( .B1(n7035), .B2(n6298), .A(n6297), .ZN(n7166) );
  NAND2_X2 U6312 ( .A1(n6395), .A2(n6394), .ZN(n8848) );
  NAND2_X1 U6313 ( .A1(n6108), .A2(n4839), .ZN(n6109) );
  NAND2_X1 U6314 ( .A1(n6108), .A2(n4838), .ZN(n6158) );
  NOR2_X1 U6315 ( .A1(n4840), .A2(n4355), .ZN(n5732) );
  NAND2_X1 U6316 ( .A1(n8555), .A2(n4356), .ZN(n4843) );
  NAND2_X1 U6317 ( .A1(n7345), .A2(n4856), .ZN(n4855) );
  NAND3_X1 U6318 ( .A1(n4860), .A2(n5661), .A3(n8072), .ZN(n4858) );
  NAND2_X1 U6319 ( .A1(n4863), .A2(n4862), .ZN(n7581) );
  NAND2_X1 U6320 ( .A1(n7511), .A2(n5364), .ZN(n4863) );
  XNOR2_X1 U6321 ( .A(n6207), .B(n6206), .ZN(n8221) );
  NAND2_X1 U6322 ( .A1(n7734), .A2(n7725), .ZN(n7823) );
  NAND2_X1 U6323 ( .A1(n7759), .A2(n9115), .ZN(n7763) );
  NAND2_X1 U6324 ( .A1(n9720), .A2(n6943), .ZN(n9713) );
  NAND2_X1 U6325 ( .A1(n5144), .A2(n5143), .ZN(n5160) );
  CLKBUF_X1 U6326 ( .A(n7266), .Z(n7268) );
  NAND2_X1 U6327 ( .A1(n5138), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5106) );
  INV_X1 U6328 ( .A(n5146), .ZN(n5143) );
  OAI21_X1 U6329 ( .B1(n6514), .B2(n6528), .A(n5210), .ZN(n5211) );
  NAND2_X1 U6330 ( .A1(n6514), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6331 ( .A1(n5819), .A2(n5818), .ZN(n5825) );
  OR2_X1 U6332 ( .A1(n5819), .A2(n5808), .ZN(n5809) );
  NAND2_X1 U6333 ( .A1(n5820), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6334 ( .A1(n5645), .A2(n5644), .ZN(n7399) );
  NAND2_X1 U6335 ( .A1(n7970), .A2(n7969), .ZN(n6897) );
  NAND2_X1 U6336 ( .A1(n9128), .A2(n6104), .ZN(n9150) );
  INV_X1 U6337 ( .A(n8220), .ZN(n5760) );
  OR2_X1 U6338 ( .A1(n6103), .A2(n7801), .ZN(n6104) );
  XNOR2_X1 U6339 ( .A(n7919), .B(n8105), .ZN(n8480) );
  CLKBUF_X1 U6340 ( .A(n7031), .Z(n7035) );
  INV_X1 U6341 ( .A(n8310), .ZN(n8312) );
  NAND2_X1 U6342 ( .A1(n7984), .A2(n7992), .ZN(n7933) );
  OR2_X1 U6343 ( .A1(n6860), .A2(n7296), .ZN(n6851) );
  AOI21_X1 U6344 ( .B1(n7043), .B2(n6448), .A(n6237), .ZN(n6241) );
  INV_X1 U6345 ( .A(n5096), .ZN(n5094) );
  XNOR2_X1 U6346 ( .A(n7101), .B(n7102), .ZN(n7610) );
  AND2_X1 U6347 ( .A1(n5727), .A2(n5726), .ZN(n9936) );
  INV_X1 U6348 ( .A(n9954), .ZN(n5718) );
  INV_X1 U6349 ( .A(n7101), .ZN(n6763) );
  AND3_X1 U6350 ( .A1(n6107), .A2(n6106), .A3(n6105), .ZN(n4870) );
  INV_X1 U6351 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5690) );
  AND2_X1 U6352 ( .A1(n7987), .A2(n7985), .ZN(n4871) );
  OR2_X1 U6353 ( .A1(n9145), .A2(n9414), .ZN(n4872) );
  AND2_X1 U6354 ( .A1(n6454), .A2(n9531), .ZN(n4874) );
  NOR2_X1 U6355 ( .A1(n5659), .A2(n5658), .ZN(n4875) );
  AND2_X1 U6356 ( .A1(n6455), .A2(n4874), .ZN(n4876) );
  INV_X1 U6357 ( .A(n9353), .ZN(n6220) );
  INV_X1 U6358 ( .A(n8040), .ZN(n5378) );
  INV_X1 U6359 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8294) );
  AND2_X1 U6360 ( .A1(n6531), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4878) );
  INV_X1 U6361 ( .A(n9142), .ZN(n6152) );
  INV_X1 U6362 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5137) );
  INV_X1 U6363 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5109) );
  AND2_X2 U6364 ( .A1(n6185), .A2(n6844), .ZN(n9753) );
  INV_X1 U6365 ( .A(n8222), .ZN(n9476) );
  OR2_X1 U6366 ( .A1(n5663), .A2(n8328), .ZN(n4879) );
  NAND2_X1 U6367 ( .A1(n8602), .A2(n5655), .ZN(n4880) );
  NAND2_X1 U6368 ( .A1(n5135), .A2(n5134), .ZN(n5145) );
  OR2_X1 U6369 ( .A1(n8169), .A2(n8604), .ZN(n4881) );
  OR2_X1 U6370 ( .A1(n5416), .A2(SI_16_), .ZN(n4882) );
  OR2_X1 U6371 ( .A1(n8377), .A2(n7257), .ZN(n4883) );
  OR2_X1 U6372 ( .A1(n5493), .A2(SI_21_), .ZN(n4884) );
  NAND2_X1 U6373 ( .A1(n7568), .A2(n8372), .ZN(n4885) );
  INV_X1 U6374 ( .A(n7460), .ZN(n8958) );
  INV_X1 U6375 ( .A(n7965), .ZN(n7958) );
  NOR2_X1 U6376 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4896) );
  NAND2_X1 U6377 ( .A1(n4958), .A2(n5157), .ZN(n4959) );
  INV_X1 U6378 ( .A(n9115), .ZN(n7761) );
  INV_X1 U6379 ( .A(n8620), .ZN(n8165) );
  NOR2_X1 U6380 ( .A1(n8278), .A2(n8634), .ZN(n8154) );
  INV_X1 U6381 ( .A(n8912), .ZN(n6417) );
  INV_X1 U6382 ( .A(n8926), .ZN(n6396) );
  INV_X1 U6383 ( .A(SI_20_), .ZN(n5479) );
  NAND2_X1 U6384 ( .A1(n8164), .A2(n8165), .ZN(n8166) );
  OR2_X1 U6385 ( .A1(n4284), .A2(n5097), .ZN(n5098) );
  NAND2_X1 U6386 ( .A1(n6544), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4983) );
  INV_X1 U6387 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8253) );
  INV_X1 U6388 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5283) );
  AOI22_X1 U6389 ( .A1(n8490), .A2(n8491), .B1(n8369), .B2(n8495), .ZN(n5671)
         );
  INV_X1 U6390 ( .A(n9858), .ZN(n9865) );
  INV_X1 U6391 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4923) );
  INV_X1 U6392 ( .A(n6039), .ZN(n5737) );
  INV_X1 U6393 ( .A(SI_22_), .ZN(n5496) );
  INV_X1 U6394 ( .A(SI_19_), .ZN(n5452) );
  INV_X1 U6395 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5741) );
  OR2_X1 U6396 ( .A1(n5439), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5459) );
  AND2_X1 U6397 ( .A1(n5013), .A2(n9816), .ZN(n5014) );
  INV_X1 U6398 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7412) );
  INV_X1 U6399 ( .A(n5556), .ZN(n5555) );
  NAND2_X1 U6400 ( .A1(n5356), .A2(n5355), .ZN(n5371) );
  OR2_X1 U6401 ( .A1(n8799), .A2(n8647), .ZN(n8061) );
  OR2_X1 U6402 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  INV_X1 U6403 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5916) );
  INV_X1 U6404 ( .A(n7742), .ZN(n6212) );
  NOR2_X1 U6405 ( .A1(n9151), .A2(n9157), .ZN(n9154) );
  OR2_X1 U6406 ( .A1(n9399), .A2(n9311), .ZN(n6033) );
  INV_X1 U6407 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U6408 ( .A1(n5163), .A2(n5162), .ZN(n5165) );
  INV_X1 U6409 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5241) );
  INV_X1 U6410 ( .A(n8604), .ZN(n8336) );
  XNOR2_X1 U6411 ( .A(n7100), .B(n7099), .ZN(n7102) );
  NAND2_X1 U6412 ( .A1(n8190), .A2(n5631), .ZN(n8191) );
  INV_X1 U6413 ( .A(n7137), .ZN(n5504) );
  OR2_X1 U6414 ( .A1(n5608), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U6415 ( .A1(n5485), .A2(n5484), .ZN(n5502) );
  NAND2_X1 U6416 ( .A1(n7093), .A2(n7095), .ZN(n6813) );
  INV_X1 U6417 ( .A(n8372), .ZN(n7563) );
  INV_X1 U6418 ( .A(n9933), .ZN(n9911) );
  OR2_X1 U6419 ( .A1(n4932), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U6420 ( .A1(n6255), .A2(n6254), .ZN(n6713) );
  INV_X1 U6421 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U6422 ( .A1(n6660), .A2(n6245), .ZN(n6629) );
  OR2_X1 U6423 ( .A1(n9677), .A2(n9638), .ZN(n6848) );
  INV_X1 U6424 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6184) );
  OAI21_X1 U6425 ( .B1(n6905), .B2(n6906), .A(n5873), .ZN(n6850) );
  INV_X1 U6426 ( .A(n9345), .ZN(n9723) );
  NAND2_X1 U6427 ( .A1(n5790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  INV_X1 U6428 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10000) );
  INV_X1 U6429 ( .A(n5193), .ZN(n5190) );
  AND2_X1 U6430 ( .A1(n5562), .A2(n5561), .ZN(n5631) );
  INV_X1 U6431 ( .A(n9835), .ZN(n9817) );
  INV_X1 U6432 ( .A(n9826), .ZN(n9843) );
  INV_X1 U6433 ( .A(n8661), .ZN(n8613) );
  INV_X1 U6434 ( .A(n8481), .ZN(n8658) );
  INV_X1 U6435 ( .A(n8670), .ZN(n8714) );
  AND2_X1 U6436 ( .A1(n9954), .A2(n9933), .ZN(n8715) );
  AND2_X1 U6437 ( .A1(n7451), .A2(n9873), .ZN(n9926) );
  NAND2_X1 U6438 ( .A1(n7451), .A2(n7958), .ZN(n9928) );
  AND2_X1 U6439 ( .A1(n4995), .A2(n4933), .ZN(n5403) );
  INV_X1 U6440 ( .A(n9535), .ZN(n8955) );
  OR2_X1 U6441 ( .A1(n6089), .A2(n6088), .ZN(n9134) );
  OR2_X1 U6442 ( .A1(n9236), .A2(n6081), .ZN(n5766) );
  INV_X1 U6443 ( .A(n9620), .ZN(n9595) );
  AND2_X1 U6444 ( .A1(n6615), .A2(n8994), .ZN(n9623) );
  OR2_X1 U6445 ( .A1(n7907), .A2(n7484), .ZN(n6552) );
  AND2_X1 U6446 ( .A1(n7701), .A2(n7878), .ZN(n9294) );
  INV_X1 U6447 ( .A(n9341), .ZN(n9334) );
  AND2_X1 U6448 ( .A1(n6146), .A2(n6138), .ZN(n9345) );
  INV_X1 U6449 ( .A(n9655), .ZN(n10148) );
  INV_X1 U6450 ( .A(n10140), .ZN(n9652) );
  AOI21_X1 U6451 ( .B1(n6536), .B2(n6184), .A(n6542), .ZN(n6464) );
  AND2_X1 U6452 ( .A1(n9687), .A2(n6232), .ZN(n9416) );
  NAND2_X1 U6453 ( .A1(n9638), .A2(n9689), .ZN(n9750) );
  AND2_X1 U6454 ( .A1(n6115), .A2(n7840), .ZN(n9687) );
  XNOR2_X1 U6455 ( .A(n6162), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6180) );
  AND2_X1 U6456 ( .A1(n5912), .A2(n5902), .ZN(n6612) );
  INV_X1 U6457 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5842) );
  INV_X1 U6458 ( .A(n8362), .ZN(n8339) );
  INV_X1 U6459 ( .A(n8350), .ZN(n8365) );
  INV_X1 U6460 ( .A(n8635), .ZN(n8605) );
  OR2_X1 U6461 ( .A1(n8381), .A2(n5676), .ZN(n9826) );
  INV_X1 U6462 ( .A(n9821), .ZN(n9852) );
  OR2_X1 U6463 ( .A1(n6572), .A2(n5675), .ZN(n9848) );
  INV_X2 U6464 ( .A(n9881), .ZN(n9878) );
  OR2_X1 U6465 ( .A1(n6820), .A2(n8532), .ZN(n8481) );
  INV_X1 U6466 ( .A(n8715), .ZN(n8693) );
  AND3_X2 U6467 ( .A1(n6814), .A2(n5714), .A3(n5720), .ZN(n9954) );
  INV_X1 U6468 ( .A(n8807), .ZN(n8787) );
  AND3_X1 U6469 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(n9945) );
  INV_X2 U6470 ( .A(n9936), .ZN(n9934) );
  NAND2_X1 U6471 ( .A1(n5697), .A2(n5696), .ZN(n6812) );
  NAND2_X1 U6472 ( .A1(n5693), .A2(n6761), .ZN(n6565) );
  INV_X1 U6473 ( .A(n6226), .ZN(n6495) );
  INV_X1 U6474 ( .A(n7275), .ZN(n9739) );
  INV_X1 U6475 ( .A(n9531), .ZN(n8945) );
  NAND2_X1 U6476 ( .A1(n6102), .A2(n6101), .ZN(n8961) );
  OAI21_X1 U6477 ( .B1(n9288), .B2(n6081), .A(n5789), .ZN(n9311) );
  NAND2_X1 U6478 ( .A1(n6552), .A2(n6550), .ZN(n9635) );
  OR2_X1 U6479 ( .A1(n9677), .A2(n6851), .ZN(n10140) );
  NAND2_X1 U6480 ( .A1(n6845), .A2(n9326), .ZN(n10141) );
  NAND2_X1 U6481 ( .A1(n9770), .A2(n9416), .ZN(n9414) );
  INV_X1 U6482 ( .A(n9770), .ZN(n9768) );
  INV_X1 U6483 ( .A(n9753), .ZN(n9752) );
  AND2_X1 U6484 ( .A1(n6537), .A2(n7907), .ZN(n9678) );
  AND2_X1 U6485 ( .A1(n7532), .A2(n7606), .ZN(n6542) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7626) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7453) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7009) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10109) );
  INV_X1 U6490 ( .A(n8381), .ZN(P2_U3893) );
  OAI21_X1 U6491 ( .B1(n5082), .B2(n9848), .A(n5081), .ZN(P2_U3200) );
  AND2_X2 U6492 ( .A1(n6496), .A2(n6495), .ZN(P1_U3973) );
  AOI21_X1 U6493 ( .B1(n9537), .B2(n9753), .A(n6224), .ZN(P1_U3521) );
  NAND2_X1 U6494 ( .A1(n4935), .A2(n4892), .ZN(n4930) );
  INV_X1 U6495 ( .A(n4930), .ZN(n4899) );
  INV_X1 U6496 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4895) );
  INV_X1 U6497 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U6498 ( .A1(n4920), .A2(n4921), .ZN(n4902) );
  NAND2_X1 U6499 ( .A1(n4908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4907) );
  MUX2_X1 U6500 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4907), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n4909) );
  INV_X1 U6501 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6502 ( .A1(n4911), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U6503 ( .A1(n4915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4916) );
  INV_X1 U6504 ( .A(n4917), .ZN(n4918) );
  NAND2_X1 U6505 ( .A1(n4918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U6506 ( .A1(n5721), .A2(n8127), .ZN(n4922) );
  NAND2_X1 U6507 ( .A1(n4922), .A2(n7090), .ZN(n5074) );
  NAND2_X1 U6508 ( .A1(n4925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4926) );
  NAND2_X1 U6509 ( .A1(n5074), .A2(n5685), .ZN(n4928) );
  NAND2_X1 U6510 ( .A1(n4928), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U6511 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U6512 ( .A1(n4929), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U6513 ( .A1(n4946), .A2(n4894), .ZN(n4941) );
  OAI21_X1 U6514 ( .B1(n4939), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4936) );
  NAND2_X1 U6515 ( .A1(n4930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U6516 ( .A1(n4936), .A2(n4931), .ZN(n4932) );
  NAND2_X1 U6517 ( .A1(n4932), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6518 ( .A1(n4936), .A2(n4935), .ZN(n4938) );
  NAND2_X1 U6519 ( .A1(n4938), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4934) );
  XNOR2_X1 U6520 ( .A(n4934), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6521 ( .A1(n4936), .A2(n4935), .ZN(n4937) );
  NAND2_X1 U6522 ( .A1(n4939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U6523 ( .A(n4940), .B(P2_IR_REG_13__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6524 ( .A1(n4941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4942) );
  XNOR2_X1 U6525 ( .A(n4942), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7420) );
  INV_X1 U6526 ( .A(n7420), .ZN(n6626) );
  OR2_X1 U6527 ( .A1(n4946), .A2(n5090), .ZN(n4943) );
  XNOR2_X1 U6528 ( .A(n4943), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7476) );
  NOR2_X1 U6529 ( .A1(n4944), .A2(n5090), .ZN(n4945) );
  MUX2_X1 U6530 ( .A(n5090), .B(n4945), .S(P2_IR_REG_10__SCAN_IN), .Z(n4947)
         );
  INV_X1 U6531 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9793) );
  INV_X1 U6532 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9880) );
  INV_X1 U6533 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U6534 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4950) );
  INV_X1 U6535 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U6536 ( .A1(n5004), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4951) );
  INV_X1 U6537 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U6538 ( .A1(n6645), .A2(n4951), .ZN(n9773) );
  OR2_X1 U6539 ( .A1(n9771), .A2(n9880), .ZN(n4952) );
  NAND2_X1 U6540 ( .A1(n9772), .A2(n4952), .ZN(n4957) );
  NAND2_X1 U6541 ( .A1(n4955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4954) );
  INV_X1 U6542 ( .A(n4957), .ZN(n4958) );
  INV_X1 U6543 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6701) );
  INV_X1 U6544 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U6545 ( .A1(n4961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4960) );
  MUX2_X1 U6546 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4960), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n4964) );
  INV_X1 U6547 ( .A(n4961), .ZN(n4963) );
  INV_X1 U6548 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6549 ( .A1(n4963), .A2(n4962), .ZN(n4972) );
  NAND2_X1 U6550 ( .A1(n4964), .A2(n4972), .ZN(n6520) );
  MUX2_X1 U6551 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n4965), .S(n6520), .Z(n6672)
         );
  NAND2_X1 U6552 ( .A1(n6520), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4966) );
  INV_X1 U6553 ( .A(n4969), .ZN(n4968) );
  NAND2_X1 U6554 ( .A1(n4972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4967) );
  XNOR2_X1 U6555 ( .A(n4967), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6556 ( .A1(n4969), .A2(n6527), .ZN(n6723) );
  INV_X1 U6557 ( .A(n6501), .ZN(n4971) );
  INV_X1 U6558 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U6559 ( .A1(n4975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4974) );
  MUX2_X1 U6560 ( .A(n4974), .B(P2_IR_REG_31__SCAN_IN), .S(n4973), .Z(n4977)
         );
  INV_X1 U6561 ( .A(n4975), .ZN(n4976) );
  NAND2_X1 U6562 ( .A1(n4976), .A2(n4973), .ZN(n4980) );
  XNOR2_X1 U6563 ( .A(n6531), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U6564 ( .A1(n4980), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4978) );
  INV_X1 U6565 ( .A(n4982), .ZN(n6877) );
  OAI21_X1 U6566 ( .B1(n4980), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4981) );
  XNOR2_X1 U6567 ( .A(n6882), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U6568 ( .A1(n4929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4984) );
  XNOR2_X1 U6569 ( .A(n4984), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9816) );
  INV_X1 U6570 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U6571 ( .A1(n4986), .A2(n9812), .ZN(n7370) );
  NAND2_X1 U6572 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6568), .ZN(n4987) );
  OAI21_X1 U6573 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6568), .A(n4987), .ZN(
        n7369) );
  NOR2_X1 U6574 ( .A1(n7476), .A2(n4988), .ZN(n4989) );
  INV_X1 U6575 ( .A(n7476), .ZN(n6622) );
  INV_X1 U6576 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n4990) );
  AOI22_X1 U6577 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7420), .B1(n6626), .B2(
        n4990), .ZN(n7410) );
  NOR2_X1 U6578 ( .A1(n7411), .A2(n7410), .ZN(n7409) );
  NOR2_X1 U6579 ( .A1(n5352), .A2(n4991), .ZN(n4992) );
  INV_X1 U6580 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8384) );
  INV_X1 U6581 ( .A(n5352), .ZN(n8394) );
  INV_X1 U6582 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7585) );
  AOI22_X1 U6583 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n5368), .B1(n8408), .B2(
        n7585), .ZN(n8400) );
  NOR2_X1 U6584 ( .A1(n5383), .A2(n4993), .ZN(n4994) );
  INV_X1 U6585 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8656) );
  INV_X1 U6586 ( .A(n5383), .ZN(n8425) );
  INV_X1 U6587 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8639) );
  AOI22_X1 U6588 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n5403), .B1(n8443), .B2(
        n8639), .ZN(n8435) );
  NOR2_X1 U6589 ( .A1(n8436), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U6590 ( .A1(n4995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4996) );
  XNOR2_X1 U6591 ( .A(n4996), .B(P2_IR_REG_17__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U6592 ( .A(n4997), .B(n5423), .ZN(n9846) );
  NAND2_X1 U6593 ( .A1(n4998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4999) );
  XNOR2_X1 U6594 ( .A(n4999), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8461) );
  INV_X1 U6595 ( .A(n8461), .ZN(n7163) );
  NAND2_X1 U6596 ( .A1(n7163), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8452) );
  OAI21_X1 U6597 ( .B1(n7163), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8452), .ZN(
        n5000) );
  AOI21_X1 U6598 ( .B1(n5001), .B2(n5000), .A(n8453), .ZN(n5082) );
  NOR2_X1 U6599 ( .A1(n5002), .A2(P2_U3151), .ZN(n8822) );
  AND2_X1 U6600 ( .A1(n5074), .A2(n8822), .ZN(n5027) );
  INV_X1 U6601 ( .A(n5027), .ZN(n6572) );
  INV_X1 U6602 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9937) );
  INV_X1 U6603 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U6604 ( .A1(n5116), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6605 ( .A1(n5004), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5006) );
  OAI21_X1 U6606 ( .B1(n6523), .B2(n5005), .A(n5006), .ZN(n6637) );
  INV_X1 U6607 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6921) );
  OR2_X1 U6608 ( .A1(n9771), .A2(n9937), .ZN(n5007) );
  INV_X1 U6609 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U6610 ( .A1(n6698), .A2(n6679), .ZN(n5008) );
  INV_X1 U6611 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9941) );
  MUX2_X1 U6612 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9941), .S(n6520), .Z(n6678)
         );
  NAND2_X1 U6613 ( .A1(n6520), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U6614 ( .A1(n6682), .A2(n5009), .ZN(n5010) );
  OAI21_X1 U6615 ( .B1(n5010), .B2(n6527), .A(n6729), .ZN(n6503) );
  INV_X1 U6616 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9943) );
  XNOR2_X1 U6617 ( .A(n6531), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6730) );
  INV_X1 U6618 ( .A(n6885), .ZN(n5012) );
  INV_X1 U6619 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5264) );
  XNOR2_X1 U6620 ( .A(n6882), .B(n5264), .ZN(n6883) );
  INV_X1 U6621 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U6622 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6568), .ZN(n5016) );
  OAI21_X1 U6623 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6568), .A(n5016), .ZN(
        n7379) );
  NOR2_X1 U6624 ( .A1(n7476), .A2(n5017), .ZN(n5018) );
  INV_X1 U6625 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9952) );
  XOR2_X1 U6626 ( .A(n6622), .B(n5017), .Z(n7472) );
  NOR2_X1 U6627 ( .A1(n9952), .A2(n7472), .ZN(n7471) );
  INV_X1 U6628 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10079) );
  XNOR2_X1 U6629 ( .A(n7420), .B(n10079), .ZN(n7415) );
  NOR2_X1 U6630 ( .A1(n7416), .A2(n7415), .ZN(n7414) );
  NOR2_X1 U6631 ( .A1(n5352), .A2(n5019), .ZN(n5020) );
  INV_X1 U6632 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10050) );
  INV_X1 U6633 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5373) );
  AOI22_X1 U6634 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n5368), .B1(n8408), .B2(
        n5373), .ZN(n8410) );
  NOR2_X1 U6635 ( .A1(n5383), .A2(n5021), .ZN(n5022) );
  INV_X1 U6636 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8713) );
  INV_X1 U6637 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8710) );
  AOI22_X1 U6638 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n5403), .B1(n8443), .B2(
        n8710), .ZN(n8445) );
  INV_X1 U6639 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9839) );
  INV_X1 U6640 ( .A(n5423), .ZN(n9834) );
  NAND2_X1 U6641 ( .A1(n7163), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8454) );
  OAI21_X1 U6642 ( .B1(n7163), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8454), .ZN(
        n5025) );
  MUX2_X1 U6643 ( .A(n9847), .B(n9839), .S(n5675), .Z(n5028) );
  NAND2_X1 U6644 ( .A1(n5028), .A2(n5423), .ZN(n5063) );
  XNOR2_X1 U6645 ( .A(n5028), .B(n9834), .ZN(n9842) );
  MUX2_X1 U6646 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4287), .Z(n5029) );
  OR2_X1 U6647 ( .A1(n5029), .A2(n8443), .ZN(n5062) );
  XNOR2_X1 U6648 ( .A(n5029), .B(n5403), .ZN(n8439) );
  MUX2_X1 U6649 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5675), .Z(n5030) );
  OR2_X1 U6650 ( .A1(n5030), .A2(n8425), .ZN(n5061) );
  XNOR2_X1 U6651 ( .A(n5030), .B(n5383), .ZN(n8421) );
  MUX2_X1 U6652 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4287), .Z(n5031) );
  OR2_X1 U6653 ( .A1(n5031), .A2(n8408), .ZN(n5060) );
  XNOR2_X1 U6654 ( .A(n5031), .B(n5368), .ZN(n8404) );
  MUX2_X1 U6655 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n5675), .Z(n5058) );
  OR2_X1 U6656 ( .A1(n5058), .A2(n8394), .ZN(n5059) );
  INV_X1 U6657 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5315) );
  MUX2_X1 U6658 ( .A(n5315), .B(n9952), .S(n5675), .Z(n5053) );
  NAND2_X1 U6659 ( .A1(n5053), .A2(n7476), .ZN(n5052) );
  INV_X1 U6660 ( .A(n5052), .ZN(n5054) );
  INV_X1 U6661 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7404) );
  INV_X1 U6662 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U6663 ( .A(n7404), .B(n9950), .S(n4287), .Z(n5050) );
  INV_X1 U6664 ( .A(n6568), .ZN(n7384) );
  NAND2_X1 U6665 ( .A1(n5050), .A2(n7384), .ZN(n5049) );
  INV_X1 U6666 ( .A(n5049), .ZN(n5051) );
  MUX2_X1 U6667 ( .A(n9813), .B(n9948), .S(n5675), .Z(n5047) );
  NAND2_X1 U6668 ( .A1(n5047), .A2(n9816), .ZN(n5046) );
  INV_X1 U6669 ( .A(n5046), .ZN(n5048) );
  MUX2_X1 U6670 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n4287), .Z(n5044) );
  INV_X1 U6671 ( .A(n5044), .ZN(n5045) );
  INV_X1 U6672 ( .A(n6520), .ZN(n6688) );
  MUX2_X1 U6673 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4287), .Z(n5036) );
  INV_X1 U6674 ( .A(n5036), .ZN(n5037) );
  MUX2_X1 U6675 ( .A(n6642), .B(n6921), .S(n5675), .Z(n5032) );
  INV_X1 U6676 ( .A(n6523), .ZN(n6650) );
  XNOR2_X1 U6677 ( .A(n5032), .B(n6650), .ZN(n6636) );
  MUX2_X1 U6678 ( .A(n6822), .B(n5116), .S(n4287), .Z(n6574) );
  NAND2_X1 U6679 ( .A1(n6574), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6573) );
  INV_X1 U6680 ( .A(n6573), .ZN(n6635) );
  OAI22_X1 U6681 ( .A1(n6636), .A2(n6635), .B1(n6650), .B2(n5032), .ZN(n9787)
         );
  MUX2_X1 U6682 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4287), .Z(n5033) );
  XNOR2_X1 U6683 ( .A(n5033), .B(n9771), .ZN(n9788) );
  INV_X1 U6684 ( .A(n9771), .ZN(n6512) );
  AOI22_X1 U6685 ( .A1(n9787), .A2(n9788), .B1(n5033), .B2(n6512), .ZN(n6694)
         );
  MUX2_X1 U6686 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5675), .Z(n5034) );
  XNOR2_X1 U6687 ( .A(n5034), .B(n5157), .ZN(n6693) );
  NAND2_X1 U6688 ( .A1(n6694), .A2(n6693), .ZN(n6692) );
  INV_X1 U6689 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6690 ( .A1(n5035), .A2(n5157), .ZN(n6669) );
  XNOR2_X1 U6691 ( .A(n5036), .B(n6688), .ZN(n6668) );
  NAND3_X1 U6692 ( .A1(n6692), .A2(n6669), .A3(n6668), .ZN(n6667) );
  OAI21_X1 U6693 ( .B1(n6688), .B2(n5037), .A(n6667), .ZN(n6498) );
  MUX2_X1 U6694 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n5675), .Z(n5038) );
  XNOR2_X1 U6695 ( .A(n5038), .B(n5207), .ZN(n6497) );
  AOI22_X1 U6696 ( .A1(n6498), .A2(n6497), .B1(n5038), .B2(n6527), .ZN(n6721)
         );
  MUX2_X1 U6697 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4287), .Z(n5039) );
  INV_X1 U6698 ( .A(n6531), .ZN(n6738) );
  XNOR2_X1 U6699 ( .A(n5039), .B(n6738), .ZN(n6722) );
  INV_X1 U6700 ( .A(n5039), .ZN(n5040) );
  AOI22_X1 U6701 ( .A1(n6721), .A2(n6722), .B1(n6738), .B2(n5040), .ZN(n9800)
         );
  INV_X1 U6702 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5240) );
  MUX2_X1 U6703 ( .A(n9793), .B(n5240), .S(n5675), .Z(n5041) );
  NAND2_X1 U6704 ( .A1(n5041), .A2(n5249), .ZN(n5042) );
  OAI21_X1 U6705 ( .B1(n5041), .B2(n5249), .A(n5042), .ZN(n9799) );
  NOR2_X1 U6706 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  INV_X1 U6707 ( .A(n5042), .ZN(n5043) );
  NOR2_X1 U6708 ( .A1(n9798), .A2(n5043), .ZN(n6870) );
  XOR2_X1 U6709 ( .A(n6882), .B(n5044), .Z(n6869) );
  NOR2_X1 U6710 ( .A1(n6870), .A2(n6869), .ZN(n6868) );
  AOI21_X1 U6711 ( .B1(n6882), .B2(n5045), .A(n6868), .ZN(n9825) );
  OAI21_X1 U6712 ( .B1(n5047), .B2(n9816), .A(n5046), .ZN(n9824) );
  NOR2_X1 U6713 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  NOR2_X1 U6714 ( .A1(n5048), .A2(n9823), .ZN(n7372) );
  OAI21_X1 U6715 ( .B1(n5050), .B2(n7384), .A(n5049), .ZN(n7373) );
  NOR2_X1 U6716 ( .A1(n7372), .A2(n7373), .ZN(n7371) );
  NOR2_X1 U6717 ( .A1(n5051), .A2(n7371), .ZN(n7466) );
  OAI21_X1 U6718 ( .B1(n5053), .B2(n7476), .A(n5052), .ZN(n7467) );
  NOR2_X1 U6719 ( .A1(n7466), .A2(n7467), .ZN(n7465) );
  NOR2_X1 U6720 ( .A1(n5054), .A2(n7465), .ZN(n7424) );
  MUX2_X1 U6721 ( .A(n4990), .B(n10079), .S(n4287), .Z(n5055) );
  NAND2_X1 U6722 ( .A1(n5055), .A2(n7420), .ZN(n7421) );
  INV_X1 U6723 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6724 ( .A1(n5056), .A2(n6626), .ZN(n7422) );
  INV_X1 U6725 ( .A(n7422), .ZN(n5057) );
  AOI21_X1 U6726 ( .B1(n7424), .B2(n7421), .A(n5057), .ZN(n8387) );
  XNOR2_X1 U6727 ( .A(n5058), .B(n5352), .ZN(n8386) );
  NAND2_X1 U6728 ( .A1(n8387), .A2(n8386), .ZN(n8385) );
  NAND2_X1 U6729 ( .A1(n5059), .A2(n8385), .ZN(n8403) );
  NAND2_X1 U6730 ( .A1(n8404), .A2(n8403), .ZN(n8402) );
  NAND2_X1 U6731 ( .A1(n5060), .A2(n8402), .ZN(n8420) );
  NAND2_X1 U6732 ( .A1(n8421), .A2(n8420), .ZN(n8419) );
  NAND2_X1 U6733 ( .A1(n5061), .A2(n8419), .ZN(n8438) );
  NAND2_X1 U6734 ( .A1(n8439), .A2(n8438), .ZN(n8437) );
  NAND2_X1 U6735 ( .A1(n5062), .A2(n8437), .ZN(n9841) );
  NAND2_X1 U6736 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  NAND2_X1 U6737 ( .A1(n5063), .A2(n9840), .ZN(n5064) );
  INV_X1 U6738 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8609) );
  INV_X1 U6739 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5442) );
  MUX2_X1 U6740 ( .A(n8609), .B(n5442), .S(n4287), .Z(n5065) );
  AND2_X1 U6741 ( .A1(n5064), .A2(n5065), .ZN(n8462) );
  INV_X1 U6742 ( .A(n8462), .ZN(n5068) );
  INV_X1 U6743 ( .A(n5064), .ZN(n5067) );
  INV_X1 U6744 ( .A(n5065), .ZN(n5066) );
  NAND2_X1 U6745 ( .A1(n5067), .A2(n5066), .ZN(n8460) );
  NAND2_X1 U6746 ( .A1(n5068), .A2(n8460), .ZN(n5076) );
  INV_X1 U6747 ( .A(n6562), .ZN(n6754) );
  INV_X1 U6748 ( .A(n5002), .ZN(n5676) );
  NAND3_X1 U6749 ( .A1(n5076), .A2(n9843), .A3(n7163), .ZN(n5073) );
  INV_X1 U6750 ( .A(n7090), .ZN(n5069) );
  NOR2_X1 U6751 ( .A1(n5721), .A2(n5069), .ZN(n5070) );
  OR2_X1 U6752 ( .A1(P2_U3150), .A2(n5070), .ZN(n9832) );
  INV_X1 U6753 ( .A(n9832), .ZN(n9797) );
  INV_X1 U6754 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8335) );
  NOR2_X1 U6755 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8335), .ZN(n5071) );
  AOI21_X1 U6756 ( .B1(n9797), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n5071), .ZN(
        n5072) );
  NAND2_X1 U6757 ( .A1(n5073), .A2(n5072), .ZN(n5079) );
  NOR2_X1 U6758 ( .A1(n4287), .A2(P2_U3151), .ZN(n7608) );
  NAND2_X1 U6759 ( .A1(n5074), .A2(n7608), .ZN(n5075) );
  MUX2_X1 U6760 ( .A(n8381), .B(n5075), .S(n5002), .Z(n9835) );
  OAI21_X1 U6761 ( .B1(n5076), .B2(n8381), .A(n9835), .ZN(n5077) );
  NAND2_X1 U6762 ( .A1(n4345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6763 ( .A1(n5085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6764 ( .A1(n5091), .A2(n5092), .ZN(n8814) );
  INV_X1 U6765 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5090) );
  INV_X1 U6766 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6900) );
  OR2_X1 U6767 ( .A1(n5177), .A2(n6900), .ZN(n5101) );
  OR2_X1 U6768 ( .A1(n5179), .A2(n6921), .ZN(n5099) );
  INV_X1 U6769 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6770 ( .A1(n7076), .A2(n5102), .ZN(n5105) );
  AND2_X2 U6771 ( .A1(n5128), .A2(n6514), .ZN(n5155) );
  NAND2_X1 U6772 ( .A1(n5155), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6773 ( .A(n5131), .B(SI_1_), .ZN(n5111) );
  OAI21_X1 U6774 ( .B1(n5138), .B2(n5109), .A(n5108), .ZN(n5110) );
  NAND2_X1 U6775 ( .A1(n5110), .A2(SI_0_), .ZN(n5129) );
  XNOR2_X1 U6776 ( .A(n5111), .B(n5129), .ZN(n6522) );
  NAND2_X1 U6777 ( .A1(n4330), .A2(n5685), .ZN(n5113) );
  INV_X1 U6778 ( .A(n5128), .ZN(n5127) );
  NAND2_X1 U6779 ( .A1(n5127), .A2(n6650), .ZN(n5112) );
  INV_X1 U6780 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6768) );
  OR2_X1 U6781 ( .A1(n5177), .A2(n6768), .ZN(n5120) );
  INV_X1 U6782 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5115) );
  OR2_X1 U6783 ( .A1(n5179), .A2(n5116), .ZN(n5117) );
  NAND4_X2 U6784 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n7098)
         );
  NAND2_X1 U6785 ( .A1(n5774), .A2(SI_0_), .ZN(n5121) );
  XNOR2_X1 U6786 ( .A(n5121), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U6787 ( .A1(n7101), .A2(n7099), .ZN(n7969) );
  OR2_X1 U6788 ( .A1(n7134), .A2(n9880), .ZN(n5126) );
  INV_X1 U6789 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6790 ( .A1(n4284), .A2(n5122), .ZN(n5125) );
  INV_X1 U6791 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7620) );
  OR2_X1 U6792 ( .A1(n5177), .A2(n7620), .ZN(n5124) );
  OR2_X1 U6793 ( .A1(n4290), .A2(n9937), .ZN(n5123) );
  NAND4_X4 U6794 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n8380)
         );
  NAND2_X1 U6795 ( .A1(n5155), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6796 ( .A1(n5131), .A2(SI_1_), .ZN(n5130) );
  NAND2_X1 U6797 ( .A1(n5130), .A2(n5129), .ZN(n5135) );
  INV_X1 U6798 ( .A(n5131), .ZN(n5133) );
  INV_X1 U6799 ( .A(SI_1_), .ZN(n5132) );
  NAND2_X1 U6800 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  INV_X1 U6801 ( .A(n5145), .ZN(n5144) );
  NAND2_X1 U6802 ( .A1(n5139), .A2(SI_2_), .ZN(n5159) );
  INV_X1 U6803 ( .A(n5139), .ZN(n5141) );
  INV_X1 U6804 ( .A(SI_2_), .ZN(n5140) );
  NAND2_X1 U6805 ( .A1(n5141), .A2(n5140), .ZN(n5142) );
  NAND2_X1 U6806 ( .A1(n5159), .A2(n5142), .ZN(n5146) );
  NAND2_X1 U6807 ( .A1(n5145), .A2(n5146), .ZN(n5147) );
  NAND2_X1 U6808 ( .A1(n5160), .A2(n5147), .ZN(n6515) );
  OR2_X1 U6809 ( .A1(n8380), .A2(n9871), .ZN(n7974) );
  INV_X4 U6810 ( .A(n4284), .ZN(n5678) );
  NAND2_X1 U6811 ( .A1(n5678), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5154) );
  OR2_X1 U6812 ( .A1(n5175), .A2(n6701), .ZN(n5153) );
  OR2_X1 U6813 ( .A1(n5177), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5152) );
  OR2_X1 U6814 ( .A1(n4290), .A2(n9939), .ZN(n5151) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6816 ( .A1(n5206), .A2(n5156), .ZN(n5173) );
  NAND2_X1 U6817 ( .A1(n4289), .A2(n5157), .ZN(n5172) );
  INV_X1 U6818 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5161) );
  INV_X1 U6819 ( .A(n5164), .ZN(n5163) );
  INV_X1 U6820 ( .A(SI_3_), .ZN(n5162) );
  NAND2_X1 U6821 ( .A1(n5165), .A2(n5184), .ZN(n5167) );
  NAND2_X1 U6822 ( .A1(n5166), .A2(n5167), .ZN(n5170) );
  INV_X1 U6823 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6824 ( .A1(n5170), .A2(n5185), .ZN(n6518) );
  OR2_X1 U6825 ( .A1(n5158), .A2(n6518), .ZN(n5171) );
  NAND2_X1 U6826 ( .A1(n9861), .A2(n8215), .ZN(n7983) );
  NAND2_X1 U6827 ( .A1(n7991), .A2(n7983), .ZN(n5633) );
  INV_X1 U6828 ( .A(n5633), .ZN(n7936) );
  NAND2_X1 U6829 ( .A1(n7004), .A2(n7936), .ZN(n5174) );
  NAND2_X1 U6830 ( .A1(n5174), .A2(n7991), .ZN(n7081) );
  INV_X2 U6831 ( .A(n7134), .ZN(n5219) );
  INV_X1 U6832 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6833 ( .A1(n4284), .A2(n5176), .ZN(n5182) );
  NAND2_X1 U6834 ( .A1(n6699), .A2(n6676), .ZN(n5200) );
  NAND2_X1 U6835 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5178) );
  AND2_X1 U6836 ( .A1(n5200), .A2(n5178), .ZN(n7086) );
  OR2_X1 U6837 ( .A1(n5438), .A2(n7086), .ZN(n5181) );
  OR2_X1 U6838 ( .A1(n4290), .A2(n9941), .ZN(n5180) );
  NAND2_X1 U6839 ( .A1(n7915), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6840 ( .A1(n4289), .A2(n6688), .ZN(n5196) );
  MUX2_X1 U6841 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5325), .Z(n5186) );
  NAND2_X1 U6842 ( .A1(n5186), .A2(SI_4_), .ZN(n5208) );
  INV_X1 U6843 ( .A(n5186), .ZN(n5188) );
  INV_X1 U6844 ( .A(SI_4_), .ZN(n5187) );
  NAND2_X1 U6845 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  NAND2_X1 U6846 ( .A1(n5208), .A2(n5189), .ZN(n5191) );
  NAND2_X1 U6847 ( .A1(n5190), .A2(n5191), .ZN(n5194) );
  INV_X1 U6848 ( .A(n5191), .ZN(n5192) );
  NAND2_X1 U6849 ( .A1(n5193), .A2(n5192), .ZN(n5209) );
  NAND2_X1 U6850 ( .A1(n5194), .A2(n5209), .ZN(n6519) );
  OR2_X1 U6851 ( .A1(n5158), .A2(n6519), .ZN(n5195) );
  OR2_X1 U6852 ( .A1(n7143), .A2(n8204), .ZN(n7984) );
  NAND2_X1 U6853 ( .A1(n7143), .A2(n8204), .ZN(n7992) );
  INV_X1 U6854 ( .A(n7933), .ZN(n7981) );
  NAND2_X1 U6855 ( .A1(n7081), .A2(n7981), .ZN(n7080) );
  NAND2_X1 U6856 ( .A1(n7080), .A2(n7984), .ZN(n7142) );
  NAND2_X1 U6857 ( .A1(n5678), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6858 ( .A1(n7134), .A2(n6500), .ZN(n5204) );
  INV_X1 U6859 ( .A(n5200), .ZN(n5199) );
  NAND2_X1 U6860 ( .A1(n5199), .A2(n5198), .ZN(n5221) );
  NAND2_X1 U6861 ( .A1(n5200), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5201) );
  AND2_X1 U6862 ( .A1(n5221), .A2(n5201), .ZN(n7148) );
  OR2_X1 U6863 ( .A1(n5438), .A2(n7148), .ZN(n5203) );
  OR2_X1 U6864 ( .A1(n4290), .A2(n9943), .ZN(n5202) );
  NAND4_X1 U6865 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n8379)
         );
  INV_X1 U6866 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U6867 ( .A1(n4289), .A2(n5207), .ZN(n5218) );
  NAND2_X1 U6868 ( .A1(n5209), .A2(n5208), .ZN(n5215) );
  NAND2_X1 U6869 ( .A1(n5211), .A2(SI_5_), .ZN(n5228) );
  INV_X1 U6870 ( .A(n5211), .ZN(n5212) );
  INV_X1 U6871 ( .A(SI_5_), .ZN(n10081) );
  NAND2_X1 U6872 ( .A1(n5212), .A2(n10081), .ZN(n5213) );
  NAND2_X1 U6873 ( .A1(n5215), .A2(n5214), .ZN(n5229) );
  OR2_X1 U6874 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  NAND2_X1 U6875 ( .A1(n5229), .A2(n5216), .ZN(n6526) );
  OR2_X1 U6876 ( .A1(n5158), .A2(n6526), .ZN(n5217) );
  OAI211_X1 U6877 ( .C1(n5206), .C2(n6528), .A(n5218), .B(n5217), .ZN(n5638)
         );
  NAND2_X1 U6878 ( .A1(n8379), .A2(n9895), .ZN(n7993) );
  NAND2_X1 U6879 ( .A1(n7142), .A2(n7993), .ZN(n7209) );
  NAND2_X1 U6880 ( .A1(n5219), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5227) );
  INV_X1 U6881 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6882 ( .A1(n4284), .A2(n5220), .ZN(n5226) );
  NAND2_X1 U6883 ( .A1(n5221), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5222) );
  AND2_X1 U6884 ( .A1(n5243), .A2(n5222), .ZN(n7251) );
  OR2_X1 U6885 ( .A1(n5438), .A2(n7251), .ZN(n5225) );
  INV_X1 U6886 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5223) );
  OR2_X1 U6887 ( .A1(n4290), .A2(n5223), .ZN(n5224) );
  NAND4_X1 U6888 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n8378)
         );
  NAND2_X1 U6889 ( .A1(n7915), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6890 ( .A1(n4289), .A2(n6738), .ZN(n5237) );
  NAND2_X1 U6891 ( .A1(n5229), .A2(n5228), .ZN(n5234) );
  MUX2_X1 U6892 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6514), .Z(n5230) );
  NAND2_X1 U6893 ( .A1(n5230), .A2(SI_6_), .ZN(n5250) );
  INV_X1 U6894 ( .A(n5230), .ZN(n5231) );
  INV_X1 U6895 ( .A(SI_6_), .ZN(n10049) );
  NAND2_X1 U6896 ( .A1(n5231), .A2(n10049), .ZN(n5232) );
  NAND2_X1 U6897 ( .A1(n5234), .A2(n5233), .ZN(n5251) );
  OR2_X1 U6898 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6899 ( .A1(n5251), .A2(n5235), .ZN(n6530) );
  OR2_X1 U6900 ( .A1(n5158), .A2(n6530), .ZN(n5236) );
  OR2_X1 U6901 ( .A1(n8378), .A2(n7246), .ZN(n7987) );
  OR2_X1 U6902 ( .A1(n8379), .A2(n9895), .ZN(n7985) );
  NAND2_X1 U6903 ( .A1(n7209), .A2(n4871), .ZN(n5239) );
  NAND2_X1 U6904 ( .A1(n8378), .A2(n7246), .ZN(n7996) );
  NAND2_X1 U6905 ( .A1(n5239), .A2(n7996), .ZN(n7220) );
  NAND2_X1 U6906 ( .A1(n5678), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5248) );
  OR2_X1 U6907 ( .A1(n4290), .A2(n5240), .ZN(n5247) );
  NAND2_X1 U6908 ( .A1(n5242), .A2(n5241), .ZN(n5262) );
  NAND2_X1 U6909 ( .A1(n5243), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5244) );
  AND2_X1 U6910 ( .A1(n5262), .A2(n5244), .ZN(n7265) );
  OR2_X1 U6911 ( .A1(n5438), .A2(n7265), .ZN(n5246) );
  OR2_X1 U6912 ( .A1(n7134), .A2(n9793), .ZN(n5245) );
  NAND4_X1 U6913 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n8377)
         );
  NAND2_X1 U6914 ( .A1(n4289), .A2(n5249), .ZN(n5260) );
  NAND2_X1 U6915 ( .A1(n5252), .A2(SI_7_), .ZN(n5269) );
  INV_X1 U6916 ( .A(n5252), .ZN(n5254) );
  INV_X1 U6917 ( .A(SI_7_), .ZN(n5253) );
  NAND2_X1 U6918 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  OR2_X1 U6919 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6920 ( .A1(n5270), .A2(n5258), .ZN(n6533) );
  OR2_X1 U6921 ( .A1(n5158), .A2(n6533), .ZN(n5259) );
  NAND2_X1 U6922 ( .A1(n8377), .A2(n9905), .ZN(n7311) );
  NAND2_X1 U6923 ( .A1(n7220), .A2(n8004), .ZN(n7219) );
  NAND2_X1 U6924 ( .A1(n5219), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5268) );
  INV_X1 U6925 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5261) );
  OR2_X1 U6926 ( .A1(n4284), .A2(n5261), .ZN(n5267) );
  NAND2_X1 U6927 ( .A1(n5262), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5263) );
  AND2_X1 U6928 ( .A1(n5285), .A2(n5263), .ZN(n7331) );
  OR2_X1 U6929 ( .A1(n5438), .A2(n7331), .ZN(n5266) );
  OR2_X1 U6930 ( .A1(n4290), .A2(n5264), .ZN(n5265) );
  NAND4_X1 U6931 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8376)
         );
  MUX2_X1 U6932 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6514), .Z(n5274) );
  XNOR2_X1 U6933 ( .A(n5274), .B(SI_8_), .ZN(n5278) );
  NAND2_X1 U6934 ( .A1(n6543), .A2(n7914), .ZN(n5272) );
  AOI22_X1 U6935 ( .A1(n7915), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4289), .B2(
        n6882), .ZN(n5271) );
  NAND2_X1 U6936 ( .A1(n8376), .A2(n9910), .ZN(n8001) );
  AND2_X1 U6937 ( .A1(n7311), .A2(n8001), .ZN(n8009) );
  NAND2_X1 U6938 ( .A1(n7219), .A2(n8009), .ZN(n5273) );
  NAND2_X1 U6939 ( .A1(n5273), .A2(n8011), .ZN(n7345) );
  INV_X1 U6940 ( .A(n5274), .ZN(n5276) );
  INV_X1 U6941 ( .A(SI_8_), .ZN(n5275) );
  NAND2_X1 U6942 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5280) );
  MUX2_X1 U6944 ( .A(n5280), .B(n10109), .S(n6514), .Z(n5291) );
  XNOR2_X1 U6945 ( .A(n5291), .B(SI_9_), .ZN(n5294) );
  XNOR2_X1 U6946 ( .A(n5295), .B(n5294), .ZN(n6563) );
  NAND2_X1 U6947 ( .A1(n6563), .A2(n7914), .ZN(n5282) );
  AOI22_X1 U6948 ( .A1(n7915), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4289), .B2(
        n9816), .ZN(n5281) );
  NAND2_X1 U6949 ( .A1(n5678), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5290) );
  OR2_X1 U6950 ( .A1(n4290), .A2(n9948), .ZN(n5289) );
  NAND2_X1 U6951 ( .A1(n5285), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5286) );
  AND2_X1 U6952 ( .A1(n5305), .A2(n5286), .ZN(n7361) );
  OR2_X1 U6953 ( .A1(n5438), .A2(n7361), .ZN(n5288) );
  OR2_X1 U6954 ( .A1(n7134), .A2(n9813), .ZN(n5287) );
  NAND4_X1 U6955 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n8375)
         );
  NAND2_X1 U6956 ( .A1(n9919), .A2(n7487), .ZN(n8012) );
  NAND2_X1 U6957 ( .A1(n8008), .A2(n8012), .ZN(n7943) );
  INV_X1 U6958 ( .A(n5291), .ZN(n5292) );
  NOR2_X1 U6959 ( .A1(n5292), .A2(SI_9_), .ZN(n5293) );
  MUX2_X1 U6960 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6514), .Z(n5296) );
  NAND2_X1 U6961 ( .A1(n5296), .A2(SI_10_), .ZN(n5311) );
  INV_X1 U6962 ( .A(n5296), .ZN(n5298) );
  INV_X1 U6963 ( .A(SI_10_), .ZN(n5297) );
  NAND2_X1 U6964 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6965 ( .A1(n5312), .A2(n5302), .ZN(n6570) );
  AOI22_X1 U6966 ( .A1(n7915), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4289), .B2(
        n7384), .ZN(n5303) );
  INV_X1 U6967 ( .A(n7496), .ZN(n9922) );
  NAND2_X1 U6968 ( .A1(n5678), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5310) );
  OR2_X1 U6969 ( .A1(n4290), .A2(n9950), .ZN(n5309) );
  NAND2_X1 U6970 ( .A1(n5305), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5306) );
  AND2_X1 U6971 ( .A1(n5316), .A2(n5306), .ZN(n7493) );
  OR2_X1 U6972 ( .A1(n5438), .A2(n7493), .ZN(n5308) );
  OR2_X1 U6973 ( .A1(n7134), .A2(n7404), .ZN(n5307) );
  NAND4_X1 U6974 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n8374)
         );
  INV_X1 U6975 ( .A(n8374), .ZN(n7553) );
  NAND2_X1 U6976 ( .A1(n7496), .A2(n7553), .ZN(n8023) );
  MUX2_X1 U6977 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6514), .Z(n5322) );
  XNOR2_X1 U6978 ( .A(n5322), .B(SI_11_), .ZN(n5323) );
  XNOR2_X1 U6979 ( .A(n5324), .B(n5323), .ZN(n6580) );
  NAND2_X1 U6980 ( .A1(n6580), .A2(n7914), .ZN(n5314) );
  AOI22_X1 U6981 ( .A1(n7915), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4289), .B2(
        n7476), .ZN(n5313) );
  NAND2_X1 U6982 ( .A1(n5314), .A2(n5313), .ZN(n7507) );
  NAND2_X1 U6983 ( .A1(n5678), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6984 ( .A1(n7134), .A2(n5315), .ZN(n5320) );
  NAND2_X1 U6985 ( .A1(n5316), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5317) );
  AND2_X1 U6986 ( .A1(n5336), .A2(n5317), .ZN(n7445) );
  OR2_X1 U6987 ( .A1(n5438), .A2(n7445), .ZN(n5319) );
  OR2_X1 U6988 ( .A1(n4290), .A2(n9952), .ZN(n5318) );
  OR2_X1 U6989 ( .A1(n7507), .A2(n7556), .ZN(n8026) );
  NAND2_X1 U6990 ( .A1(n7507), .A2(n7556), .ZN(n8021) );
  NAND2_X1 U6991 ( .A1(n8026), .A2(n8021), .ZN(n7944) );
  INV_X1 U6992 ( .A(n7944), .ZN(n7555) );
  NAND2_X1 U6993 ( .A1(n7444), .A2(n7555), .ZN(n7443) );
  MUX2_X1 U6994 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6513), .Z(n5326) );
  NAND2_X1 U6995 ( .A1(n5326), .A2(SI_12_), .ZN(n5343) );
  INV_X1 U6996 ( .A(n5326), .ZN(n5328) );
  INV_X1 U6997 ( .A(SI_12_), .ZN(n5327) );
  NAND2_X1 U6998 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  NAND2_X1 U6999 ( .A1(n5343), .A2(n5329), .ZN(n5330) );
  NAND2_X1 U7000 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  NAND2_X1 U7001 ( .A1(n5332), .A2(n5344), .ZN(n6628) );
  OR2_X1 U7002 ( .A1(n6628), .A2(n5158), .ZN(n5334) );
  AOI22_X1 U7003 ( .A1(n7915), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4289), .B2(
        n7420), .ZN(n5333) );
  NAND2_X1 U7004 ( .A1(n5219), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5341) );
  INV_X1 U7005 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7517) );
  OR2_X1 U7006 ( .A1(n4284), .A2(n7517), .ZN(n5340) );
  NAND2_X1 U7007 ( .A1(n5336), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5337) );
  AND2_X1 U7008 ( .A1(n5357), .A2(n5337), .ZN(n7550) );
  OR2_X1 U7009 ( .A1(n5438), .A2(n7550), .ZN(n5339) );
  OR2_X1 U7010 ( .A1(n7137), .A2(n10079), .ZN(n5338) );
  NAND4_X1 U7011 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n8372)
         );
  NAND2_X1 U7012 ( .A1(n7568), .A2(n7563), .ZN(n8030) );
  NAND2_X1 U7013 ( .A1(n8031), .A2(n8030), .ZN(n8034) );
  INV_X1 U7014 ( .A(n8021), .ZN(n8025) );
  NOR2_X1 U7015 ( .A1(n8034), .A2(n8025), .ZN(n5342) );
  NAND2_X1 U7016 ( .A1(n7443), .A2(n5342), .ZN(n7511) );
  MUX2_X1 U7017 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6514), .Z(n5345) );
  NAND2_X1 U7018 ( .A1(n5345), .A2(SI_13_), .ZN(n5365) );
  INV_X1 U7019 ( .A(n5345), .ZN(n5347) );
  INV_X1 U7020 ( .A(SI_13_), .ZN(n5346) );
  NAND2_X1 U7021 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  OR2_X1 U7022 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  AND2_X1 U7023 ( .A1(n5366), .A2(n5351), .ZN(n6711) );
  NAND2_X1 U7024 ( .A1(n6711), .A2(n7914), .ZN(n5354) );
  AOI22_X1 U7025 ( .A1(n5155), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4289), .B2(
        n5352), .ZN(n5353) );
  NAND2_X1 U7026 ( .A1(n5678), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5362) );
  OR2_X1 U7027 ( .A1(n7134), .A2(n8384), .ZN(n5361) );
  NAND2_X1 U7028 ( .A1(n5357), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5358) );
  AND2_X1 U7029 ( .A1(n5371), .A2(n5358), .ZN(n7593) );
  OR2_X1 U7030 ( .A1(n5438), .A2(n7593), .ZN(n5360) );
  OR2_X1 U7031 ( .A1(n7137), .A2(n10050), .ZN(n5359) );
  NAND4_X1 U7032 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n8371)
         );
  INV_X1 U7033 ( .A(n8371), .ZN(n7547) );
  NOR2_X1 U7034 ( .A1(n7589), .A2(n7547), .ZN(n8038) );
  INV_X1 U7035 ( .A(n8038), .ZN(n5363) );
  AND2_X1 U7036 ( .A1(n5363), .A2(n8031), .ZN(n5364) );
  NAND2_X1 U7037 ( .A1(n7589), .A2(n7547), .ZN(n8036) );
  MUX2_X1 U7038 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6514), .Z(n5380) );
  XNOR2_X1 U7039 ( .A(n5380), .B(SI_14_), .ZN(n5367) );
  XNOR2_X1 U7040 ( .A(n5381), .B(n5367), .ZN(n6769) );
  NAND2_X1 U7041 ( .A1(n6769), .A2(n7914), .ZN(n5370) );
  AOI22_X1 U7042 ( .A1(n5155), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4289), .B2(
        n5368), .ZN(n5369) );
  NAND2_X1 U7043 ( .A1(n5678), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5377) );
  OR2_X1 U7044 ( .A1(n7134), .A2(n7585), .ZN(n5376) );
  NAND2_X1 U7045 ( .A1(n5371), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5372) );
  AND2_X1 U7046 ( .A1(n5388), .A2(n5372), .ZN(n8238) );
  OR2_X1 U7047 ( .A1(n5438), .A2(n8238), .ZN(n5375) );
  OR2_X1 U7048 ( .A1(n7137), .A2(n5373), .ZN(n5374) );
  NAND4_X1 U7049 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n8655)
         );
  XNOR2_X1 U7050 ( .A(n8240), .B(n8153), .ZN(n8040) );
  OR2_X1 U7051 ( .A1(n8240), .A2(n8153), .ZN(n5379) );
  NAND2_X1 U7052 ( .A1(n7581), .A2(n5379), .ZN(n8645) );
  MUX2_X1 U7053 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6513), .Z(n5395) );
  XNOR2_X1 U7054 ( .A(n5395), .B(SI_15_), .ZN(n5382) );
  XNOR2_X1 U7055 ( .A(n5398), .B(n5382), .ZN(n6824) );
  NAND2_X1 U7056 ( .A1(n6824), .A2(n7914), .ZN(n5385) );
  AOI22_X1 U7057 ( .A1(n7915), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4289), .B2(
        n5383), .ZN(n5384) );
  NAND2_X1 U7058 ( .A1(n5678), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5393) );
  OR2_X1 U7059 ( .A1(n7134), .A2(n8656), .ZN(n5392) );
  NAND2_X1 U7060 ( .A1(n5388), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5389) );
  AND2_X1 U7061 ( .A1(n5406), .A2(n5389), .ZN(n8357) );
  OR2_X1 U7062 ( .A1(n5438), .A2(n8357), .ZN(n5391) );
  OR2_X1 U7063 ( .A1(n7137), .A2(n8713), .ZN(n5390) );
  INV_X1 U7064 ( .A(n8048), .ZN(n5394) );
  NAND2_X1 U7065 ( .A1(n8805), .A2(n8634), .ZN(n8059) );
  INV_X1 U7066 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U7067 ( .A1(n5397), .A2(n5396), .ZN(n5401) );
  NAND2_X1 U7068 ( .A1(n5399), .A2(n4719), .ZN(n5400) );
  NAND2_X1 U7069 ( .A1(n5401), .A2(n5400), .ZN(n5413) );
  MUX2_X1 U7070 ( .A(n6893), .B(n10111), .S(n6513), .Z(n5414) );
  XNOR2_X1 U7071 ( .A(n5414), .B(SI_16_), .ZN(n5402) );
  XNOR2_X1 U7072 ( .A(n5413), .B(n5402), .ZN(n6892) );
  NAND2_X1 U7073 ( .A1(n6892), .A2(n7914), .ZN(n5405) );
  AOI22_X1 U7074 ( .A1(n7915), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4289), .B2(
        n5403), .ZN(n5404) );
  NAND2_X1 U7075 ( .A1(n5678), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5411) );
  OR2_X1 U7076 ( .A1(n7134), .A2(n8639), .ZN(n5410) );
  NAND2_X1 U7077 ( .A1(n5406), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5407) );
  AND2_X1 U7078 ( .A1(n5427), .A2(n5407), .ZN(n8640) );
  OR2_X1 U7079 ( .A1(n5438), .A2(n8640), .ZN(n5409) );
  OR2_X1 U7080 ( .A1(n7137), .A2(n8710), .ZN(n5408) );
  NAND2_X1 U7081 ( .A1(n8799), .A2(n8647), .ZN(n8058) );
  INV_X1 U7082 ( .A(n8058), .ZN(n5412) );
  INV_X1 U7083 ( .A(n5413), .ZN(n5415) );
  NAND2_X1 U7084 ( .A1(n5415), .A2(n4882), .ZN(n5418) );
  NAND2_X1 U7085 ( .A1(n5416), .A2(SI_16_), .ZN(n5417) );
  MUX2_X1 U7086 ( .A(n10035), .B(n7009), .S(n6514), .Z(n5420) );
  INV_X1 U7087 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U7088 ( .A1(n5421), .A2(SI_17_), .ZN(n5422) );
  NAND2_X1 U7089 ( .A1(n5435), .A2(n5422), .ZN(n5434) );
  XNOR2_X1 U7090 ( .A(n5433), .B(n5434), .ZN(n7007) );
  NAND2_X1 U7091 ( .A1(n7007), .A2(n7914), .ZN(n5425) );
  AOI22_X1 U7092 ( .A1(n5155), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4289), .B2(
        n5423), .ZN(n5424) );
  NAND2_X1 U7093 ( .A1(n5678), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5432) );
  OR2_X1 U7094 ( .A1(n7134), .A2(n9847), .ZN(n5431) );
  NAND2_X1 U7095 ( .A1(n5427), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5428) );
  AND2_X1 U7096 ( .A1(n5439), .A2(n5428), .ZN(n8293) );
  OR2_X1 U7097 ( .A1(n5438), .A2(n8293), .ZN(n5430) );
  OR2_X1 U7098 ( .A1(n7137), .A2(n9839), .ZN(n5429) );
  OR2_X1 U7099 ( .A1(n8793), .A2(n8635), .ZN(n7929) );
  NAND2_X1 U7100 ( .A1(n8793), .A2(n8635), .ZN(n7930) );
  NAND2_X1 U7101 ( .A1(n7929), .A2(n7930), .ZN(n8618) );
  MUX2_X1 U7102 ( .A(n7162), .B(n7165), .S(n6513), .Z(n5448) );
  XNOR2_X1 U7103 ( .A(n5448), .B(SI_18_), .ZN(n5447) );
  XNOR2_X1 U7104 ( .A(n5451), .B(n5447), .ZN(n7161) );
  NAND2_X1 U7105 ( .A1(n7161), .A2(n7914), .ZN(n5437) );
  AOI22_X1 U7106 ( .A1(n5155), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4289), .B2(
        n8461), .ZN(n5436) );
  NAND2_X1 U7107 ( .A1(n5439), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U7108 ( .A1(n5459), .A2(n5440), .ZN(n8334) );
  NAND2_X1 U7109 ( .A1(n5625), .A2(n8334), .ZN(n5446) );
  INV_X1 U7110 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5441) );
  OR2_X1 U7111 ( .A1(n4284), .A2(n5441), .ZN(n5445) );
  OR2_X1 U7112 ( .A1(n7134), .A2(n8609), .ZN(n5444) );
  OR2_X1 U7113 ( .A1(n7137), .A2(n5442), .ZN(n5443) );
  NAND4_X1 U7114 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n8620)
         );
  NAND2_X1 U7115 ( .A1(n8702), .A2(n8165), .ZN(n7931) );
  NAND2_X1 U7116 ( .A1(n8053), .A2(n7931), .ZN(n8611) );
  INV_X1 U7117 ( .A(n5447), .ZN(n5450) );
  INV_X1 U7118 ( .A(n5448), .ZN(n5449) );
  MUX2_X1 U7119 ( .A(n7253), .B(n7254), .S(n6514), .Z(n5453) );
  NAND2_X1 U7120 ( .A1(n5453), .A2(n5452), .ZN(n5465) );
  INV_X1 U7121 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U7122 ( .A1(n5454), .A2(SI_19_), .ZN(n5455) );
  NAND2_X1 U7123 ( .A1(n5465), .A2(n5455), .ZN(n5466) );
  XNOR2_X1 U7124 ( .A(n5467), .B(n5466), .ZN(n7252) );
  NAND2_X1 U7125 ( .A1(n7252), .A2(n7914), .ZN(n5457) );
  AOI22_X1 U7126 ( .A1(n7915), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5673), .B2(
        n5127), .ZN(n5456) );
  NAND2_X1 U7127 ( .A1(n5459), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7128 ( .A1(n5471), .A2(n5460), .ZN(n8252) );
  NAND2_X1 U7129 ( .A1(n5625), .A2(n8252), .ZN(n5464) );
  NAND2_X1 U7130 ( .A1(n5504), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5463) );
  INV_X1 U7131 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8594) );
  OR2_X1 U7132 ( .A1(n7134), .A2(n8594), .ZN(n5462) );
  INV_X1 U7133 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10017) );
  OR2_X1 U7134 ( .A1(n4284), .A2(n10017), .ZN(n5461) );
  NAND4_X1 U7135 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n8604)
         );
  XNOR2_X1 U7136 ( .A(n8695), .B(n8336), .ZN(n5661) );
  NOR2_X1 U7137 ( .A1(n8695), .A2(n8336), .ZN(n7960) );
  INV_X1 U7138 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7282) );
  MUX2_X1 U7139 ( .A(n7282), .B(n10016), .S(n6513), .Z(n5478) );
  XNOR2_X1 U7140 ( .A(n5478), .B(SI_20_), .ZN(n5468) );
  NAND2_X1 U7141 ( .A1(n7281), .A2(n7914), .ZN(n5470) );
  NAND2_X1 U7142 ( .A1(n7915), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7143 ( .A1(n5471), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7144 ( .A1(n5486), .A2(n5472), .ZN(n8586) );
  NAND2_X1 U7145 ( .A1(n8586), .A2(n5625), .ZN(n5477) );
  INV_X1 U7146 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10123) );
  OR2_X1 U7147 ( .A1(n7134), .A2(n10123), .ZN(n5474) );
  INV_X1 U7148 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8783) );
  OR2_X1 U7149 ( .A1(n4284), .A2(n8783), .ZN(n5473) );
  AND2_X1 U7150 ( .A1(n5474), .A2(n5473), .ZN(n5476) );
  NAND2_X1 U7151 ( .A1(n5504), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7152 ( .A1(n8784), .A2(n8590), .ZN(n8073) );
  INV_X1 U7153 ( .A(n8073), .ZN(n7963) );
  MUX2_X1 U7154 ( .A(n7344), .B(n7387), .S(n6514), .Z(n5492) );
  XNOR2_X1 U7155 ( .A(n5492), .B(SI_21_), .ZN(n5481) );
  NAND2_X1 U7156 ( .A1(n7343), .A2(n7914), .ZN(n5483) );
  NAND2_X1 U7157 ( .A1(n5155), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5482) );
  INV_X1 U7158 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7159 ( .A1(n5486), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7160 ( .A1(n5502), .A2(n5487), .ZN(n8577) );
  NAND2_X1 U7161 ( .A1(n8577), .A2(n5625), .ZN(n5490) );
  AOI22_X1 U7162 ( .A1(n5219), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5678), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7163 ( .A1(n5504), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7164 ( .A1(n8778), .A2(n8315), .ZN(n8078) );
  INV_X1 U7165 ( .A(n8071), .ZN(n8080) );
  NAND2_X1 U7166 ( .A1(n5493), .A2(SI_21_), .ZN(n5494) );
  MUX2_X1 U7167 ( .A(n7452), .B(n7453), .S(n6513), .Z(n5497) );
  NAND2_X1 U7168 ( .A1(n5497), .A2(n5496), .ZN(n5509) );
  INV_X1 U7169 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U7170 ( .A1(n5498), .A2(SI_22_), .ZN(n5499) );
  NAND2_X1 U7171 ( .A1(n5509), .A2(n5499), .ZN(n5510) );
  NAND2_X1 U7172 ( .A1(n7450), .A2(n7914), .ZN(n5501) );
  NAND2_X1 U7173 ( .A1(n7915), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7174 ( .A1(n5502), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7175 ( .A1(n5519), .A2(n5503), .ZN(n8563) );
  NAND2_X1 U7176 ( .A1(n8563), .A2(n5625), .ZN(n5507) );
  AOI22_X1 U7177 ( .A1(n5219), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n5678), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7178 ( .A1(n5504), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7179 ( .A1(n8772), .A2(n8180), .ZN(n8082) );
  INV_X1 U7180 ( .A(n8082), .ZN(n5508) );
  OR2_X1 U7181 ( .A1(n8772), .A2(n8180), .ZN(n5662) );
  OAI21_X2 U7182 ( .B1(n5511), .B2(n5510), .A(n5509), .ZN(n5527) );
  INV_X1 U7183 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5512) );
  MUX2_X1 U7184 ( .A(n5512), .B(n7486), .S(n6514), .Z(n5514) );
  INV_X1 U7185 ( .A(SI_23_), .ZN(n5513) );
  NAND2_X1 U7186 ( .A1(n5514), .A2(n5513), .ZN(n5528) );
  INV_X1 U7187 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U7188 ( .A1(n5515), .A2(SI_23_), .ZN(n5516) );
  NAND2_X1 U7189 ( .A1(n7483), .A2(n7914), .ZN(n5518) );
  NAND2_X1 U7190 ( .A1(n7915), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7191 ( .A1(n5519), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7192 ( .A1(n5537), .A2(n5520), .ZN(n8552) );
  NAND2_X1 U7193 ( .A1(n8552), .A2(n5625), .ZN(n5525) );
  INV_X1 U7194 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U7195 ( .A1(n5678), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7196 ( .A1(n5219), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5521) );
  OAI211_X1 U7197 ( .C1(n10120), .C2(n7137), .A(n5522), .B(n5521), .ZN(n5523)
         );
  INV_X1 U7198 ( .A(n5523), .ZN(n5524) );
  INV_X2 U7199 ( .A(n8328), .ZN(n8560) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7529) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7530) );
  MUX2_X1 U7202 ( .A(n7529), .B(n7530), .S(n6513), .Z(n5530) );
  INV_X1 U7203 ( .A(SI_24_), .ZN(n5529) );
  NAND2_X1 U7204 ( .A1(n5530), .A2(n5529), .ZN(n5546) );
  INV_X1 U7205 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7206 ( .A1(n5531), .A2(SI_24_), .ZN(n5532) );
  NAND2_X1 U7207 ( .A1(n7527), .A2(n7914), .ZN(n5534) );
  NAND2_X1 U7208 ( .A1(n7915), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5533) );
  INV_X1 U7209 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7210 ( .A1(n5537), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7211 ( .A1(n5556), .A2(n5538), .ZN(n8539) );
  NAND2_X1 U7212 ( .A1(n8539), .A2(n5625), .ZN(n5543) );
  INV_X1 U7213 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U7214 ( .A1(n5678), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7215 ( .A1(n5219), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U7216 ( .C1(n8679), .C2(n7137), .A(n5540), .B(n5539), .ZN(n5541)
         );
  INV_X1 U7217 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7218 ( .A1(n8760), .A2(n8246), .ZN(n8085) );
  NAND2_X1 U7219 ( .A1(n8766), .A2(n8328), .ZN(n8083) );
  NAND2_X1 U7220 ( .A1(n8085), .A2(n8083), .ZN(n8095) );
  INV_X1 U7221 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5547) );
  INV_X1 U7222 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7599) );
  MUX2_X1 U7223 ( .A(n5547), .B(n7599), .S(n6514), .Z(n5549) );
  INV_X1 U7224 ( .A(SI_25_), .ZN(n5548) );
  NAND2_X1 U7225 ( .A1(n5549), .A2(n5548), .ZN(n5565) );
  INV_X1 U7226 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U7227 ( .A1(n5550), .A2(SI_25_), .ZN(n5551) );
  XNOR2_X1 U7228 ( .A(n5564), .B(n5563), .ZN(n7570) );
  NAND2_X1 U7229 ( .A1(n7570), .A2(n7914), .ZN(n5553) );
  NAND2_X1 U7230 ( .A1(n7915), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5552) );
  INV_X1 U7231 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7232 ( .A1(n5556), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7233 ( .A1(n5574), .A2(n5557), .ZN(n8527) );
  NAND2_X1 U7234 ( .A1(n8527), .A2(n5625), .ZN(n5562) );
  INV_X1 U7235 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U7236 ( .A1(n5678), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7237 ( .A1(n5219), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5558) );
  OAI211_X1 U7238 ( .C1(n10029), .C2(n7137), .A(n5559), .B(n5558), .ZN(n5560)
         );
  INV_X1 U7239 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7240 ( .A1(n8754), .A2(n5631), .ZN(n8087) );
  NAND2_X1 U7241 ( .A1(n5564), .A2(n5563), .ZN(n5566) );
  INV_X1 U7242 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5567) );
  INV_X1 U7243 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U7244 ( .A(n5567), .B(n10108), .S(n6513), .Z(n5569) );
  INV_X1 U7245 ( .A(SI_26_), .ZN(n5568) );
  NAND2_X1 U7246 ( .A1(n5569), .A2(n5568), .ZN(n5583) );
  INV_X1 U7247 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7248 ( .A1(n5570), .A2(SI_26_), .ZN(n5571) );
  NAND2_X1 U7249 ( .A1(n7602), .A2(n7914), .ZN(n5573) );
  NAND2_X1 U7250 ( .A1(n5155), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7251 ( .A1(n5574), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7252 ( .A1(n8517), .A2(n5625), .ZN(n5580) );
  INV_X1 U7253 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U7254 ( .A1(n5219), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7255 ( .A1(n5678), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U7256 ( .C1(n8674), .C2(n7137), .A(n5577), .B(n5576), .ZN(n5578)
         );
  INV_X1 U7257 ( .A(n5578), .ZN(n5579) );
  OAI21_X1 U7258 ( .B1(n8511), .B2(n7927), .A(n8101), .ZN(n8500) );
  NAND2_X1 U7259 ( .A1(n5582), .A2(n5581), .ZN(n5584) );
  INV_X1 U7260 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5585) );
  MUX2_X1 U7261 ( .A(n5585), .B(n7626), .S(n6513), .Z(n5587) );
  INV_X1 U7262 ( .A(SI_27_), .ZN(n5586) );
  NAND2_X1 U7263 ( .A1(n5587), .A2(n5586), .ZN(n5603) );
  INV_X1 U7264 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7265 ( .A1(n5588), .A2(SI_27_), .ZN(n5589) );
  NAND2_X1 U7266 ( .A1(n7607), .A2(n7914), .ZN(n5591) );
  NAND2_X1 U7267 ( .A1(n7915), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5590) );
  INV_X1 U7268 ( .A(n5594), .ZN(n5593) );
  INV_X1 U7269 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7270 ( .A1(n5593), .A2(n5592), .ZN(n5608) );
  NAND2_X1 U7271 ( .A1(n5594), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7272 ( .A1(n5608), .A2(n5595), .ZN(n8195) );
  NAND2_X1 U7273 ( .A1(n8195), .A2(n5625), .ZN(n5600) );
  INV_X1 U7274 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U7275 ( .A1(n5678), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7276 ( .A1(n5219), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U7277 ( .C1(n7137), .C2(n10055), .A(n5597), .B(n5596), .ZN(n5598)
         );
  INV_X1 U7278 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U7279 ( .A1(n8672), .A2(n8348), .ZN(n8107) );
  NOR2_X1 U7280 ( .A1(n8672), .A2(n8348), .ZN(n8106) );
  NAND2_X1 U7281 ( .A1(n5602), .A2(n5601), .ZN(n5604) );
  INV_X1 U7282 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5605) );
  INV_X1 U7283 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7632) );
  MUX2_X1 U7284 ( .A(n5605), .B(n7632), .S(n6514), .Z(n5619) );
  XNOR2_X1 U7285 ( .A(n5619), .B(SI_28_), .ZN(n5616) );
  NAND2_X1 U7286 ( .A1(n7631), .A2(n7914), .ZN(n5607) );
  NAND2_X1 U7287 ( .A1(n5155), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7288 ( .A1(n5608), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7289 ( .A1(n8475), .A2(n5609), .ZN(n8494) );
  NAND2_X1 U7290 ( .A1(n8494), .A2(n5625), .ZN(n5614) );
  INV_X1 U7291 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U7292 ( .A1(n5219), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7293 ( .A1(n5678), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7294 ( .C1(n10097), .C2(n7137), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U7295 ( .A(n5612), .ZN(n5613) );
  NOR2_X1 U7296 ( .A1(n8741), .A2(n8369), .ZN(n5615) );
  OAI22_X1 U7297 ( .A1(n8489), .A2(n5615), .B1(n8505), .B2(n8495), .ZN(n7919)
         );
  NAND2_X1 U7298 ( .A1(n5617), .A2(n5616), .ZN(n5621) );
  INV_X1 U7299 ( .A(SI_28_), .ZN(n5618) );
  NAND2_X1 U7300 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  INV_X1 U7301 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5622) );
  INV_X1 U7302 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7629) );
  MUX2_X1 U7303 ( .A(n5622), .B(n7629), .S(n6513), .Z(n6188) );
  NAND2_X1 U7304 ( .A1(n7628), .A2(n7914), .ZN(n5624) );
  NAND2_X1 U7305 ( .A1(n7915), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5623) );
  INV_X1 U7306 ( .A(n8475), .ZN(n5626) );
  NAND2_X1 U7307 ( .A1(n5626), .A2(n5625), .ZN(n7140) );
  INV_X1 U7308 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U7309 ( .A1(n5678), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7310 ( .A1(n5219), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7311 ( .C1(n7137), .C2(n10127), .A(n5628), .B(n5627), .ZN(n5629)
         );
  INV_X1 U7312 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7313 ( .A1(n5715), .A2(n8368), .ZN(n7920) );
  INV_X1 U7314 ( .A(n8672), .ZN(n8200) );
  NAND2_X1 U7315 ( .A1(n6897), .A2(n6898), .ZN(n6896) );
  INV_X1 U7316 ( .A(n7099), .ZN(n6902) );
  OR2_X1 U7317 ( .A1(n7101), .A2(n6902), .ZN(n5632) );
  NAND2_X1 U7318 ( .A1(n6896), .A2(n5632), .ZN(n9864) );
  NAND2_X1 U7319 ( .A1(n9864), .A2(n9865), .ZN(n9863) );
  OR2_X1 U7320 ( .A1(n8380), .A2(n5149), .ZN(n6998) );
  NAND2_X1 U7321 ( .A1(n9863), .A2(n6998), .ZN(n5634) );
  NAND2_X1 U7322 ( .A1(n5634), .A2(n5633), .ZN(n6997) );
  OR2_X1 U7323 ( .A1(n9861), .A2(n9886), .ZN(n7082) );
  NAND2_X1 U7324 ( .A1(n6997), .A2(n7082), .ZN(n5635) );
  INV_X1 U7325 ( .A(n8204), .ZN(n9891) );
  OR2_X1 U7326 ( .A1(n7143), .A2(n9891), .ZN(n5636) );
  NAND2_X1 U7327 ( .A1(n8379), .A2(n5638), .ZN(n5637) );
  NAND2_X1 U7328 ( .A1(n7987), .A2(n7996), .ZN(n7932) );
  NAND2_X1 U7329 ( .A1(n7211), .A2(n7932), .ZN(n5640) );
  INV_X1 U7330 ( .A(n7246), .ZN(n9901) );
  OR2_X1 U7331 ( .A1(n8378), .A2(n9901), .ZN(n5639) );
  NAND2_X1 U7332 ( .A1(n5640), .A2(n5639), .ZN(n7222) );
  NAND2_X1 U7333 ( .A1(n8377), .A2(n7257), .ZN(n7313) );
  INV_X1 U7334 ( .A(n9910), .ZN(n7325) );
  NAND2_X1 U7335 ( .A1(n8376), .A2(n7325), .ZN(n5641) );
  INV_X1 U7336 ( .A(n5641), .ZN(n5642) );
  NAND2_X1 U7337 ( .A1(n8011), .A2(n8001), .ZN(n7938) );
  OR2_X1 U7338 ( .A1(n9919), .A2(n8375), .ZN(n5643) );
  NAND2_X1 U7339 ( .A1(n9919), .A2(n8375), .ZN(n5644) );
  OR2_X1 U7340 ( .A1(n7496), .A2(n8374), .ZN(n5646) );
  NAND2_X1 U7341 ( .A1(n7399), .A2(n5646), .ZN(n5647) );
  NAND2_X1 U7342 ( .A1(n7496), .A2(n8374), .ZN(n7558) );
  INV_X1 U7343 ( .A(n7556), .ZN(n8373) );
  NAND2_X1 U7344 ( .A1(n7507), .A2(n8373), .ZN(n7513) );
  INV_X1 U7345 ( .A(n7568), .ZN(n5648) );
  NAND2_X1 U7346 ( .A1(n7589), .A2(n8371), .ZN(n7573) );
  NAND2_X1 U7347 ( .A1(n8240), .A2(n8655), .ZN(n5649) );
  AND2_X1 U7348 ( .A1(n7573), .A2(n5649), .ZN(n5651) );
  INV_X1 U7349 ( .A(n5649), .ZN(n5650) );
  OR2_X1 U7350 ( .A1(n7589), .A2(n8371), .ZN(n7575) );
  AOI21_X1 U7351 ( .B1(n7574), .B2(n5651), .A(n4327), .ZN(n5653) );
  OR2_X1 U7352 ( .A1(n8240), .A2(n8655), .ZN(n5652) );
  NAND2_X1 U7353 ( .A1(n8805), .A2(n8370), .ZN(n5654) );
  NAND2_X1 U7354 ( .A1(n8061), .A2(n8058), .ZN(n8630) );
  INV_X1 U7355 ( .A(n8647), .ZN(n8621) );
  NAND2_X1 U7356 ( .A1(n8799), .A2(n8621), .ZN(n8601) );
  OR2_X1 U7357 ( .A1(n8702), .A2(n8620), .ZN(n5657) );
  NAND2_X1 U7358 ( .A1(n8793), .A2(n8605), .ZN(n8602) );
  NAND2_X1 U7359 ( .A1(n8702), .A2(n8620), .ZN(n5655) );
  AND2_X1 U7360 ( .A1(n8601), .A2(n5656), .ZN(n5660) );
  INV_X1 U7361 ( .A(n5656), .ZN(n5659) );
  AND2_X1 U7362 ( .A1(n8618), .A2(n5657), .ZN(n5658) );
  INV_X1 U7363 ( .A(n8784), .ZN(n8321) );
  NAND2_X1 U7364 ( .A1(n8321), .A2(n8590), .ZN(n8569) );
  NOR2_X1 U7365 ( .A1(n8778), .A2(n8584), .ZN(n8557) );
  NAND2_X1 U7366 ( .A1(n5662), .A2(n8082), .ZN(n8556) );
  OAI21_X1 U7367 ( .B1(n8573), .B2(n8772), .A(n8559), .ZN(n8548) );
  NAND2_X1 U7368 ( .A1(n8548), .A2(n4879), .ZN(n5665) );
  NAND2_X1 U7369 ( .A1(n5665), .A2(n5664), .ZN(n8534) );
  NAND2_X1 U7370 ( .A1(n5666), .A2(n8087), .ZN(n8528) );
  NAND2_X1 U7371 ( .A1(n8748), .A2(n8523), .ZN(n5668) );
  INV_X1 U7372 ( .A(n8748), .ZN(n5667) );
  NAND2_X1 U7373 ( .A1(n8502), .A2(n5669), .ZN(n5670) );
  OAI21_X1 U7374 ( .B1(n8348), .B2(n8200), .A(n5670), .ZN(n8490) );
  NAND2_X1 U7375 ( .A1(n8144), .A2(n5673), .ZN(n5722) );
  INV_X1 U7376 ( .A(n7283), .ZN(n8135) );
  NAND2_X1 U7377 ( .A1(n7965), .A2(n8135), .ZN(n5672) );
  AOI21_X1 U7378 ( .B1(n7451), .B2(n8135), .A(n5673), .ZN(n5674) );
  INV_X1 U7379 ( .A(n5675), .ZN(n8142) );
  NAND2_X1 U7380 ( .A1(n5676), .A2(n8142), .ZN(n5677) );
  NAND2_X1 U7381 ( .A1(n5685), .A2(n5677), .ZN(n5684) );
  INV_X1 U7382 ( .A(n5684), .ZN(n7109) );
  INV_X1 U7383 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7384 ( .A1(n5219), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7385 ( .A1(n5678), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5679) );
  OAI211_X1 U7386 ( .C1(n5681), .C2(n7137), .A(n5680), .B(n5679), .ZN(n5682)
         );
  INV_X1 U7387 ( .A(n5682), .ZN(n5683) );
  NAND2_X1 U7388 ( .A1(n7140), .A2(n5683), .ZN(n8367) );
  AOI21_X1 U7389 ( .B1(P2_B_REG_SCAN_IN), .B2(n5685), .A(n8646), .ZN(n8472) );
  AOI22_X1 U7390 ( .A1(n9862), .A2(n8369), .B1(n8367), .B2(n8472), .ZN(n5686)
         );
  NAND2_X1 U7391 ( .A1(n5694), .A2(n5687), .ZN(n7093) );
  XNOR2_X1 U7392 ( .A(n5687), .B(P2_B_REG_SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7393 ( .A1(n5688), .A2(n5695), .ZN(n5689) );
  NAND3_X1 U7394 ( .A1(n8144), .A2(n8135), .A3(n8468), .ZN(n5692) );
  NAND2_X1 U7395 ( .A1(n8127), .A2(n5692), .ZN(n5698) );
  OR2_X1 U7396 ( .A1(n6813), .A2(n5698), .ZN(n5701) );
  OR2_X1 U7397 ( .A1(n5693), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7398 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  INV_X1 U7399 ( .A(n5698), .ZN(n5699) );
  OR2_X1 U7400 ( .A1(n6812), .A2(n5699), .ZN(n5700) );
  NAND2_X1 U7401 ( .A1(n5701), .A2(n5700), .ZN(n6814) );
  NOR2_X1 U7402 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n9999) );
  NOR4_X1 U7403 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5704) );
  NOR4_X1 U7404 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5703) );
  NOR4_X1 U7405 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5702) );
  NAND4_X1 U7406 ( .A1(n9999), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n5710)
         );
  NOR4_X1 U7407 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5708) );
  NOR4_X1 U7408 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5707) );
  NOR4_X1 U7409 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5706) );
  NOR4_X1 U7410 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5705) );
  NAND4_X1 U7411 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n5709)
         );
  NOR2_X1 U7412 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  OR2_X1 U7413 ( .A1(n8127), .A2(n5712), .ZN(n5713) );
  AND2_X1 U7414 ( .A1(n5721), .A2(n5713), .ZN(n6743) );
  NAND3_X1 U7415 ( .A1(n5724), .A2(n6562), .A3(n6743), .ZN(n6811) );
  AND2_X1 U7416 ( .A1(n9926), .A2(n7958), .ZN(n6760) );
  NOR2_X1 U7417 ( .A1(n6811), .A2(n6760), .ZN(n5714) );
  NAND2_X1 U7418 ( .A1(n9954), .A2(n9920), .ZN(n8670) );
  INV_X1 U7419 ( .A(n5716), .ZN(n5717) );
  OAI21_X1 U7420 ( .B1(n5732), .B2(n5718), .A(n5717), .ZN(P2_U3488) );
  INV_X1 U7421 ( .A(n5724), .ZN(n5719) );
  NAND2_X1 U7422 ( .A1(n6747), .A2(n6761), .ZN(n6759) );
  OR3_X1 U7423 ( .A1(n5722), .A2(n7965), .A3(n7283), .ZN(n6742) );
  AND2_X1 U7424 ( .A1(n6749), .A2(n6742), .ZN(n5723) );
  OR2_X1 U7425 ( .A1(n6759), .A2(n5723), .ZN(n5727) );
  NAND3_X1 U7426 ( .A1(n6813), .A2(n6812), .A3(n5724), .ZN(n6751) );
  INV_X1 U7427 ( .A(n6761), .ZN(n6535) );
  AND2_X1 U7428 ( .A1(n8127), .A2(n9928), .ZN(n5725) );
  NAND2_X1 U7429 ( .A1(n5725), .A2(n6742), .ZN(n6755) );
  NAND2_X1 U7430 ( .A1(n6755), .A2(n8532), .ZN(n6741) );
  NAND2_X1 U7431 ( .A1(n6764), .A2(n6741), .ZN(n5726) );
  INV_X1 U7432 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5729) );
  OAI21_X1 U7433 ( .B1(n5732), .B2(n9936), .A(n5731), .ZN(P2_U3456) );
  NAND2_X1 U7434 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5862) );
  NAND2_X1 U7435 ( .A1(n5881), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7436 ( .A1(n5933), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5945) );
  INV_X1 U7437 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5783) );
  INV_X1 U7438 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6047) );
  INV_X1 U7439 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U7440 ( .A1(n6050), .A2(n10032), .ZN(n5739) );
  NAND2_X1 U7441 ( .A1(n6058), .A2(n5739), .ZN(n9236) );
  INV_X2 U7442 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5875) );
  NOR2_X1 U7443 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5746) );
  NOR2_X1 U7444 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5745) );
  NOR2_X1 U7445 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5743) );
  NOR2_X1 U7446 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5749) );
  NOR2_X1 U7447 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5748) );
  NOR2_X1 U7448 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5747) );
  NAND4_X1 U7449 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n5751)
         );
  INV_X1 U7450 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7451 ( .A1(n5769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5753) );
  INV_X1 U7452 ( .A(n5756), .ZN(n9474) );
  INV_X1 U7453 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5763) );
  INV_X4 U7454 ( .A(n5852), .ZN(n7753) );
  NAND2_X1 U7455 ( .A1(n7753), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7456 ( .A1(n6140), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5761) );
  OAI211_X1 U7457 ( .C1(n5763), .C2(n6099), .A(n5762), .B(n5761), .ZN(n5764)
         );
  INV_X1 U7458 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U7459 ( .A1(n7483), .A2(n6210), .ZN(n5776) );
  OR2_X1 U7460 ( .A1(n5844), .A2(n7486), .ZN(n5775) );
  NAND2_X1 U7461 ( .A1(n7281), .A2(n6210), .ZN(n5778) );
  OR2_X1 U7462 ( .A1(n5844), .A2(n10016), .ZN(n5777) );
  AND2_X2 U7463 ( .A1(n5778), .A2(n5777), .ZN(n6035) );
  INV_X1 U7464 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U7465 ( .A1(n5785), .A2(n8920), .ZN(n5779) );
  AND2_X1 U7466 ( .A1(n6039), .A2(n5779), .ZN(n9280) );
  INV_X1 U7467 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U7468 ( .A1(n6140), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7469 ( .A1(n7753), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5780) );
  OAI211_X1 U7470 ( .C1(n6099), .C2(n9397), .A(n5781), .B(n5780), .ZN(n5782)
         );
  AOI21_X1 U7471 ( .B1(n9280), .B2(n4285), .A(n5782), .ZN(n8871) );
  NAND2_X1 U7472 ( .A1(n5796), .A2(n5783), .ZN(n5784) );
  NAND2_X1 U7473 ( .A1(n5785), .A2(n5784), .ZN(n9288) );
  INV_X1 U7474 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U7475 ( .A1(n7753), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7476 ( .A1(n6140), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5786) );
  OAI211_X1 U7477 ( .C1(n6099), .C2(n9097), .A(n5787), .B(n5786), .ZN(n5788)
         );
  INV_X1 U7478 ( .A(n5788), .ZN(n5789) );
  INV_X1 U7479 ( .A(n9311), .ZN(n6134) );
  NAND2_X1 U7480 ( .A1(n7252), .A2(n6210), .ZN(n5794) );
  INV_X1 U7481 ( .A(n6108), .ZN(n5790) );
  NAND2_X1 U7482 ( .A1(n6021), .A2(n6106), .ZN(n5791) );
  NAND2_X1 U7483 ( .A1(n5791), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7484 ( .A1(n5800), .A2(n6107), .ZN(n5802) );
  XNOR2_X2 U7485 ( .A(n5792), .B(n6105), .ZN(n7900) );
  AOI22_X1 U7486 ( .A1(n6023), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9103), .B2(
        n6022), .ZN(n5793) );
  INV_X1 U7487 ( .A(n9399), .ZN(n9291) );
  INV_X1 U7488 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7489 ( .A1(n6029), .A2(n8936), .ZN(n5795) );
  NAND2_X1 U7490 ( .A1(n5796), .A2(n5795), .ZN(n9304) );
  OR2_X1 U7491 ( .A1(n9304), .A2(n6081), .ZN(n5798) );
  AOI22_X1 U7492 ( .A1(n6140), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n7753), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5797) );
  OAI211_X1 U7493 ( .C1(n6099), .C2(n5799), .A(n5798), .B(n5797), .ZN(n9295)
         );
  NAND2_X1 U7494 ( .A1(n7161), .A2(n6210), .ZN(n5804) );
  OR2_X1 U7495 ( .A1(n5800), .A2(n6107), .ZN(n5801) );
  AND2_X1 U7496 ( .A1(n5802), .A2(n5801), .ZN(n9094) );
  AOI22_X1 U7497 ( .A1(n6023), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6022), .B2(
        n9094), .ZN(n5803) );
  NAND2_X1 U7498 ( .A1(n5821), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7499 ( .A1(n5837), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5806) );
  INV_X1 U7500 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7501 ( .A1(n5810), .A2(n5809), .ZN(n6225) );
  INV_X1 U7502 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7503 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5811) );
  XNOR2_X1 U7504 ( .A(n5812), .B(n5811), .ZN(n6599) );
  INV_X1 U7505 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7506 ( .A1(n6139), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7507 ( .A1(n5837), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7508 ( .A1(n5821), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7509 ( .A1(n5820), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7510 ( .A1(n6514), .A2(SI_0_), .ZN(n5817) );
  XNOR2_X1 U7511 ( .A(n5817), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9480) );
  MUX2_X1 U7512 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9480), .S(n6548), .Z(n9686) );
  AND2_X1 U7513 ( .A1(n7043), .A2(n9686), .ZN(n7040) );
  OAI22_X1 U7514 ( .A1(n6117), .A2(n7040), .B1(n8983), .B2(n7053), .ZN(n9670)
         );
  INV_X1 U7515 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7516 ( .A1(n5820), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7517 ( .A1(n5837), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7518 ( .A1(n5821), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U7519 ( .A1(n5826), .A2(n9473), .ZN(n5827) );
  MUX2_X1 U7520 ( .A(n9473), .B(n5827), .S(P1_IR_REG_2__SCAN_IN), .Z(n5828) );
  INV_X1 U7521 ( .A(n5828), .ZN(n5831) );
  BUF_X1 U7522 ( .A(n5829), .Z(n5830) );
  NAND2_X1 U7523 ( .A1(n5831), .A2(n5830), .ZN(n9003) );
  INV_X1 U7524 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6516) );
  OR2_X1 U7525 ( .A1(n5844), .A2(n6516), .ZN(n5833) );
  OR2_X1 U7526 ( .A1(n5845), .A2(n6515), .ZN(n5832) );
  OAI211_X1 U7527 ( .C1(n6548), .C2(n9003), .A(n5833), .B(n5832), .ZN(n6249)
         );
  NAND2_X1 U7528 ( .A1(n6941), .A2(n6249), .ZN(n6119) );
  NAND2_X1 U7529 ( .A1(n8982), .A2(n5834), .ZN(n7838) );
  NAND2_X1 U7530 ( .A1(n6119), .A2(n7838), .ZN(n9669) );
  NAND2_X1 U7531 ( .A1(n9670), .A2(n9669), .ZN(n5836) );
  NAND2_X1 U7532 ( .A1(n6941), .A2(n5834), .ZN(n5835) );
  NAND2_X1 U7533 ( .A1(n5836), .A2(n5835), .ZN(n6938) );
  NAND2_X1 U7534 ( .A1(n7752), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7535 ( .A1(n7751), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7536 ( .A1(n5837), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5839) );
  INV_X1 U7537 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U7538 ( .A1(n6139), .A2(n6944), .ZN(n5838) );
  NAND4_X2 U7539 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n8981)
         );
  NAND2_X1 U7540 ( .A1(n5830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U7541 ( .A(n5843), .B(n5842), .ZN(n9019) );
  OR2_X1 U7542 ( .A1(n5844), .A2(n5161), .ZN(n5847) );
  OR2_X1 U7543 ( .A1(n5845), .A2(n6518), .ZN(n5846) );
  OAI211_X1 U7544 ( .C1(n6548), .C2(n9019), .A(n5847), .B(n5846), .ZN(n6943)
         );
  AND2_X1 U7545 ( .A1(n8981), .A2(n9703), .ZN(n7645) );
  NAND2_X1 U7546 ( .A1(n6938), .A2(n7775), .ZN(n5849) );
  NAND2_X1 U7547 ( .A1(n9720), .A2(n9703), .ZN(n5848) );
  NAND2_X1 U7548 ( .A1(n5849), .A2(n5848), .ZN(n9708) );
  NAND2_X1 U7549 ( .A1(n7751), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5856) );
  INV_X1 U7550 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7551 ( .A1(n6944), .A2(n5850), .ZN(n5851) );
  AND2_X1 U7552 ( .A1(n5851), .A2(n5862), .ZN(n10145) );
  NAND2_X1 U7553 ( .A1(n6139), .A2(n10145), .ZN(n5855) );
  NAND2_X1 U7554 ( .A1(n7753), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7555 ( .A1(n7752), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7556 ( .A1(n5830), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7557 ( .A1(n5877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  XNOR2_X1 U7558 ( .A(n5868), .B(n5875), .ZN(n9030) );
  OR2_X1 U7559 ( .A1(n5845), .A2(n6519), .ZN(n5859) );
  INV_X1 U7560 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7561 ( .A1(n5844), .A2(n5857), .ZN(n5858) );
  OAI211_X1 U7562 ( .C1(n6548), .C2(n9030), .A(n5859), .B(n5858), .ZN(n6267)
         );
  NOR2_X1 U7563 ( .A1(n8980), .A2(n6267), .ZN(n5861) );
  NAND2_X1 U7564 ( .A1(n8980), .A2(n6267), .ZN(n5860) );
  AND2_X1 U7565 ( .A1(n5862), .A2(n6777), .ZN(n5863) );
  NOR2_X1 U7566 ( .A1(n5881), .A2(n5863), .ZN(n6951) );
  NAND2_X1 U7567 ( .A1(n4285), .A2(n6951), .ZN(n5867) );
  NAND2_X1 U7568 ( .A1(n7751), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7569 ( .A1(n7753), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7570 ( .A1(n7752), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5864) );
  NAND4_X1 U7571 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n8979)
         );
  INV_X1 U7572 ( .A(n8979), .ZN(n9722) );
  NOR2_X1 U7573 ( .A1(n6526), .A2(n5845), .ZN(n5872) );
  INV_X1 U7574 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7575 ( .A1(n5868), .A2(n5875), .ZN(n5869) );
  NAND2_X1 U7576 ( .A1(n5869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U7577 ( .A(n5870), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9542) );
  INV_X1 U7578 ( .A(n9542), .ZN(n6525) );
  OAI22_X1 U7579 ( .A1(n5844), .A2(n6524), .B1(n6548), .B2(n6525), .ZN(n5871)
         );
  NAND2_X1 U7580 ( .A1(n9722), .A2(n6952), .ZN(n7650) );
  INV_X1 U7581 ( .A(n6952), .ZN(n6915) );
  NAND2_X1 U7582 ( .A1(n6915), .A2(n8979), .ZN(n7852) );
  NAND2_X1 U7583 ( .A1(n7650), .A2(n7852), .ZN(n7774) );
  INV_X1 U7584 ( .A(n7774), .ZN(n6906) );
  NAND2_X1 U7585 ( .A1(n9722), .A2(n6915), .ZN(n5873) );
  OR2_X1 U7586 ( .A1(n6530), .A2(n5845), .ZN(n5880) );
  INV_X1 U7587 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7588 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  OR2_X1 U7589 ( .A1(n5980), .A2(n9473), .ZN(n5878) );
  XNOR2_X1 U7590 ( .A(n5878), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6607) );
  AOI22_X1 U7591 ( .A1(n6023), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6022), .B2(
        n6607), .ZN(n5879) );
  NAND2_X1 U7592 ( .A1(n5880), .A2(n5879), .ZN(n6852) );
  INV_X1 U7593 ( .A(n6852), .ZN(n6934) );
  NAND2_X1 U7594 ( .A1(n7751), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7595 ( .A1(n5881), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5882) );
  AND2_X1 U7596 ( .A1(n5893), .A2(n5882), .ZN(n6853) );
  NAND2_X1 U7597 ( .A1(n4285), .A2(n6853), .ZN(n5885) );
  NAND2_X1 U7598 ( .A1(n7753), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7599 ( .A1(n7752), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5883) );
  NAND4_X1 U7600 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n8978)
         );
  NAND2_X1 U7601 ( .A1(n6934), .A2(n8978), .ZN(n7648) );
  INV_X1 U7602 ( .A(n8978), .ZN(n6778) );
  NAND2_X1 U7603 ( .A1(n6778), .A2(n6852), .ZN(n7654) );
  NAND2_X1 U7604 ( .A1(n7648), .A2(n7654), .ZN(n7773) );
  NAND2_X1 U7605 ( .A1(n6850), .A2(n7773), .ZN(n6849) );
  NAND2_X1 U7606 ( .A1(n6934), .A2(n6778), .ZN(n5887) );
  NAND2_X1 U7607 ( .A1(n6849), .A2(n5887), .ZN(n7011) );
  OR2_X1 U7608 ( .A1(n6533), .A2(n5845), .ZN(n5891) );
  INV_X1 U7609 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7610 ( .A1(n5980), .A2(n5888), .ZN(n5900) );
  NAND2_X1 U7611 ( .A1(n5900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7612 ( .A(n5889), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6610) );
  AOI22_X1 U7613 ( .A1(n6023), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6022), .B2(
        n6610), .ZN(n5890) );
  NAND2_X1 U7614 ( .A1(n5891), .A2(n5890), .ZN(n9651) );
  NAND2_X1 U7615 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  AND2_X1 U7616 ( .A1(n5906), .A2(n5894), .ZN(n9650) );
  NAND2_X1 U7617 ( .A1(n4285), .A2(n9650), .ZN(n5898) );
  NAND2_X1 U7618 ( .A1(n7751), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7619 ( .A1(n7753), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7620 ( .A1(n6140), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5895) );
  NAND4_X1 U7621 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n8977)
         );
  NAND2_X1 U7622 ( .A1(n7025), .A2(n8977), .ZN(n6127) );
  INV_X1 U7623 ( .A(n8977), .ZN(n7176) );
  NAND2_X1 U7624 ( .A1(n9651), .A2(n7176), .ZN(n6963) );
  NAND2_X1 U7625 ( .A1(n7025), .A2(n7176), .ZN(n5899) );
  NAND2_X1 U7626 ( .A1(n6543), .A2(n6210), .ZN(n5904) );
  NAND2_X1 U7627 ( .A1(n5927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7628 ( .A1(n5901), .A2(n5925), .ZN(n5912) );
  OR2_X1 U7629 ( .A1(n5901), .A2(n5925), .ZN(n5902) );
  AOI22_X1 U7630 ( .A1(n6023), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6022), .B2(
        n6612), .ZN(n5903) );
  NAND2_X1 U7631 ( .A1(n7751), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7632 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7633 ( .A1(n5917), .A2(n5907), .ZN(n7173) );
  INV_X1 U7634 ( .A(n7173), .ZN(n6974) );
  NAND2_X1 U7635 ( .A1(n4285), .A2(n6974), .ZN(n5910) );
  NAND2_X1 U7636 ( .A1(n7753), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7637 ( .A1(n6140), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5908) );
  NAND4_X1 U7638 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n8976)
         );
  INV_X1 U7639 ( .A(n8976), .ZN(n7203) );
  OR2_X1 U7640 ( .A1(n7178), .A2(n7203), .ZN(n6980) );
  NAND2_X1 U7641 ( .A1(n7178), .A2(n7203), .ZN(n7661) );
  NAND2_X1 U7642 ( .A1(n6980), .A2(n7661), .ZN(n6966) );
  NAND2_X1 U7643 ( .A1(n6563), .A2(n6210), .ZN(n5915) );
  NAND2_X1 U7644 ( .A1(n5912), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5913) );
  XNOR2_X1 U7645 ( .A(n5913), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7646 ( .A1(n6023), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6022), .B2(
        n6790), .ZN(n5914) );
  NAND2_X1 U7647 ( .A1(n7751), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5922) );
  AND2_X1 U7648 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NOR2_X1 U7649 ( .A1(n5933), .A2(n5918), .ZN(n7206) );
  NAND2_X1 U7650 ( .A1(n4285), .A2(n7206), .ZN(n5921) );
  NAND2_X1 U7651 ( .A1(n7753), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7652 ( .A1(n6140), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5919) );
  NAND4_X1 U7653 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n8975)
         );
  INV_X1 U7654 ( .A(n8975), .ZN(n6968) );
  OR2_X1 U7655 ( .A1(n6992), .A2(n6968), .ZN(n7783) );
  NAND2_X1 U7656 ( .A1(n6992), .A2(n6968), .ZN(n7671) );
  NAND2_X1 U7657 ( .A1(n7783), .A2(n7671), .ZN(n6986) );
  NAND2_X1 U7658 ( .A1(n6987), .A2(n6986), .ZN(n6989) );
  OR2_X1 U7659 ( .A1(n6570), .A2(n5845), .ZN(n5932) );
  INV_X1 U7660 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7661 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NOR2_X1 U7662 ( .A1(n5927), .A2(n5926), .ZN(n5929) );
  OR2_X1 U7663 ( .A1(n5929), .A2(n9473), .ZN(n5928) );
  MUX2_X1 U7664 ( .A(n5928), .B(P1_IR_REG_31__SCAN_IN), .S(n10000), .Z(n5930)
         );
  NAND2_X1 U7665 ( .A1(n5929), .A2(n10000), .ZN(n5953) );
  NAND2_X1 U7666 ( .A1(n5930), .A2(n5953), .ZN(n6791) );
  INV_X1 U7667 ( .A(n6791), .ZN(n9489) );
  AOI22_X1 U7668 ( .A1(n6023), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6022), .B2(
        n9489), .ZN(n5931) );
  NAND2_X1 U7669 ( .A1(n7751), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5940) );
  INV_X1 U7670 ( .A(n5933), .ZN(n5935) );
  INV_X1 U7671 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7672 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7673 ( .A1(n5945), .A2(n5936), .ZN(n9534) );
  INV_X1 U7674 ( .A(n9534), .ZN(n7128) );
  NAND2_X1 U7675 ( .A1(n4285), .A2(n7128), .ZN(n5939) );
  NAND2_X1 U7676 ( .A1(n7753), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7677 ( .A1(n6140), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5937) );
  NAND4_X1 U7678 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n8974)
         );
  INV_X1 U7679 ( .A(n8974), .ZN(n7289) );
  OR2_X1 U7680 ( .A1(n7158), .A2(n7289), .ZN(n7853) );
  NAND2_X1 U7681 ( .A1(n7158), .A2(n7289), .ZN(n7665) );
  NAND2_X1 U7682 ( .A1(n6580), .A2(n6210), .ZN(n5943) );
  NAND2_X1 U7683 ( .A1(n5953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5941) );
  XNOR2_X1 U7684 ( .A(n5941), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U7685 ( .A1(n6023), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6022), .B2(
        n9575), .ZN(n5942) );
  INV_X1 U7686 ( .A(n7233), .ZN(n7294) );
  NAND2_X1 U7687 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  AND2_X1 U7688 ( .A1(n5960), .A2(n5946), .ZN(n7291) );
  NAND2_X1 U7689 ( .A1(n4285), .A2(n7291), .ZN(n5950) );
  NAND2_X1 U7690 ( .A1(n7751), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7691 ( .A1(n7753), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7692 ( .A1(n6140), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5947) );
  NAND4_X1 U7693 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n8973)
         );
  INV_X1 U7694 ( .A(n8973), .ZN(n7338) );
  NAND2_X1 U7695 ( .A1(n7294), .A2(n7338), .ZN(n5951) );
  NAND2_X1 U7696 ( .A1(n5952), .A2(n5951), .ZN(n7266) );
  OR2_X1 U7697 ( .A1(n6628), .A2(n5845), .ZN(n5958) );
  NAND2_X1 U7698 ( .A1(n5954), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5955) );
  INV_X1 U7699 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U7700 ( .A1(n5955), .A2(n10091), .ZN(n5967) );
  OR2_X1 U7701 ( .A1(n5955), .A2(n10091), .ZN(n5956) );
  AOI22_X1 U7702 ( .A1(n6023), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6022), .B2(
        n9060), .ZN(n5957) );
  NAND2_X1 U7703 ( .A1(n7751), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5965) );
  INV_X1 U7704 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7705 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  AND2_X1 U7706 ( .A1(n5972), .A2(n5961), .ZN(n7340) );
  NAND2_X1 U7707 ( .A1(n4285), .A2(n7340), .ZN(n5964) );
  NAND2_X1 U7708 ( .A1(n7753), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7709 ( .A1(n6140), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5962) );
  NAND4_X1 U7710 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n8972)
         );
  INV_X1 U7711 ( .A(n8972), .ZN(n7186) );
  AND2_X1 U7712 ( .A1(n7275), .A2(n7186), .ZN(n7677) );
  INV_X1 U7713 ( .A(n7677), .ZN(n7860) );
  INV_X1 U7714 ( .A(n7270), .ZN(n7267) );
  INV_X1 U7715 ( .A(n9739), .ZN(n5966) );
  NAND2_X1 U7716 ( .A1(n6711), .A2(n6210), .ZN(n5970) );
  NAND2_X1 U7717 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  AOI22_X1 U7718 ( .A1(n9587), .A2(n6022), .B1(n6023), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7719 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  AND2_X1 U7720 ( .A1(n5989), .A2(n5973), .ZN(n7395) );
  NAND2_X1 U7721 ( .A1(n4285), .A2(n7395), .ZN(n5977) );
  NAND2_X1 U7722 ( .A1(n7751), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7723 ( .A1(n7753), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7724 ( .A1(n6140), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U7725 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8971)
         );
  INV_X1 U7726 ( .A(n8971), .ZN(n5978) );
  NOR2_X1 U7727 ( .A1(n6339), .A2(n5978), .ZN(n7687) );
  INV_X1 U7728 ( .A(n7687), .ZN(n7640) );
  NAND2_X1 U7729 ( .A1(n6339), .A2(n5978), .ZN(n7685) );
  NAND2_X1 U7730 ( .A1(n6769), .A2(n6210), .ZN(n5987) );
  AND2_X1 U7731 ( .A1(n5980), .A2(n5979), .ZN(n5983) );
  NOR2_X1 U7732 ( .A1(n5983), .A2(n9473), .ZN(n5981) );
  MUX2_X1 U7733 ( .A(n9473), .B(n5981), .S(P1_IR_REG_14__SCAN_IN), .Z(n5985)
         );
  NAND2_X1 U7734 ( .A1(n5983), .A2(n5982), .ZN(n5995) );
  INV_X1 U7735 ( .A(n5995), .ZN(n5984) );
  OR2_X1 U7736 ( .A1(n5985), .A2(n5984), .ZN(n9602) );
  INV_X1 U7737 ( .A(n9602), .ZN(n9062) );
  AOI22_X1 U7738 ( .A1(n6023), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6022), .B2(
        n9062), .ZN(n5986) );
  NAND2_X1 U7739 ( .A1(n7751), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7740 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  AND2_X1 U7741 ( .A1(n6002), .A2(n5990), .ZN(n9640) );
  NAND2_X1 U7742 ( .A1(n4285), .A2(n9640), .ZN(n5993) );
  NAND2_X1 U7743 ( .A1(n7753), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7744 ( .A1(n6140), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5991) );
  NAND4_X1 U7745 ( .A1(n5994), .A2(n5993), .A3(n5992), .A4(n5991), .ZN(n8970)
         );
  INV_X1 U7746 ( .A(n8970), .ZN(n6347) );
  NOR2_X1 U7747 ( .A1(n9430), .A2(n6347), .ZN(n7691) );
  INV_X1 U7748 ( .A(n7691), .ZN(n7641) );
  NAND2_X1 U7749 ( .A1(n9430), .A2(n6347), .ZN(n7686) );
  NAND2_X1 U7750 ( .A1(n7641), .A2(n7686), .ZN(n9422) );
  NAND2_X1 U7751 ( .A1(n6824), .A2(n6210), .ZN(n6000) );
  NAND2_X1 U7752 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  MUX2_X1 U7753 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5996), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5998) );
  NAND2_X1 U7754 ( .A1(n5998), .A2(n5997), .ZN(n9064) );
  INV_X1 U7755 ( .A(n9064), .ZN(n9615) );
  AOI22_X1 U7756 ( .A1(n6023), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6022), .B2(
        n9615), .ZN(n5999) );
  INV_X1 U7757 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7758 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  AND2_X1 U7759 ( .A1(n6014), .A2(n6003), .ZN(n8954) );
  NAND2_X1 U7760 ( .A1(n4285), .A2(n8954), .ZN(n6007) );
  NAND2_X1 U7761 ( .A1(n7751), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7762 ( .A1(n7753), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7763 ( .A1(n6140), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6004) );
  NAND4_X1 U7764 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n9344)
         );
  INV_X1 U7765 ( .A(n9344), .ZN(n6132) );
  NAND2_X1 U7766 ( .A1(n6892), .A2(n6210), .ZN(n6012) );
  NAND2_X1 U7767 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7768 ( .A(n6010), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9075) );
  AOI22_X1 U7769 ( .A1(n6023), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6022), .B2(
        n9075), .ZN(n6011) );
  NAND2_X1 U7770 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  NAND2_X1 U7771 ( .A1(n6027), .A2(n6015), .ZN(n9338) );
  NAND2_X1 U7772 ( .A1(n7751), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7773 ( .A1(n7753), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6016) );
  AND2_X1 U7774 ( .A1(n6017), .A2(n6016), .ZN(n6019) );
  NAND2_X1 U7775 ( .A1(n6140), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6018) );
  OAI211_X1 U7776 ( .C1(n9338), .C2(n6081), .A(n6019), .B(n6018), .ZN(n8969)
         );
  INV_X1 U7777 ( .A(n8969), .ZN(n6020) );
  NAND2_X1 U7778 ( .A1(n9415), .A2(n6020), .ZN(n7868) );
  NAND2_X1 U7779 ( .A1(n7007), .A2(n6210), .ZN(n6025) );
  XNOR2_X1 U7780 ( .A(n6021), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9085) );
  AOI22_X1 U7781 ( .A1(n6023), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6022), .B2(
        n9085), .ZN(n6024) );
  INV_X1 U7782 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9328) );
  INV_X1 U7783 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7784 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  NAND2_X1 U7785 ( .A1(n6029), .A2(n6028), .ZN(n9327) );
  OR2_X1 U7786 ( .A1(n9327), .A2(n6081), .ZN(n6031) );
  AOI22_X1 U7787 ( .A1(n7751), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7753), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6030) );
  OAI211_X1 U7788 ( .C1(n6032), .C2(n9328), .A(n6031), .B(n6030), .ZN(n9346)
         );
  INV_X1 U7789 ( .A(n9346), .ZN(n8937) );
  INV_X1 U7790 ( .A(n9405), .ZN(n9307) );
  INV_X1 U7791 ( .A(n9295), .ZN(n8862) );
  OAI21_X1 U7792 ( .B1(n6134), .B2(n9291), .A(n6034), .ZN(n9274) );
  INV_X1 U7793 ( .A(n8871), .ZN(n9296) );
  NAND2_X1 U7794 ( .A1(n6035), .A2(n9296), .ZN(n9256) );
  NAND2_X1 U7795 ( .A1(n9258), .A2(n9256), .ZN(n9275) );
  NAND2_X1 U7796 ( .A1(n7343), .A2(n6210), .ZN(n6037) );
  OR2_X1 U7797 ( .A1(n5844), .A2(n7387), .ZN(n6036) );
  INV_X1 U7798 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7799 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U7800 ( .A1(n6048), .A2(n6040), .ZN(n9266) );
  OR2_X1 U7801 ( .A1(n9266), .A2(n6081), .ZN(n6045) );
  INV_X1 U7802 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U7803 ( .A1(n7753), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7804 ( .A1(n6140), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6041) );
  OAI211_X1 U7805 ( .C1(n6099), .C2(n9391), .A(n6042), .B(n6041), .ZN(n6043)
         );
  INV_X1 U7806 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7807 ( .A1(n6045), .A2(n6044), .ZN(n8968) );
  INV_X1 U7808 ( .A(n8968), .ZN(n7769) );
  NOR2_X1 U7809 ( .A1(n9457), .A2(n7769), .ZN(n6046) );
  INV_X1 U7810 ( .A(n9453), .ZN(n9248) );
  NAND2_X1 U7811 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  AND2_X1 U7812 ( .A1(n6050), .A2(n6049), .ZN(n9249) );
  INV_X1 U7813 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U7814 ( .A1(n7753), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7815 ( .A1(n6140), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7816 ( .C1(n9386), .C2(n6099), .A(n6052), .B(n6051), .ZN(n6053)
         );
  INV_X1 U7817 ( .A(n4292), .ZN(n8967) );
  NAND2_X1 U7818 ( .A1(n9248), .A2(n8967), .ZN(n6054) );
  NOR2_X1 U7819 ( .A1(n9380), .A2(n8966), .ZN(n9218) );
  NAND2_X1 U7820 ( .A1(n7527), .A2(n6210), .ZN(n6056) );
  OR2_X1 U7821 ( .A1(n5844), .A2(n7530), .ZN(n6055) );
  INV_X1 U7822 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6057) );
  OR2_X2 U7823 ( .A1(n6058), .A2(n6057), .ZN(n6067) );
  NAND2_X1 U7824 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  AND2_X1 U7825 ( .A1(n6067), .A2(n6059), .ZN(n9212) );
  NAND2_X1 U7826 ( .A1(n9212), .A2(n4285), .ZN(n6064) );
  INV_X1 U7827 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U7828 ( .A1(n7751), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7829 ( .A1(n7752), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6060) );
  OAI211_X1 U7830 ( .C1(n5852), .C2(n10125), .A(n6061), .B(n6060), .ZN(n6062)
         );
  INV_X1 U7831 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7832 ( .A1(n6064), .A2(n6063), .ZN(n8965) );
  INV_X1 U7833 ( .A(n8965), .ZN(n9235) );
  NAND2_X1 U7834 ( .A1(n7570), .A2(n6210), .ZN(n6066) );
  OR2_X1 U7835 ( .A1(n5844), .A2(n7599), .ZN(n6065) );
  INV_X1 U7836 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10031) );
  OR2_X2 U7837 ( .A1(n6067), .A2(n10031), .ZN(n6079) );
  NAND2_X1 U7838 ( .A1(n6067), .A2(n10031), .ZN(n6068) );
  NAND2_X1 U7839 ( .A1(n9195), .A2(n4285), .ZN(n6073) );
  INV_X1 U7840 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U7841 ( .A1(n7753), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7842 ( .A1(n7752), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6069) );
  OAI211_X1 U7843 ( .C1(n6099), .C2(n9371), .A(n6070), .B(n6069), .ZN(n6071)
         );
  INV_X1 U7844 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7845 ( .A1(n9194), .A2(n8964), .ZN(n6075) );
  NOR2_X1 U7846 ( .A1(n9194), .A2(n8964), .ZN(n6074) );
  NAND2_X1 U7847 ( .A1(n7602), .A2(n6210), .ZN(n6077) );
  OR2_X1 U7848 ( .A1(n5844), .A2(n10108), .ZN(n6076) );
  INV_X1 U7849 ( .A(n6079), .ZN(n6078) );
  NAND2_X1 U7850 ( .A1(n6078), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6089) );
  INV_X1 U7851 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7852 ( .A1(n6079), .A2(n6488), .ZN(n6080) );
  NAND2_X1 U7853 ( .A1(n6089), .A2(n6080), .ZN(n9178) );
  INV_X1 U7854 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U7855 ( .A1(n7751), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7856 ( .A1(n6140), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6082) );
  OAI211_X1 U7857 ( .C1(n5852), .C2(n10014), .A(n6083), .B(n6082), .ZN(n6084)
         );
  INV_X1 U7858 ( .A(n6084), .ZN(n6085) );
  NAND2_X1 U7859 ( .A1(n9442), .A2(n7724), .ZN(n6087) );
  INV_X1 U7860 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7861 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  INV_X1 U7862 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U7863 ( .A1(n6140), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7864 ( .A1(n7753), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6091) );
  OAI211_X1 U7865 ( .C1(n6099), .C2(n9361), .A(n6092), .B(n6091), .ZN(n6093)
         );
  AOI21_X2 U7866 ( .B1(n9163), .B2(n6139), .A(n6093), .ZN(n6485) );
  INV_X1 U7867 ( .A(n6485), .ZN(n8962) );
  OR2_X1 U7868 ( .A1(n9439), .A2(n8962), .ZN(n7732) );
  NAND2_X1 U7869 ( .A1(n7732), .A2(n7734), .ZN(n9157) );
  INV_X1 U7870 ( .A(n9439), .ZN(n9162) );
  NAND2_X1 U7871 ( .A1(n7631), .A2(n6210), .ZN(n6095) );
  OR2_X1 U7872 ( .A1(n5844), .A2(n7632), .ZN(n6094) );
  XNOR2_X1 U7873 ( .A(n9134), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U7874 ( .A1(n9143), .A2(n4285), .ZN(n6102) );
  INV_X1 U7875 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7876 ( .A1(n6140), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7877 ( .A1(n7753), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7878 ( .C1(n6099), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6100)
         );
  INV_X1 U7879 ( .A(n6100), .ZN(n6101) );
  NAND2_X1 U7880 ( .A1(n6474), .A2(n9127), .ZN(n7743) );
  NAND2_X1 U7881 ( .A1(n7828), .A2(n7743), .ZN(n7801) );
  NAND2_X1 U7882 ( .A1(n6112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6114) );
  NOR2_X1 U7883 ( .A1(n6229), .A2(n6231), .ZN(n7906) );
  NAND2_X1 U7884 ( .A1(n7900), .A2(n7296), .ZN(n6232) );
  AND2_X1 U7885 ( .A1(n6229), .A2(n6232), .ZN(n6116) );
  OR3_X1 U7886 ( .A1(n7906), .A2(n9687), .A3(n6116), .ZN(n9638) );
  INV_X1 U7887 ( .A(n7296), .ZN(n7905) );
  OR2_X1 U7888 ( .A1(n7760), .A2(n7905), .ZN(n9689) );
  XNOR2_X1 U7889 ( .A(n9380), .B(n8966), .ZN(n9219) );
  INV_X1 U7890 ( .A(n9219), .ZN(n9232) );
  NAND2_X1 U7891 ( .A1(n9453), .A2(n8967), .ZN(n7715) );
  OR2_X1 U7892 ( .A1(n9405), .A2(n8862), .ZN(n7874) );
  NAND2_X1 U7893 ( .A1(n9405), .A2(n8862), .ZN(n7638) );
  INV_X1 U7894 ( .A(n9686), .ZN(n7052) );
  NOR2_X1 U7895 ( .A1(n7043), .A2(n7052), .ZN(n7042) );
  INV_X1 U7896 ( .A(n8983), .ZN(n6656) );
  NAND2_X1 U7897 ( .A1(n6656), .A2(n7053), .ZN(n6118) );
  NAND2_X1 U7898 ( .A1(n6120), .A2(n7838), .ZN(n7646) );
  OR2_X1 U7899 ( .A1(n7646), .A2(n7775), .ZN(n9715) );
  NAND2_X1 U7900 ( .A1(n9715), .A2(n9713), .ZN(n6122) );
  INV_X1 U7901 ( .A(n8980), .ZN(n6942) );
  NAND2_X1 U7902 ( .A1(n6942), .A2(n6267), .ZN(n7651) );
  INV_X1 U7903 ( .A(n6267), .ZN(n10139) );
  NAND2_X1 U7904 ( .A1(n8980), .A2(n10139), .ZN(n7647) );
  NAND2_X1 U7905 ( .A1(n7651), .A2(n7647), .ZN(n9714) );
  INV_X1 U7906 ( .A(n9714), .ZN(n6121) );
  NAND2_X1 U7907 ( .A1(n6122), .A2(n6121), .ZN(n9717) );
  NAND2_X1 U7908 ( .A1(n9717), .A2(n7651), .ZN(n6907) );
  INV_X1 U7909 ( .A(n7650), .ZN(n6123) );
  NAND2_X1 U7910 ( .A1(n7661), .A2(n6963), .ZN(n7660) );
  INV_X1 U7911 ( .A(n7660), .ZN(n6124) );
  OR2_X1 U7912 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND3_X1 U7913 ( .A1(n6961), .A2(n7848), .A3(n7654), .ZN(n6129) );
  AND2_X1 U7914 ( .A1(n6980), .A2(n6127), .ZN(n7771) );
  NAND3_X1 U7915 ( .A1(n7783), .A2(n7771), .A3(n7648), .ZN(n6128) );
  NAND2_X1 U7916 ( .A1(n7848), .A2(n6128), .ZN(n7858) );
  NAND2_X1 U7917 ( .A1(n7233), .A2(n7338), .ZN(n7668) );
  AND2_X1 U7918 ( .A1(n7668), .A2(n7665), .ZN(n7856) );
  OR2_X1 U7919 ( .A1(n7233), .A2(n7338), .ZN(n7674) );
  NAND2_X1 U7920 ( .A1(n6130), .A2(n7674), .ZN(n7269) );
  INV_X1 U7921 ( .A(n7790), .ZN(n7298) );
  INV_X1 U7922 ( .A(n7675), .ZN(n7669) );
  NOR2_X1 U7923 ( .A1(n7298), .A2(n7669), .ZN(n6131) );
  OR2_X1 U7924 ( .A1(n7460), .A2(n6132), .ZN(n7689) );
  AND2_X1 U7925 ( .A1(n7460), .A2(n6132), .ZN(n7864) );
  INV_X1 U7926 ( .A(n7864), .ZN(n6133) );
  NAND2_X1 U7927 ( .A1(n7689), .A2(n6133), .ZN(n7791) );
  NAND2_X1 U7928 ( .A1(n7431), .A2(n7432), .ZN(n7430) );
  OR2_X1 U7929 ( .A1(n9325), .A2(n8937), .ZN(n7698) );
  NAND2_X1 U7930 ( .A1(n9325), .A2(n8937), .ZN(n7697) );
  NAND2_X1 U7931 ( .A1(n9310), .A2(n9309), .ZN(n9308) );
  NAND2_X1 U7932 ( .A1(n9308), .A2(n7638), .ZN(n9293) );
  NOR2_X1 U7933 ( .A1(n9399), .A2(n6134), .ZN(n7876) );
  INV_X1 U7934 ( .A(n7876), .ZN(n7701) );
  NAND2_X1 U7935 ( .A1(n9399), .A2(n6134), .ZN(n7878) );
  NAND2_X1 U7936 ( .A1(n9265), .A2(n7769), .ZN(n7711) );
  NAND2_X1 U7937 ( .A1(n7711), .A2(n9258), .ZN(n7704) );
  NAND2_X1 U7938 ( .A1(n7704), .A2(n7712), .ZN(n7815) );
  OR2_X2 U7939 ( .A1(n9232), .A2(n9231), .ZN(n9229) );
  NAND2_X1 U7940 ( .A1(n9211), .A2(n9235), .ZN(n7817) );
  NAND2_X1 U7941 ( .A1(n7809), .A2(n7817), .ZN(n9202) );
  INV_X1 U7942 ( .A(n8966), .ZN(n7714) );
  NAND2_X1 U7943 ( .A1(n9380), .A2(n7714), .ZN(n9201) );
  NAND3_X1 U7944 ( .A1(n9229), .A2(n9208), .A3(n9201), .ZN(n9205) );
  NAND2_X1 U7945 ( .A1(n9205), .A2(n7809), .ZN(n9186) );
  INV_X1 U7946 ( .A(n8964), .ZN(n6135) );
  NAND2_X1 U7947 ( .A1(n9194), .A2(n6135), .ZN(n7729) );
  NAND2_X1 U7948 ( .A1(n9186), .A2(n9190), .ZN(n9185) );
  XNOR2_X1 U7949 ( .A(n9177), .B(n7724), .ZN(n9175) );
  NAND2_X1 U7950 ( .A1(n9177), .A2(n7724), .ZN(n7733) );
  INV_X1 U7951 ( .A(n7734), .ZN(n6136) );
  NOR2_X1 U7952 ( .A1(n6115), .A2(n7900), .ZN(n7768) );
  NOR2_X1 U7953 ( .A1(n7840), .A2(n7296), .ZN(n7899) );
  AOI211_X1 U7954 ( .C1(n6137), .C2(n7801), .A(n9719), .B(n9121), .ZN(n6150)
         );
  NAND2_X1 U7955 ( .A1(n7909), .A2(n7776), .ZN(n7805) );
  INV_X1 U7956 ( .A(n7805), .ZN(n6146) );
  INV_X1 U7957 ( .A(n6138), .ZN(n8995) );
  INV_X1 U7958 ( .A(n9343), .ZN(n9721) );
  OR2_X1 U7959 ( .A1(n6485), .A2(n9721), .ZN(n6148) );
  NAND2_X1 U7960 ( .A1(n6139), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7961 ( .A1(n7751), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7962 ( .A1(n6140), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7963 ( .A1(n7753), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6141) );
  AND3_X1 U7964 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n6144) );
  OAI21_X1 U7965 ( .B1(n9134), .B2(n6145), .A(n6144), .ZN(n8960) );
  NAND2_X1 U7966 ( .A1(n8960), .A2(n9345), .ZN(n6147) );
  AND2_X1 U7967 ( .A1(n6148), .A2(n6147), .ZN(n6472) );
  INV_X1 U7968 ( .A(n6472), .ZN(n6149) );
  NOR2_X1 U7969 ( .A1(n6150), .A2(n6149), .ZN(n9146) );
  AND2_X1 U7970 ( .A1(n9671), .A2(n5834), .ZN(n9672) );
  NAND2_X1 U7971 ( .A1(n9672), .A2(n9703), .ZN(n9709) );
  OR2_X1 U7972 ( .A1(n9710), .A2(n6952), .ZN(n6909) );
  AND2_X1 U7973 ( .A1(n7019), .A2(n7025), .ZN(n7017) );
  INV_X1 U7974 ( .A(n7178), .ZN(n9727) );
  INV_X1 U7975 ( .A(n6992), .ZN(n9733) );
  INV_X1 U7976 ( .A(n7158), .ZN(n9529) );
  NAND3_X1 U7977 ( .A1(n7125), .A2(n9733), .A3(n9529), .ZN(n7188) );
  OR2_X1 U7978 ( .A1(n7188), .A2(n7233), .ZN(n7187) );
  NOR2_X2 U7979 ( .A1(n7187), .A2(n7275), .ZN(n7305) );
  NAND2_X1 U7980 ( .A1(n9466), .A2(n9336), .ZN(n9322) );
  NAND2_X1 U7981 ( .A1(n6035), .A2(n9287), .ZN(n9279) );
  NAND2_X1 U7982 ( .A1(n9439), .A2(n9176), .ZN(n9159) );
  NAND2_X1 U7983 ( .A1(n9687), .A2(n7296), .ZN(n9740) );
  NAND2_X1 U7984 ( .A1(n6474), .A2(n9159), .ZN(n6151) );
  NAND3_X1 U7985 ( .A1(n9131), .A2(n9711), .A3(n6151), .ZN(n9142) );
  OAI21_X1 U7986 ( .B1(n9150), .B2(n9683), .A(n6153), .ZN(n6186) );
  NAND2_X1 U7987 ( .A1(n4666), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7988 ( .A1(n7601), .A2(P1_B_REG_SCAN_IN), .ZN(n6160) );
  MUX2_X1 U7989 ( .A(n6160), .B(P1_B_REG_SCAN_IN), .S(n6181), .Z(n6163) );
  NAND2_X1 U7990 ( .A1(n6161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  INV_X1 U7991 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6538) );
  INV_X1 U7992 ( .A(n6180), .ZN(n7606) );
  AND2_X1 U7993 ( .A1(n7606), .A2(n7601), .ZN(n6540) );
  INV_X1 U7994 ( .A(n9687), .ZN(n6860) );
  NAND2_X1 U7995 ( .A1(n9416), .A2(n6851), .ZN(n6465) );
  OR2_X1 U7996 ( .A1(n6842), .A2(n6460), .ZN(n6183) );
  NOR2_X1 U7997 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6167) );
  NOR4_X1 U7998 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6166) );
  NOR4_X1 U7999 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6165) );
  NOR4_X1 U8000 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U8001 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n6173)
         );
  NOR4_X1 U8002 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6171) );
  NOR4_X1 U8003 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U8004 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6169) );
  NOR4_X1 U8005 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6168) );
  NAND4_X1 U8006 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n6172)
         );
  OAI21_X1 U8007 ( .B1(n6173), .B2(n6172), .A(n6536), .ZN(n6463) );
  NAND2_X1 U8008 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  NAND2_X1 U8009 ( .A1(n6176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6177) );
  INV_X1 U8010 ( .A(n6547), .ZN(n6178) );
  INV_X1 U8011 ( .A(n7601), .ZN(n6179) );
  INV_X1 U8012 ( .A(n6232), .ZN(n7896) );
  OR2_X1 U8013 ( .A1(n7805), .A2(n7896), .ZN(n6467) );
  AND2_X1 U8014 ( .A1(n7907), .A2(n6467), .ZN(n6182) );
  NAND2_X1 U8015 ( .A1(n6463), .A2(n6182), .ZN(n6841) );
  INV_X1 U8016 ( .A(n6181), .ZN(n7532) );
  INV_X1 U8017 ( .A(n6464), .ZN(n6844) );
  NAND2_X1 U8018 ( .A1(n6187), .A2(n4872), .ZN(P1_U3550) );
  INV_X1 U8019 ( .A(SI_29_), .ZN(n6191) );
  INV_X1 U8020 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6193) );
  INV_X1 U8021 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8223) );
  MUX2_X1 U8022 ( .A(n6193), .B(n8223), .S(n6514), .Z(n6195) );
  INV_X1 U8023 ( .A(SI_30_), .ZN(n6194) );
  NAND2_X1 U8024 ( .A1(n6195), .A2(n6194), .ZN(n6198) );
  INV_X1 U8025 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U8026 ( .A1(n6196), .A2(SI_30_), .ZN(n6197) );
  NAND2_X1 U8027 ( .A1(n6198), .A2(n6197), .ZN(n6206) );
  INV_X1 U8028 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6199) );
  INV_X1 U8029 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6203) );
  MUX2_X1 U8030 ( .A(n6199), .B(n6203), .S(n6513), .Z(n6200) );
  XNOR2_X1 U8031 ( .A(n6200), .B(SI_31_), .ZN(n6201) );
  NAND2_X1 U8032 ( .A1(n8813), .A2(n6210), .ZN(n6205) );
  OR2_X1 U8033 ( .A1(n5844), .A2(n6203), .ZN(n6204) );
  NAND2_X1 U8034 ( .A1(n8221), .A2(n6210), .ZN(n6209) );
  OR2_X1 U8035 ( .A1(n5844), .A2(n8223), .ZN(n6208) );
  OR2_X1 U8036 ( .A1(n5844), .A2(n7629), .ZN(n6211) );
  NOR2_X2 U8037 ( .A1(n9115), .A2(n9132), .ZN(n9114) );
  XOR2_X1 U8038 ( .A(n9109), .B(n9114), .Z(n9113) );
  NOR2_X1 U8039 ( .A1(n9113), .A2(n9740), .ZN(n6223) );
  NAND2_X1 U8040 ( .A1(n7751), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U8041 ( .A1(n7752), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U8042 ( .A1(n7753), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6214) );
  AND3_X1 U8043 ( .A1(n6216), .A2(n6215), .A3(n6214), .ZN(n7758) );
  INV_X1 U8044 ( .A(P1_B_REG_SCAN_IN), .ZN(n6218) );
  OR2_X1 U8045 ( .A1(n8994), .A2(n6218), .ZN(n6219) );
  NAND2_X1 U8046 ( .A1(n9345), .A2(n6219), .ZN(n9124) );
  NOR2_X1 U8047 ( .A1(n7758), .A2(n9124), .ZN(n9353) );
  NOR2_X1 U8048 ( .A1(n9753), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U8049 ( .A1(n6225), .A2(n4288), .ZN(n6228) );
  AND2_X4 U8050 ( .A1(n6226), .A2(n6231), .ZN(n6449) );
  NAND2_X1 U8051 ( .A1(n6235), .A2(n6449), .ZN(n6227) );
  NAND2_X1 U8052 ( .A1(n6228), .A2(n6227), .ZN(n6230) );
  NAND2_X4 U8053 ( .A1(n6229), .A2(n6231), .ZN(n6446) );
  NAND2_X1 U8054 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  NAND2_X1 U8055 ( .A1(n6229), .A2(n6233), .ZN(n6234) );
  AND2_X4 U8056 ( .A1(n6234), .A2(n6226), .ZN(n6443) );
  AOI21_X2 U8057 ( .B1(n8983), .B2(n6443), .A(n6236), .ZN(n6243) );
  NAND2_X1 U8058 ( .A1(n6495), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U8059 ( .A1(n6241), .A2(n6238), .ZN(n6655) );
  NAND2_X1 U8060 ( .A1(n7043), .A2(n6443), .ZN(n6240) );
  AOI22_X1 U8061 ( .A1(n9686), .A2(n6442), .B1(n6495), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U8062 ( .A1(n6240), .A2(n6239), .ZN(n6654) );
  AOI22_X1 U8063 ( .A1(n6655), .A2(n6654), .B1(n6409), .B2(n6241), .ZN(n6661)
         );
  INV_X1 U8064 ( .A(n6242), .ZN(n6244) );
  NAND2_X1 U8065 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  NAND2_X1 U8066 ( .A1(n8982), .A2(n6442), .ZN(n6247) );
  NAND2_X1 U8067 ( .A1(n6249), .A2(n6449), .ZN(n6246) );
  AND2_X1 U8068 ( .A1(n6249), .A2(n6442), .ZN(n6250) );
  AOI21_X1 U8069 ( .B1(n8982), .B2(n6443), .A(n6250), .ZN(n6252) );
  XNOR2_X1 U8070 ( .A(n6251), .B(n6252), .ZN(n6630) );
  NAND2_X1 U8071 ( .A1(n6629), .A2(n6630), .ZN(n6255) );
  INV_X1 U8072 ( .A(n6251), .ZN(n6253) );
  NAND2_X1 U8073 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  INV_X4 U8074 ( .A(n6433), .ZN(n6442) );
  NAND2_X1 U8075 ( .A1(n8981), .A2(n6442), .ZN(n6257) );
  NAND2_X1 U8076 ( .A1(n6943), .A2(n6449), .ZN(n6256) );
  NAND2_X1 U8077 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  XNOR2_X1 U8078 ( .A(n6258), .B(n6446), .ZN(n6260) );
  AND2_X1 U8079 ( .A1(n6943), .A2(n6442), .ZN(n6259) );
  AOI21_X1 U8080 ( .B1(n8981), .B2(n6443), .A(n6259), .ZN(n6261) );
  INV_X1 U8081 ( .A(n6260), .ZN(n6262) );
  NAND2_X1 U8082 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U8083 ( .A1(n8980), .A2(n6442), .ZN(n6265) );
  NAND2_X1 U8084 ( .A1(n6267), .A2(n6449), .ZN(n6264) );
  NAND2_X1 U8085 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U8086 ( .A1(n8980), .A2(n6443), .ZN(n6269) );
  NAND2_X1 U8087 ( .A1(n6267), .A2(n6442), .ZN(n6268) );
  NAND2_X1 U8088 ( .A1(n6269), .A2(n6268), .ZN(n6271) );
  INV_X1 U8089 ( .A(n6270), .ZN(n6273) );
  INV_X1 U8090 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U8091 ( .A1(n8979), .A2(n6442), .ZN(n6275) );
  NAND2_X1 U8092 ( .A1(n6952), .A2(n6449), .ZN(n6274) );
  NAND2_X1 U8093 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  XNOR2_X1 U8094 ( .A(n6276), .B(n6446), .ZN(n6279) );
  AOI22_X1 U8095 ( .A1(n8979), .A2(n6443), .B1(n6952), .B2(n6448), .ZN(n6775)
         );
  INV_X1 U8096 ( .A(n6277), .ZN(n6278) );
  NOR2_X1 U8097 ( .A1(n6279), .A2(n6278), .ZN(n6281) );
  NAND2_X1 U8098 ( .A1(n6282), .A2(n6773), .ZN(n6828) );
  NAND2_X1 U8099 ( .A1(n6852), .A2(n6449), .ZN(n6284) );
  NAND2_X1 U8100 ( .A1(n8978), .A2(n6442), .ZN(n6283) );
  NAND2_X1 U8101 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  XNOR2_X1 U8102 ( .A(n6285), .B(n6446), .ZN(n6286) );
  AOI22_X1 U8103 ( .A1(n6852), .A2(n6442), .B1(n8978), .B2(n6443), .ZN(n6287)
         );
  XNOR2_X1 U8104 ( .A(n6286), .B(n6287), .ZN(n6829) );
  NAND2_X1 U8105 ( .A1(n6828), .A2(n6829), .ZN(n6290) );
  INV_X1 U8106 ( .A(n6286), .ZN(n6288) );
  NAND2_X1 U8107 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  NAND2_X1 U8108 ( .A1(n9651), .A2(n6449), .ZN(n6292) );
  NAND2_X1 U8109 ( .A1(n8977), .A2(n6442), .ZN(n6291) );
  NAND2_X1 U8110 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  XNOR2_X1 U8111 ( .A(n6293), .B(n6409), .ZN(n7033) );
  AND2_X1 U8112 ( .A1(n8977), .A2(n6443), .ZN(n6294) );
  AOI21_X1 U8113 ( .B1(n9651), .B2(n6442), .A(n6294), .ZN(n7032) );
  AND2_X1 U8114 ( .A1(n7033), .A2(n7032), .ZN(n6298) );
  INV_X1 U8115 ( .A(n7033), .ZN(n6296) );
  INV_X1 U8116 ( .A(n7032), .ZN(n6295) );
  NAND2_X1 U8117 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  NAND2_X1 U8118 ( .A1(n7178), .A2(n6449), .ZN(n6300) );
  NAND2_X1 U8119 ( .A1(n8976), .A2(n6442), .ZN(n6299) );
  NAND2_X1 U8120 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  XNOR2_X1 U8121 ( .A(n6301), .B(n6446), .ZN(n7167) );
  NAND2_X1 U8122 ( .A1(n7178), .A2(n6442), .ZN(n6303) );
  NAND2_X1 U8123 ( .A1(n8976), .A2(n6443), .ZN(n6302) );
  NAND2_X1 U8124 ( .A1(n6303), .A2(n6302), .ZN(n7171) );
  AND2_X1 U8125 ( .A1(n7167), .A2(n7171), .ZN(n6311) );
  NAND2_X1 U8126 ( .A1(n6992), .A2(n6449), .ZN(n6305) );
  NAND2_X1 U8127 ( .A1(n8975), .A2(n6442), .ZN(n6304) );
  NAND2_X1 U8128 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  XNOR2_X1 U8129 ( .A(n6306), .B(n6446), .ZN(n7198) );
  NAND2_X1 U8130 ( .A1(n6992), .A2(n6442), .ZN(n6308) );
  NAND2_X1 U8131 ( .A1(n8975), .A2(n6443), .ZN(n6307) );
  NAND2_X1 U8132 ( .A1(n6308), .A2(n6307), .ZN(n6312) );
  OAI22_X1 U8133 ( .A1(n7198), .A2(n6312), .B1(n7171), .B2(n7167), .ZN(n6309)
         );
  INV_X1 U8134 ( .A(n6309), .ZN(n6310) );
  INV_X1 U8135 ( .A(n6312), .ZN(n7197) );
  AOI22_X1 U8136 ( .A1(n7158), .A2(n6449), .B1(n6448), .B2(n8974), .ZN(n6313)
         );
  XOR2_X1 U8137 ( .A(n6446), .B(n6313), .Z(n6314) );
  AOI22_X1 U8138 ( .A1(n7158), .A2(n6448), .B1(n6443), .B2(n8974), .ZN(n9522)
         );
  INV_X1 U8139 ( .A(n6315), .ZN(n7286) );
  NAND2_X1 U8140 ( .A1(n7233), .A2(n6449), .ZN(n6317) );
  NAND2_X1 U8141 ( .A1(n8973), .A2(n6442), .ZN(n6316) );
  NAND2_X1 U8142 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  XNOR2_X1 U8143 ( .A(n6318), .B(n6409), .ZN(n6320) );
  AND2_X1 U8144 ( .A1(n8973), .A2(n6443), .ZN(n6319) );
  AOI21_X1 U8145 ( .B1(n7233), .B2(n6442), .A(n6319), .ZN(n6321) );
  NAND2_X1 U8146 ( .A1(n6320), .A2(n6321), .ZN(n6325) );
  INV_X1 U8147 ( .A(n6320), .ZN(n6323) );
  INV_X1 U8148 ( .A(n6321), .ZN(n6322) );
  NAND2_X1 U8149 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U8150 ( .A1(n6325), .A2(n6324), .ZN(n7285) );
  INV_X1 U8151 ( .A(n6325), .ZN(n7333) );
  NAND2_X1 U8152 ( .A1(n7275), .A2(n6449), .ZN(n6327) );
  NAND2_X1 U8153 ( .A1(n8972), .A2(n6448), .ZN(n6326) );
  NAND2_X1 U8154 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  XNOR2_X1 U8155 ( .A(n6328), .B(n6409), .ZN(n6330) );
  AND2_X1 U8156 ( .A1(n8972), .A2(n6443), .ZN(n6329) );
  AOI21_X1 U8157 ( .B1(n5966), .B2(n6442), .A(n6329), .ZN(n6331) );
  NAND2_X1 U8158 ( .A1(n6330), .A2(n6331), .ZN(n6335) );
  INV_X1 U8159 ( .A(n6330), .ZN(n6333) );
  INV_X1 U8160 ( .A(n6331), .ZN(n6332) );
  NAND2_X1 U8161 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  AND2_X1 U8162 ( .A1(n6335), .A2(n6334), .ZN(n7332) );
  NAND2_X1 U8163 ( .A1(n6339), .A2(n6449), .ZN(n6337) );
  NAND2_X1 U8164 ( .A1(n8971), .A2(n6442), .ZN(n6336) );
  NAND2_X1 U8165 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  XNOR2_X1 U8166 ( .A(n6338), .B(n6446), .ZN(n6340) );
  AOI22_X1 U8167 ( .A1(n6339), .A2(n6442), .B1(n6443), .B2(n8971), .ZN(n6341)
         );
  XNOR2_X1 U8168 ( .A(n6340), .B(n6341), .ZN(n7391) );
  INV_X1 U8169 ( .A(n6340), .ZN(n6342) );
  NAND2_X1 U8170 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  NAND2_X1 U8171 ( .A1(n7389), .A2(n6343), .ZN(n6346) );
  AOI22_X1 U8172 ( .A1(n9430), .A2(n6449), .B1(n6442), .B2(n8970), .ZN(n6344)
         );
  XNOR2_X1 U8173 ( .A(n6344), .B(n6446), .ZN(n6345) );
  INV_X1 U8174 ( .A(n6443), .ZN(n6432) );
  OAI22_X1 U8175 ( .A1(n9642), .A2(n6433), .B1(n6347), .B2(n6432), .ZN(n8840)
         );
  INV_X1 U8176 ( .A(n6348), .ZN(n6349) );
  AOI22_X1 U8177 ( .A1(n7460), .A2(n6449), .B1(n6442), .B2(n9344), .ZN(n6350)
         );
  XOR2_X1 U8178 ( .A(n6446), .B(n6350), .Z(n6351) );
  AOI22_X1 U8179 ( .A1(n7460), .A2(n6448), .B1(n6443), .B2(n9344), .ZN(n8948)
         );
  NAND2_X1 U8180 ( .A1(n8947), .A2(n4338), .ZN(n8889) );
  NAND2_X1 U8181 ( .A1(n9415), .A2(n6449), .ZN(n6353) );
  NAND2_X1 U8182 ( .A1(n8969), .A2(n6448), .ZN(n6352) );
  NAND2_X1 U8183 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  XNOR2_X1 U8184 ( .A(n6354), .B(n6446), .ZN(n6357) );
  AOI22_X1 U8185 ( .A1(n9415), .A2(n4288), .B1(n6443), .B2(n8969), .ZN(n6355)
         );
  XNOR2_X1 U8186 ( .A(n6357), .B(n6355), .ZN(n8890) );
  NAND2_X1 U8187 ( .A1(n8889), .A2(n8890), .ZN(n8888) );
  INV_X1 U8188 ( .A(n6355), .ZN(n6356) );
  NAND2_X1 U8189 ( .A1(n8888), .A2(n6358), .ZN(n8899) );
  NAND2_X1 U8190 ( .A1(n9325), .A2(n6449), .ZN(n6360) );
  NAND2_X1 U8191 ( .A1(n9346), .A2(n4288), .ZN(n6359) );
  NAND2_X1 U8192 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  XNOR2_X1 U8193 ( .A(n6361), .B(n6446), .ZN(n6364) );
  NAND2_X1 U8194 ( .A1(n9325), .A2(n6442), .ZN(n6363) );
  NAND2_X1 U8195 ( .A1(n9346), .A2(n6443), .ZN(n6362) );
  NAND2_X1 U8196 ( .A1(n6363), .A2(n6362), .ZN(n6365) );
  NAND2_X1 U8197 ( .A1(n6364), .A2(n6365), .ZN(n8900) );
  INV_X1 U8198 ( .A(n6364), .ZN(n6367) );
  INV_X1 U8199 ( .A(n6365), .ZN(n6366) );
  NAND2_X1 U8200 ( .A1(n6367), .A2(n6366), .ZN(n8902) );
  NAND2_X1 U8201 ( .A1(n9405), .A2(n6449), .ZN(n6369) );
  NAND2_X1 U8202 ( .A1(n9295), .A2(n6442), .ZN(n6368) );
  NAND2_X1 U8203 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  XNOR2_X1 U8204 ( .A(n6370), .B(n6446), .ZN(n8933) );
  NAND2_X1 U8205 ( .A1(n9405), .A2(n6448), .ZN(n6372) );
  NAND2_X1 U8206 ( .A1(n9295), .A2(n6443), .ZN(n6371) );
  NAND2_X1 U8207 ( .A1(n6372), .A2(n6371), .ZN(n8932) );
  INV_X1 U8208 ( .A(n8933), .ZN(n6374) );
  INV_X1 U8209 ( .A(n8932), .ZN(n6373) );
  NAND2_X1 U8210 ( .A1(n9399), .A2(n6449), .ZN(n6376) );
  NAND2_X1 U8211 ( .A1(n9311), .A2(n6448), .ZN(n6375) );
  NAND2_X1 U8212 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  XNOR2_X1 U8213 ( .A(n6377), .B(n6409), .ZN(n8858) );
  AND2_X1 U8214 ( .A1(n9311), .A2(n6443), .ZN(n6378) );
  AOI21_X1 U8215 ( .B1(n9399), .B2(n6448), .A(n6378), .ZN(n8859) );
  NAND2_X1 U8216 ( .A1(n8858), .A2(n8859), .ZN(n6379) );
  INV_X1 U8217 ( .A(n6449), .ZN(n6430) );
  OAI22_X1 U8218 ( .A1(n6035), .A2(n6430), .B1(n8871), .B2(n6433), .ZN(n6380)
         );
  XNOR2_X1 U8219 ( .A(n6380), .B(n6446), .ZN(n6382) );
  OAI22_X1 U8220 ( .A1(n6035), .A2(n6433), .B1(n8871), .B2(n6432), .ZN(n6381)
         );
  NOR2_X1 U8221 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  AOI21_X1 U8222 ( .B1(n6382), .B2(n6381), .A(n6383), .ZN(n8917) );
  NAND2_X1 U8223 ( .A1(n9265), .A2(n6449), .ZN(n6385) );
  NAND2_X1 U8224 ( .A1(n8968), .A2(n6442), .ZN(n6384) );
  NAND2_X1 U8225 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  XNOR2_X1 U8226 ( .A(n6386), .B(n6446), .ZN(n6387) );
  AOI22_X1 U8227 ( .A1(n9265), .A2(n6442), .B1(n6443), .B2(n8968), .ZN(n6388)
         );
  XNOR2_X1 U8228 ( .A(n6387), .B(n6388), .ZN(n8870) );
  INV_X1 U8229 ( .A(n6387), .ZN(n6389) );
  NAND2_X1 U8230 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U8231 ( .A1(n8868), .A2(n6390), .ZN(n6395) );
  INV_X1 U8232 ( .A(n6395), .ZN(n6393) );
  OAI22_X1 U8233 ( .A1(n9453), .A2(n6430), .B1(n4292), .B2(n6433), .ZN(n6391)
         );
  XOR2_X1 U8234 ( .A(n6446), .B(n6391), .Z(n6394) );
  INV_X1 U8235 ( .A(n6394), .ZN(n6392) );
  OAI22_X1 U8236 ( .A1(n9453), .A2(n6433), .B1(n4292), .B2(n6432), .ZN(n8926)
         );
  NAND2_X1 U8237 ( .A1(n9380), .A2(n6449), .ZN(n6398) );
  NAND2_X1 U8238 ( .A1(n8966), .A2(n4288), .ZN(n6397) );
  NAND2_X1 U8239 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  XNOR2_X1 U8240 ( .A(n6399), .B(n6409), .ZN(n6401) );
  AND2_X1 U8241 ( .A1(n8966), .A2(n6443), .ZN(n6400) );
  AOI21_X1 U8242 ( .B1(n9380), .B2(n6442), .A(n6400), .ZN(n6402) );
  NAND2_X1 U8243 ( .A1(n6401), .A2(n6402), .ZN(n8913) );
  INV_X1 U8244 ( .A(n6401), .ZN(n6404) );
  INV_X1 U8245 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U8246 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U8247 ( .A1(n9211), .A2(n6449), .ZN(n6408) );
  NAND2_X1 U8248 ( .A1(n8965), .A2(n6448), .ZN(n6407) );
  NAND2_X1 U8249 ( .A1(n6408), .A2(n6407), .ZN(n6410) );
  XNOR2_X1 U8250 ( .A(n6410), .B(n6409), .ZN(n6412) );
  AND2_X1 U8251 ( .A1(n8965), .A2(n6443), .ZN(n6411) );
  AOI21_X1 U8252 ( .B1(n9211), .B2(n6442), .A(n6411), .ZN(n6413) );
  NAND2_X1 U8253 ( .A1(n6412), .A2(n6413), .ZN(n6418) );
  INV_X1 U8254 ( .A(n6412), .ZN(n6415) );
  INV_X1 U8255 ( .A(n6413), .ZN(n6414) );
  NAND2_X1 U8256 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  AND2_X1 U8257 ( .A1(n6418), .A2(n6416), .ZN(n8912) );
  NAND2_X1 U8258 ( .A1(n9194), .A2(n6449), .ZN(n6420) );
  NAND2_X1 U8259 ( .A1(n8964), .A2(n6448), .ZN(n6419) );
  NAND2_X1 U8260 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  XNOR2_X1 U8261 ( .A(n6421), .B(n6446), .ZN(n6426) );
  AOI22_X1 U8262 ( .A1(n9194), .A2(n4288), .B1(n6443), .B2(n8964), .ZN(n6427)
         );
  NAND2_X1 U8263 ( .A1(n9177), .A2(n6449), .ZN(n6423) );
  NAND2_X1 U8264 ( .A1(n8963), .A2(n4288), .ZN(n6422) );
  NAND2_X1 U8265 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  XNOR2_X1 U8266 ( .A(n6424), .B(n6446), .ZN(n6438) );
  AND2_X1 U8267 ( .A1(n8963), .A2(n6443), .ZN(n6425) );
  AOI21_X1 U8268 ( .B1(n9177), .B2(n6442), .A(n6425), .ZN(n6436) );
  XNOR2_X1 U8269 ( .A(n6438), .B(n6436), .ZN(n6483) );
  INV_X1 U8270 ( .A(n6426), .ZN(n6428) );
  NAND2_X1 U8271 ( .A1(n6428), .A2(n6427), .ZN(n6482) );
  NAND2_X2 U8272 ( .A1(n6481), .A2(n6429), .ZN(n8830) );
  OAI22_X1 U8273 ( .A1(n9439), .A2(n6430), .B1(n6485), .B2(n6433), .ZN(n6431)
         );
  XNOR2_X1 U8274 ( .A(n6431), .B(n6446), .ZN(n6435) );
  OAI22_X1 U8275 ( .A1(n9439), .A2(n6433), .B1(n6485), .B2(n6432), .ZN(n6434)
         );
  NOR2_X1 U8276 ( .A1(n6435), .A2(n6434), .ZN(n6457) );
  AOI21_X1 U8277 ( .B1(n6435), .B2(n6434), .A(n6457), .ZN(n8828) );
  INV_X1 U8278 ( .A(n8828), .ZN(n6440) );
  INV_X1 U8279 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U8280 ( .A1(n6438), .A2(n6437), .ZN(n8829) );
  INV_X1 U8281 ( .A(n8829), .ZN(n6439) );
  NOR2_X1 U8282 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  AND2_X2 U8283 ( .A1(n8830), .A2(n6441), .ZN(n8832) );
  INV_X1 U8284 ( .A(n8832), .ZN(n6456) );
  NAND2_X1 U8285 ( .A1(n6474), .A2(n4288), .ZN(n6445) );
  NAND2_X1 U8286 ( .A1(n8961), .A2(n6443), .ZN(n6444) );
  NAND2_X1 U8287 ( .A1(n6445), .A2(n6444), .ZN(n6447) );
  XNOR2_X1 U8288 ( .A(n6447), .B(n6446), .ZN(n6451) );
  AOI22_X1 U8289 ( .A1(n6474), .A2(n6449), .B1(n6442), .B2(n8961), .ZN(n6450)
         );
  XNOR2_X1 U8290 ( .A(n6451), .B(n6450), .ZN(n6458) );
  INV_X1 U8291 ( .A(n6458), .ZN(n6455) );
  INV_X1 U8292 ( .A(n6457), .ZN(n6454) );
  AND2_X1 U8293 ( .A1(n6463), .A2(n7907), .ZN(n6452) );
  AND3_X1 U8294 ( .A1(n6452), .A2(n6464), .A3(n6842), .ZN(n6462) );
  INV_X1 U8295 ( .A(n9416), .ZN(n9748) );
  AND2_X1 U8296 ( .A1(n9748), .A2(n7805), .ZN(n6453) );
  NAND2_X1 U8297 ( .A1(n6456), .A2(n4876), .ZN(n6480) );
  NAND3_X1 U8298 ( .A1(n6458), .A2(n9531), .A3(n6457), .ZN(n6476) );
  INV_X1 U8299 ( .A(n6851), .ZN(n6459) );
  NAND2_X1 U8300 ( .A1(n6462), .A2(n6459), .ZN(n6461) );
  NAND2_X1 U8301 ( .A1(n6462), .A2(n7896), .ZN(n8952) );
  NAND3_X1 U8302 ( .A1(n6842), .A2(n6464), .A3(n6463), .ZN(n6466) );
  NAND2_X1 U8303 ( .A1(n6466), .A2(n6465), .ZN(n6469) );
  AND2_X1 U8304 ( .A1(n6467), .A2(n6226), .ZN(n6468) );
  NAND2_X1 U8305 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  AND2_X1 U8306 ( .A1(n6547), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7484) );
  AOI21_X2 U8307 ( .B1(n6470), .B2(P1_STATE_REG_SCAN_IN), .A(n7484), .ZN(n9535) );
  AOI22_X1 U8308 ( .A1(n9143), .A2(n8955), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6471) );
  OAI21_X1 U8309 ( .B1(n6472), .B2(n8952), .A(n6471), .ZN(n6473) );
  AOI21_X1 U8310 ( .B1(n6474), .B2(n8943), .A(n6473), .ZN(n6475) );
  NAND2_X1 U8311 ( .A1(n6480), .A2(n6479), .ZN(P1_U3220) );
  AND2_X1 U8312 ( .A1(n6481), .A2(n6482), .ZN(n6484) );
  NAND2_X1 U8313 ( .A1(n8830), .A2(n9531), .ZN(n6493) );
  OR2_X1 U8314 ( .A1(n6485), .A2(n9723), .ZN(n6487) );
  NAND2_X1 U8315 ( .A1(n8964), .A2(n9343), .ZN(n6486) );
  NAND2_X1 U8316 ( .A1(n6487), .A2(n6486), .ZN(n9171) );
  INV_X1 U8317 ( .A(n8952), .ZN(n9526) );
  OAI22_X1 U8318 ( .A1(n9178), .A2(n9535), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6488), .ZN(n6489) );
  AOI21_X1 U8319 ( .B1(n9171), .B2(n9526), .A(n6489), .ZN(n6490) );
  INV_X1 U8320 ( .A(n6491), .ZN(n6492) );
  OAI21_X1 U8321 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(P1_U3240) );
  XNOR2_X1 U8322 ( .A(n6498), .B(n6497), .ZN(n6499) );
  NOR2_X1 U8323 ( .A1(n6499), .A2(n9826), .ZN(n6511) );
  NOR2_X1 U8324 ( .A1(n9835), .A2(n6527), .ZN(n6510) );
  INV_X1 U8325 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10001) );
  NOR2_X1 U8326 ( .A1(n9832), .A2(n10001), .ZN(n6509) );
  NAND2_X1 U8327 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  AND2_X1 U8328 ( .A1(n6725), .A2(n6502), .ZN(n6507) );
  NAND2_X1 U8329 ( .A1(n6503), .A2(n9943), .ZN(n6504) );
  NAND2_X1 U8330 ( .A1(n6731), .A2(n6504), .ZN(n6505) );
  NAND2_X1 U8331 ( .A1(n9821), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U8332 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7111) );
  OAI211_X1 U8333 ( .C1(n6507), .C2(n9848), .A(n6506), .B(n7111), .ZN(n6508)
         );
  OR4_X1 U8334 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(P2_U3187)
         );
  XNOR2_X1 U8335 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U8336 ( .A(n8823), .ZN(n7528) );
  OR2_X2 U8337 ( .A1(n6513), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8825) );
  OAI222_X1 U8338 ( .A1(n7528), .A2(n5137), .B1(n6512), .B2(P2_U3151), .C1(
        n8825), .C2(n6515), .ZN(P2_U3293) );
  OR2_X2 U8339 ( .A1(n6513), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8222) );
  AND2_X1 U8340 ( .A1(n6514), .A2(P1_U3086), .ZN(n7482) );
  INV_X2 U8341 ( .A(n7482), .ZN(n9478) );
  OAI222_X1 U8342 ( .A1(n8222), .A2(n6516), .B1(n9478), .B2(n6515), .C1(
        P1_U3086), .C2(n9003), .ZN(P1_U3353) );
  OAI222_X1 U8343 ( .A1(n8222), .A2(n6517), .B1(n9478), .B2(n6522), .C1(
        P1_U3086), .C2(n6599), .ZN(P1_U3354) );
  OAI222_X1 U8344 ( .A1(n8222), .A2(n5161), .B1(n9478), .B2(n6518), .C1(
        P1_U3086), .C2(n9019), .ZN(P1_U3352) );
  OAI222_X1 U8345 ( .A1(n7528), .A2(n5156), .B1(n6695), .B2(P2_U3151), .C1(
        n8825), .C2(n6518), .ZN(P2_U3292) );
  OAI222_X1 U8346 ( .A1(n9030), .A2(P1_U3086), .B1(n8222), .B2(n5857), .C1(
        n6519), .C2(n9478), .ZN(P1_U3351) );
  INV_X1 U8347 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6521) );
  OAI222_X1 U8348 ( .A1(n7528), .A2(n6521), .B1(n6520), .B2(P2_U3151), .C1(
        n8825), .C2(n6519), .ZN(P2_U3291) );
  OAI222_X1 U8349 ( .A1(n7528), .A2(n5107), .B1(n6523), .B2(P2_U3151), .C1(
        n8825), .C2(n6522), .ZN(P2_U3294) );
  OAI222_X1 U8350 ( .A1(P1_U3086), .A2(n6525), .B1(n9478), .B2(n6526), .C1(
        n6524), .C2(n8222), .ZN(P1_U3350) );
  OAI222_X1 U8351 ( .A1(n7528), .A2(n6528), .B1(n6527), .B2(P2_U3151), .C1(
        n8825), .C2(n6526), .ZN(P2_U3290) );
  INV_X1 U8352 ( .A(n6607), .ZN(n9562) );
  INV_X1 U8353 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6529) );
  OAI222_X1 U8354 ( .A1(P1_U3086), .A2(n9562), .B1(n9478), .B2(n6530), .C1(
        n6529), .C2(n8222), .ZN(P1_U3349) );
  INV_X1 U8355 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6532) );
  OAI222_X1 U8356 ( .A1(n7528), .A2(n6532), .B1(n6531), .B2(P2_U3151), .C1(
        n8825), .C2(n6530), .ZN(P2_U3289) );
  OAI222_X1 U8357 ( .A1(n8825), .A2(n6533), .B1(n4587), .B2(P2_U3151), .C1(
        n4417), .C2(n7528), .ZN(P2_U3288) );
  INV_X1 U8358 ( .A(n6610), .ZN(n9502) );
  INV_X1 U8359 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10092) );
  OAI222_X1 U8360 ( .A1(P1_U3086), .A2(n9502), .B1(n9478), .B2(n6533), .C1(
        n10092), .C2(n8222), .ZN(P1_U3348) );
  NAND2_X1 U8361 ( .A1(n6535), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6534) );
  OAI21_X1 U8362 ( .B1(n6812), .B2(n6535), .A(n6534), .ZN(P2_U3377) );
  INV_X1 U8363 ( .A(n6536), .ZN(n6537) );
  OR2_X1 U8364 ( .A1(n9678), .A2(n6538), .ZN(n6539) );
  OAI21_X1 U8365 ( .B1(n9679), .B2(n6540), .A(n6539), .ZN(P1_U3440) );
  NAND2_X1 U8366 ( .A1(n9679), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U8367 ( .B1(n9679), .B2(n6542), .A(n6541), .ZN(P1_U3439) );
  INV_X1 U8368 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10121) );
  INV_X1 U8369 ( .A(n6543), .ZN(n6546) );
  OAI222_X1 U8370 ( .A1(n7528), .A2(n10121), .B1(n8825), .B2(n6546), .C1(
        P2_U3151), .C2(n6544), .ZN(P2_U3287) );
  INV_X1 U8371 ( .A(n6612), .ZN(n9516) );
  INV_X1 U8372 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6545) );
  OAI222_X1 U8373 ( .A1(n9516), .A2(P1_U3086), .B1(n9478), .B2(n6546), .C1(
        n6545), .C2(n8222), .ZN(P1_U3347) );
  OR2_X1 U8374 ( .A1(n6547), .A2(n7805), .ZN(n6549) );
  AND2_X1 U8375 ( .A1(n6549), .A2(n6548), .ZN(n6551) );
  INV_X1 U8376 ( .A(n6551), .ZN(n6550) );
  INV_X1 U8377 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6558) );
  AND2_X1 U8378 ( .A1(n6552), .A2(n6551), .ZN(n6615) );
  INV_X1 U8379 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6554) );
  NOR2_X1 U8380 ( .A1(n8994), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6553) );
  OR2_X1 U8381 ( .A1(n6138), .A2(n6553), .ZN(n8996) );
  AOI21_X1 U8382 ( .B1(n8994), .B2(n6554), .A(n8996), .ZN(n6555) );
  INV_X1 U8383 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8997) );
  XNOR2_X1 U8384 ( .A(n6555), .B(n8997), .ZN(n6556) );
  AOI22_X1 U8385 ( .A1(n6615), .A2(n6556), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6557) );
  OAI21_X1 U8386 ( .B1(n9635), .B2(n6558), .A(n6557), .ZN(P1_U3243) );
  INV_X1 U8387 ( .A(n9635), .ZN(n9076) );
  NOR2_X1 U8388 ( .A1(n9076), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8389 ( .A1(n7043), .A2(P1_U3973), .ZN(n6559) );
  OAI21_X1 U8390 ( .B1(P1_U3973), .B2(n5109), .A(n6559), .ZN(P1_U3554) );
  INV_X1 U8391 ( .A(n7758), .ZN(n7757) );
  NAND2_X1 U8392 ( .A1(n7757), .A2(P1_U3973), .ZN(n6560) );
  OAI21_X1 U8393 ( .B1(P1_U3973), .B2(n6199), .A(n6560), .ZN(P1_U3585) );
  INV_X1 U8394 ( .A(n7093), .ZN(n6561) );
  AOI22_X1 U8395 ( .A1(n6565), .A2(n5690), .B1(n6562), .B2(n6561), .ZN(
        P2_U3376) );
  AND2_X1 U8396 ( .A1(n6565), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8397 ( .A1(n6565), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8398 ( .A1(n6565), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8399 ( .A1(n6565), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8400 ( .A1(n6565), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8401 ( .A1(n6565), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8402 ( .A1(n6565), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8403 ( .A1(n6565), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8404 ( .A1(n6565), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8405 ( .A1(n6565), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8406 ( .A1(n6565), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8407 ( .A1(n6565), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8408 ( .A1(n6565), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8409 ( .A1(n6565), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8410 ( .A1(n6565), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8411 ( .A1(n6565), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8412 ( .A1(n6565), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8413 ( .A1(n6565), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8414 ( .A1(n6565), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8415 ( .A1(n6565), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8416 ( .A1(n6565), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8417 ( .A1(n6565), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8418 ( .A1(n6565), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8419 ( .A1(n6565), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8420 ( .A1(n6565), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8421 ( .A1(n6565), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  INV_X1 U8422 ( .A(n6563), .ZN(n6571) );
  AOI22_X1 U8423 ( .A1(n9816), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8823), .ZN(n6564) );
  OAI21_X1 U8424 ( .B1(n6571), .B2(n8825), .A(n6564), .ZN(P2_U3286) );
  INV_X1 U8425 ( .A(n6565), .ZN(n6566) );
  INV_X1 U8426 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U8427 ( .A1(n6566), .A2(n10066), .ZN(P2_U3248) );
  INV_X1 U8428 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U8429 ( .A1(n6566), .A2(n10067), .ZN(P2_U3253) );
  INV_X1 U8430 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U8431 ( .A1(n6566), .A2(n10040), .ZN(P2_U3245) );
  INV_X1 U8432 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U8433 ( .A1(n6566), .A2(n10128), .ZN(P2_U3255) );
  INV_X1 U8434 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6567) );
  OAI222_X1 U8435 ( .A1(n8825), .A2(n6570), .B1(n6568), .B2(P2_U3151), .C1(
        n6567), .C2(n7528), .ZN(P2_U3285) );
  INV_X1 U8436 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6569) );
  OAI222_X1 U8437 ( .A1(P1_U3086), .A2(n6791), .B1(n9478), .B2(n6570), .C1(
        n6569), .C2(n8222), .ZN(P1_U3345) );
  INV_X1 U8438 ( .A(n6790), .ZN(n6617) );
  OAI222_X1 U8439 ( .A1(P1_U3086), .A2(n6617), .B1(n9478), .B2(n6571), .C1(
        n10109), .C2(n8222), .ZN(P1_U3346) );
  INV_X1 U8440 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U8441 ( .A1(n6572), .A2(n9826), .ZN(n6576) );
  OAI21_X1 U8442 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6574), .A(n6573), .ZN(n6575) );
  AOI22_X1 U8443 ( .A1(n6576), .A2(n6575), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6578) );
  NAND2_X1 U8444 ( .A1(n9817), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6577) );
  OAI211_X1 U8445 ( .C1(n9832), .C2(n6579), .A(n6578), .B(n6577), .ZN(P2_U3182) );
  INV_X1 U8446 ( .A(n6580), .ZN(n6623) );
  AOI22_X1 U8447 ( .A1(n9575), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9476), .ZN(n6581) );
  OAI21_X1 U8448 ( .B1(n6623), .B2(n9478), .A(n6581), .ZN(P1_U3344) );
  NOR2_X1 U8449 ( .A1(n6790), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6582) );
  AOI21_X1 U8450 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6790), .A(n6582), .ZN(
        n6597) );
  XNOR2_X1 U8451 ( .A(n9003), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9012) );
  INV_X1 U8452 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6583) );
  MUX2_X1 U8453 ( .A(n6583), .B(P1_REG2_REG_1__SCAN_IN), .S(n6599), .Z(n8989)
         );
  AND2_X1 U8454 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8998) );
  NAND2_X1 U8455 ( .A1(n8989), .A2(n8998), .ZN(n8988) );
  INV_X1 U8456 ( .A(n6599), .ZN(n8987) );
  NAND2_X1 U8457 ( .A1(n8987), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6584) );
  INV_X1 U8458 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6585) );
  OR2_X1 U8459 ( .A1(n9003), .A2(n6585), .ZN(n6586) );
  NAND2_X1 U8460 ( .A1(n9010), .A2(n6586), .ZN(n9025) );
  XNOR2_X1 U8461 ( .A(n9019), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U8462 ( .A1(n9025), .A2(n9026), .ZN(n9024) );
  INV_X1 U8463 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6587) );
  OR2_X1 U8464 ( .A1(n9019), .A2(n6587), .ZN(n6588) );
  NAND2_X1 U8465 ( .A1(n9024), .A2(n6588), .ZN(n9036) );
  INV_X1 U8466 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6589) );
  MUX2_X1 U8467 ( .A(n6589), .B(P1_REG2_REG_4__SCAN_IN), .S(n9030), .Z(n9037)
         );
  NAND2_X1 U8468 ( .A1(n9036), .A2(n9037), .ZN(n9035) );
  OR2_X1 U8469 ( .A1(n9030), .A2(n6589), .ZN(n6590) );
  NAND2_X1 U8470 ( .A1(n9035), .A2(n6590), .ZN(n9540) );
  OR2_X1 U8471 ( .A1(n9542), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8472 ( .A1(n9542), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6591) );
  AND2_X1 U8473 ( .A1(n6592), .A2(n6591), .ZN(n9541) );
  AND2_X1 U8474 ( .A1(n9540), .A2(n9541), .ZN(n9538) );
  INV_X1 U8475 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U8476 ( .A1(n6607), .A2(n6593), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9562), .ZN(n9554) );
  NOR2_X1 U8477 ( .A1(n9553), .A2(n9554), .ZN(n9552) );
  AOI21_X1 U8478 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6607), .A(n9552), .ZN(
        n9493) );
  NAND2_X1 U8479 ( .A1(n6610), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6594) );
  OAI21_X1 U8480 ( .B1(n6610), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6594), .ZN(
        n9494) );
  NOR2_X1 U8481 ( .A1(n9493), .A2(n9494), .ZN(n9492) );
  NAND2_X1 U8482 ( .A1(n6612), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U8483 ( .B1(n6612), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6595), .ZN(
        n9508) );
  NOR2_X1 U8484 ( .A1(n9507), .A2(n9508), .ZN(n9506) );
  AOI21_X1 U8485 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6612), .A(n9506), .ZN(
        n6596) );
  NAND2_X1 U8486 ( .A1(n6597), .A2(n6596), .ZN(n6784) );
  OAI21_X1 U8487 ( .B1(n6597), .B2(n6596), .A(n6784), .ZN(n6598) );
  NOR2_X1 U8488 ( .A1(n6138), .A2(n8994), .ZN(n8999) );
  NAND2_X1 U8489 ( .A1(n6615), .A2(n8999), .ZN(n9620) );
  NAND2_X1 U8490 ( .A1(n6598), .A2(n9595), .ZN(n6621) );
  INV_X1 U8491 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U8492 ( .A1(n6790), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n9764), .B2(
        n6617), .ZN(n6614) );
  XNOR2_X1 U8493 ( .A(n9003), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9009) );
  INV_X1 U8494 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9755) );
  MUX2_X1 U8495 ( .A(n9755), .B(P1_REG1_REG_1__SCAN_IN), .S(n6599), .Z(n8986)
         );
  AND2_X1 U8496 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8985) );
  NAND2_X1 U8497 ( .A1(n8986), .A2(n8985), .ZN(n8984) );
  NAND2_X1 U8498 ( .A1(n8987), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8499 ( .A1(n8984), .A2(n6600), .ZN(n9008) );
  NAND2_X1 U8500 ( .A1(n9009), .A2(n9008), .ZN(n9007) );
  INV_X1 U8501 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10096) );
  OR2_X1 U8502 ( .A1(n9003), .A2(n10096), .ZN(n6601) );
  NAND2_X1 U8503 ( .A1(n9007), .A2(n6601), .ZN(n9017) );
  XNOR2_X1 U8504 ( .A(n9019), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U8505 ( .A1(n9017), .A2(n9018), .ZN(n9016) );
  OR2_X1 U8506 ( .A1(n9019), .A2(n9758), .ZN(n6602) );
  NAND2_X1 U8507 ( .A1(n9016), .A2(n6602), .ZN(n9039) );
  INV_X1 U8508 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U8509 ( .A(n9760), .B(P1_REG1_REG_4__SCAN_IN), .S(n9030), .Z(n9040)
         );
  NAND2_X1 U8510 ( .A1(n9039), .A2(n9040), .ZN(n9038) );
  OR2_X1 U8511 ( .A1(n9030), .A2(n9760), .ZN(n6603) );
  NAND2_X1 U8512 ( .A1(n9038), .A2(n6603), .ZN(n9544) );
  OR2_X1 U8513 ( .A1(n9542), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U8514 ( .A1(n9542), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6605) );
  AND2_X1 U8515 ( .A1(n6604), .A2(n6605), .ZN(n9545) );
  NAND2_X1 U8516 ( .A1(n9544), .A2(n9545), .ZN(n9543) );
  AND2_X1 U8517 ( .A1(n9543), .A2(n6605), .ZN(n9558) );
  INV_X1 U8518 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6606) );
  MUX2_X1 U8519 ( .A(n6606), .B(P1_REG1_REG_6__SCAN_IN), .S(n6607), .Z(n9557)
         );
  NOR2_X1 U8520 ( .A1(n9558), .A2(n9557), .ZN(n9556) );
  AOI21_X1 U8521 ( .B1(n6607), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9556), .ZN(
        n9497) );
  OR2_X1 U8522 ( .A1(n6610), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U8523 ( .A1(n6610), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8524 ( .A1(n6609), .A2(n6608), .ZN(n9498) );
  NOR2_X1 U8525 ( .A1(n9497), .A2(n9498), .ZN(n9496) );
  AOI21_X1 U8526 ( .B1(n6610), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9496), .ZN(
        n9511) );
  NAND2_X1 U8527 ( .A1(n6612), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6611) );
  OAI21_X1 U8528 ( .B1(n6612), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6611), .ZN(
        n9512) );
  NOR2_X1 U8529 ( .A1(n9511), .A2(n9512), .ZN(n9510) );
  AOI21_X1 U8530 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6612), .A(n9510), .ZN(
        n6613) );
  NAND2_X1 U8531 ( .A1(n6614), .A2(n6613), .ZN(n6789) );
  OAI21_X1 U8532 ( .B1(n6614), .B2(n6613), .A(n6789), .ZN(n6619) );
  NAND2_X1 U8533 ( .A1(n6615), .A2(n6138), .ZN(n9629) );
  NAND2_X1 U8534 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U8535 ( .A1(n9076), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6616) );
  OAI211_X1 U8536 ( .C1(n9629), .C2(n6617), .A(n7201), .B(n6616), .ZN(n6618)
         );
  AOI21_X1 U8537 ( .B1(n6619), .B2(n9623), .A(n6618), .ZN(n6620) );
  NAND2_X1 U8538 ( .A1(n6621), .A2(n6620), .ZN(P1_U3252) );
  INV_X1 U8539 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6624) );
  OAI222_X1 U8540 ( .A1(n7528), .A2(n6624), .B1(n8825), .B2(n6623), .C1(
        P2_U3151), .C2(n6622), .ZN(P2_U3284) );
  INV_X1 U8541 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6625) );
  OAI222_X1 U8542 ( .A1(n8825), .A2(n6628), .B1(n6626), .B2(P2_U3151), .C1(
        n6625), .C2(n7528), .ZN(P2_U3283) );
  INV_X1 U8543 ( .A(n9060), .ZN(n6799) );
  INV_X1 U8544 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6627) );
  OAI222_X1 U8545 ( .A1(P1_U3086), .A2(n6799), .B1(n9478), .B2(n6628), .C1(
        n6627), .C2(n8222), .ZN(P1_U3343) );
  XOR2_X1 U8546 ( .A(n6630), .B(n6629), .Z(n6633) );
  NAND2_X1 U8547 ( .A1(n9535), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6653) );
  AOI22_X1 U8548 ( .A1(n9343), .A2(n8983), .B1(n8981), .B2(n9345), .ZN(n9663)
         );
  OAI22_X1 U8549 ( .A1(n9528), .A2(n5834), .B1(n9663), .B2(n8952), .ZN(n6631)
         );
  AOI21_X1 U8550 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6653), .A(n6631), .ZN(
        n6632) );
  OAI21_X1 U8551 ( .B1(n6633), .B2(n8945), .A(n6632), .ZN(P1_U3237) );
  NAND2_X1 U8552 ( .A1(n7143), .A2(P2_U3893), .ZN(n6634) );
  OAI21_X1 U8553 ( .B1(P2_U3893), .B2(n5857), .A(n6634), .ZN(P2_U3495) );
  XNOR2_X1 U8554 ( .A(n6636), .B(n6635), .ZN(n6652) );
  INV_X1 U8555 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U8556 ( .A1(n6637), .A2(n6921), .ZN(n6638) );
  NAND2_X1 U8557 ( .A1(n6639), .A2(n6638), .ZN(n6641) );
  NOR2_X1 U8558 ( .A1(n6900), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6640) );
  AOI21_X1 U8559 ( .B1(n9821), .B2(n6641), .A(n6640), .ZN(n6648) );
  INV_X1 U8560 ( .A(n9848), .ZN(n9777) );
  NAND2_X1 U8561 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  NAND2_X1 U8562 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  NAND2_X1 U8563 ( .A1(n9777), .A2(n6646), .ZN(n6647) );
  OAI211_X1 U8564 ( .C1(n9959), .C2(n9832), .A(n6648), .B(n6647), .ZN(n6649)
         );
  AOI21_X1 U8565 ( .B1(n6650), .B2(n9817), .A(n6649), .ZN(n6651) );
  OAI21_X1 U8566 ( .B1(n6652), .B2(n9826), .A(n6651), .ZN(P2_U3183) );
  INV_X1 U8567 ( .A(n6653), .ZN(n6666) );
  INV_X1 U8568 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6863) );
  XOR2_X1 U8569 ( .A(n6655), .B(n6654), .Z(n9002) );
  NOR2_X1 U8570 ( .A1(n8952), .A2(n9723), .ZN(n8940) );
  INV_X1 U8571 ( .A(n8940), .ZN(n8892) );
  OAI22_X1 U8572 ( .A1(n8892), .A2(n6656), .B1(n9528), .B2(n7052), .ZN(n6657)
         );
  AOI21_X1 U8573 ( .B1(n9531), .B2(n9002), .A(n6657), .ZN(n6658) );
  OAI21_X1 U8574 ( .B1(n6666), .B2(n6863), .A(n6658), .ZN(P1_U3232) );
  NAND2_X1 U8575 ( .A1(n9526), .A2(n9343), .ZN(n8938) );
  INV_X1 U8576 ( .A(n8938), .ZN(n8895) );
  INV_X1 U8577 ( .A(n7053), .ZN(n9691) );
  OAI22_X1 U8578 ( .A1(n8892), .A2(n6941), .B1(n9691), .B2(n9528), .ZN(n6659)
         );
  AOI21_X1 U8579 ( .B1(n8895), .B2(n7043), .A(n6659), .ZN(n6665) );
  OAI21_X1 U8580 ( .B1(n6662), .B2(n6661), .A(n6660), .ZN(n6663) );
  NAND2_X1 U8581 ( .A1(n6663), .A2(n9531), .ZN(n6664) );
  OAI211_X1 U8582 ( .C1(n6666), .C2(n5808), .A(n6665), .B(n6664), .ZN(P1_U3222) );
  NAND2_X1 U8583 ( .A1(n6667), .A2(n9843), .ZN(n6691) );
  AOI21_X1 U8584 ( .B1(n6692), .B2(n6669), .A(n6668), .ZN(n6690) );
  INV_X1 U8585 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6686) );
  INV_X1 U8586 ( .A(n6672), .ZN(n6674) );
  NAND3_X1 U8587 ( .A1(n6671), .A2(n6674), .A3(n6673), .ZN(n6675) );
  NAND2_X1 U8588 ( .A1(n6670), .A2(n6675), .ZN(n6677) );
  NOR2_X1 U8589 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6676), .ZN(n8206) );
  AOI21_X1 U8590 ( .B1(n9777), .B2(n6677), .A(n8206), .ZN(n6685) );
  INV_X1 U8591 ( .A(n6678), .ZN(n6680) );
  NAND3_X1 U8592 ( .A1(n6698), .A2(n6680), .A3(n6679), .ZN(n6681) );
  NAND2_X1 U8593 ( .A1(n6682), .A2(n6681), .ZN(n6683) );
  NAND2_X1 U8594 ( .A1(n9821), .A2(n6683), .ZN(n6684) );
  OAI211_X1 U8595 ( .C1(n6686), .C2(n9832), .A(n6685), .B(n6684), .ZN(n6687)
         );
  AOI21_X1 U8596 ( .B1(n6688), .B2(n9817), .A(n6687), .ZN(n6689) );
  OAI21_X1 U8597 ( .B1(n6691), .B2(n6690), .A(n6689), .ZN(P2_U3186) );
  OAI21_X1 U8598 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6709) );
  NOR2_X1 U8599 ( .A1(n9835), .A2(n6695), .ZN(n6708) );
  INV_X1 U8600 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U8601 ( .A1(n6696), .A2(n9939), .ZN(n6697) );
  NAND2_X1 U8602 ( .A1(n6698), .A2(n6697), .ZN(n6700) );
  NOR2_X1 U8603 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6699), .ZN(n8217) );
  AOI21_X1 U8604 ( .B1(n9821), .B2(n6700), .A(n8217), .ZN(n6706) );
  NAND2_X1 U8605 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U8606 ( .A1(n6671), .A2(n6703), .ZN(n6704) );
  NAND2_X1 U8607 ( .A1(n9777), .A2(n6704), .ZN(n6705) );
  OAI211_X1 U8608 ( .C1(n10027), .C2(n9832), .A(n6706), .B(n6705), .ZN(n6707)
         );
  AOI211_X1 U8609 ( .C1(n6709), .C2(n9843), .A(n6708), .B(n6707), .ZN(n6710)
         );
  INV_X1 U8610 ( .A(n6710), .ZN(P2_U3185) );
  INV_X1 U8611 ( .A(n6711), .ZN(n6720) );
  AOI22_X1 U8612 ( .A1(n9587), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9476), .ZN(n6712) );
  OAI21_X1 U8613 ( .B1(n6720), .B2(n9478), .A(n6712), .ZN(P1_U3342) );
  XOR2_X1 U8614 ( .A(n6714), .B(n6713), .Z(n6718) );
  MUX2_X1 U8615 ( .A(P1_U3086), .B(n8955), .S(n6944), .Z(n6716) );
  OAI22_X1 U8616 ( .A1(n8892), .A2(n6942), .B1(n9703), .B2(n9528), .ZN(n6715)
         );
  AOI211_X1 U8617 ( .C1(n8895), .C2(n8982), .A(n6716), .B(n6715), .ZN(n6717)
         );
  OAI21_X1 U8618 ( .B1(n6718), .B2(n8945), .A(n6717), .ZN(P1_U3218) );
  INV_X1 U8619 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6719) );
  OAI222_X1 U8620 ( .A1(n8825), .A2(n6720), .B1(n8394), .B2(P2_U3151), .C1(
        n6719), .C2(n7528), .ZN(P2_U3282) );
  XOR2_X1 U8621 ( .A(n6722), .B(n6721), .Z(n6740) );
  AND3_X1 U8622 ( .A1(n6725), .A2(n6724), .A3(n6723), .ZN(n6726) );
  NOR2_X1 U8623 ( .A1(n6727), .A2(n6726), .ZN(n6736) );
  INV_X1 U8624 ( .A(n6728), .ZN(n6733) );
  NAND3_X1 U8625 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n6732) );
  AOI21_X1 U8626 ( .B1(n6733), .B2(n6732), .A(n9852), .ZN(n6734) );
  AOI21_X1 U8627 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n9797), .A(n6734), .ZN(
        n6735) );
  NAND2_X1 U8628 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7245) );
  OAI211_X1 U8629 ( .C1(n6736), .C2(n9848), .A(n6735), .B(n7245), .ZN(n6737)
         );
  AOI21_X1 U8630 ( .B1(n6738), .B2(n9817), .A(n6737), .ZN(n6739) );
  OAI21_X1 U8631 ( .B1(n6740), .B2(n9826), .A(n6739), .ZN(P2_U3188) );
  INV_X1 U8632 ( .A(n6741), .ZN(n6746) );
  INV_X1 U8633 ( .A(n6742), .ZN(n6756) );
  INV_X1 U8634 ( .A(n6743), .ZN(n6744) );
  AOI21_X1 U8635 ( .B1(n6751), .B2(n6756), .A(n6744), .ZN(n6745) );
  OAI21_X1 U8636 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(n6748) );
  NAND2_X1 U8637 ( .A1(n6748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6753) );
  INV_X1 U8638 ( .A(n6749), .ZN(n6817) );
  NAND2_X1 U8639 ( .A1(n6761), .A2(n6817), .ZN(n8143) );
  INV_X1 U8640 ( .A(n8143), .ZN(n6750) );
  NAND2_X1 U8641 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  NAND2_X1 U8642 ( .A1(n6753), .A2(n6752), .ZN(n7091) );
  NOR2_X1 U8643 ( .A1(n7091), .A2(n6754), .ZN(n7621) );
  NAND2_X1 U8644 ( .A1(n7098), .A2(n8726), .ZN(n7968) );
  NAND2_X1 U8645 ( .A1(n6894), .A2(n7968), .ZN(n8723) );
  OR2_X1 U8646 ( .A1(n6759), .A2(n6755), .ZN(n6758) );
  NAND2_X1 U8647 ( .A1(n6764), .A2(n6756), .ZN(n6757) );
  OR2_X1 U8648 ( .A1(n6759), .A2(n9928), .ZN(n6762) );
  AND2_X1 U8649 ( .A1(n6764), .A2(n6817), .ZN(n7110) );
  INV_X1 U8650 ( .A(n7110), .ZN(n6765) );
  OR2_X2 U8651 ( .A1(n6765), .A2(n7109), .ZN(n8360) );
  OAI22_X1 U8652 ( .A1(n8365), .A2(n8726), .B1(n6763), .B2(n8360), .ZN(n6766)
         );
  AOI21_X1 U8653 ( .B1(n8723), .B2(n8354), .A(n6766), .ZN(n6767) );
  OAI21_X1 U8654 ( .B1(n7621), .B2(n6768), .A(n6767), .ZN(P2_U3172) );
  INV_X1 U8655 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6770) );
  INV_X1 U8656 ( .A(n6769), .ZN(n6771) );
  OAI222_X1 U8657 ( .A1(n7528), .A2(n6770), .B1(n8825), .B2(n6771), .C1(
        P2_U3151), .C2(n8408), .ZN(P2_U3281) );
  INV_X1 U8658 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6772) );
  OAI222_X1 U8659 ( .A1(n8222), .A2(n6772), .B1(n9478), .B2(n6771), .C1(n9602), 
        .C2(P1_U3086), .ZN(P1_U3341) );
  NAND2_X1 U8660 ( .A1(n6774), .A2(n6773), .ZN(n6776) );
  XNOR2_X1 U8661 ( .A(n6776), .B(n6775), .ZN(n6782) );
  OAI22_X1 U8662 ( .A1(n9528), .A2(n6915), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6777), .ZN(n6780) );
  OAI22_X1 U8663 ( .A1(n8892), .A2(n6778), .B1(n6942), .B2(n8938), .ZN(n6779)
         );
  AOI211_X1 U8664 ( .C1(n6951), .C2(n8955), .A(n6780), .B(n6779), .ZN(n6781)
         );
  OAI21_X1 U8665 ( .B1(n6782), .B2(n8945), .A(n6781), .ZN(P1_U3227) );
  NOR2_X1 U8666 ( .A1(n9060), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6783) );
  AOI21_X1 U8667 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9060), .A(n6783), .ZN(
        n6788) );
  OAI21_X1 U8668 ( .B1(n6790), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6784), .ZN(
        n9486) );
  INV_X1 U8669 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6785) );
  XNOR2_X1 U8670 ( .A(n6791), .B(n6785), .ZN(n9485) );
  NOR2_X1 U8671 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  NAND2_X1 U8672 ( .A1(n9575), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6786) );
  OAI21_X1 U8673 ( .B1(n9575), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6786), .ZN(
        n9568) );
  NOR2_X1 U8674 ( .A1(n9569), .A2(n9568), .ZN(n9567) );
  AOI21_X1 U8675 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9575), .A(n9567), .ZN(
        n6787) );
  NAND2_X1 U8676 ( .A1(n6788), .A2(n6787), .ZN(n9059) );
  OAI21_X1 U8677 ( .B1(n6788), .B2(n6787), .A(n9059), .ZN(n6801) );
  OAI21_X1 U8678 ( .B1(n6790), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6789), .ZN(
        n9482) );
  INV_X1 U8679 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6792) );
  MUX2_X1 U8680 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6792), .S(n6791), .Z(n9483)
         );
  NOR2_X1 U8681 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  AOI21_X1 U8682 ( .B1(n9489), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9481), .ZN(
        n9572) );
  INV_X1 U8683 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6793) );
  MUX2_X1 U8684 ( .A(n6793), .B(P1_REG1_REG_11__SCAN_IN), .S(n9575), .Z(n9571)
         );
  NOR2_X1 U8685 ( .A1(n9572), .A2(n9571), .ZN(n9570) );
  AOI21_X1 U8686 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9575), .A(n9570), .ZN(
        n6795) );
  INV_X1 U8687 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U8688 ( .A1(n9060), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9766), .B2(
        n6799), .ZN(n6794) );
  NAND2_X1 U8689 ( .A1(n6795), .A2(n6794), .ZN(n9046) );
  OAI21_X1 U8690 ( .B1(n6795), .B2(n6794), .A(n9046), .ZN(n6796) );
  NAND2_X1 U8691 ( .A1(n6796), .A2(n9623), .ZN(n6798) );
  AND2_X1 U8692 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7336) );
  AOI21_X1 U8693 ( .B1(n9076), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7336), .ZN(
        n6797) );
  OAI211_X1 U8694 ( .C1(n9629), .C2(n6799), .A(n6798), .B(n6797), .ZN(n6800)
         );
  AOI21_X1 U8695 ( .B1(n9595), .B2(n6801), .A(n6800), .ZN(n6802) );
  INV_X1 U8696 ( .A(n6802), .ZN(P1_U3255) );
  AOI22_X1 U8697 ( .A1(n8895), .A2(n8981), .B1(n8940), .B2(n8979), .ZN(n6803)
         );
  NAND2_X1 U8698 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U8699 ( .C1(n10139), .C2(n9528), .A(n6803), .B(n9031), .ZN(n6809)
         );
  INV_X1 U8700 ( .A(n6805), .ZN(n6806) );
  AOI211_X1 U8701 ( .C1(n6807), .C2(n6804), .A(n8945), .B(n6806), .ZN(n6808)
         );
  AOI211_X1 U8702 ( .C1(n10145), .C2(n8955), .A(n6809), .B(n6808), .ZN(n6810)
         );
  INV_X1 U8703 ( .A(n6810), .ZN(P1_U3230) );
  AOI21_X1 U8704 ( .B1(n6813), .B2(n6812), .A(n6811), .ZN(n6816) );
  INV_X1 U8705 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8706 ( .A1(n6816), .A2(n6815), .ZN(n6820) );
  NOR2_X1 U8707 ( .A1(n6763), .A2(n8646), .ZN(n8722) );
  INV_X1 U8708 ( .A(n8723), .ZN(n6818) );
  NOR3_X1 U8709 ( .A1(n6818), .A2(n6817), .A3(n9920), .ZN(n6819) );
  AOI211_X1 U8710 ( .C1(n9877), .C2(P2_REG3_REG_0__SCAN_IN), .A(n8722), .B(
        n6819), .ZN(n6821) );
  MUX2_X1 U8711 ( .A(n6822), .B(n6821), .S(n9878), .Z(n6823) );
  OAI21_X1 U8712 ( .B1(n8481), .B2(n8726), .A(n6823), .ZN(P2_U3233) );
  INV_X1 U8713 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6825) );
  INV_X1 U8714 ( .A(n6824), .ZN(n6827) );
  OAI222_X1 U8715 ( .A1(n7528), .A2(n6825), .B1(n8825), .B2(n6827), .C1(
        P2_U3151), .C2(n8425), .ZN(P2_U3280) );
  INV_X1 U8716 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6826) );
  OAI222_X1 U8717 ( .A1(n9064), .A2(P1_U3086), .B1(n9478), .B2(n6827), .C1(
        n6826), .C2(n8222), .ZN(P1_U3340) );
  XNOR2_X1 U8718 ( .A(n6828), .B(n6829), .ZN(n6836) );
  INV_X1 U8719 ( .A(n6853), .ZN(n6834) );
  NAND2_X1 U8720 ( .A1(n8979), .A2(n9343), .ZN(n6831) );
  NAND2_X1 U8721 ( .A1(n8977), .A2(n9345), .ZN(n6830) );
  NAND2_X1 U8722 ( .A1(n6831), .A2(n6830), .ZN(n6838) );
  AOI22_X1 U8723 ( .A1(n9526), .A2(n6838), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6833) );
  NAND2_X1 U8724 ( .A1(n8943), .A2(n6852), .ZN(n6832) );
  OAI211_X1 U8725 ( .C1(n9535), .C2(n6834), .A(n6833), .B(n6832), .ZN(n6835)
         );
  AOI21_X1 U8726 ( .B1(n6836), .B2(n9531), .A(n6835), .ZN(n6837) );
  INV_X1 U8727 ( .A(n6837), .ZN(P1_U3239) );
  XOR2_X1 U8728 ( .A(n7773), .B(n6961), .Z(n6840) );
  INV_X1 U8729 ( .A(n6838), .ZN(n6839) );
  OAI21_X1 U8730 ( .B1(n6840), .B2(n9719), .A(n6839), .ZN(n6928) );
  INV_X1 U8731 ( .A(n6928), .ZN(n6858) );
  INV_X1 U8732 ( .A(n6841), .ZN(n6843) );
  NAND3_X1 U8733 ( .A1(n6844), .A2(n6843), .A3(n6842), .ZN(n6845) );
  NAND2_X1 U8734 ( .A1(n9103), .A2(n6846), .ZN(n6847) );
  OR2_X1 U8735 ( .A1(n9677), .A2(n6847), .ZN(n6972) );
  OAI21_X1 U8736 ( .B1(n6850), .B2(n7773), .A(n6849), .ZN(n6930) );
  AOI211_X1 U8737 ( .C1(n6852), .C2(n6909), .A(n9740), .B(n7019), .ZN(n6929)
         );
  NAND2_X1 U8738 ( .A1(n6929), .A2(n10148), .ZN(n6855) );
  INV_X2 U8739 ( .A(n9326), .ZN(n10146) );
  AOI22_X1 U8740 ( .A1(n9677), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6853), .B2(
        n10146), .ZN(n6854) );
  OAI211_X1 U8741 ( .C1(n6934), .C2(n10140), .A(n6855), .B(n6854), .ZN(n6856)
         );
  AOI21_X1 U8742 ( .B1(n10150), .B2(n6930), .A(n6856), .ZN(n6857) );
  OAI21_X1 U8743 ( .B1(n6858), .B2(n9677), .A(n6857), .ZN(P1_U3287) );
  INV_X1 U8744 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U8745 ( .A1(n10148), .A2(n9711), .ZN(n9112) );
  INV_X1 U8746 ( .A(n9112), .ZN(n9350) );
  OAI21_X1 U8747 ( .B1(n9350), .B2(n9652), .A(n9686), .ZN(n6866) );
  INV_X1 U8748 ( .A(n7042), .ZN(n6859) );
  NAND2_X1 U8749 ( .A1(n7043), .A2(n7052), .ZN(n7837) );
  NAND2_X1 U8750 ( .A1(n6859), .A2(n7837), .ZN(n9681) );
  INV_X1 U8751 ( .A(n7906), .ZN(n6861) );
  NAND3_X1 U8752 ( .A1(n9681), .A2(n6861), .A3(n6860), .ZN(n6862) );
  NAND2_X1 U8753 ( .A1(n8983), .A2(n9345), .ZN(n9680) );
  OAI211_X1 U8754 ( .C1(n9326), .C2(n6863), .A(n6862), .B(n9680), .ZN(n6864)
         );
  NAND2_X1 U8755 ( .A1(n10141), .A2(n6864), .ZN(n6865) );
  OAI211_X1 U8756 ( .C1(n6867), .C2(n10141), .A(n6866), .B(n6865), .ZN(
        P1_U3293) );
  AOI21_X1 U8757 ( .B1(n6870), .B2(n6869), .A(n6868), .ZN(n6891) );
  INV_X1 U8758 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6873) );
  INV_X1 U8759 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6871) );
  NOR2_X1 U8760 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6871), .ZN(n7328) );
  INV_X1 U8761 ( .A(n7328), .ZN(n6872) );
  OAI21_X1 U8762 ( .B1(n9832), .B2(n6873), .A(n6872), .ZN(n6881) );
  INV_X1 U8763 ( .A(n6874), .ZN(n6876) );
  INV_X1 U8764 ( .A(n9792), .ZN(n6875) );
  NAND3_X1 U8765 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n6878) );
  AOI21_X1 U8766 ( .B1(n6879), .B2(n6878), .A(n9848), .ZN(n6880) );
  AOI211_X1 U8767 ( .C1(n9817), .C2(n6882), .A(n6881), .B(n6880), .ZN(n6890)
         );
  INV_X1 U8768 ( .A(n9802), .ZN(n6886) );
  INV_X1 U8769 ( .A(n6883), .ZN(n6884) );
  NOR3_X1 U8770 ( .A1(n6886), .A2(n6885), .A3(n6884), .ZN(n6887) );
  OAI21_X1 U8771 ( .B1(n6888), .B2(n6887), .A(n9821), .ZN(n6889) );
  OAI211_X1 U8772 ( .C1(n6891), .C2(n9826), .A(n6890), .B(n6889), .ZN(P2_U3190) );
  INV_X1 U8773 ( .A(n6892), .ZN(n6927) );
  OAI222_X1 U8774 ( .A1(n8825), .A2(n6927), .B1(n8443), .B2(P2_U3151), .C1(
        n6893), .C2(n7528), .ZN(P2_U3279) );
  INV_X1 U8775 ( .A(n6897), .ZN(n7935) );
  XNOR2_X1 U8776 ( .A(n7935), .B(n6894), .ZN(n6920) );
  AND2_X1 U8777 ( .A1(n9873), .A2(n7965), .ZN(n7226) );
  OR2_X1 U8778 ( .A1(n7401), .A2(n7226), .ZN(n6895) );
  OAI21_X1 U8779 ( .B1(n6898), .B2(n6897), .A(n6896), .ZN(n6899) );
  AOI222_X1 U8780 ( .A1(n9866), .A2(n6899), .B1(n8380), .B2(n9860), .C1(n7098), 
        .C2(n9862), .ZN(n6919) );
  OAI21_X1 U8781 ( .B1(n6900), .B2(n8607), .A(n6919), .ZN(n6901) );
  NAND2_X1 U8782 ( .A1(n6901), .A2(n9878), .ZN(n6904) );
  AOI22_X1 U8783 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n9881), .B1(n8658), .B2(
        n6902), .ZN(n6903) );
  OAI211_X1 U8784 ( .C1(n6920), .C2(n8661), .A(n6904), .B(n6903), .ZN(P2_U3232) );
  XNOR2_X1 U8785 ( .A(n6905), .B(n7774), .ZN(n6950) );
  XNOR2_X1 U8786 ( .A(n6907), .B(n6906), .ZN(n6908) );
  AOI222_X1 U8787 ( .A1(n9665), .A2(n6908), .B1(n8980), .B2(n9343), .C1(n8978), 
        .C2(n9345), .ZN(n6959) );
  AOI21_X1 U8788 ( .B1(n9710), .B2(n6952), .A(n9740), .ZN(n6910) );
  NAND2_X1 U8789 ( .A1(n6910), .A2(n6909), .ZN(n6955) );
  OAI211_X1 U8790 ( .C1(n9683), .C2(n6950), .A(n6959), .B(n6955), .ZN(n6917)
         );
  INV_X1 U8791 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6911) );
  OAI22_X1 U8792 ( .A1(n9469), .A2(n6915), .B1(n9753), .B2(n6911), .ZN(n6912)
         );
  AOI21_X1 U8793 ( .B1(n6917), .B2(n9753), .A(n6912), .ZN(n6913) );
  INV_X1 U8794 ( .A(n6913), .ZN(P1_U3468) );
  INV_X1 U8795 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6914) );
  OAI22_X1 U8796 ( .A1(n9414), .A2(n6915), .B1(n9770), .B2(n6914), .ZN(n6916)
         );
  AOI21_X1 U8797 ( .B1(n6917), .B2(n9770), .A(n6916), .ZN(n6918) );
  INV_X1 U8798 ( .A(n6918), .ZN(P1_U3527) );
  OAI21_X1 U8799 ( .B1(n9911), .B2(n6920), .A(n6919), .ZN(n6925) );
  OAI22_X1 U8800 ( .A1(n8670), .A2(n7099), .B1(n9954), .B2(n6921), .ZN(n6922)
         );
  AOI21_X1 U8801 ( .B1(n6925), .B2(n9954), .A(n6922), .ZN(n6923) );
  INV_X1 U8802 ( .A(n6923), .ZN(P2_U3460) );
  OAI22_X1 U8803 ( .A1(n7099), .A2(n8740), .B1(n9934), .B2(n5097), .ZN(n6924)
         );
  AOI21_X1 U8804 ( .B1(n6925), .B2(n9934), .A(n6924), .ZN(n6926) );
  INV_X1 U8805 ( .A(n6926), .ZN(P2_U3393) );
  INV_X1 U8806 ( .A(n9075), .ZN(n9057) );
  OAI222_X1 U8807 ( .A1(P1_U3086), .A2(n9057), .B1(n9478), .B2(n6927), .C1(
        n10111), .C2(n8222), .ZN(P1_U3339) );
  AOI211_X1 U8808 ( .C1(n9750), .C2(n6930), .A(n6929), .B(n6928), .ZN(n6937)
         );
  OAI22_X1 U8809 ( .A1(n9414), .A2(n6934), .B1(n9770), .B2(n6606), .ZN(n6931)
         );
  INV_X1 U8810 ( .A(n6931), .ZN(n6932) );
  OAI21_X1 U8811 ( .B1(n6937), .B2(n9768), .A(n6932), .ZN(P1_U3528) );
  INV_X1 U8812 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6933) );
  OAI22_X1 U8813 ( .A1(n9469), .A2(n6934), .B1(n9753), .B2(n6933), .ZN(n6935)
         );
  INV_X1 U8814 ( .A(n6935), .ZN(n6936) );
  OAI21_X1 U8815 ( .B1(n6937), .B2(n9752), .A(n6936), .ZN(P1_U3471) );
  INV_X1 U8816 ( .A(n10150), .ZN(n9352) );
  XNOR2_X1 U8817 ( .A(n6938), .B(n7775), .ZN(n9706) );
  INV_X1 U8818 ( .A(n9706), .ZN(n6949) );
  INV_X1 U8819 ( .A(n9715), .ZN(n6939) );
  AOI21_X1 U8820 ( .B1(n7775), .B2(n7646), .A(n6939), .ZN(n6940) );
  OAI222_X1 U8821 ( .A1(n9723), .A2(n6942), .B1(n9721), .B2(n6941), .C1(n9719), 
        .C2(n6940), .ZN(n9704) );
  OAI211_X1 U8822 ( .C1(n9672), .C2(n9703), .A(n9711), .B(n9709), .ZN(n9702)
         );
  NAND2_X1 U8823 ( .A1(n9652), .A2(n6943), .ZN(n6946) );
  AOI22_X1 U8824 ( .A1(n9677), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10146), .B2(
        n6944), .ZN(n6945) );
  OAI211_X1 U8825 ( .C1(n9702), .C2(n9655), .A(n6946), .B(n6945), .ZN(n6947)
         );
  AOI21_X1 U8826 ( .B1(n9704), .B2(n10141), .A(n6947), .ZN(n6948) );
  OAI21_X1 U8827 ( .B1(n9352), .B2(n6949), .A(n6948), .ZN(P1_U3290) );
  INV_X1 U8828 ( .A(n6950), .ZN(n6957) );
  AOI22_X1 U8829 ( .A1(n9677), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6951), .B2(
        n10146), .ZN(n6954) );
  NAND2_X1 U8830 ( .A1(n9652), .A2(n6952), .ZN(n6953) );
  OAI211_X1 U8831 ( .C1(n6955), .C2(n9655), .A(n6954), .B(n6953), .ZN(n6956)
         );
  AOI21_X1 U8832 ( .B1(n6957), .B2(n10150), .A(n6956), .ZN(n6958) );
  OAI21_X1 U8833 ( .B1(n6959), .B2(n9677), .A(n6958), .ZN(P1_U3288) );
  INV_X1 U8834 ( .A(n7648), .ZN(n6960) );
  OR2_X1 U8835 ( .A1(n6961), .A2(n6960), .ZN(n6962) );
  NAND2_X1 U8836 ( .A1(n6962), .A2(n7654), .ZN(n7012) );
  NAND2_X1 U8837 ( .A1(n7012), .A2(n7658), .ZN(n6964) );
  NAND2_X1 U8838 ( .A1(n6964), .A2(n6963), .ZN(n6982) );
  XNOR2_X1 U8839 ( .A(n6982), .B(n6966), .ZN(n6971) );
  OAI21_X1 U8840 ( .B1(n6967), .B2(n6966), .A(n6965), .ZN(n9730) );
  INV_X1 U8841 ( .A(n9638), .ZN(n7048) );
  OAI22_X1 U8842 ( .A1(n6968), .A2(n9723), .B1(n7176), .B2(n9721), .ZN(n6969)
         );
  AOI21_X1 U8843 ( .B1(n9730), .B2(n7048), .A(n6969), .ZN(n6970) );
  OAI21_X1 U8844 ( .B1(n9719), .B2(n6971), .A(n6970), .ZN(n9728) );
  INV_X1 U8845 ( .A(n9728), .ZN(n6979) );
  INV_X1 U8846 ( .A(n6972), .ZN(n9658) );
  INV_X1 U8847 ( .A(n7125), .ZN(n6973) );
  OAI211_X1 U8848 ( .C1(n9727), .C2(n7017), .A(n6973), .B(n9711), .ZN(n9726)
         );
  AOI22_X1 U8849 ( .A1(n9677), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6974), .B2(
        n10146), .ZN(n6976) );
  NAND2_X1 U8850 ( .A1(n9652), .A2(n7178), .ZN(n6975) );
  OAI211_X1 U8851 ( .C1(n9726), .C2(n9655), .A(n6976), .B(n6975), .ZN(n6977)
         );
  AOI21_X1 U8852 ( .B1(n9730), .B2(n9658), .A(n6977), .ZN(n6978) );
  OAI21_X1 U8853 ( .B1(n6979), .B2(n9677), .A(n6978), .ZN(P1_U3285) );
  INV_X1 U8854 ( .A(n7661), .ZN(n6981) );
  OAI21_X1 U8855 ( .B1(n6982), .B2(n6981), .A(n6980), .ZN(n6983) );
  XNOR2_X1 U8856 ( .A(n6983), .B(n6986), .ZN(n6985) );
  AND2_X1 U8857 ( .A1(n8976), .A2(n9343), .ZN(n6984) );
  AOI21_X1 U8858 ( .B1(n6985), .B2(n9665), .A(n6984), .ZN(n9737) );
  OR2_X1 U8859 ( .A1(n6987), .A2(n6986), .ZN(n6988) );
  NAND2_X1 U8860 ( .A1(n6989), .A2(n6988), .ZN(n9735) );
  XNOR2_X1 U8861 ( .A(n7125), .B(n6992), .ZN(n6991) );
  AND2_X1 U8862 ( .A1(n8974), .A2(n9345), .ZN(n6990) );
  AOI21_X1 U8863 ( .B1(n6991), .B2(n9711), .A(n6990), .ZN(n9732) );
  AOI22_X1 U8864 ( .A1(n9677), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7206), .B2(
        n10146), .ZN(n6994) );
  NAND2_X1 U8865 ( .A1(n6992), .A2(n9652), .ZN(n6993) );
  OAI211_X1 U8866 ( .C1(n9732), .C2(n9655), .A(n6994), .B(n6993), .ZN(n6995)
         );
  AOI21_X1 U8867 ( .B1(n9735), .B2(n10150), .A(n6995), .ZN(n6996) );
  OAI21_X1 U8868 ( .B1(n9737), .B2(n9677), .A(n6996), .ZN(P1_U3284) );
  NAND3_X1 U8869 ( .A1(n9863), .A2(n7936), .A3(n6998), .ZN(n6999) );
  NAND2_X1 U8870 ( .A1(n6997), .A2(n6999), .ZN(n7000) );
  NAND2_X1 U8871 ( .A1(n7000), .A2(n9866), .ZN(n7002) );
  AOI22_X1 U8872 ( .A1(n9860), .A2(n7143), .B1(n8380), .B2(n9862), .ZN(n7001)
         );
  AND2_X1 U8873 ( .A1(n7002), .A2(n7001), .ZN(n9889) );
  OAI22_X1 U8874 ( .A1(n8481), .A2(n8215), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8607), .ZN(n7003) );
  AOI21_X1 U8875 ( .B1(n9881), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7003), .ZN(
        n7006) );
  XNOR2_X1 U8876 ( .A(n7004), .B(n7936), .ZN(n9885) );
  NAND2_X1 U8877 ( .A1(n9885), .A2(n8613), .ZN(n7005) );
  OAI211_X1 U8878 ( .C1(n9889), .C2(n9881), .A(n7006), .B(n7005), .ZN(P2_U3230) );
  INV_X1 U8879 ( .A(n7007), .ZN(n7008) );
  OAI222_X1 U8880 ( .A1(n7528), .A2(n10035), .B1(n8825), .B2(n7008), .C1(
        P2_U3151), .C2(n9834), .ZN(P2_U3278) );
  INV_X1 U8881 ( .A(n9085), .ZN(n9091) );
  OAI222_X1 U8882 ( .A1(n8222), .A2(n7009), .B1(n9478), .B2(n7008), .C1(n9091), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  OAI21_X1 U8883 ( .B1(n7011), .B2(n4477), .A(n7010), .ZN(n9659) );
  INV_X1 U8884 ( .A(n9659), .ZN(n7020) );
  XNOR2_X1 U8885 ( .A(n7012), .B(n7658), .ZN(n7016) );
  NAND2_X1 U8886 ( .A1(n8978), .A2(n9343), .ZN(n7014) );
  NAND2_X1 U8887 ( .A1(n8976), .A2(n9345), .ZN(n7013) );
  AND2_X1 U8888 ( .A1(n7014), .A2(n7013), .ZN(n7030) );
  OAI21_X1 U8889 ( .B1(n7020), .B2(n9638), .A(n7030), .ZN(n7015) );
  AOI21_X1 U8890 ( .B1(n7016), .B2(n9665), .A(n7015), .ZN(n9661) );
  INV_X1 U8891 ( .A(n7017), .ZN(n7018) );
  OAI211_X1 U8892 ( .C1(n7025), .C2(n7019), .A(n7018), .B(n9711), .ZN(n9656)
         );
  OAI211_X1 U8893 ( .C1(n7020), .C2(n9689), .A(n9661), .B(n9656), .ZN(n7027)
         );
  INV_X1 U8894 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7021) );
  OAI22_X1 U8895 ( .A1(n9414), .A2(n7025), .B1(n9770), .B2(n7021), .ZN(n7022)
         );
  AOI21_X1 U8896 ( .B1(n7027), .B2(n9770), .A(n7022), .ZN(n7023) );
  INV_X1 U8897 ( .A(n7023), .ZN(P1_U3529) );
  INV_X1 U8898 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7024) );
  OAI22_X1 U8899 ( .A1(n9469), .A2(n7025), .B1(n9753), .B2(n7024), .ZN(n7026)
         );
  AOI21_X1 U8900 ( .B1(n7027), .B2(n9753), .A(n7026), .ZN(n7028) );
  INV_X1 U8901 ( .A(n7028), .ZN(P1_U3474) );
  NAND2_X1 U8902 ( .A1(n8943), .A2(n9651), .ZN(n7029) );
  NAND2_X1 U8903 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9504) );
  OAI211_X1 U8904 ( .C1(n7030), .C2(n8952), .A(n7029), .B(n9504), .ZN(n7038)
         );
  XNOR2_X1 U8905 ( .A(n7033), .B(n7032), .ZN(n7034) );
  XNOR2_X1 U8906 ( .A(n7035), .B(n7034), .ZN(n7036) );
  NOR2_X1 U8907 ( .A1(n7036), .A2(n8945), .ZN(n7037) );
  AOI211_X1 U8908 ( .C1(n9650), .C2(n8955), .A(n7038), .B(n7037), .ZN(n7039)
         );
  INV_X1 U8909 ( .A(n7039), .ZN(P1_U3213) );
  NAND2_X1 U8910 ( .A1(n7043), .A2(n9343), .ZN(n7045) );
  NAND2_X1 U8911 ( .A1(n8982), .A2(n9345), .ZN(n7044) );
  NAND2_X1 U8912 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  AOI21_X1 U8913 ( .B1(n7047), .B2(n9665), .A(n7046), .ZN(n7050) );
  NAND2_X1 U8914 ( .A1(n9694), .A2(n7048), .ZN(n7049) );
  NAND2_X1 U8915 ( .A1(n7050), .A2(n7049), .ZN(n9692) );
  MUX2_X1 U8916 ( .A(n9692), .B(P1_REG2_REG_1__SCAN_IN), .S(n9677), .Z(n7056)
         );
  INV_X1 U8917 ( .A(n9671), .ZN(n7051) );
  OAI211_X1 U8918 ( .C1(n9691), .C2(n7052), .A(n7051), .B(n9711), .ZN(n9690)
         );
  AOI22_X1 U8919 ( .A1(n9652), .A2(n7053), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n10146), .ZN(n7054) );
  OAI21_X1 U8920 ( .B1(n9655), .B2(n9690), .A(n7054), .ZN(n7055) );
  AOI211_X1 U8921 ( .C1(n9694), .C2(n9658), .A(n7056), .B(n7055), .ZN(n7057)
         );
  INV_X1 U8922 ( .A(n7057), .ZN(P1_U3292) );
  INV_X1 U8923 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9961) );
  NOR2_X1 U8924 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7058) );
  AOI21_X1 U8925 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7058), .ZN(n9966) );
  NOR2_X1 U8926 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7059) );
  AOI21_X1 U8927 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7059), .ZN(n9969) );
  NOR2_X1 U8928 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7060) );
  AOI21_X1 U8929 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7060), .ZN(n9972) );
  NOR2_X1 U8930 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7061) );
  AOI21_X1 U8931 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7061), .ZN(n9975) );
  NOR2_X1 U8932 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7062) );
  AOI21_X1 U8933 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7062), .ZN(n9978) );
  NOR2_X1 U8934 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7063) );
  AOI21_X1 U8935 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7063), .ZN(n9981) );
  NOR2_X1 U8936 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7064) );
  AOI21_X1 U8937 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7064), .ZN(n9984) );
  NOR2_X1 U8938 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7065) );
  AOI21_X1 U8939 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7065), .ZN(n9987) );
  NOR2_X1 U8940 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7066) );
  AOI21_X1 U8941 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7066), .ZN(n10166) );
  NOR2_X1 U8942 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7067) );
  AOI21_X1 U8943 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7067), .ZN(n10172) );
  NOR2_X1 U8944 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7068) );
  AOI21_X1 U8945 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7068), .ZN(n10169) );
  NOR2_X1 U8946 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7069) );
  AOI21_X1 U8947 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7069), .ZN(n10160) );
  NOR2_X1 U8948 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7070) );
  AOI21_X1 U8949 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7070), .ZN(n10163) );
  AND2_X1 U8950 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7071) );
  NOR2_X1 U8951 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7071), .ZN(n9956) );
  INV_X1 U8952 ( .A(n9956), .ZN(n9957) );
  NAND3_X1 U8953 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U8954 ( .A1(n9959), .A2(n9958), .ZN(n9955) );
  NAND2_X1 U8955 ( .A1(n9957), .A2(n9955), .ZN(n10175) );
  NAND2_X1 U8956 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7072) );
  OAI21_X1 U8957 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7072), .ZN(n10174) );
  NOR2_X1 U8958 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  AOI21_X1 U8959 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10173), .ZN(n10178) );
  NAND2_X1 U8960 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7073) );
  OAI21_X1 U8961 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7073), .ZN(n10177) );
  NOR2_X1 U8962 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  AOI21_X1 U8963 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10176), .ZN(n10181) );
  NOR2_X1 U8964 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7074) );
  AOI21_X1 U8965 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7074), .ZN(n10180) );
  NAND2_X1 U8966 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  OAI21_X1 U8967 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10179), .ZN(n10162) );
  NAND2_X1 U8968 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  OAI21_X1 U8969 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10161), .ZN(n10159) );
  NAND2_X1 U8970 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  OAI21_X1 U8971 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10158), .ZN(n10168) );
  NAND2_X1 U8972 ( .A1(n10169), .A2(n10168), .ZN(n10167) );
  OAI21_X1 U8973 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10167), .ZN(n10171) );
  NAND2_X1 U8974 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  OAI21_X1 U8975 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10170), .ZN(n10165) );
  NAND2_X1 U8976 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  OAI21_X1 U8977 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10164), .ZN(n9986) );
  NAND2_X1 U8978 ( .A1(n9987), .A2(n9986), .ZN(n9985) );
  OAI21_X1 U8979 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9985), .ZN(n9983) );
  NAND2_X1 U8980 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  OAI21_X1 U8981 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9982), .ZN(n9980) );
  NAND2_X1 U8982 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  OAI21_X1 U8983 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9979), .ZN(n9977) );
  NAND2_X1 U8984 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  OAI21_X1 U8985 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9976), .ZN(n9974) );
  NAND2_X1 U8986 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  OAI21_X1 U8987 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9973), .ZN(n9971) );
  NAND2_X1 U8988 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  OAI21_X1 U8989 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9970), .ZN(n9968) );
  NAND2_X1 U8990 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  OAI21_X1 U8991 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9967), .ZN(n9965) );
  NAND2_X1 U8992 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  OAI21_X1 U8993 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9964), .ZN(n9962) );
  NOR2_X1 U8994 ( .A1(n9961), .A2(n9962), .ZN(n7075) );
  NAND2_X1 U8995 ( .A1(n9961), .A2(n9962), .ZN(n9960) );
  OAI21_X1 U8996 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7075), .A(n9960), .ZN(
        n7079) );
  NOR2_X1 U8997 ( .A1(n7076), .A2(n7077), .ZN(n7078) );
  XNOR2_X1 U8998 ( .A(n7079), .B(n7078), .ZN(ADD_1068_U4) );
  OAI21_X1 U8999 ( .B1(n7081), .B2(n7981), .A(n7080), .ZN(n9892) );
  INV_X1 U9000 ( .A(n9892), .ZN(n7089) );
  NAND3_X1 U9001 ( .A1(n6997), .A2(n7981), .A3(n7082), .ZN(n7083) );
  NAND2_X1 U9002 ( .A1(n7084), .A2(n7083), .ZN(n7085) );
  AOI222_X1 U9003 ( .A1(n9866), .A2(n7085), .B1(n9861), .B2(n9862), .C1(n8379), 
        .C2(n9860), .ZN(n9894) );
  MUX2_X1 U9004 ( .A(n4965), .B(n9894), .S(n9878), .Z(n7088) );
  INV_X1 U9005 ( .A(n7086), .ZN(n8207) );
  AOI22_X1 U9006 ( .A1(n8658), .A2(n9891), .B1(n9877), .B2(n8207), .ZN(n7087)
         );
  OAI211_X1 U9007 ( .C1(n7089), .C2(n8661), .A(n7088), .B(n7087), .ZN(P2_U3229) );
  OR2_X1 U9008 ( .A1(n7090), .A2(P2_U3151), .ZN(n8147) );
  INV_X1 U9009 ( .A(n8147), .ZN(n7479) );
  INV_X1 U9010 ( .A(n7143), .ZN(n8214) );
  XNOR2_X1 U9011 ( .A(n7965), .B(n7283), .ZN(n7092) );
  AND2_X1 U9012 ( .A1(n7093), .A2(n7092), .ZN(n7094) );
  NAND2_X1 U9013 ( .A1(n7095), .A2(n7094), .ZN(n7097) );
  XNOR2_X1 U9014 ( .A(n8204), .B(n4291), .ZN(n7106) );
  INV_X1 U9015 ( .A(n7106), .ZN(n7107) );
  INV_X1 U9016 ( .A(n9861), .ZN(n7619) );
  XNOR2_X1 U9017 ( .A(n9886), .B(n7100), .ZN(n7105) );
  MUX2_X1 U9018 ( .A(n7098), .B(n7100), .S(n8726), .Z(n7611) );
  XNOR2_X1 U9019 ( .A(n9871), .B(n8184), .ZN(n7103) );
  XNOR2_X1 U9020 ( .A(n7103), .B(n8380), .ZN(n7617) );
  INV_X1 U9021 ( .A(n8380), .ZN(n7104) );
  AOI22_X1 U9022 ( .A1(n7618), .A2(n7617), .B1(n7104), .B2(n7103), .ZN(n8213)
         );
  XNOR2_X1 U9023 ( .A(n7105), .B(n9861), .ZN(n8212) );
  NAND2_X1 U9024 ( .A1(n8213), .A2(n8212), .ZN(n8211) );
  OAI21_X1 U9025 ( .B1(n7619), .B2(n7105), .A(n8211), .ZN(n8202) );
  XNOR2_X1 U9026 ( .A(n7106), .B(n7143), .ZN(n8203) );
  AOI21_X1 U9027 ( .B1(n8214), .B2(n7107), .A(n8201), .ZN(n7241) );
  XNOR2_X1 U9028 ( .A(n9895), .B(n4291), .ZN(n7239) );
  XNOR2_X1 U9029 ( .A(n7239), .B(n8379), .ZN(n7240) );
  XNOR2_X1 U9030 ( .A(n7241), .B(n7240), .ZN(n7108) );
  NAND2_X1 U9031 ( .A1(n7108), .A2(n8354), .ZN(n7116) );
  INV_X1 U9032 ( .A(n7111), .ZN(n7114) );
  INV_X1 U9033 ( .A(n8378), .ZN(n7112) );
  OAI22_X1 U9034 ( .A1(n8365), .A2(n9895), .B1(n7112), .B2(n8360), .ZN(n7113)
         );
  AOI211_X1 U9035 ( .C1(n8358), .C2(n7143), .A(n7114), .B(n7113), .ZN(n7115)
         );
  OAI211_X1 U9036 ( .C1(n7148), .C2(n8339), .A(n7116), .B(n7115), .ZN(P2_U3167) );
  OAI21_X1 U9037 ( .B1(n7118), .B2(n4691), .A(n7117), .ZN(n7154) );
  INV_X1 U9038 ( .A(n7154), .ZN(n7133) );
  INV_X1 U9039 ( .A(n7182), .ZN(n7119) );
  AOI21_X1 U9040 ( .B1(n4691), .B2(n7120), .A(n7119), .ZN(n7124) );
  NAND2_X1 U9041 ( .A1(n8975), .A2(n9343), .ZN(n7122) );
  NAND2_X1 U9042 ( .A1(n8973), .A2(n9345), .ZN(n7121) );
  NAND2_X1 U9043 ( .A1(n7122), .A2(n7121), .ZN(n9525) );
  INV_X1 U9044 ( .A(n9525), .ZN(n7123) );
  OAI21_X1 U9045 ( .B1(n7124), .B2(n9719), .A(n7123), .ZN(n7152) );
  INV_X1 U9046 ( .A(n7188), .ZN(n7127) );
  AOI21_X1 U9047 ( .B1(n7125), .B2(n9733), .A(n9529), .ZN(n7126) );
  NOR3_X1 U9048 ( .A1(n7127), .A2(n7126), .A3(n9740), .ZN(n7153) );
  NAND2_X1 U9049 ( .A1(n7153), .A2(n10148), .ZN(n7130) );
  AOI22_X1 U9050 ( .A1(n9677), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7128), .B2(
        n10146), .ZN(n7129) );
  OAI211_X1 U9051 ( .C1(n9529), .C2(n10140), .A(n7130), .B(n7129), .ZN(n7131)
         );
  AOI21_X1 U9052 ( .B1(n7152), .B2(n10141), .A(n7131), .ZN(n7132) );
  OAI21_X1 U9053 ( .B1(n7133), .B2(n9352), .A(n7132), .ZN(P1_U3283) );
  INV_X1 U9054 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U9055 ( .A1(n5678), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7136) );
  INV_X1 U9056 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8477) );
  OR2_X1 U9057 ( .A1(n7134), .A2(n8477), .ZN(n7135) );
  OAI211_X1 U9058 ( .C1(n8664), .C2(n7137), .A(n7136), .B(n7135), .ZN(n7138)
         );
  INV_X1 U9059 ( .A(n7138), .ZN(n7139) );
  NAND2_X1 U9060 ( .A1(n8381), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U9061 ( .B1(n8474), .B2(n8381), .A(n7141), .ZN(P2_U3522) );
  XNOR2_X1 U9062 ( .A(n8379), .B(n9895), .ZN(n7940) );
  XNOR2_X1 U9063 ( .A(n7142), .B(n7940), .ZN(n9896) );
  NAND2_X1 U9064 ( .A1(n9878), .A2(n7226), .ZN(n8487) );
  INV_X1 U9065 ( .A(n7401), .ZN(n9870) );
  AOI22_X1 U9066 ( .A1(n9862), .A2(n7143), .B1(n8378), .B2(n9860), .ZN(n7147)
         );
  XNOR2_X1 U9067 ( .A(n7144), .B(n7940), .ZN(n7145) );
  NAND2_X1 U9068 ( .A1(n7145), .A2(n9866), .ZN(n7146) );
  OAI211_X1 U9069 ( .C1(n9896), .C2(n9870), .A(n7147), .B(n7146), .ZN(n9898)
         );
  NAND2_X1 U9070 ( .A1(n9898), .A2(n9878), .ZN(n7151) );
  OAI22_X1 U9071 ( .A1(n8481), .A2(n9895), .B1(n7148), .B2(n8607), .ZN(n7149)
         );
  AOI21_X1 U9072 ( .B1(n9881), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7149), .ZN(
        n7150) );
  OAI211_X1 U9073 ( .C1(n9896), .C2(n8487), .A(n7151), .B(n7150), .ZN(P2_U3228) );
  AOI211_X1 U9074 ( .C1(n9750), .C2(n7154), .A(n7153), .B(n7152), .ZN(n7160)
         );
  INV_X1 U9075 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7155) );
  OAI22_X1 U9076 ( .A1(n9529), .A2(n9469), .B1(n9753), .B2(n7155), .ZN(n7156)
         );
  INV_X1 U9077 ( .A(n7156), .ZN(n7157) );
  OAI21_X1 U9078 ( .B1(n7160), .B2(n9752), .A(n7157), .ZN(P1_U3483) );
  INV_X1 U9079 ( .A(n9414), .ZN(n9429) );
  AOI22_X1 U9080 ( .A1(n7158), .A2(n9429), .B1(n9768), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7159) );
  OAI21_X1 U9081 ( .B1(n7160), .B2(n9768), .A(n7159), .ZN(P1_U3532) );
  INV_X1 U9082 ( .A(n7161), .ZN(n7164) );
  OAI222_X1 U9083 ( .A1(n8825), .A2(n7164), .B1(n7163), .B2(P2_U3151), .C1(
        n7162), .C2(n7528), .ZN(P2_U3277) );
  INV_X1 U9084 ( .A(n9094), .ZN(n9628) );
  OAI222_X1 U9085 ( .A1(n8222), .A2(n7165), .B1(n9478), .B2(n7164), .C1(
        P1_U3086), .C2(n9628), .ZN(P1_U3337) );
  INV_X1 U9086 ( .A(n7167), .ZN(n7169) );
  INV_X1 U9087 ( .A(n7166), .ZN(n7168) );
  OR2_X1 U9088 ( .A1(n7166), .A2(n7167), .ZN(n7194) );
  OAI21_X1 U9089 ( .B1(n7169), .B2(n7168), .A(n7194), .ZN(n7170) );
  NOR2_X1 U9090 ( .A1(n7170), .A2(n7171), .ZN(n7196) );
  AOI21_X1 U9091 ( .B1(n7171), .B2(n7170), .A(n7196), .ZN(n7180) );
  NAND2_X1 U9092 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9518) );
  INV_X1 U9093 ( .A(n9518), .ZN(n7172) );
  AOI21_X1 U9094 ( .B1(n8940), .B2(n8975), .A(n7172), .ZN(n7175) );
  OR2_X1 U9095 ( .A1(n9535), .A2(n7173), .ZN(n7174) );
  OAI211_X1 U9096 ( .C1(n7176), .C2(n8938), .A(n7175), .B(n7174), .ZN(n7177)
         );
  AOI21_X1 U9097 ( .B1(n7178), .B2(n8943), .A(n7177), .ZN(n7179) );
  OAI21_X1 U9098 ( .B1(n7180), .B2(n8945), .A(n7179), .ZN(P1_U3221) );
  XNOR2_X1 U9099 ( .A(n7233), .B(n7338), .ZN(n7183) );
  XNOR2_X1 U9100 ( .A(n7181), .B(n7183), .ZN(n7232) );
  INV_X1 U9101 ( .A(n7232), .ZN(n7193) );
  NAND2_X1 U9102 ( .A1(n7182), .A2(n7665), .ZN(n7184) );
  XNOR2_X1 U9103 ( .A(n7184), .B(n7183), .ZN(n7185) );
  OAI222_X1 U9104 ( .A1(n9723), .A2(n7186), .B1(n9721), .B2(n7289), .C1(n9719), 
        .C2(n7185), .ZN(n7230) );
  INV_X1 U9105 ( .A(n7187), .ZN(n7274) );
  AOI211_X1 U9106 ( .C1(n7233), .C2(n7188), .A(n9740), .B(n7274), .ZN(n7231)
         );
  NAND2_X1 U9107 ( .A1(n7231), .A2(n10148), .ZN(n7190) );
  AOI22_X1 U9108 ( .A1(n9677), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7291), .B2(
        n10146), .ZN(n7189) );
  OAI211_X1 U9109 ( .C1(n7294), .C2(n10140), .A(n7190), .B(n7189), .ZN(n7191)
         );
  AOI21_X1 U9110 ( .B1(n7230), .B2(n10141), .A(n7191), .ZN(n7192) );
  OAI21_X1 U9111 ( .B1(n7193), .B2(n9352), .A(n7192), .ZN(P1_U3282) );
  INV_X1 U9112 ( .A(n7194), .ZN(n7195) );
  NOR2_X1 U9113 ( .A1(n7196), .A2(n7195), .ZN(n7200) );
  XNOR2_X1 U9114 ( .A(n7198), .B(n7197), .ZN(n7199) );
  XNOR2_X1 U9115 ( .A(n7200), .B(n7199), .ZN(n7208) );
  NAND2_X1 U9116 ( .A1(n8940), .A2(n8974), .ZN(n7202) );
  OAI211_X1 U9117 ( .C1(n8938), .C2(n7203), .A(n7202), .B(n7201), .ZN(n7205)
         );
  NOR2_X1 U9118 ( .A1(n9733), .A2(n9528), .ZN(n7204) );
  AOI211_X1 U9119 ( .C1(n7206), .C2(n8955), .A(n7205), .B(n7204), .ZN(n7207)
         );
  OAI21_X1 U9120 ( .B1(n7208), .B2(n8945), .A(n7207), .ZN(P1_U3231) );
  NAND2_X1 U9121 ( .A1(n7209), .A2(n7985), .ZN(n7210) );
  XNOR2_X1 U9122 ( .A(n7210), .B(n7932), .ZN(n9900) );
  INV_X1 U9123 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7215) );
  XNOR2_X1 U9124 ( .A(n7211), .B(n7932), .ZN(n7212) );
  NAND2_X1 U9125 ( .A1(n7212), .A2(n9866), .ZN(n7214) );
  AOI22_X1 U9126 ( .A1(n9862), .A2(n8379), .B1(n8377), .B2(n9860), .ZN(n7213)
         );
  AND2_X1 U9127 ( .A1(n7214), .A2(n7213), .ZN(n9904) );
  MUX2_X1 U9128 ( .A(n7215), .B(n9904), .S(n9878), .Z(n7218) );
  INV_X1 U9129 ( .A(n7251), .ZN(n7216) );
  AOI22_X1 U9130 ( .A1(n8658), .A2(n9901), .B1(n9877), .B2(n7216), .ZN(n7217)
         );
  OAI211_X1 U9131 ( .C1(n8661), .C2(n9900), .A(n7218), .B(n7217), .ZN(P2_U3227) );
  OR2_X1 U9132 ( .A1(n7220), .A2(n8004), .ZN(n7221) );
  NAND2_X1 U9133 ( .A1(n7219), .A2(n7221), .ZN(n9906) );
  INV_X1 U9134 ( .A(n8004), .ZN(n7934) );
  XNOR2_X1 U9135 ( .A(n7222), .B(n7934), .ZN(n7223) );
  NAND2_X1 U9136 ( .A1(n7223), .A2(n9866), .ZN(n7225) );
  AOI22_X1 U9137 ( .A1(n9862), .A2(n8378), .B1(n8376), .B2(n9860), .ZN(n7224)
         );
  OAI211_X1 U9138 ( .C1(n9870), .C2(n9906), .A(n7225), .B(n7224), .ZN(n9908)
         );
  INV_X1 U9139 ( .A(n7226), .ZN(n9874) );
  OAI22_X1 U9140 ( .A1(n9906), .A2(n9874), .B1(n7265), .B2(n8607), .ZN(n7227)
         );
  OAI21_X1 U9141 ( .B1(n9908), .B2(n7227), .A(n9878), .ZN(n7229) );
  NAND2_X1 U9142 ( .A1(n8658), .A2(n7257), .ZN(n7228) );
  OAI211_X1 U9143 ( .C1(n9793), .C2(n9878), .A(n7229), .B(n7228), .ZN(P2_U3226) );
  AOI211_X1 U9144 ( .C1(n7232), .C2(n9750), .A(n7231), .B(n7230), .ZN(n7238)
         );
  AOI22_X1 U9145 ( .A1(n7233), .A2(n9429), .B1(n9768), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7234) );
  OAI21_X1 U9146 ( .B1(n7238), .B2(n9768), .A(n7234), .ZN(P1_U3533) );
  INV_X1 U9147 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7235) );
  OAI22_X1 U9148 ( .A1(n7294), .A2(n9469), .B1(n9753), .B2(n7235), .ZN(n7236)
         );
  INV_X1 U9149 ( .A(n7236), .ZN(n7237) );
  OAI21_X1 U9150 ( .B1(n7238), .B2(n9752), .A(n7237), .ZN(P1_U3486) );
  XNOR2_X1 U9151 ( .A(n7246), .B(n4291), .ZN(n7256) );
  XNOR2_X1 U9152 ( .A(n7256), .B(n8378), .ZN(n7243) );
  AOI211_X1 U9153 ( .C1(n7243), .C2(n7242), .A(n8352), .B(n4372), .ZN(n7244)
         );
  INV_X1 U9154 ( .A(n7244), .ZN(n7250) );
  INV_X1 U9155 ( .A(n7245), .ZN(n7248) );
  INV_X1 U9156 ( .A(n8377), .ZN(n7317) );
  OAI22_X1 U9157 ( .A1(n8365), .A2(n7246), .B1(n7317), .B2(n8360), .ZN(n7247)
         );
  AOI211_X1 U9158 ( .C1(n8358), .C2(n8379), .A(n7248), .B(n7247), .ZN(n7249)
         );
  OAI211_X1 U9159 ( .C1(n7251), .C2(n8339), .A(n7250), .B(n7249), .ZN(P2_U3179) );
  INV_X1 U9160 ( .A(n7252), .ZN(n7255) );
  OAI222_X1 U9161 ( .A1(n7528), .A2(n7253), .B1(n8825), .B2(n7255), .C1(
        P2_U3151), .C2(n8468), .ZN(P2_U3276) );
  OAI222_X1 U9162 ( .A1(n7900), .A2(P1_U3086), .B1(n9478), .B2(n7255), .C1(
        n7254), .C2(n8222), .ZN(P1_U3336) );
  XNOR2_X1 U9163 ( .A(n7257), .B(n4291), .ZN(n7322) );
  XNOR2_X1 U9164 ( .A(n7322), .B(n8377), .ZN(n7258) );
  OAI21_X1 U9165 ( .B1(n7259), .B2(n7258), .A(n7323), .ZN(n7260) );
  NAND2_X1 U9166 ( .A1(n7260), .A2(n8354), .ZN(n7264) );
  NAND2_X1 U9167 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9807) );
  INV_X1 U9168 ( .A(n9807), .ZN(n7262) );
  INV_X1 U9169 ( .A(n8376), .ZN(n7356) );
  OAI22_X1 U9170 ( .A1(n8365), .A2(n9905), .B1(n7356), .B2(n8360), .ZN(n7261)
         );
  AOI211_X1 U9171 ( .C1(n8358), .C2(n8378), .A(n7262), .B(n7261), .ZN(n7263)
         );
  OAI211_X1 U9172 ( .C1(n7265), .C2(n8339), .A(n7264), .B(n7263), .ZN(P2_U3153) );
  XNOR2_X1 U9173 ( .A(n7267), .B(n7268), .ZN(n9744) );
  INV_X1 U9174 ( .A(n9744), .ZN(n7280) );
  OAI211_X1 U9175 ( .C1(n7270), .C2(n7269), .A(n7297), .B(n9665), .ZN(n7272)
         );
  AOI22_X1 U9176 ( .A1(n9343), .A2(n8973), .B1(n8971), .B2(n9345), .ZN(n7271)
         );
  NAND2_X1 U9177 ( .A1(n7272), .A2(n7271), .ZN(n9743) );
  INV_X1 U9178 ( .A(n7305), .ZN(n7273) );
  OAI21_X1 U9179 ( .B1(n9739), .B2(n7274), .A(n7273), .ZN(n9741) );
  AOI22_X1 U9180 ( .A1(n9677), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7340), .B2(
        n10146), .ZN(n7277) );
  NAND2_X1 U9181 ( .A1(n7275), .A2(n9652), .ZN(n7276) );
  OAI211_X1 U9182 ( .C1(n9741), .C2(n9112), .A(n7277), .B(n7276), .ZN(n7278)
         );
  AOI21_X1 U9183 ( .B1(n9743), .B2(n10141), .A(n7278), .ZN(n7279) );
  OAI21_X1 U9184 ( .B1(n7280), .B2(n9352), .A(n7279), .ZN(P1_U3281) );
  INV_X1 U9185 ( .A(n7281), .ZN(n7295) );
  OAI222_X1 U9186 ( .A1(n8825), .A2(n7295), .B1(n7283), .B2(P2_U3151), .C1(
        n7282), .C2(n7528), .ZN(P2_U3275) );
  AND3_X1 U9187 ( .A1(n7284), .A2(n7286), .A3(n7285), .ZN(n7287) );
  OAI21_X1 U9188 ( .B1(n7334), .B2(n7287), .A(n9531), .ZN(n7293) );
  NAND2_X1 U9189 ( .A1(n8940), .A2(n8972), .ZN(n7288) );
  NAND2_X1 U9190 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9576) );
  OAI211_X1 U9191 ( .C1(n8938), .C2(n7289), .A(n7288), .B(n9576), .ZN(n7290)
         );
  AOI21_X1 U9192 ( .B1(n7291), .B2(n8955), .A(n7290), .ZN(n7292) );
  OAI211_X1 U9193 ( .C1(n7294), .C2(n9528), .A(n7293), .B(n7292), .ZN(P1_U3236) );
  OAI222_X1 U9194 ( .A1(P1_U3086), .A2(n7296), .B1(n9478), .B2(n7295), .C1(
        n10016), .C2(n8222), .ZN(P1_U3335) );
  NAND2_X1 U9195 ( .A1(n7297), .A2(n7675), .ZN(n7299) );
  XNOR2_X1 U9196 ( .A(n7299), .B(n7298), .ZN(n7303) );
  NAND2_X1 U9197 ( .A1(n8972), .A2(n9343), .ZN(n7301) );
  NAND2_X1 U9198 ( .A1(n8970), .A2(n9345), .ZN(n7300) );
  AND2_X1 U9199 ( .A1(n7301), .A2(n7300), .ZN(n7393) );
  INV_X1 U9200 ( .A(n7393), .ZN(n7302) );
  AOI21_X1 U9201 ( .B1(n7303), .B2(n9665), .A(n7302), .ZN(n9747) );
  XNOR2_X1 U9202 ( .A(n7304), .B(n7790), .ZN(n9751) );
  NAND2_X1 U9203 ( .A1(n9751), .A2(n10150), .ZN(n7310) );
  OAI211_X1 U9204 ( .C1(n4772), .C2(n7305), .A(n9711), .B(n9426), .ZN(n9746)
         );
  INV_X1 U9205 ( .A(n9746), .ZN(n7308) );
  AOI22_X1 U9206 ( .A1(n9677), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7395), .B2(
        n10146), .ZN(n7306) );
  OAI21_X1 U9207 ( .B1(n4772), .B2(n10140), .A(n7306), .ZN(n7307) );
  AOI21_X1 U9208 ( .B1(n7308), .B2(n10148), .A(n7307), .ZN(n7309) );
  OAI211_X1 U9209 ( .C1(n9677), .C2(n9747), .A(n7310), .B(n7309), .ZN(P1_U3280) );
  NAND2_X1 U9210 ( .A1(n7219), .A2(n7311), .ZN(n7312) );
  XOR2_X1 U9211 ( .A(n7938), .B(n7312), .Z(n9912) );
  NAND2_X1 U9212 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  XNOR2_X1 U9213 ( .A(n7315), .B(n7938), .ZN(n7316) );
  OAI222_X1 U9214 ( .A1(n8633), .A2(n7317), .B1(n8646), .B2(n7487), .C1(n7316), 
        .C2(n8650), .ZN(n9914) );
  NAND2_X1 U9215 ( .A1(n9914), .A2(n9878), .ZN(n7321) );
  INV_X1 U9216 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7318) );
  OAI22_X1 U9217 ( .A1(n9878), .A2(n7318), .B1(n7331), .B2(n8607), .ZN(n7319)
         );
  AOI21_X1 U9218 ( .B1(n8658), .B2(n7325), .A(n7319), .ZN(n7320) );
  OAI211_X1 U9219 ( .C1(n9912), .C2(n8661), .A(n7321), .B(n7320), .ZN(P2_U3225) );
  INV_X1 U9220 ( .A(n7322), .ZN(n7324) );
  OAI21_X1 U9221 ( .B1(n7324), .B2(n8377), .A(n7323), .ZN(n7358) );
  XNOR2_X1 U9222 ( .A(n7325), .B(n4291), .ZN(n7355) );
  XNOR2_X1 U9223 ( .A(n7355), .B(n8376), .ZN(n7357) );
  XNOR2_X1 U9224 ( .A(n7358), .B(n7357), .ZN(n7326) );
  NAND2_X1 U9225 ( .A1(n7326), .A2(n8354), .ZN(n7330) );
  OAI22_X1 U9226 ( .A1(n8365), .A2(n9910), .B1(n7487), .B2(n8360), .ZN(n7327)
         );
  AOI211_X1 U9227 ( .C1(n8358), .C2(n8377), .A(n7328), .B(n7327), .ZN(n7329)
         );
  OAI211_X1 U9228 ( .C1(n7331), .C2(n8339), .A(n7330), .B(n7329), .ZN(P2_U3161) );
  NOR3_X1 U9229 ( .A1(n7334), .A2(n7333), .A3(n7332), .ZN(n7335) );
  OAI21_X1 U9230 ( .B1(n4367), .B2(n7335), .A(n9531), .ZN(n7342) );
  AOI21_X1 U9231 ( .B1(n8940), .B2(n8971), .A(n7336), .ZN(n7337) );
  OAI21_X1 U9232 ( .B1(n7338), .B2(n8938), .A(n7337), .ZN(n7339) );
  AOI21_X1 U9233 ( .B1(n7340), .B2(n8955), .A(n7339), .ZN(n7341) );
  OAI211_X1 U9234 ( .C1(n9739), .C2(n9528), .A(n7342), .B(n7341), .ZN(P1_U3224) );
  INV_X1 U9235 ( .A(n7343), .ZN(n7388) );
  OAI222_X1 U9236 ( .A1(n8825), .A2(n7388), .B1(n7958), .B2(P2_U3151), .C1(
        n7344), .C2(n7528), .ZN(P2_U3274) );
  NAND2_X1 U9237 ( .A1(n7345), .A2(n7943), .ZN(n7346) );
  NAND2_X1 U9238 ( .A1(n7347), .A2(n7346), .ZN(n9916) );
  XOR2_X1 U9239 ( .A(n7348), .B(n7943), .Z(n7349) );
  NAND2_X1 U9240 ( .A1(n7349), .A2(n9866), .ZN(n7351) );
  AOI22_X1 U9241 ( .A1(n9862), .A2(n8376), .B1(n8374), .B2(n9860), .ZN(n7350)
         );
  OAI211_X1 U9242 ( .C1(n9870), .C2(n9916), .A(n7351), .B(n7350), .ZN(n9917)
         );
  NAND2_X1 U9243 ( .A1(n9917), .A2(n9878), .ZN(n7354) );
  OAI22_X1 U9244 ( .A1(n9878), .A2(n9813), .B1(n7361), .B2(n8607), .ZN(n7352)
         );
  AOI21_X1 U9245 ( .B1(n8658), .B2(n9919), .A(n7352), .ZN(n7353) );
  OAI211_X1 U9246 ( .C1(n9916), .C2(n8487), .A(n7354), .B(n7353), .ZN(P2_U3224) );
  XNOR2_X1 U9247 ( .A(n9919), .B(n4291), .ZN(n7488) );
  XNOR2_X1 U9248 ( .A(n7488), .B(n8375), .ZN(n7359) );
  NAND2_X1 U9249 ( .A1(n7360), .A2(n7359), .ZN(n7490) );
  OAI211_X1 U9250 ( .C1(n7360), .C2(n7359), .A(n7490), .B(n8354), .ZN(n7367)
         );
  INV_X1 U9251 ( .A(n7361), .ZN(n7362) );
  NAND2_X1 U9252 ( .A1(n8362), .A2(n7362), .ZN(n7364) );
  NOR2_X1 U9253 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5283), .ZN(n9815) );
  AOI21_X1 U9254 ( .B1(n8358), .B2(n8376), .A(n9815), .ZN(n7363) );
  OAI211_X1 U9255 ( .C1(n7553), .C2(n8360), .A(n7364), .B(n7363), .ZN(n7365)
         );
  AOI21_X1 U9256 ( .B1(n9919), .B2(n8350), .A(n7365), .ZN(n7366) );
  NAND2_X1 U9257 ( .A1(n7367), .A2(n7366), .ZN(P2_U3171) );
  AOI21_X1 U9258 ( .B1(n7370), .B2(n7369), .A(n7368), .ZN(n7386) );
  AOI21_X1 U9259 ( .B1(n7373), .B2(n7372), .A(n7371), .ZN(n7377) );
  INV_X1 U9260 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7374) );
  OR2_X1 U9261 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7374), .ZN(n7491) );
  INV_X1 U9262 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7375) );
  OR2_X1 U9263 ( .A1(n9832), .A2(n7375), .ZN(n7376) );
  OAI211_X1 U9264 ( .C1(n7377), .C2(n9826), .A(n7491), .B(n7376), .ZN(n7383)
         );
  AOI21_X1 U9265 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7381) );
  NOR2_X1 U9266 ( .A1(n7381), .A2(n9852), .ZN(n7382) );
  AOI211_X1 U9267 ( .C1(n9817), .C2(n7384), .A(n7383), .B(n7382), .ZN(n7385)
         );
  OAI21_X1 U9268 ( .B1(n7386), .B2(n9848), .A(n7385), .ZN(P2_U3192) );
  OAI21_X1 U9269 ( .B1(n7391), .B2(n7390), .A(n7389), .ZN(n7392) );
  NAND2_X1 U9270 ( .A1(n7392), .A2(n9531), .ZN(n7397) );
  NAND2_X1 U9271 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9588) );
  OAI21_X1 U9272 ( .B1(n8952), .B2(n7393), .A(n9588), .ZN(n7394) );
  AOI21_X1 U9273 ( .B1(n8955), .B2(n7395), .A(n7394), .ZN(n7396) );
  OAI211_X1 U9274 ( .C1(n4772), .C2(n9528), .A(n7397), .B(n7396), .ZN(P1_U3234) );
  NOR2_X1 U9275 ( .A1(n8007), .A2(n4854), .ZN(n7941) );
  XOR2_X1 U9276 ( .A(n7398), .B(n7941), .Z(n9925) );
  INV_X1 U9277 ( .A(n9925), .ZN(n7408) );
  XOR2_X1 U9278 ( .A(n7941), .B(n7399), .Z(n7403) );
  OAI22_X1 U9279 ( .A1(n7487), .A2(n8633), .B1(n7556), .B2(n8646), .ZN(n7400)
         );
  AOI21_X1 U9280 ( .B1(n9925), .B2(n7401), .A(n7400), .ZN(n7402) );
  OAI21_X1 U9281 ( .B1(n8650), .B2(n7403), .A(n7402), .ZN(n9923) );
  NAND2_X1 U9282 ( .A1(n9923), .A2(n9878), .ZN(n7407) );
  OAI22_X1 U9283 ( .A1(n9878), .A2(n7404), .B1(n7493), .B2(n8607), .ZN(n7405)
         );
  AOI21_X1 U9284 ( .B1(n8658), .B2(n7496), .A(n7405), .ZN(n7406) );
  OAI211_X1 U9285 ( .C1(n7408), .C2(n8487), .A(n7407), .B(n7406), .ZN(P2_U3223) );
  AOI21_X1 U9286 ( .B1(n7411), .B2(n7410), .A(n7409), .ZN(n7428) );
  INV_X1 U9287 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7413) );
  OR2_X1 U9288 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7412), .ZN(n7546) );
  OAI21_X1 U9289 ( .B1(n9832), .B2(n7413), .A(n7546), .ZN(n7419) );
  AOI21_X1 U9290 ( .B1(n7416), .B2(n7415), .A(n7414), .ZN(n7417) );
  NOR2_X1 U9291 ( .A1(n7417), .A2(n9852), .ZN(n7418) );
  AOI211_X1 U9292 ( .C1(n9817), .C2(n7420), .A(n7419), .B(n7418), .ZN(n7427)
         );
  NAND2_X1 U9293 ( .A1(n7422), .A2(n7421), .ZN(n7423) );
  XNOR2_X1 U9294 ( .A(n7424), .B(n7423), .ZN(n7425) );
  NAND2_X1 U9295 ( .A1(n7425), .A2(n9843), .ZN(n7426) );
  OAI211_X1 U9296 ( .C1(n7428), .C2(n9848), .A(n7427), .B(n7426), .ZN(P2_U3194) );
  XNOR2_X1 U9297 ( .A(n7429), .B(n7432), .ZN(n7457) );
  INV_X1 U9298 ( .A(n7457), .ZN(n7440) );
  OAI21_X1 U9299 ( .B1(n7432), .B2(n7431), .A(n7430), .ZN(n7433) );
  NAND2_X1 U9300 ( .A1(n7433), .A2(n9665), .ZN(n7434) );
  AOI22_X1 U9301 ( .A1(n8969), .A2(n9345), .B1(n8970), .B2(n9343), .ZN(n8951)
         );
  NAND2_X1 U9302 ( .A1(n7434), .A2(n8951), .ZN(n7455) );
  INV_X1 U9303 ( .A(n9337), .ZN(n7435) );
  AOI211_X1 U9304 ( .C1(n7460), .C2(n4366), .A(n9740), .B(n7435), .ZN(n7456)
         );
  NAND2_X1 U9305 ( .A1(n7456), .A2(n10148), .ZN(n7437) );
  AOI22_X1 U9306 ( .A1(n9677), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8954), .B2(
        n10146), .ZN(n7436) );
  OAI211_X1 U9307 ( .C1(n8958), .C2(n10140), .A(n7437), .B(n7436), .ZN(n7438)
         );
  AOI21_X1 U9308 ( .B1(n10141), .B2(n7455), .A(n7438), .ZN(n7439) );
  OAI21_X1 U9309 ( .B1(n7440), .B2(n9352), .A(n7439), .ZN(P1_U3278) );
  XNOR2_X1 U9310 ( .A(n7441), .B(n7944), .ZN(n7442) );
  OAI222_X1 U9311 ( .A1(n8633), .A2(n7553), .B1(n8646), .B2(n7563), .C1(n7442), 
        .C2(n8650), .ZN(n9930) );
  INV_X1 U9312 ( .A(n9930), .ZN(n7449) );
  OAI21_X1 U9313 ( .B1(n7444), .B2(n7555), .A(n7443), .ZN(n9932) );
  INV_X1 U9314 ( .A(n7507), .ZN(n9929) );
  INV_X1 U9315 ( .A(n7445), .ZN(n7502) );
  AOI22_X1 U9316 ( .A1(n9881), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9877), .B2(
        n7502), .ZN(n7446) );
  OAI21_X1 U9317 ( .B1(n9929), .B2(n8481), .A(n7446), .ZN(n7447) );
  AOI21_X1 U9318 ( .B1(n9932), .B2(n8613), .A(n7447), .ZN(n7448) );
  OAI21_X1 U9319 ( .B1(n7449), .B2(n9881), .A(n7448), .ZN(P2_U3222) );
  INV_X1 U9320 ( .A(n7450), .ZN(n7454) );
  OAI222_X1 U9321 ( .A1(n7528), .A2(n7452), .B1(n8825), .B2(n7454), .C1(
        P2_U3151), .C2(n7451), .ZN(P2_U3273) );
  OAI222_X1 U9322 ( .A1(n6115), .A2(P1_U3086), .B1(n9478), .B2(n7454), .C1(
        n7453), .C2(n8222), .ZN(P1_U3333) );
  AOI211_X1 U9323 ( .C1(n7457), .C2(n9750), .A(n7456), .B(n7455), .ZN(n7462)
         );
  INV_X1 U9324 ( .A(n9469), .ZN(n7458) );
  AOI22_X1 U9325 ( .A1(n7460), .A2(n7458), .B1(n9752), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n7459) );
  OAI21_X1 U9326 ( .B1(n7462), .B2(n9752), .A(n7459), .ZN(P1_U3498) );
  AOI22_X1 U9327 ( .A1(n7460), .A2(n9429), .B1(n9768), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n7461) );
  OAI21_X1 U9328 ( .B1(n7462), .B2(n9768), .A(n7461), .ZN(P1_U3537) );
  AOI21_X1 U9329 ( .B1(n5315), .B2(n7464), .A(n7463), .ZN(n7478) );
  AOI21_X1 U9330 ( .B1(n7467), .B2(n7466), .A(n7465), .ZN(n7470) );
  AND2_X1 U9331 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7503) );
  INV_X1 U9332 ( .A(n7503), .ZN(n7469) );
  INV_X1 U9333 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10013) );
  OR2_X1 U9334 ( .A1(n9832), .A2(n10013), .ZN(n7468) );
  OAI211_X1 U9335 ( .C1(n7470), .C2(n9826), .A(n7469), .B(n7468), .ZN(n7475)
         );
  AOI21_X1 U9336 ( .B1(n9952), .B2(n7472), .A(n7471), .ZN(n7473) );
  NOR2_X1 U9337 ( .A1(n7473), .A2(n9852), .ZN(n7474) );
  AOI211_X1 U9338 ( .C1(n9817), .C2(n7476), .A(n7475), .B(n7474), .ZN(n7477)
         );
  OAI21_X1 U9339 ( .B1(n7478), .B2(n9848), .A(n7477), .ZN(P2_U3193) );
  INV_X1 U9340 ( .A(n7483), .ZN(n7481) );
  AOI21_X1 U9341 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8823), .A(n7479), .ZN(
        n7480) );
  OAI21_X1 U9342 ( .B1(n7481), .B2(n8825), .A(n7480), .ZN(P2_U3272) );
  NAND2_X1 U9343 ( .A1(n7483), .A2(n7482), .ZN(n7485) );
  INV_X1 U9344 ( .A(n7484), .ZN(n7911) );
  OAI211_X1 U9345 ( .C1(n7486), .C2(n8222), .A(n7485), .B(n7911), .ZN(P1_U3332) );
  XNOR2_X1 U9346 ( .A(n7562), .B(n8374), .ZN(n7500) );
  XNOR2_X1 U9347 ( .A(n7496), .B(n4291), .ZN(n7552) );
  XNOR2_X1 U9348 ( .A(n7500), .B(n7552), .ZN(n7498) );
  NAND2_X1 U9349 ( .A1(n8358), .A2(n8375), .ZN(n7492) );
  OAI211_X1 U9350 ( .C1(n7556), .C2(n8360), .A(n7492), .B(n7491), .ZN(n7495)
         );
  NOR2_X1 U9351 ( .A1(n8339), .A2(n7493), .ZN(n7494) );
  AOI211_X1 U9352 ( .C1(n7496), .C2(n8350), .A(n7495), .B(n7494), .ZN(n7497)
         );
  OAI21_X1 U9353 ( .B1(n7498), .B2(n8352), .A(n7497), .ZN(P2_U3157) );
  INV_X1 U9354 ( .A(n7552), .ZN(n7499) );
  OAI22_X1 U9355 ( .A1(n7500), .A2(n7499), .B1(n8374), .B2(n7562), .ZN(n7501)
         );
  XNOR2_X1 U9356 ( .A(n7944), .B(n4291), .ZN(n7551) );
  XNOR2_X1 U9357 ( .A(n7501), .B(n7551), .ZN(n7509) );
  NAND2_X1 U9358 ( .A1(n8362), .A2(n7502), .ZN(n7505) );
  AOI21_X1 U9359 ( .B1(n8358), .B2(n8374), .A(n7503), .ZN(n7504) );
  OAI211_X1 U9360 ( .C1(n7563), .C2(n8360), .A(n7505), .B(n7504), .ZN(n7506)
         );
  AOI21_X1 U9361 ( .B1(n7507), .B2(n8350), .A(n7506), .ZN(n7508) );
  OAI21_X1 U9362 ( .B1(n7509), .B2(n8352), .A(n7508), .ZN(P2_U3176) );
  INV_X1 U9363 ( .A(n7443), .ZN(n7510) );
  OAI21_X1 U9364 ( .B1(n7510), .B2(n8025), .A(n8034), .ZN(n7512) );
  NAND2_X1 U9365 ( .A1(n7512), .A2(n7511), .ZN(n7526) );
  NAND2_X1 U9366 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  XOR2_X1 U9367 ( .A(n8034), .B(n7515), .Z(n7516) );
  AOI222_X1 U9368 ( .A1(n9866), .A2(n7516), .B1(n8373), .B2(n9862), .C1(n8371), 
        .C2(n9860), .ZN(n7522) );
  MUX2_X1 U9369 ( .A(n7517), .B(n7522), .S(n9934), .Z(n7519) );
  NAND2_X1 U9370 ( .A1(n7568), .A2(n8806), .ZN(n7518) );
  OAI211_X1 U9371 ( .C1(n7526), .C2(n8787), .A(n7519), .B(n7518), .ZN(P2_U3426) );
  MUX2_X1 U9372 ( .A(n10079), .B(n7522), .S(n9954), .Z(n7521) );
  NAND2_X1 U9373 ( .A1(n7568), .A2(n8714), .ZN(n7520) );
  OAI211_X1 U9374 ( .C1(n8693), .C2(n7526), .A(n7521), .B(n7520), .ZN(P2_U3471) );
  MUX2_X1 U9375 ( .A(n4990), .B(n7522), .S(n9878), .Z(n7525) );
  INV_X1 U9376 ( .A(n7550), .ZN(n7523) );
  AOI22_X1 U9377 ( .A1(n7568), .A2(n8658), .B1(n9877), .B2(n7523), .ZN(n7524)
         );
  OAI211_X1 U9378 ( .C1(n7526), .C2(n8661), .A(n7525), .B(n7524), .ZN(P2_U3221) );
  INV_X1 U9379 ( .A(n7527), .ZN(n7531) );
  OAI222_X1 U9380 ( .A1(n8825), .A2(n7531), .B1(P2_U3151), .B2(n5687), .C1(
        n7529), .C2(n7528), .ZN(P2_U3271) );
  OAI222_X1 U9381 ( .A1(n7532), .A2(P1_U3086), .B1(n9478), .B2(n7531), .C1(
        n7530), .C2(n8222), .ZN(P1_U3331) );
  NAND2_X1 U9382 ( .A1(n7575), .A2(n7573), .ZN(n8033) );
  XOR2_X1 U9383 ( .A(n7574), .B(n8033), .Z(n7533) );
  AOI222_X1 U9384 ( .A1(n9866), .A2(n7533), .B1(n8372), .B2(n9862), .C1(n8655), 
        .C2(n9860), .ZN(n7542) );
  INV_X1 U9385 ( .A(n7542), .ZN(n7535) );
  INV_X1 U9386 ( .A(n7589), .ZN(n7598) );
  OAI22_X1 U9387 ( .A1(n7598), .A2(n8532), .B1(n7593), .B2(n8607), .ZN(n7534)
         );
  OAI21_X1 U9388 ( .B1(n7535), .B2(n7534), .A(n9878), .ZN(n7538) );
  NAND2_X1 U9389 ( .A1(n7511), .A2(n8031), .ZN(n7536) );
  XOR2_X1 U9390 ( .A(n8033), .B(n7536), .Z(n7543) );
  AOI22_X1 U9391 ( .A1(n7543), .A2(n8613), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9881), .ZN(n7537) );
  NAND2_X1 U9392 ( .A1(n7538), .A2(n7537), .ZN(P2_U3220) );
  INV_X1 U9393 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7539) );
  MUX2_X1 U9394 ( .A(n7539), .B(n7542), .S(n9934), .Z(n7541) );
  AOI22_X1 U9395 ( .A1(n7543), .A2(n8807), .B1(n8806), .B2(n7589), .ZN(n7540)
         );
  NAND2_X1 U9396 ( .A1(n7541), .A2(n7540), .ZN(P2_U3429) );
  MUX2_X1 U9397 ( .A(n10050), .B(n7542), .S(n9954), .Z(n7545) );
  AOI22_X1 U9398 ( .A1(n7543), .A2(n8715), .B1(n8714), .B2(n7589), .ZN(n7544)
         );
  NAND2_X1 U9399 ( .A1(n7545), .A2(n7544), .ZN(P2_U3472) );
  OAI21_X1 U9400 ( .B1(n8360), .B2(n7547), .A(n7546), .ZN(n7548) );
  AOI21_X1 U9401 ( .B1(n8358), .B2(n8373), .A(n7548), .ZN(n7549) );
  OAI21_X1 U9402 ( .B1(n7550), .B2(n8339), .A(n7549), .ZN(n7567) );
  AOI21_X1 U9403 ( .B1(n7553), .B2(n7552), .A(n7551), .ZN(n7561) );
  NAND2_X1 U9404 ( .A1(n8007), .A2(n4291), .ZN(n7554) );
  OAI211_X1 U9405 ( .C1(n7556), .C2(n4291), .A(n7555), .B(n7554), .ZN(n7560)
         );
  NAND2_X1 U9406 ( .A1(n8373), .A2(n4291), .ZN(n7557) );
  OAI211_X1 U9407 ( .C1(n4291), .C2(n7558), .A(n7944), .B(n7557), .ZN(n7559)
         );
  XNOR2_X1 U9408 ( .A(n7568), .B(n4291), .ZN(n7586) );
  XNOR2_X1 U9409 ( .A(n7586), .B(n7563), .ZN(n7564) );
  AOI211_X1 U9410 ( .C1(n7565), .C2(n7564), .A(n8352), .B(n7587), .ZN(n7566)
         );
  AOI211_X1 U9411 ( .C1(n7568), .C2(n8350), .A(n7567), .B(n7566), .ZN(n7569)
         );
  INV_X1 U9412 ( .A(n7569), .ZN(P2_U3164) );
  INV_X1 U9413 ( .A(n7570), .ZN(n7600) );
  AOI22_X1 U9414 ( .A1(n7571), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8823), .ZN(n7572) );
  OAI21_X1 U9415 ( .B1(n7600), .B2(n8825), .A(n7572), .ZN(P2_U3270) );
  NAND2_X1 U9416 ( .A1(n7574), .A2(n7573), .ZN(n7576) );
  NAND2_X1 U9417 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  XNOR2_X1 U9418 ( .A(n7577), .B(n8040), .ZN(n7578) );
  AOI222_X1 U9419 ( .A1(n9866), .A2(n7578), .B1(n8371), .B2(n9862), .C1(n8370), 
        .C2(n9860), .ZN(n8720) );
  INV_X1 U9420 ( .A(n8720), .ZN(n7580) );
  INV_X1 U9421 ( .A(n8240), .ZN(n8721) );
  OAI22_X1 U9422 ( .A1(n8721), .A2(n8532), .B1(n8238), .B2(n8607), .ZN(n7579)
         );
  OAI21_X1 U9423 ( .B1(n7580), .B2(n7579), .A(n9878), .ZN(n7584) );
  NAND2_X1 U9424 ( .A1(n7582), .A2(n8040), .ZN(n8718) );
  NAND3_X1 U9425 ( .A1(n7581), .A2(n8718), .A3(n8613), .ZN(n7583) );
  OAI211_X1 U9426 ( .C1(n9878), .C2(n7585), .A(n7584), .B(n7583), .ZN(P2_U3219) );
  INV_X1 U9427 ( .A(n7586), .ZN(n7588) );
  XNOR2_X1 U9428 ( .A(n7589), .B(n4291), .ZN(n8149) );
  XNOR2_X1 U9429 ( .A(n8149), .B(n8371), .ZN(n7590) );
  NAND2_X1 U9430 ( .A1(n7591), .A2(n7590), .ZN(n8150) );
  OAI21_X1 U9431 ( .B1(n7591), .B2(n7590), .A(n8150), .ZN(n7592) );
  NAND2_X1 U9432 ( .A1(n7592), .A2(n8354), .ZN(n7597) );
  NAND2_X1 U9433 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8390) );
  OAI21_X1 U9434 ( .B1(n8360), .B2(n8153), .A(n8390), .ZN(n7595) );
  NOR2_X1 U9435 ( .A1(n8339), .A2(n7593), .ZN(n7594) );
  AOI211_X1 U9436 ( .C1(n8358), .C2(n8372), .A(n7595), .B(n7594), .ZN(n7596)
         );
  OAI211_X1 U9437 ( .C1(n7598), .C2(n8365), .A(n7597), .B(n7596), .ZN(P2_U3174) );
  OAI222_X1 U9438 ( .A1(n7601), .A2(P1_U3086), .B1(n9478), .B2(n7600), .C1(
        n7599), .C2(n8222), .ZN(P1_U3330) );
  INV_X1 U9439 ( .A(n7602), .ZN(n7605) );
  AOI22_X1 U9440 ( .A1(n7603), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8823), .ZN(n7604) );
  OAI21_X1 U9441 ( .B1(n7605), .B2(n8825), .A(n7604), .ZN(P2_U3269) );
  OAI222_X1 U9442 ( .A1(n7606), .A2(P1_U3086), .B1(n9478), .B2(n7605), .C1(
        n10108), .C2(n8222), .ZN(P1_U3329) );
  INV_X1 U9443 ( .A(n7607), .ZN(n7627) );
  AOI21_X1 U9444 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8823), .A(n7608), .ZN(
        n7609) );
  OAI21_X1 U9445 ( .B1(n7627), .B2(n8825), .A(n7609), .ZN(P2_U3268) );
  AOI21_X1 U9446 ( .B1(n7610), .B2(n7611), .A(n4305), .ZN(n7616) );
  INV_X1 U9447 ( .A(n7621), .ZN(n7614) );
  INV_X1 U9448 ( .A(n8360), .ZN(n8305) );
  AOI22_X1 U9449 ( .A1(n8305), .A2(n8380), .B1(n8358), .B2(n7098), .ZN(n7612)
         );
  OAI21_X1 U9450 ( .B1(n7099), .B2(n8365), .A(n7612), .ZN(n7613) );
  AOI21_X1 U9451 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7614), .A(n7613), .ZN(
        n7615) );
  OAI21_X1 U9452 ( .B1(n8352), .B2(n7616), .A(n7615), .ZN(P2_U3162) );
  XOR2_X1 U9453 ( .A(n7618), .B(n7617), .Z(n7625) );
  INV_X1 U9454 ( .A(n8358), .ZN(n8316) );
  OAI22_X1 U9455 ( .A1(n8316), .A2(n6763), .B1(n7619), .B2(n8360), .ZN(n7623)
         );
  NOR2_X1 U9456 ( .A1(n7621), .A2(n7620), .ZN(n7622) );
  AOI211_X1 U9457 ( .C1(n5149), .C2(n8350), .A(n7623), .B(n7622), .ZN(n7624)
         );
  OAI21_X1 U9458 ( .B1(n8352), .B2(n7625), .A(n7624), .ZN(P2_U3177) );
  OAI222_X1 U9459 ( .A1(P1_U3086), .A2(n8994), .B1(n9478), .B2(n7627), .C1(
        n7626), .C2(n8222), .ZN(P1_U3328) );
  INV_X1 U9460 ( .A(n7628), .ZN(n8821) );
  OAI222_X1 U9461 ( .A1(P1_U3086), .A2(n7630), .B1(n9478), .B2(n8821), .C1(
        n7629), .C2(n8222), .ZN(P1_U3326) );
  INV_X1 U9462 ( .A(n7631), .ZN(n8826) );
  OAI222_X1 U9463 ( .A1(P1_U3086), .A2(n6138), .B1(n9478), .B2(n8826), .C1(
        n7632), .C2(n8222), .ZN(P1_U3327) );
  NAND2_X1 U9464 ( .A1(n9201), .A2(n7633), .ZN(n7814) );
  AND2_X1 U9465 ( .A1(n7874), .A2(n7698), .ZN(n7873) );
  INV_X1 U9466 ( .A(n7760), .ZN(n7897) );
  AOI22_X1 U9467 ( .A1(n7634), .A2(n9291), .B1(n7897), .B2(n9256), .ZN(n7637)
         );
  INV_X1 U9468 ( .A(n9258), .ZN(n7636) );
  NAND2_X1 U9469 ( .A1(n9311), .A2(n7760), .ZN(n7635) );
  OAI22_X1 U9470 ( .A1(n7637), .A2(n7876), .B1(n7636), .B2(n7635), .ZN(n7707)
         );
  NAND2_X1 U9471 ( .A1(n7638), .A2(n7697), .ZN(n7871) );
  NAND2_X1 U9472 ( .A1(n7871), .A2(n7760), .ZN(n7639) );
  OAI211_X1 U9473 ( .C1(n7873), .C2(n7760), .A(n7707), .B(n7639), .ZN(n7710)
         );
  INV_X1 U9474 ( .A(n7690), .ZN(n7684) );
  AND2_X1 U9475 ( .A1(n7641), .A2(n7640), .ZN(n7867) );
  INV_X1 U9476 ( .A(n7867), .ZN(n7642) );
  OR2_X1 U9477 ( .A1(n7642), .A2(n7685), .ZN(n7643) );
  AND2_X1 U9478 ( .A1(n7643), .A2(n7686), .ZN(n7863) );
  AND2_X1 U9479 ( .A1(n7647), .A2(n7644), .ZN(n7843) );
  AND2_X1 U9480 ( .A1(n7648), .A2(n7852), .ZN(n7652) );
  INV_X1 U9481 ( .A(n7654), .ZN(n7850) );
  AOI21_X1 U9482 ( .B1(n7649), .B2(n7652), .A(n7850), .ZN(n7657) );
  NAND2_X1 U9483 ( .A1(n7651), .A2(n7650), .ZN(n7844) );
  OAI21_X1 U9484 ( .B1(n7653), .B2(n7844), .A(n7652), .ZN(n7655) );
  NAND2_X1 U9485 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  MUX2_X1 U9486 ( .A(n7657), .B(n7656), .S(n7760), .Z(n7659) );
  NAND2_X1 U9487 ( .A1(n7671), .A2(n7661), .ZN(n7663) );
  AOI21_X1 U9488 ( .B1(n4475), .B2(n7771), .A(n7664), .ZN(n7673) );
  INV_X1 U9489 ( .A(n7783), .ZN(n7666) );
  OAI21_X1 U9490 ( .B1(n7673), .B2(n7666), .A(n7665), .ZN(n7667) );
  NAND3_X1 U9491 ( .A1(n7667), .A2(n7674), .A3(n7853), .ZN(n7670) );
  AND2_X1 U9492 ( .A1(n7860), .A2(n7668), .ZN(n7770) );
  AOI21_X1 U9493 ( .B1(n7670), .B2(n7770), .A(n7669), .ZN(n7680) );
  INV_X1 U9494 ( .A(n7671), .ZN(n7672) );
  OAI21_X1 U9495 ( .B1(n7673), .B2(n7672), .A(n7853), .ZN(n7676) );
  NAND2_X1 U9496 ( .A1(n7675), .A2(n7674), .ZN(n7861) );
  AOI21_X1 U9497 ( .B1(n7676), .B2(n7856), .A(n7861), .ZN(n7678) );
  NOR2_X1 U9498 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  MUX2_X1 U9499 ( .A(n7680), .B(n7679), .S(n7760), .Z(n7688) );
  NAND3_X1 U9500 ( .A1(n7688), .A2(n7867), .A3(n7690), .ZN(n7683) );
  NAND2_X1 U9501 ( .A1(n7690), .A2(n7864), .ZN(n7681) );
  NAND2_X1 U9502 ( .A1(n7681), .A2(n7868), .ZN(n7692) );
  INV_X1 U9503 ( .A(n7692), .ZN(n7682) );
  OAI211_X1 U9504 ( .C1(n7684), .C2(n7863), .A(n7683), .B(n7682), .ZN(n7696)
         );
  OAI211_X1 U9505 ( .C1(n7688), .C2(n7687), .A(n7686), .B(n7685), .ZN(n7694)
         );
  NAND2_X1 U9506 ( .A1(n7690), .A2(n7689), .ZN(n7869) );
  NOR2_X1 U9507 ( .A1(n7869), .A2(n7691), .ZN(n7693) );
  AOI21_X1 U9508 ( .B1(n7694), .B2(n7693), .A(n7692), .ZN(n7695) );
  MUX2_X1 U9509 ( .A(n7696), .B(n7695), .S(n7760), .Z(n7700) );
  NAND4_X1 U9510 ( .A1(n7868), .A2(n8958), .A3(n7897), .A4(n9344), .ZN(n7699)
         );
  NAND2_X1 U9511 ( .A1(n7698), .A2(n7697), .ZN(n9320) );
  AOI21_X1 U9512 ( .B1(n7700), .B2(n7699), .A(n9320), .ZN(n7709) );
  AOI21_X1 U9513 ( .B1(n8862), .B2(n7897), .A(n9307), .ZN(n7703) );
  AOI21_X1 U9514 ( .B1(n9295), .B2(n7760), .A(n9405), .ZN(n7702) );
  OAI211_X1 U9515 ( .C1(n7703), .C2(n7702), .A(n7878), .B(n7701), .ZN(n7706)
         );
  MUX2_X1 U9516 ( .A(n7712), .B(n7711), .S(n7760), .Z(n7713) );
  OR2_X1 U9517 ( .A1(n9380), .A2(n7714), .ZN(n7716) );
  INV_X1 U9518 ( .A(n7716), .ZN(n7717) );
  AND2_X1 U9519 ( .A1(n7716), .A2(n7715), .ZN(n7806) );
  INV_X1 U9520 ( .A(n9201), .ZN(n7718) );
  AOI21_X1 U9521 ( .B1(n7897), .B2(n7718), .A(n9202), .ZN(n7722) );
  INV_X1 U9522 ( .A(n7809), .ZN(n7720) );
  INV_X1 U9523 ( .A(n7817), .ZN(n7719) );
  AOI21_X1 U9524 ( .B1(n7723), .B2(n7722), .A(n7721), .ZN(n7730) );
  NAND2_X1 U9525 ( .A1(n7733), .A2(n7729), .ZN(n7821) );
  AOI21_X1 U9526 ( .B1(n7730), .B2(n7812), .A(n7821), .ZN(n7726) );
  OR2_X1 U9527 ( .A1(n9177), .A2(n7724), .ZN(n7725) );
  NOR2_X1 U9528 ( .A1(n7726), .A2(n7823), .ZN(n7727) );
  NAND2_X1 U9529 ( .A1(n7743), .A2(n7732), .ZN(n7824) );
  OAI21_X1 U9530 ( .B1(n7727), .B2(n7824), .A(n7828), .ZN(n7740) );
  INV_X1 U9531 ( .A(n7812), .ZN(n7728) );
  INV_X1 U9532 ( .A(n7731), .ZN(n7738) );
  INV_X1 U9533 ( .A(n7732), .ZN(n7736) );
  INV_X1 U9534 ( .A(n7733), .ZN(n7735) );
  OAI21_X1 U9535 ( .B1(n7736), .B2(n7735), .A(n7734), .ZN(n7737) );
  INV_X1 U9536 ( .A(n7828), .ZN(n9120) );
  AOI21_X1 U9537 ( .B1(n7738), .B2(n7737), .A(n9120), .ZN(n7739) );
  INV_X1 U9538 ( .A(n8960), .ZN(n7741) );
  NAND2_X1 U9539 ( .A1(n7742), .A2(n7741), .ZN(n7746) );
  NAND2_X1 U9540 ( .A1(n7827), .A2(n7746), .ZN(n9122) );
  INV_X1 U9541 ( .A(n7743), .ZN(n7744) );
  INV_X1 U9542 ( .A(n7746), .ZN(n7885) );
  INV_X1 U9543 ( .A(n7827), .ZN(n7747) );
  INV_X1 U9544 ( .A(n7759), .ZN(n7750) );
  MUX2_X1 U9545 ( .A(n7750), .B(n7760), .S(n9115), .Z(n7767) );
  NAND2_X1 U9546 ( .A1(n7751), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9547 ( .A1(n7752), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U9548 ( .A1(n7753), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7754) );
  NAND3_X1 U9549 ( .A1(n7756), .A2(n7755), .A3(n7754), .ZN(n8959) );
  NAND2_X1 U9550 ( .A1(n7757), .A2(n8959), .ZN(n7829) );
  NAND2_X1 U9551 ( .A1(n7901), .A2(n7829), .ZN(n7766) );
  NAND2_X1 U9552 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  NAND3_X1 U9553 ( .A1(n7764), .A2(n9109), .A3(n8959), .ZN(n7765) );
  INV_X1 U9554 ( .A(n9122), .ZN(n9129) );
  INV_X1 U9555 ( .A(n8959), .ZN(n9123) );
  NOR2_X1 U9556 ( .A1(n9115), .A2(n9123), .ZN(n7889) );
  INV_X1 U9557 ( .A(n7889), .ZN(n7803) );
  XNOR2_X1 U9558 ( .A(n9265), .B(n7769), .ZN(n9260) );
  INV_X1 U9559 ( .A(n7871), .ZN(n7796) );
  INV_X1 U9560 ( .A(n7873), .ZN(n7794) );
  INV_X1 U9561 ( .A(n7861), .ZN(n7789) );
  INV_X1 U9562 ( .A(n7770), .ZN(n7787) );
  INV_X1 U9563 ( .A(n7771), .ZN(n7782) );
  NOR2_X1 U9564 ( .A1(n7773), .A2(n7772), .ZN(n7780) );
  NOR2_X1 U9565 ( .A1(n9714), .A2(n7774), .ZN(n7779) );
  NOR2_X1 U9566 ( .A1(n7775), .A2(n9669), .ZN(n7778) );
  NOR2_X1 U9567 ( .A1(n9681), .A2(n7776), .ZN(n7777) );
  NAND4_X1 U9568 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n7781)
         );
  NOR2_X1 U9569 ( .A1(n7782), .A2(n7781), .ZN(n7784) );
  NAND4_X1 U9570 ( .A1(n7785), .A2(n7848), .A3(n7784), .A4(n7783), .ZN(n7786)
         );
  NOR2_X1 U9571 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  NAND3_X1 U9572 ( .A1(n7790), .A2(n7789), .A3(n7788), .ZN(n7792) );
  OR4_X1 U9573 ( .A1(n9334), .A2(n7792), .A3(n7791), .A4(n9422), .ZN(n7793) );
  NOR2_X1 U9574 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  NAND4_X1 U9575 ( .A1(n7634), .A2(n9294), .A3(n7796), .A4(n7795), .ZN(n7797)
         );
  NOR3_X1 U9576 ( .A1(n9241), .A2(n9260), .A3(n7797), .ZN(n7798) );
  NAND4_X1 U9577 ( .A1(n9190), .A2(n9208), .A3(n7798), .A4(n9219), .ZN(n7799)
         );
  OR3_X1 U9578 ( .A1(n9157), .A2(n7799), .A3(n9175), .ZN(n7800) );
  NOR2_X1 U9579 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  NAND2_X1 U9580 ( .A1(n9115), .A2(n9123), .ZN(n7888) );
  AND4_X1 U9581 ( .A1(n7803), .A2(n9129), .A3(n7802), .A4(n7888), .ZN(n7804)
         );
  AND3_X1 U9582 ( .A1(n7901), .A2(n7804), .A3(n7893), .ZN(n7835) );
  INV_X1 U9583 ( .A(n7893), .ZN(n7898) );
  AOI211_X1 U9584 ( .C1(n7889), .C2(n9109), .A(n7805), .B(n7898), .ZN(n7833)
         );
  INV_X1 U9585 ( .A(n7806), .ZN(n7807) );
  NAND2_X1 U9586 ( .A1(n7807), .A2(n9201), .ZN(n7808) );
  NAND2_X1 U9587 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  NAND2_X1 U9588 ( .A1(n7810), .A2(n7817), .ZN(n7811) );
  NAND2_X1 U9589 ( .A1(n7812), .A2(n7811), .ZN(n7819) );
  OR3_X1 U9590 ( .A1(n7823), .A2(n7813), .A3(n7819), .ZN(n7883) );
  NOR2_X1 U9591 ( .A1(n7883), .A2(n4312), .ZN(n7826) );
  INV_X1 U9592 ( .A(n7814), .ZN(n7816) );
  AND3_X1 U9593 ( .A1(n7817), .A2(n7816), .A3(n7815), .ZN(n7818) );
  NOR2_X1 U9594 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  NOR2_X1 U9595 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  NOR2_X1 U9596 ( .A1(n7823), .A2(n7822), .ZN(n7825) );
  OR2_X1 U9597 ( .A1(n7825), .A2(n7824), .ZN(n7881) );
  NOR2_X1 U9598 ( .A1(n7826), .A2(n7881), .ZN(n7831) );
  NAND2_X1 U9599 ( .A1(n7827), .A2(n7828), .ZN(n7836) );
  AOI21_X1 U9600 ( .B1(n9115), .B2(n7829), .A(n7885), .ZN(n7830) );
  OAI211_X1 U9601 ( .C1(n7831), .C2(n7836), .A(n7901), .B(n7830), .ZN(n7832)
         );
  AOI21_X1 U9602 ( .B1(n7833), .B2(n7832), .A(n7835), .ZN(n7834) );
  NOR2_X1 U9603 ( .A1(n7900), .A2(n7905), .ZN(n7895) );
  INV_X1 U9604 ( .A(n7836), .ZN(n7887) );
  NAND2_X1 U9605 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  AOI211_X1 U9606 ( .C1(n9691), .C2(n8983), .A(n7840), .B(n7839), .ZN(n7841)
         );
  NOR2_X1 U9607 ( .A1(n7842), .A2(n7841), .ZN(n7847) );
  INV_X1 U9608 ( .A(n7843), .ZN(n7846) );
  INV_X1 U9609 ( .A(n7844), .ZN(n7845) );
  OAI21_X1 U9610 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7851) );
  INV_X1 U9611 ( .A(n7848), .ZN(n7849) );
  AOI211_X1 U9612 ( .C1(n7852), .C2(n7851), .A(n7850), .B(n7849), .ZN(n7855)
         );
  INV_X1 U9613 ( .A(n7853), .ZN(n7854) );
  NOR2_X1 U9614 ( .A1(n7855), .A2(n7854), .ZN(n7859) );
  INV_X1 U9615 ( .A(n7856), .ZN(n7857) );
  AOI21_X1 U9616 ( .B1(n7859), .B2(n7858), .A(n7857), .ZN(n7862) );
  OAI21_X1 U9617 ( .B1(n7862), .B2(n7861), .A(n7860), .ZN(n7866) );
  INV_X1 U9618 ( .A(n7863), .ZN(n7865) );
  AOI211_X1 U9619 ( .C1(n7867), .C2(n7866), .A(n7865), .B(n7864), .ZN(n7870)
         );
  OAI21_X1 U9620 ( .B1(n7870), .B2(n7869), .A(n7868), .ZN(n7872) );
  AOI21_X1 U9621 ( .B1(n7873), .B2(n7872), .A(n7871), .ZN(n7877) );
  INV_X1 U9622 ( .A(n7874), .ZN(n7875) );
  NOR3_X1 U9623 ( .A1(n7877), .A2(n7876), .A3(n7875), .ZN(n7880) );
  INV_X1 U9624 ( .A(n7878), .ZN(n7879) );
  NOR2_X1 U9625 ( .A1(n7880), .A2(n7879), .ZN(n7884) );
  INV_X1 U9626 ( .A(n7881), .ZN(n7882) );
  OAI21_X1 U9627 ( .B1(n7884), .B2(n7883), .A(n7882), .ZN(n7886) );
  AOI21_X1 U9628 ( .B1(n7887), .B2(n7886), .A(n7885), .ZN(n7890) );
  OAI21_X1 U9629 ( .B1(n7890), .B2(n7889), .A(n7888), .ZN(n7892) );
  INV_X1 U9630 ( .A(n7901), .ZN(n7891) );
  MUX2_X1 U9631 ( .A(n7896), .B(n7895), .S(n7894), .Z(n7904) );
  OAI211_X1 U9632 ( .C1(n7901), .C2(n7900), .A(n7899), .B(n6115), .ZN(n7902)
         );
  NAND3_X1 U9633 ( .A1(n7907), .A2(n8999), .A3(n7906), .ZN(n7908) );
  OAI211_X1 U9634 ( .C1(n7909), .C2(n7911), .A(n7908), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7910) );
  INV_X1 U9635 ( .A(n7925), .ZN(n7918) );
  NAND2_X1 U9636 ( .A1(n8221), .A2(n7914), .ZN(n7913) );
  NAND2_X1 U9637 ( .A1(n5155), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U9638 ( .A1(n8813), .A2(n7914), .ZN(n7917) );
  NAND2_X1 U9639 ( .A1(n7915), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7916) );
  OAI22_X1 U9640 ( .A1(n7919), .A2(n7918), .B1(n8667), .B2(n8727), .ZN(n7923)
         );
  OR2_X1 U9641 ( .A1(n8727), .A2(n8474), .ZN(n8134) );
  INV_X1 U9642 ( .A(n8367), .ZN(n7921) );
  NAND2_X1 U9643 ( .A1(n8731), .A2(n7921), .ZN(n8125) );
  NAND2_X1 U9644 ( .A1(n8134), .A2(n8112), .ZN(n7924) );
  NOR2_X1 U9645 ( .A1(n8731), .A2(n7921), .ZN(n8116) );
  OAI21_X1 U9646 ( .B1(n8116), .B2(n8474), .A(n8727), .ZN(n7922) );
  OAI21_X1 U9647 ( .B1(n7923), .B2(n7924), .A(n7922), .ZN(n7959) );
  INV_X1 U9648 ( .A(n7924), .ZN(n7954) );
  INV_X1 U9649 ( .A(n8116), .ZN(n7926) );
  NAND2_X1 U9650 ( .A1(n7926), .A2(n7925), .ZN(n8120) );
  INV_X1 U9651 ( .A(n7927), .ZN(n8090) );
  INV_X1 U9652 ( .A(n8528), .ZN(n8098) );
  INV_X1 U9653 ( .A(n8107), .ZN(n7928) );
  INV_X1 U9654 ( .A(n8083), .ZN(n8540) );
  NAND2_X1 U9655 ( .A1(n8094), .A2(n8085), .ZN(n8542) );
  INV_X1 U9656 ( .A(n8582), .ZN(n7949) );
  NAND2_X1 U9657 ( .A1(n8053), .A2(n7929), .ZN(n8065) );
  NAND2_X1 U9658 ( .A1(n7931), .A2(n7930), .ZN(n8050) );
  NOR4_X1 U9659 ( .A1(n7934), .A2(n7933), .A3(n8723), .A4(n7932), .ZN(n7937)
         );
  NAND3_X1 U9660 ( .A1(n7937), .A2(n7936), .A3(n7935), .ZN(n7939) );
  NOR4_X1 U9661 ( .A1(n9865), .A2(n7940), .A3(n7939), .A4(n7938), .ZN(n7942)
         );
  NAND2_X1 U9662 ( .A1(n7942), .A2(n7941), .ZN(n7945) );
  NOR4_X1 U9663 ( .A1(n8034), .A2(n7945), .A3(n7944), .A4(n7943), .ZN(n7946)
         );
  NAND4_X1 U9664 ( .A1(n8652), .A2(n7946), .A3(n8033), .A4(n5378), .ZN(n7947)
         );
  NOR4_X1 U9665 ( .A1(n8065), .A2(n8050), .A3(n8630), .A4(n7947), .ZN(n7948)
         );
  NAND4_X1 U9666 ( .A1(n8570), .A2(n7949), .A3(n7948), .A4(n8596), .ZN(n7950)
         );
  NOR4_X1 U9667 ( .A1(n8547), .A2(n8556), .A3(n8542), .A4(n7950), .ZN(n7951)
         );
  NAND4_X1 U9668 ( .A1(n8100), .A2(n8098), .A3(n8499), .A4(n7951), .ZN(n7952)
         );
  NOR3_X1 U9669 ( .A1(n8120), .A2(n8491), .A3(n7952), .ZN(n7953) );
  NAND2_X1 U9670 ( .A1(n8727), .A2(n8474), .ZN(n8132) );
  NAND3_X1 U9671 ( .A1(n7954), .A2(n7953), .A3(n8132), .ZN(n7955) );
  MUX2_X1 U9672 ( .A(n8505), .B(n8741), .S(n8127), .Z(n8113) );
  INV_X1 U9673 ( .A(n7960), .ZN(n7961) );
  NAND2_X1 U9674 ( .A1(n8072), .A2(n7961), .ZN(n7962) );
  AND2_X1 U9675 ( .A1(n8695), .A2(n8336), .ZN(n8054) );
  MUX2_X1 U9676 ( .A(n7962), .B(n8054), .S(n8128), .Z(n7964) );
  NOR2_X1 U9677 ( .A1(n7964), .A2(n7963), .ZN(n8077) );
  AND2_X1 U9678 ( .A1(n7968), .A2(n7965), .ZN(n7967) );
  OAI21_X1 U9679 ( .B1(n7967), .B2(n7966), .A(n7969), .ZN(n7973) );
  NAND2_X1 U9680 ( .A1(n7969), .A2(n7968), .ZN(n7971) );
  NAND2_X1 U9681 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  NAND2_X1 U9682 ( .A1(n7991), .A2(n7974), .ZN(n7977) );
  NAND2_X1 U9683 ( .A1(n8380), .A2(n9871), .ZN(n7975) );
  NAND2_X1 U9684 ( .A1(n7983), .A2(n7975), .ZN(n7976) );
  INV_X1 U9685 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U9686 ( .A1(n7982), .A2(n7981), .ZN(n7995) );
  INV_X1 U9687 ( .A(n7983), .ZN(n7986) );
  OAI211_X1 U9688 ( .C1(n7995), .C2(n7986), .A(n7985), .B(n7984), .ZN(n7990)
         );
  AND2_X1 U9689 ( .A1(n7996), .A2(n7993), .ZN(n7989) );
  INV_X1 U9690 ( .A(n7987), .ZN(n7988) );
  AOI21_X1 U9691 ( .B1(n7990), .B2(n7989), .A(n7988), .ZN(n8000) );
  INV_X1 U9692 ( .A(n7991), .ZN(n7994) );
  OAI211_X1 U9693 ( .C1(n7995), .C2(n7994), .A(n7993), .B(n7992), .ZN(n7998)
         );
  INV_X1 U9694 ( .A(n7996), .ZN(n7997) );
  AOI21_X1 U9695 ( .B1(n7998), .B2(n4871), .A(n7997), .ZN(n7999) );
  NAND2_X1 U9696 ( .A1(n8008), .A2(n8001), .ZN(n8003) );
  NAND2_X1 U9697 ( .A1(n8012), .A2(n8011), .ZN(n8002) );
  INV_X1 U9698 ( .A(n8014), .ZN(n8005) );
  NAND3_X1 U9699 ( .A1(n8006), .A2(n8005), .A3(n8004), .ZN(n8019) );
  INV_X1 U9700 ( .A(n8007), .ZN(n8020) );
  OAI211_X1 U9701 ( .C1(n8014), .C2(n8009), .A(n8020), .B(n8008), .ZN(n8016)
         );
  AND2_X1 U9702 ( .A1(n8011), .A2(n8010), .ZN(n8013) );
  OAI211_X1 U9703 ( .C1(n8014), .C2(n8013), .A(n8023), .B(n8012), .ZN(n8015)
         );
  MUX2_X1 U9704 ( .A(n8016), .B(n8015), .S(n8128), .Z(n8017) );
  INV_X1 U9705 ( .A(n8017), .ZN(n8018) );
  NAND3_X1 U9706 ( .A1(n8024), .A2(n8026), .A3(n8020), .ZN(n8022) );
  NAND2_X1 U9707 ( .A1(n8022), .A2(n8021), .ZN(n8029) );
  AOI21_X1 U9708 ( .B1(n8027), .B2(n8026), .A(n8025), .ZN(n8028) );
  MUX2_X1 U9709 ( .A(n8031), .B(n8030), .S(n8127), .Z(n8032) );
  OAI211_X1 U9710 ( .C1(n8035), .C2(n8034), .A(n8033), .B(n8032), .ZN(n8042)
         );
  INV_X1 U9711 ( .A(n8036), .ZN(n8037) );
  MUX2_X1 U9712 ( .A(n8038), .B(n8037), .S(n8128), .Z(n8039) );
  NOR2_X1 U9713 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  NAND2_X1 U9714 ( .A1(n8042), .A2(n8041), .ZN(n8046) );
  NAND2_X1 U9715 ( .A1(n8240), .A2(n8127), .ZN(n8044) );
  OR2_X1 U9716 ( .A1(n8240), .A2(n8127), .ZN(n8043) );
  MUX2_X1 U9717 ( .A(n8044), .B(n8043), .S(n8655), .Z(n8045) );
  NAND2_X1 U9718 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  INV_X1 U9719 ( .A(n8618), .ZN(n8049) );
  NAND2_X1 U9720 ( .A1(n8050), .A2(n8128), .ZN(n8051) );
  NAND2_X1 U9721 ( .A1(n8052), .A2(n8051), .ZN(n8064) );
  NAND3_X1 U9722 ( .A1(n8064), .A2(n8053), .A3(n8596), .ZN(n8057) );
  INV_X1 U9723 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9724 ( .A1(n8055), .A2(n8127), .ZN(n8056) );
  NAND2_X1 U9725 ( .A1(n8057), .A2(n8056), .ZN(n8070) );
  NAND3_X1 U9726 ( .A1(n8060), .A2(n8059), .A3(n8058), .ZN(n8062) );
  NAND3_X1 U9727 ( .A1(n8062), .A2(n8127), .A3(n8061), .ZN(n8063) );
  NAND2_X1 U9728 ( .A1(n8064), .A2(n8063), .ZN(n8067) );
  INV_X1 U9729 ( .A(n8065), .ZN(n8066) );
  NAND2_X1 U9730 ( .A1(n8067), .A2(n8066), .ZN(n8069) );
  NAND3_X1 U9731 ( .A1(n8702), .A2(n8165), .A3(n8127), .ZN(n8068) );
  NAND2_X1 U9732 ( .A1(n8072), .A2(n8071), .ZN(n8075) );
  NAND2_X1 U9733 ( .A1(n8078), .A2(n8073), .ZN(n8074) );
  MUX2_X1 U9734 ( .A(n8075), .B(n8074), .S(n8127), .Z(n8076) );
  INV_X1 U9735 ( .A(n8078), .ZN(n8079) );
  MUX2_X1 U9736 ( .A(n8080), .B(n8079), .S(n8128), .Z(n8081) );
  NAND2_X1 U9737 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  OAI211_X1 U9738 ( .C1(n8093), .C2(n8084), .A(n4851), .B(n8094), .ZN(n8086)
         );
  AOI21_X1 U9739 ( .B1(n8086), .B2(n8085), .A(n8528), .ZN(n8089) );
  INV_X1 U9740 ( .A(n8087), .ZN(n8088) );
  NAND2_X1 U9741 ( .A1(n8091), .A2(n8090), .ZN(n8104) );
  NOR2_X1 U9742 ( .A1(n8093), .A2(n8092), .ZN(n8096) );
  OAI21_X1 U9743 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8099) );
  AOI21_X1 U9744 ( .B1(n8099), .B2(n8098), .A(n8097), .ZN(n8102) );
  OAI21_X1 U9745 ( .B1(n8102), .B2(n8512), .A(n8101), .ZN(n8103) );
  MUX2_X2 U9746 ( .A(n8104), .B(n8103), .S(n8128), .Z(n8111) );
  INV_X1 U9747 ( .A(n8499), .ZN(n8501) );
  INV_X1 U9748 ( .A(n8105), .ZN(n8110) );
  INV_X1 U9749 ( .A(n8106), .ZN(n8108) );
  MUX2_X1 U9750 ( .A(n8108), .B(n8107), .S(n8128), .Z(n8109) );
  INV_X1 U9751 ( .A(n8112), .ZN(n8115) );
  AOI211_X1 U9752 ( .C1(n8505), .C2(n8119), .A(n8115), .B(n8121), .ZN(n8118)
         );
  INV_X1 U9753 ( .A(n8119), .ZN(n8124) );
  INV_X1 U9754 ( .A(n8120), .ZN(n8123) );
  INV_X1 U9755 ( .A(n8121), .ZN(n8122) );
  OAI211_X1 U9756 ( .C1(n8124), .C2(n8495), .A(n8123), .B(n8122), .ZN(n8126)
         );
  NAND2_X1 U9757 ( .A1(n8126), .A2(n8125), .ZN(n8129) );
  NAND2_X1 U9758 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  NAND2_X1 U9759 ( .A1(n8131), .A2(n8130), .ZN(n8133) );
  INV_X1 U9760 ( .A(n8134), .ZN(n8136) );
  NAND2_X1 U9761 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  XNOR2_X1 U9762 ( .A(n8141), .B(n8468), .ZN(n8148) );
  NOR3_X1 U9763 ( .A1(n8143), .A2(n8142), .A3(n5002), .ZN(n8146) );
  OAI21_X1 U9764 ( .B1(n8147), .B2(n8144), .A(P2_B_REG_SCAN_IN), .ZN(n8145) );
  INV_X1 U9765 ( .A(n8149), .ZN(n8151) );
  OAI21_X1 U9766 ( .B1(n8151), .B2(n8371), .A(n8150), .ZN(n8235) );
  XNOR2_X1 U9767 ( .A(n8240), .B(n4291), .ZN(n8152) );
  XNOR2_X1 U9768 ( .A(n8152), .B(n8655), .ZN(n8234) );
  XNOR2_X1 U9769 ( .A(n8805), .B(n4291), .ZN(n8278) );
  XNOR2_X1 U9770 ( .A(n8278), .B(n8370), .ZN(n8355) );
  XNOR2_X1 U9771 ( .A(n8799), .B(n4291), .ZN(n8159) );
  XNOR2_X1 U9772 ( .A(n8159), .B(n8647), .ZN(n8280) );
  XNOR2_X1 U9773 ( .A(n8793), .B(n4291), .ZN(n8157) );
  XNOR2_X1 U9774 ( .A(n8157), .B(n8605), .ZN(n8287) );
  INV_X1 U9775 ( .A(n8287), .ZN(n8160) );
  OR2_X1 U9776 ( .A1(n8280), .A2(n8160), .ZN(n8155) );
  INV_X1 U9777 ( .A(n8157), .ZN(n8158) );
  NAND2_X1 U9778 ( .A1(n8159), .A2(n8647), .ZN(n8286) );
  OR2_X1 U9779 ( .A1(n8160), .A2(n8286), .ZN(n8290) );
  INV_X1 U9780 ( .A(n8290), .ZN(n8161) );
  XNOR2_X1 U9781 ( .A(n8702), .B(n4291), .ZN(n8164) );
  XNOR2_X1 U9782 ( .A(n8164), .B(n8620), .ZN(n8333) );
  NAND2_X1 U9783 ( .A1(n8167), .A2(n8166), .ZN(n8250) );
  INV_X1 U9784 ( .A(n8250), .ZN(n8171) );
  XOR2_X1 U9785 ( .A(n4291), .B(n8695), .Z(n8169) );
  INV_X1 U9786 ( .A(n8169), .ZN(n8168) );
  XNOR2_X1 U9787 ( .A(n8168), .B(n8604), .ZN(n8251) );
  INV_X1 U9788 ( .A(n8251), .ZN(n8170) );
  XNOR2_X1 U9789 ( .A(n8784), .B(n4291), .ZN(n8173) );
  XNOR2_X1 U9790 ( .A(n8173), .B(n8590), .ZN(n8311) );
  INV_X1 U9791 ( .A(n8311), .ZN(n8172) );
  NAND2_X1 U9792 ( .A1(n8310), .A2(n8172), .ZN(n8175) );
  NAND2_X1 U9793 ( .A1(n8173), .A2(n8590), .ZN(n8174) );
  NAND2_X1 U9794 ( .A1(n8175), .A2(n8174), .ZN(n8259) );
  XNOR2_X1 U9795 ( .A(n8778), .B(n4291), .ZN(n8176) );
  XNOR2_X1 U9796 ( .A(n8176), .B(n8584), .ZN(n8260) );
  NAND2_X1 U9797 ( .A1(n8259), .A2(n8260), .ZN(n8178) );
  NAND2_X1 U9798 ( .A1(n8176), .A2(n8315), .ZN(n8177) );
  NAND2_X1 U9799 ( .A1(n8178), .A2(n8177), .ZN(n8322) );
  XNOR2_X1 U9800 ( .A(n8184), .B(n8772), .ZN(n8179) );
  NAND2_X1 U9801 ( .A1(n8179), .A2(n8573), .ZN(n8323) );
  NAND2_X1 U9802 ( .A1(n8322), .A2(n8323), .ZN(n8182) );
  INV_X1 U9803 ( .A(n8179), .ZN(n8181) );
  NAND2_X1 U9804 ( .A1(n8181), .A2(n8180), .ZN(n8324) );
  XNOR2_X1 U9805 ( .A(n8766), .B(n4291), .ZN(n8183) );
  XNOR2_X1 U9806 ( .A(n8533), .B(n8184), .ZN(n8185) );
  INV_X1 U9807 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U9808 ( .A1(n8186), .A2(n8549), .ZN(n8187) );
  NAND2_X1 U9809 ( .A1(n8188), .A2(n8301), .ZN(n8266) );
  NAND2_X1 U9810 ( .A1(n8266), .A2(n8267), .ZN(n8189) );
  XNOR2_X1 U9811 ( .A(n8754), .B(n4291), .ZN(n8190) );
  XNOR2_X1 U9812 ( .A(n8190), .B(n8535), .ZN(n8268) );
  NAND2_X1 U9813 ( .A1(n8189), .A2(n8268), .ZN(n8270) );
  XNOR2_X1 U9814 ( .A(n8748), .B(n4291), .ZN(n8343) );
  XNOR2_X1 U9815 ( .A(n8672), .B(n4291), .ZN(n8192) );
  NOR2_X1 U9816 ( .A1(n8192), .A2(n8348), .ZN(n8224) );
  AOI21_X1 U9817 ( .B1(n8348), .B2(n8192), .A(n8224), .ZN(n8193) );
  OAI211_X1 U9818 ( .C1(n8194), .C2(n8193), .A(n8226), .B(n8354), .ZN(n8199)
         );
  INV_X1 U9819 ( .A(n8195), .ZN(n8507) );
  AOI22_X1 U9820 ( .A1(n8523), .A2(n8358), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8196) );
  OAI21_X1 U9821 ( .B1(n8507), .B2(n8339), .A(n8196), .ZN(n8197) );
  AOI21_X1 U9822 ( .B1(n8369), .B2(n8305), .A(n8197), .ZN(n8198) );
  OAI211_X1 U9823 ( .C1(n8200), .C2(n8365), .A(n8199), .B(n8198), .ZN(P2_U3154) );
  AOI21_X1 U9824 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8210) );
  OAI22_X1 U9825 ( .A1(n8365), .A2(n8204), .B1(n4610), .B2(n8360), .ZN(n8205)
         );
  AOI211_X1 U9826 ( .C1(n8358), .C2(n9861), .A(n8206), .B(n8205), .ZN(n8209)
         );
  NAND2_X1 U9827 ( .A1(n8362), .A2(n8207), .ZN(n8208) );
  OAI211_X1 U9828 ( .C1(n8210), .C2(n8352), .A(n8209), .B(n8208), .ZN(P2_U3170) );
  OAI211_X1 U9829 ( .C1(n8213), .C2(n8212), .A(n8211), .B(n8354), .ZN(n8219)
         );
  OAI22_X1 U9830 ( .A1(n8365), .A2(n8215), .B1(n8214), .B2(n8360), .ZN(n8216)
         );
  AOI211_X1 U9831 ( .C1(n8358), .C2(n8380), .A(n8217), .B(n8216), .ZN(n8218)
         );
  OAI211_X1 U9832 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8339), .A(n8219), .B(
        n8218), .ZN(P2_U3158) );
  INV_X1 U9833 ( .A(n8221), .ZN(n8818) );
  OAI222_X1 U9834 ( .A1(n8220), .A2(P1_U3086), .B1(n9478), .B2(n8818), .C1(
        n8223), .C2(n8222), .ZN(P1_U3325) );
  INV_X1 U9835 ( .A(n8224), .ZN(n8225) );
  XNOR2_X1 U9836 ( .A(n8228), .B(n8227), .ZN(n8233) );
  AOI22_X1 U9837 ( .A1(n8514), .A2(n8358), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8230) );
  NAND2_X1 U9838 ( .A1(n8494), .A2(n8362), .ZN(n8229) );
  OAI211_X1 U9839 ( .C1(n8368), .C2(n8360), .A(n8230), .B(n8229), .ZN(n8231)
         );
  AOI21_X1 U9840 ( .B1(n8495), .B2(n8350), .A(n8231), .ZN(n8232) );
  OAI21_X1 U9841 ( .B1(n8233), .B2(n8352), .A(n8232), .ZN(P2_U3160) );
  XOR2_X1 U9842 ( .A(n8235), .B(n8234), .Z(n8242) );
  NAND2_X1 U9843 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8406) );
  OAI21_X1 U9844 ( .B1(n8360), .B2(n8634), .A(n8406), .ZN(n8236) );
  AOI21_X1 U9845 ( .B1(n8358), .B2(n8371), .A(n8236), .ZN(n8237) );
  OAI21_X1 U9846 ( .B1(n8238), .B2(n8339), .A(n8237), .ZN(n8239) );
  AOI21_X1 U9847 ( .B1(n8240), .B2(n8350), .A(n8239), .ZN(n8241) );
  OAI21_X1 U9848 ( .B1(n8242), .B2(n8352), .A(n8241), .ZN(P2_U3155) );
  AOI21_X1 U9849 ( .B1(n8560), .B2(n8243), .A(n4294), .ZN(n8249) );
  AOI22_X1 U9850 ( .A1(n8573), .A2(n8358), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8245) );
  NAND2_X1 U9851 ( .A1(n8362), .A2(n8552), .ZN(n8244) );
  OAI211_X1 U9852 ( .C1(n8246), .C2(n8360), .A(n8245), .B(n8244), .ZN(n8247)
         );
  AOI21_X1 U9853 ( .B1(n8766), .B2(n8350), .A(n8247), .ZN(n8248) );
  OAI21_X1 U9854 ( .B1(n8249), .B2(n8352), .A(n8248), .ZN(P2_U3156) );
  XOR2_X1 U9855 ( .A(n8250), .B(n8251), .Z(n8258) );
  INV_X1 U9856 ( .A(n8252), .ZN(n8593) );
  OAI22_X1 U9857 ( .A1(n8360), .A2(n8590), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8253), .ZN(n8254) );
  AOI21_X1 U9858 ( .B1(n8358), .B2(n8620), .A(n8254), .ZN(n8255) );
  OAI21_X1 U9859 ( .B1(n8593), .B2(n8339), .A(n8255), .ZN(n8256) );
  AOI21_X1 U9860 ( .B1(n8695), .B2(n8350), .A(n8256), .ZN(n8257) );
  OAI21_X1 U9861 ( .B1(n8258), .B2(n8352), .A(n8257), .ZN(P2_U3159) );
  XOR2_X1 U9862 ( .A(n8259), .B(n8260), .Z(n8265) );
  AOI22_X1 U9863 ( .A1(n8573), .A2(n8305), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8262) );
  NAND2_X1 U9864 ( .A1(n8362), .A2(n8577), .ZN(n8261) );
  OAI211_X1 U9865 ( .C1(n8590), .C2(n8316), .A(n8262), .B(n8261), .ZN(n8263)
         );
  AOI21_X1 U9866 ( .B1(n8778), .B2(n8350), .A(n8263), .ZN(n8264) );
  OAI21_X1 U9867 ( .B1(n8265), .B2(n8352), .A(n8264), .ZN(P2_U3163) );
  INV_X1 U9868 ( .A(n8754), .ZN(n8520) );
  INV_X1 U9869 ( .A(n8266), .ZN(n8303) );
  INV_X1 U9870 ( .A(n8267), .ZN(n8269) );
  NOR3_X1 U9871 ( .A1(n8303), .A2(n8269), .A3(n8268), .ZN(n8272) );
  INV_X1 U9872 ( .A(n8270), .ZN(n8271) );
  OAI21_X1 U9873 ( .B1(n8272), .B2(n8271), .A(n8354), .ZN(n8276) );
  AOI22_X1 U9874 ( .A1(n8549), .A2(n8358), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8273) );
  OAI21_X1 U9875 ( .B1(n8504), .B2(n8360), .A(n8273), .ZN(n8274) );
  AOI21_X1 U9876 ( .B1(n8527), .B2(n8362), .A(n8274), .ZN(n8275) );
  OAI211_X1 U9877 ( .C1(n8520), .C2(n8365), .A(n8276), .B(n8275), .ZN(P2_U3165) );
  OAI21_X1 U9878 ( .B1(n8634), .B2(n8278), .A(n8277), .ZN(n8279) );
  NOR2_X1 U9879 ( .A1(n8279), .A2(n8280), .ZN(n8289) );
  AOI21_X1 U9880 ( .B1(n8280), .B2(n8279), .A(n8289), .ZN(n8285) );
  NAND2_X1 U9881 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8441) );
  OAI21_X1 U9882 ( .B1(n8360), .B2(n8635), .A(n8441), .ZN(n8281) );
  AOI21_X1 U9883 ( .B1(n8358), .B2(n8370), .A(n8281), .ZN(n8282) );
  OAI21_X1 U9884 ( .B1(n8640), .B2(n8339), .A(n8282), .ZN(n8283) );
  AOI21_X1 U9885 ( .B1(n8799), .B2(n8350), .A(n8283), .ZN(n8284) );
  OAI21_X1 U9886 ( .B1(n8285), .B2(n8352), .A(n8284), .ZN(P2_U3166) );
  INV_X1 U9887 ( .A(n8793), .ZN(n8299) );
  INV_X1 U9888 ( .A(n8286), .ZN(n8288) );
  NOR3_X1 U9889 ( .A1(n8289), .A2(n8288), .A3(n8287), .ZN(n8292) );
  OAI21_X1 U9890 ( .B1(n8292), .B2(n4370), .A(n8354), .ZN(n8298) );
  INV_X1 U9891 ( .A(n8293), .ZN(n8624) );
  OAI22_X1 U9892 ( .A1(n8360), .A2(n8165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8294), .ZN(n8296) );
  NOR2_X1 U9893 ( .A1(n8316), .A2(n8647), .ZN(n8295) );
  AOI211_X1 U9894 ( .C1(n8624), .C2(n8362), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI211_X1 U9895 ( .C1(n8299), .C2(n8365), .A(n8298), .B(n8297), .ZN(P2_U3168) );
  INV_X1 U9896 ( .A(n8300), .ZN(n8302) );
  NOR3_X1 U9897 ( .A1(n4294), .A2(n8302), .A3(n8301), .ZN(n8304) );
  OAI21_X1 U9898 ( .B1(n8304), .B2(n8303), .A(n8354), .ZN(n8309) );
  AOI22_X1 U9899 ( .A1(n8535), .A2(n8305), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8306) );
  OAI21_X1 U9900 ( .B1(n8328), .B2(n8316), .A(n8306), .ZN(n8307) );
  AOI21_X1 U9901 ( .B1(n8539), .B2(n8362), .A(n8307), .ZN(n8308) );
  OAI211_X1 U9902 ( .C1(n8533), .C2(n8365), .A(n8309), .B(n8308), .ZN(P2_U3169) );
  XNOR2_X1 U9903 ( .A(n8312), .B(n8311), .ZN(n8313) );
  NAND2_X1 U9904 ( .A1(n8313), .A2(n8354), .ZN(n8320) );
  INV_X1 U9905 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8314) );
  OAI22_X1 U9906 ( .A1(n8315), .A2(n8360), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8314), .ZN(n8318) );
  NOR2_X1 U9907 ( .A1(n8316), .A2(n8336), .ZN(n8317) );
  AOI211_X1 U9908 ( .C1(n8586), .C2(n8362), .A(n8318), .B(n8317), .ZN(n8319)
         );
  OAI211_X1 U9909 ( .C1(n8321), .C2(n8365), .A(n8320), .B(n8319), .ZN(P2_U3173) );
  NAND2_X1 U9910 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  XNOR2_X1 U9911 ( .A(n8322), .B(n8325), .ZN(n8331) );
  AOI22_X1 U9912 ( .A1(n8584), .A2(n8358), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8327) );
  NAND2_X1 U9913 ( .A1(n8362), .A2(n8563), .ZN(n8326) );
  OAI211_X1 U9914 ( .C1(n8328), .C2(n8360), .A(n8327), .B(n8326), .ZN(n8329)
         );
  AOI21_X1 U9915 ( .B1(n8772), .B2(n8350), .A(n8329), .ZN(n8330) );
  OAI21_X1 U9916 ( .B1(n8331), .B2(n8352), .A(n8330), .ZN(P2_U3175) );
  XOR2_X1 U9917 ( .A(n8332), .B(n8333), .Z(n8342) );
  INV_X1 U9918 ( .A(n8334), .ZN(n8608) );
  OAI22_X1 U9919 ( .A1(n8360), .A2(n8336), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8335), .ZN(n8337) );
  AOI21_X1 U9920 ( .B1(n8358), .B2(n8605), .A(n8337), .ZN(n8338) );
  OAI21_X1 U9921 ( .B1(n8608), .B2(n8339), .A(n8338), .ZN(n8340) );
  AOI21_X1 U9922 ( .B1(n8702), .B2(n8350), .A(n8340), .ZN(n8341) );
  OAI21_X1 U9923 ( .B1(n8342), .B2(n8352), .A(n8341), .ZN(P2_U3178) );
  XNOR2_X1 U9924 ( .A(n8343), .B(n8504), .ZN(n8344) );
  XNOR2_X1 U9925 ( .A(n8345), .B(n8344), .ZN(n8353) );
  AOI22_X1 U9926 ( .A1(n8535), .A2(n8358), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8347) );
  NAND2_X1 U9927 ( .A1(n8517), .A2(n8362), .ZN(n8346) );
  OAI211_X1 U9928 ( .C1(n8348), .C2(n8360), .A(n8347), .B(n8346), .ZN(n8349)
         );
  AOI21_X1 U9929 ( .B1(n8748), .B2(n8350), .A(n8349), .ZN(n8351) );
  OAI21_X1 U9930 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(P2_U3180) );
  INV_X1 U9931 ( .A(n8805), .ZN(n8366) );
  OAI211_X1 U9932 ( .C1(n8356), .C2(n8355), .A(n8277), .B(n8354), .ZN(n8364)
         );
  INV_X1 U9933 ( .A(n8357), .ZN(n8657) );
  NAND2_X1 U9934 ( .A1(n8358), .A2(n8655), .ZN(n8359) );
  NAND2_X1 U9935 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8423) );
  OAI211_X1 U9936 ( .C1(n8647), .C2(n8360), .A(n8359), .B(n8423), .ZN(n8361)
         );
  AOI21_X1 U9937 ( .B1(n8657), .B2(n8362), .A(n8361), .ZN(n8363) );
  OAI211_X1 U9938 ( .C1(n8366), .C2(n8365), .A(n8364), .B(n8363), .ZN(P2_U3181) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8367), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U9940 ( .A(n8368), .ZN(n8492) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8492), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8369), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8514), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9944 ( .A(n8523), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8381), .Z(
        P2_U3517) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8535), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8549), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9947 ( .A(n8560), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8381), .Z(
        P2_U3514) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8573), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8584), .S(P2_U3893), .Z(
        P2_U3512) );
  INV_X1 U9950 ( .A(n8590), .ZN(n8574) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8574), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9952 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8604), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9953 ( .A(n8620), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8381), .Z(
        P2_U3509) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8621), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8370), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9957 ( .A(n8655), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8381), .Z(
        P2_U3505) );
  MUX2_X1 U9958 ( .A(n8371), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8381), .Z(
        P2_U3504) );
  MUX2_X1 U9959 ( .A(n8372), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8381), .Z(
        P2_U3503) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8373), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9961 ( .A(n8374), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8381), .Z(
        P2_U3501) );
  MUX2_X1 U9962 ( .A(n8375), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8381), .Z(
        P2_U3500) );
  MUX2_X1 U9963 ( .A(n8376), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8381), .Z(
        P2_U3499) );
  MUX2_X1 U9964 ( .A(n8377), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8381), .Z(
        P2_U3498) );
  MUX2_X1 U9965 ( .A(n8378), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8381), .Z(
        P2_U3497) );
  MUX2_X1 U9966 ( .A(n8379), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8381), .Z(
        P2_U3496) );
  MUX2_X1 U9967 ( .A(n9861), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8381), .Z(
        P2_U3494) );
  MUX2_X1 U9968 ( .A(n8380), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8381), .Z(
        P2_U3493) );
  MUX2_X1 U9969 ( .A(n7101), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8381), .Z(
        P2_U3492) );
  MUX2_X1 U9970 ( .A(n7098), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8381), .Z(
        P2_U3491) );
  AOI21_X1 U9971 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8398) );
  OAI21_X1 U9972 ( .B1(n8387), .B2(n8386), .A(n8385), .ZN(n8396) );
  AOI21_X1 U9973 ( .B1(n8389), .B2(n10050), .A(n8388), .ZN(n8391) );
  OAI21_X1 U9974 ( .B1(n9852), .B2(n8391), .A(n8390), .ZN(n8392) );
  AOI21_X1 U9975 ( .B1(n9797), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8392), .ZN(
        n8393) );
  OAI21_X1 U9976 ( .B1(n8394), .B2(n9835), .A(n8393), .ZN(n8395) );
  AOI21_X1 U9977 ( .B1(n8396), .B2(n9843), .A(n8395), .ZN(n8397) );
  OAI21_X1 U9978 ( .B1(n8398), .B2(n9848), .A(n8397), .ZN(P2_U3195) );
  AOI21_X1 U9979 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8416) );
  OAI21_X1 U9980 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8414) );
  INV_X1 U9981 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8405) );
  OR2_X1 U9982 ( .A1(n9832), .A2(n8405), .ZN(n8407) );
  OAI211_X1 U9983 ( .C1(n9835), .C2(n8408), .A(n8407), .B(n8406), .ZN(n8413)
         );
  AOI21_X1 U9984 ( .B1(n4334), .B2(n8410), .A(n8409), .ZN(n8411) );
  NOR2_X1 U9985 ( .A1(n8411), .A2(n9852), .ZN(n8412) );
  AOI211_X1 U9986 ( .C1(n9843), .C2(n8414), .A(n8413), .B(n8412), .ZN(n8415)
         );
  OAI21_X1 U9987 ( .B1(n8416), .B2(n9848), .A(n8415), .ZN(P2_U3196) );
  AOI21_X1 U9988 ( .B1(n8418), .B2(n8713), .A(n8417), .ZN(n8433) );
  OAI21_X1 U9989 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(n8431) );
  INV_X1 U9990 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8422) );
  OR2_X1 U9991 ( .A1(n9832), .A2(n8422), .ZN(n8424) );
  OAI211_X1 U9992 ( .C1(n9835), .C2(n8425), .A(n8424), .B(n8423), .ZN(n8430)
         );
  AOI21_X1 U9993 ( .B1(n8656), .B2(n8427), .A(n8426), .ZN(n8428) );
  NOR2_X1 U9994 ( .A1(n8428), .A2(n9848), .ZN(n8429) );
  AOI211_X1 U9995 ( .C1(n9843), .C2(n8431), .A(n8430), .B(n8429), .ZN(n8432)
         );
  OAI21_X1 U9996 ( .B1(n8433), .B2(n9852), .A(n8432), .ZN(P2_U3197) );
  AOI21_X1 U9997 ( .B1(n8436), .B2(n8435), .A(n8434), .ZN(n8451) );
  OAI21_X1 U9998 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8449) );
  INV_X1 U9999 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8440) );
  OR2_X1 U10000 ( .A1(n9832), .A2(n8440), .ZN(n8442) );
  OAI211_X1 U10001 ( .C1(n9835), .C2(n8443), .A(n8442), .B(n8441), .ZN(n8448)
         );
  AOI21_X1 U10002 ( .B1(n4335), .B2(n8445), .A(n8444), .ZN(n8446) );
  NOR2_X1 U10003 ( .A1(n8446), .A2(n9852), .ZN(n8447) );
  AOI211_X1 U10004 ( .C1(n9843), .C2(n8449), .A(n8448), .B(n8447), .ZN(n8450)
         );
  OAI21_X1 U10005 ( .B1(n8451), .B2(n9848), .A(n8450), .ZN(P2_U3198) );
  MUX2_X1 U10006 ( .A(n8594), .B(P2_REG2_REG_19__SCAN_IN), .S(n8468), .Z(n8459) );
  INV_X1 U10007 ( .A(n8454), .ZN(n8455) );
  XNOR2_X1 U10008 ( .A(n8468), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8458) );
  MUX2_X1 U10009 ( .A(n8459), .B(n8458), .S(n4287), .Z(n8464) );
  OAI21_X1 U10010 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n8463) );
  XOR2_X1 U10011 ( .A(n8464), .B(n8463), .Z(n8465) );
  NAND2_X1 U10012 ( .A1(n9797), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10013 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8466) );
  OAI211_X1 U10014 ( .C1(n9835), .C2(n8468), .A(n8467), .B(n8466), .ZN(n8469)
         );
  OAI21_X1 U10015 ( .B1(n8471), .B2(n9848), .A(n8470), .ZN(P2_U3201) );
  NAND2_X1 U10016 ( .A1(n8727), .A2(n8658), .ZN(n8476) );
  INV_X1 U10017 ( .A(n8472), .ZN(n8473) );
  NOR2_X1 U10018 ( .A1(n8474), .A2(n8473), .ZN(n8728) );
  NOR2_X1 U10019 ( .A1(n8475), .A2(n8607), .ZN(n8484) );
  AOI21_X1 U10020 ( .B1(n8728), .B2(n9878), .A(n8484), .ZN(n8479) );
  OAI211_X1 U10021 ( .C1(n9878), .C2(n8477), .A(n8476), .B(n8479), .ZN(
        P2_U3202) );
  NAND2_X1 U10022 ( .A1(n9881), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8478) );
  OAI211_X1 U10023 ( .C1(n8667), .C2(n8481), .A(n8479), .B(n8478), .ZN(
        P2_U3203) );
  INV_X1 U10024 ( .A(n8480), .ZN(n8488) );
  NOR2_X1 U10025 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  AOI211_X1 U10026 ( .C1(n9881), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8484), .B(
        n8483), .ZN(n8485) );
  OAI211_X1 U10027 ( .C1(n8488), .C2(n8487), .A(n8486), .B(n8485), .ZN(
        P2_U3204) );
  XOR2_X1 U10028 ( .A(n8491), .B(n8489), .Z(n8737) );
  INV_X1 U10029 ( .A(n8737), .ZN(n8498) );
  INV_X1 U10030 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8493) );
  MUX2_X1 U10031 ( .A(n8493), .B(n8735), .S(n9878), .Z(n8497) );
  AOI22_X1 U10032 ( .A1(n8495), .A2(n8658), .B1(n9877), .B2(n8494), .ZN(n8496)
         );
  OAI211_X1 U10033 ( .C1(n8498), .C2(n8661), .A(n8497), .B(n8496), .ZN(
        P2_U3205) );
  XNOR2_X1 U10034 ( .A(n8500), .B(n8499), .ZN(n8745) );
  XNOR2_X1 U10035 ( .A(n8502), .B(n8501), .ZN(n8503) );
  NAND2_X1 U10036 ( .A1(n8671), .A2(n9878), .ZN(n8510) );
  INV_X1 U10037 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8506) );
  OAI22_X1 U10038 ( .A1(n8507), .A2(n8607), .B1(n9878), .B2(n8506), .ZN(n8508)
         );
  AOI21_X1 U10039 ( .B1(n8672), .B2(n8658), .A(n8508), .ZN(n8509) );
  OAI211_X1 U10040 ( .C1(n8745), .C2(n8661), .A(n8510), .B(n8509), .ZN(
        P2_U3206) );
  XNOR2_X1 U10041 ( .A(n8511), .B(n8512), .ZN(n8751) );
  INV_X1 U10042 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8516) );
  XNOR2_X1 U10043 ( .A(n8513), .B(n8512), .ZN(n8515) );
  AOI222_X1 U10044 ( .A1(n9866), .A2(n8515), .B1(n8535), .B2(n9862), .C1(n8514), .C2(n9860), .ZN(n8746) );
  MUX2_X1 U10045 ( .A(n8516), .B(n8746), .S(n9878), .Z(n8519) );
  AOI22_X1 U10046 ( .A1(n8748), .A2(n8658), .B1(n9877), .B2(n8517), .ZN(n8518)
         );
  OAI211_X1 U10047 ( .C1(n8751), .C2(n8661), .A(n8519), .B(n8518), .ZN(
        P2_U3207) );
  NOR2_X1 U10048 ( .A1(n8520), .A2(n8532), .ZN(n8526) );
  OAI21_X1 U10049 ( .B1(n8522), .B2(n8528), .A(n8521), .ZN(n8524) );
  AOI222_X1 U10050 ( .A1(n9866), .A2(n8524), .B1(n8523), .B2(n9860), .C1(n8549), .C2(n9862), .ZN(n8752) );
  INV_X1 U10051 ( .A(n8752), .ZN(n8525) );
  AOI211_X1 U10052 ( .C1(n9877), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8531)
         );
  XNOR2_X1 U10053 ( .A(n8529), .B(n8528), .ZN(n8755) );
  AOI22_X1 U10054 ( .A1(n8755), .A2(n8613), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9881), .ZN(n8530) );
  OAI21_X1 U10055 ( .B1(n8531), .B2(n9881), .A(n8530), .ZN(P2_U3208) );
  NOR2_X1 U10056 ( .A1(n8533), .A2(n8532), .ZN(n8538) );
  XNOR2_X1 U10057 ( .A(n8534), .B(n8542), .ZN(n8536) );
  AOI222_X1 U10058 ( .A1(n9866), .A2(n8536), .B1(n8535), .B2(n9860), .C1(n8560), .C2(n9862), .ZN(n8758) );
  INV_X1 U10059 ( .A(n8758), .ZN(n8537) );
  AOI211_X1 U10060 ( .C1(n9877), .C2(n8539), .A(n8538), .B(n8537), .ZN(n8545)
         );
  NOR2_X1 U10061 ( .A1(n8541), .A2(n8540), .ZN(n8543) );
  XNOR2_X1 U10062 ( .A(n8543), .B(n8542), .ZN(n8761) );
  AOI22_X1 U10063 ( .A1(n8761), .A2(n8613), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9881), .ZN(n8544) );
  OAI21_X1 U10064 ( .B1(n8545), .B2(n9881), .A(n8544), .ZN(P2_U3209) );
  XOR2_X1 U10065 ( .A(n8547), .B(n8546), .Z(n8769) );
  INV_X1 U10066 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U10067 ( .A(n8548), .B(n8547), .ZN(n8550) );
  AOI222_X1 U10068 ( .A1(n9866), .A2(n8550), .B1(n8549), .B2(n9860), .C1(n8573), .C2(n9862), .ZN(n8764) );
  MUX2_X1 U10069 ( .A(n8551), .B(n8764), .S(n9878), .Z(n8554) );
  AOI22_X1 U10070 ( .A1(n8766), .A2(n8658), .B1(n9877), .B2(n8552), .ZN(n8553)
         );
  OAI211_X1 U10071 ( .C1(n8769), .C2(n8661), .A(n8554), .B(n8553), .ZN(
        P2_U3210) );
  XOR2_X1 U10072 ( .A(n8555), .B(n8556), .Z(n8773) );
  INV_X1 U10073 ( .A(n8773), .ZN(n8566) );
  INV_X1 U10074 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8562) );
  OR3_X1 U10075 ( .A1(n8568), .A2(n8557), .A3(n8556), .ZN(n8558) );
  NAND2_X1 U10076 ( .A1(n8559), .A2(n8558), .ZN(n8561) );
  AOI222_X1 U10077 ( .A1(n9866), .A2(n8561), .B1(n8584), .B2(n9862), .C1(n8560), .C2(n9860), .ZN(n8770) );
  MUX2_X1 U10078 ( .A(n8562), .B(n8770), .S(n9878), .Z(n8565) );
  AOI22_X1 U10079 ( .A1(n8772), .A2(n8658), .B1(n9877), .B2(n8563), .ZN(n8564)
         );
  OAI211_X1 U10080 ( .C1(n8566), .C2(n8661), .A(n8565), .B(n8564), .ZN(
        P2_U3211) );
  XOR2_X1 U10081 ( .A(n8567), .B(n8570), .Z(n8779) );
  INV_X1 U10082 ( .A(n8779), .ZN(n8580) );
  INV_X1 U10083 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8576) );
  INV_X1 U10084 ( .A(n8568), .ZN(n8572) );
  NAND3_X1 U10085 ( .A1(n8581), .A2(n8570), .A3(n8569), .ZN(n8571) );
  NAND2_X1 U10086 ( .A1(n8572), .A2(n8571), .ZN(n8575) );
  AOI222_X1 U10087 ( .A1(n9866), .A2(n8575), .B1(n8574), .B2(n9862), .C1(n8573), .C2(n9860), .ZN(n8776) );
  MUX2_X1 U10088 ( .A(n8576), .B(n8776), .S(n9878), .Z(n8579) );
  AOI22_X1 U10089 ( .A1(n8778), .A2(n8658), .B1(n9877), .B2(n8577), .ZN(n8578)
         );
  OAI211_X1 U10090 ( .C1(n8580), .C2(n8661), .A(n8579), .B(n8578), .ZN(
        P2_U3212) );
  XNOR2_X1 U10091 ( .A(n4365), .B(n8582), .ZN(n8788) );
  OAI21_X1 U10092 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8585) );
  AOI222_X1 U10093 ( .A1(n9866), .A2(n8585), .B1(n8584), .B2(n9860), .C1(n8604), .C2(n9862), .ZN(n8782) );
  MUX2_X1 U10094 ( .A(n10123), .B(n8782), .S(n9878), .Z(n8588) );
  AOI22_X1 U10095 ( .A1(n8784), .A2(n8658), .B1(n9877), .B2(n8586), .ZN(n8587)
         );
  OAI211_X1 U10096 ( .C1(n8788), .C2(n8661), .A(n8588), .B(n8587), .ZN(
        P2_U3213) );
  XNOR2_X1 U10097 ( .A(n8589), .B(n8596), .ZN(n8592) );
  OAI22_X1 U10098 ( .A1(n8590), .A2(n8646), .B1(n8165), .B2(n8633), .ZN(n8591)
         );
  AOI21_X1 U10099 ( .B1(n8592), .B2(n9866), .A(n8591), .ZN(n8701) );
  OAI22_X1 U10100 ( .A1(n9878), .A2(n8594), .B1(n8593), .B2(n8607), .ZN(n8595)
         );
  AOI21_X1 U10101 ( .B1(n8695), .B2(n8658), .A(n8595), .ZN(n8600) );
  INV_X1 U10102 ( .A(n8697), .ZN(n8598) );
  OR2_X1 U10103 ( .A1(n8597), .A2(n8596), .ZN(n8694) );
  NAND3_X1 U10104 ( .A1(n8598), .A2(n8613), .A3(n8694), .ZN(n8599) );
  OAI211_X1 U10105 ( .C1(n8701), .C2(n9881), .A(n8600), .B(n8599), .ZN(
        P2_U3214) );
  NAND2_X1 U10106 ( .A1(n8637), .A2(n8601), .ZN(n8619) );
  NAND2_X1 U10107 ( .A1(n8619), .A2(n8618), .ZN(n8617) );
  NAND2_X1 U10108 ( .A1(n8617), .A2(n8602), .ZN(n8603) );
  XOR2_X1 U10109 ( .A(n8611), .B(n8603), .Z(n8606) );
  AOI222_X1 U10110 ( .A1(n9866), .A2(n8606), .B1(n8605), .B2(n9862), .C1(n8604), .C2(n9860), .ZN(n8706) );
  OAI22_X1 U10111 ( .A1(n9878), .A2(n8609), .B1(n8608), .B2(n8607), .ZN(n8610)
         );
  AOI21_X1 U10112 ( .B1(n8702), .B2(n8658), .A(n8610), .ZN(n8615) );
  NAND2_X1 U10113 ( .A1(n8612), .A2(n8611), .ZN(n8703) );
  NAND3_X1 U10114 ( .A1(n8704), .A2(n8703), .A3(n8613), .ZN(n8614) );
  OAI211_X1 U10115 ( .C1(n8706), .C2(n9881), .A(n8615), .B(n8614), .ZN(
        P2_U3215) );
  XNOR2_X1 U10116 ( .A(n8616), .B(n8618), .ZN(n8794) );
  INV_X1 U10117 ( .A(n8794), .ZN(n8627) );
  OAI211_X1 U10118 ( .C1(n8619), .C2(n8618), .A(n8617), .B(n9866), .ZN(n8623)
         );
  AOI22_X1 U10119 ( .A1(n8621), .A2(n9862), .B1(n9860), .B2(n8620), .ZN(n8622)
         );
  AND2_X1 U10120 ( .A1(n8623), .A2(n8622), .ZN(n8791) );
  MUX2_X1 U10121 ( .A(n9847), .B(n8791), .S(n9878), .Z(n8626) );
  AOI22_X1 U10122 ( .A1(n8793), .A2(n8658), .B1(n9877), .B2(n8624), .ZN(n8625)
         );
  OAI211_X1 U10123 ( .C1(n8627), .C2(n8661), .A(n8626), .B(n8625), .ZN(
        P2_U3216) );
  XOR2_X1 U10124 ( .A(n8630), .B(n8628), .Z(n8800) );
  INV_X1 U10125 ( .A(n8800), .ZN(n8644) );
  INV_X1 U10126 ( .A(n8629), .ZN(n8632) );
  INV_X1 U10127 ( .A(n8630), .ZN(n8631) );
  AOI21_X1 U10128 ( .B1(n8632), .B2(n8631), .A(n8650), .ZN(n8638) );
  OAI22_X1 U10129 ( .A1(n8635), .A2(n8646), .B1(n8634), .B2(n8633), .ZN(n8636)
         );
  AOI21_X1 U10130 ( .B1(n8638), .B2(n8637), .A(n8636), .ZN(n8797) );
  MUX2_X1 U10131 ( .A(n8639), .B(n8797), .S(n9878), .Z(n8643) );
  INV_X1 U10132 ( .A(n8640), .ZN(n8641) );
  AOI22_X1 U10133 ( .A1(n8799), .A2(n8658), .B1(n9877), .B2(n8641), .ZN(n8642)
         );
  OAI211_X1 U10134 ( .C1(n8644), .C2(n8661), .A(n8643), .B(n8642), .ZN(
        P2_U3217) );
  XOR2_X1 U10135 ( .A(n8652), .B(n8645), .Z(n8808) );
  INV_X1 U10136 ( .A(n8808), .ZN(n8662) );
  NOR2_X1 U10137 ( .A1(n8647), .A2(n8646), .ZN(n8654) );
  INV_X1 U10138 ( .A(n8648), .ZN(n8649) );
  AOI211_X1 U10139 ( .C1(n8652), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8653)
         );
  AOI211_X1 U10140 ( .C1(n9862), .C2(n8655), .A(n8654), .B(n8653), .ZN(n8803)
         );
  MUX2_X1 U10141 ( .A(n8656), .B(n8803), .S(n9878), .Z(n8660) );
  AOI22_X1 U10142 ( .A1(n8805), .A2(n8658), .B1(n9877), .B2(n8657), .ZN(n8659)
         );
  OAI211_X1 U10143 ( .C1(n8662), .C2(n8661), .A(n8660), .B(n8659), .ZN(
        P2_U3218) );
  NAND2_X1 U10144 ( .A1(n8727), .A2(n8714), .ZN(n8663) );
  NAND2_X1 U10145 ( .A1(n8728), .A2(n9954), .ZN(n8665) );
  OAI211_X1 U10146 ( .C1(n9954), .C2(n8664), .A(n8663), .B(n8665), .ZN(
        P2_U3490) );
  NAND2_X1 U10147 ( .A1(n5718), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8666) );
  OAI211_X1 U10148 ( .C1(n8667), .C2(n8670), .A(n8666), .B(n8665), .ZN(
        P2_U3489) );
  MUX2_X1 U10149 ( .A(n10097), .B(n8735), .S(n9954), .Z(n8669) );
  NAND2_X1 U10150 ( .A1(n8737), .A2(n8715), .ZN(n8668) );
  OAI211_X1 U10151 ( .C1(n8741), .C2(n8670), .A(n8669), .B(n8668), .ZN(
        P2_U3487) );
  AOI21_X1 U10152 ( .B1(n9920), .B2(n8672), .A(n8671), .ZN(n8742) );
  MUX2_X1 U10153 ( .A(n10055), .B(n8742), .S(n9954), .Z(n8673) );
  OAI21_X1 U10154 ( .B1(n8745), .B2(n8693), .A(n8673), .ZN(P2_U3486) );
  MUX2_X1 U10155 ( .A(n8674), .B(n8746), .S(n9954), .Z(n8676) );
  NAND2_X1 U10156 ( .A1(n8748), .A2(n8714), .ZN(n8675) );
  OAI211_X1 U10157 ( .C1(n8693), .C2(n8751), .A(n8676), .B(n8675), .ZN(
        P2_U3485) );
  MUX2_X1 U10158 ( .A(n10029), .B(n8752), .S(n9954), .Z(n8678) );
  AOI22_X1 U10159 ( .A1(n8755), .A2(n8715), .B1(n8714), .B2(n8754), .ZN(n8677)
         );
  NAND2_X1 U10160 ( .A1(n8678), .A2(n8677), .ZN(P2_U3484) );
  MUX2_X1 U10161 ( .A(n8679), .B(n8758), .S(n9954), .Z(n8681) );
  AOI22_X1 U10162 ( .A1(n8761), .A2(n8715), .B1(n8714), .B2(n8760), .ZN(n8680)
         );
  NAND2_X1 U10163 ( .A1(n8681), .A2(n8680), .ZN(P2_U3483) );
  MUX2_X1 U10164 ( .A(n10120), .B(n8764), .S(n9954), .Z(n8683) );
  NAND2_X1 U10165 ( .A1(n8766), .A2(n8714), .ZN(n8682) );
  OAI211_X1 U10166 ( .C1(n8769), .C2(n8693), .A(n8683), .B(n8682), .ZN(
        P2_U3482) );
  INV_X1 U10167 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8684) );
  MUX2_X1 U10168 ( .A(n8684), .B(n8770), .S(n9954), .Z(n8686) );
  AOI22_X1 U10169 ( .A1(n8773), .A2(n8715), .B1(n8714), .B2(n8772), .ZN(n8685)
         );
  NAND2_X1 U10170 ( .A1(n8686), .A2(n8685), .ZN(P2_U3481) );
  INV_X1 U10171 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8687) );
  MUX2_X1 U10172 ( .A(n8687), .B(n8776), .S(n9954), .Z(n8689) );
  AOI22_X1 U10173 ( .A1(n8779), .A2(n8715), .B1(n8714), .B2(n8778), .ZN(n8688)
         );
  NAND2_X1 U10174 ( .A1(n8689), .A2(n8688), .ZN(P2_U3480) );
  INV_X1 U10175 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8690) );
  MUX2_X1 U10176 ( .A(n8690), .B(n8782), .S(n9954), .Z(n8692) );
  NAND2_X1 U10177 ( .A1(n8784), .A2(n8714), .ZN(n8691) );
  OAI211_X1 U10178 ( .C1(n8788), .C2(n8693), .A(n8692), .B(n8691), .ZN(
        P2_U3479) );
  NAND2_X1 U10179 ( .A1(n8694), .A2(n9933), .ZN(n8698) );
  INV_X1 U10180 ( .A(n8695), .ZN(n8696) );
  OAI22_X1 U10181 ( .A1(n8698), .A2(n8697), .B1(n8696), .B2(n9928), .ZN(n8699)
         );
  INV_X1 U10182 ( .A(n8699), .ZN(n8700) );
  NAND2_X1 U10183 ( .A1(n8701), .A2(n8700), .ZN(n8789) );
  MUX2_X1 U10184 ( .A(n8789), .B(P2_REG1_REG_19__SCAN_IN), .S(n5718), .Z(
        P2_U3478) );
  INV_X1 U10185 ( .A(n8702), .ZN(n8707) );
  NAND3_X1 U10186 ( .A1(n8704), .A2(n8703), .A3(n9933), .ZN(n8705) );
  OAI211_X1 U10187 ( .C1(n8707), .C2(n9928), .A(n8706), .B(n8705), .ZN(n8790)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8790), .S(n9954), .Z(
        P2_U3477) );
  MUX2_X1 U10189 ( .A(n9839), .B(n8791), .S(n9954), .Z(n8709) );
  AOI22_X1 U10190 ( .A1(n8794), .A2(n8715), .B1(n8714), .B2(n8793), .ZN(n8708)
         );
  NAND2_X1 U10191 ( .A1(n8709), .A2(n8708), .ZN(P2_U3476) );
  MUX2_X1 U10192 ( .A(n8710), .B(n8797), .S(n9954), .Z(n8712) );
  AOI22_X1 U10193 ( .A1(n8800), .A2(n8715), .B1(n8714), .B2(n8799), .ZN(n8711)
         );
  NAND2_X1 U10194 ( .A1(n8712), .A2(n8711), .ZN(P2_U3475) );
  MUX2_X1 U10195 ( .A(n8713), .B(n8803), .S(n9954), .Z(n8717) );
  AOI22_X1 U10196 ( .A1(n8808), .A2(n8715), .B1(n8714), .B2(n8805), .ZN(n8716)
         );
  NAND2_X1 U10197 ( .A1(n8717), .A2(n8716), .ZN(P2_U3474) );
  NAND3_X1 U10198 ( .A1(n7581), .A2(n9933), .A3(n8718), .ZN(n8719) );
  OAI211_X1 U10199 ( .C1(n8721), .C2(n9928), .A(n8720), .B(n8719), .ZN(n8811)
         );
  MUX2_X1 U10200 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8811), .S(n9954), .Z(
        P2_U3473) );
  INV_X1 U10201 ( .A(n8722), .ZN(n8725) );
  OAI21_X1 U10202 ( .B1(n9866), .B2(n9933), .A(n8723), .ZN(n8724) );
  OAI211_X1 U10203 ( .C1(n9928), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8812)
         );
  MUX2_X1 U10204 ( .A(n8812), .B(P2_REG1_REG_0__SCAN_IN), .S(n5718), .Z(
        P2_U3459) );
  INV_X1 U10205 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U10206 ( .A1(n8727), .A2(n8806), .ZN(n8729) );
  NAND2_X1 U10207 ( .A1(n8728), .A2(n9934), .ZN(n8732) );
  OAI211_X1 U10208 ( .C1(n8730), .C2(n9934), .A(n8729), .B(n8732), .ZN(
        P2_U3458) );
  INV_X1 U10209 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10210 ( .A1(n8731), .A2(n8806), .ZN(n8733) );
  OAI211_X1 U10211 ( .C1(n8734), .C2(n9934), .A(n8733), .B(n8732), .ZN(
        P2_U3457) );
  INV_X1 U10212 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8736) );
  MUX2_X1 U10213 ( .A(n8736), .B(n8735), .S(n9934), .Z(n8739) );
  NAND2_X1 U10214 ( .A1(n8737), .A2(n8807), .ZN(n8738) );
  OAI211_X1 U10215 ( .C1(n8741), .C2(n8740), .A(n8739), .B(n8738), .ZN(
        P2_U3455) );
  INV_X1 U10216 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8743) );
  MUX2_X1 U10217 ( .A(n8743), .B(n8742), .S(n9934), .Z(n8744) );
  OAI21_X1 U10218 ( .B1(n8745), .B2(n8787), .A(n8744), .ZN(P2_U3454) );
  INV_X1 U10219 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8747) );
  MUX2_X1 U10220 ( .A(n8747), .B(n8746), .S(n9934), .Z(n8750) );
  NAND2_X1 U10221 ( .A1(n8748), .A2(n8806), .ZN(n8749) );
  OAI211_X1 U10222 ( .C1(n8751), .C2(n8787), .A(n8750), .B(n8749), .ZN(
        P2_U3453) );
  INV_X1 U10223 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8753) );
  MUX2_X1 U10224 ( .A(n8753), .B(n8752), .S(n9934), .Z(n8757) );
  AOI22_X1 U10225 ( .A1(n8755), .A2(n8807), .B1(n8806), .B2(n8754), .ZN(n8756)
         );
  NAND2_X1 U10226 ( .A1(n8757), .A2(n8756), .ZN(P2_U3452) );
  INV_X1 U10227 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8759) );
  MUX2_X1 U10228 ( .A(n8759), .B(n8758), .S(n9934), .Z(n8763) );
  AOI22_X1 U10229 ( .A1(n8761), .A2(n8807), .B1(n8806), .B2(n8760), .ZN(n8762)
         );
  NAND2_X1 U10230 ( .A1(n8763), .A2(n8762), .ZN(P2_U3451) );
  INV_X1 U10231 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8765) );
  MUX2_X1 U10232 ( .A(n8765), .B(n8764), .S(n9934), .Z(n8768) );
  NAND2_X1 U10233 ( .A1(n8766), .A2(n8806), .ZN(n8767) );
  OAI211_X1 U10234 ( .C1(n8769), .C2(n8787), .A(n8768), .B(n8767), .ZN(
        P2_U3450) );
  INV_X1 U10235 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8771) );
  MUX2_X1 U10236 ( .A(n8771), .B(n8770), .S(n9934), .Z(n8775) );
  AOI22_X1 U10237 ( .A1(n8773), .A2(n8807), .B1(n8806), .B2(n8772), .ZN(n8774)
         );
  NAND2_X1 U10238 ( .A1(n8775), .A2(n8774), .ZN(P2_U3449) );
  INV_X1 U10239 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8777) );
  MUX2_X1 U10240 ( .A(n8777), .B(n8776), .S(n9934), .Z(n8781) );
  AOI22_X1 U10241 ( .A1(n8779), .A2(n8807), .B1(n8806), .B2(n8778), .ZN(n8780)
         );
  NAND2_X1 U10242 ( .A1(n8781), .A2(n8780), .ZN(P2_U3448) );
  MUX2_X1 U10243 ( .A(n8783), .B(n8782), .S(n9934), .Z(n8786) );
  NAND2_X1 U10244 ( .A1(n8784), .A2(n8806), .ZN(n8785) );
  OAI211_X1 U10245 ( .C1(n8788), .C2(n8787), .A(n8786), .B(n8785), .ZN(
        P2_U3447) );
  MUX2_X1 U10246 ( .A(n8789), .B(P2_REG0_REG_19__SCAN_IN), .S(n9936), .Z(
        P2_U3446) );
  MUX2_X1 U10247 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8790), .S(n9934), .Z(
        P2_U3444) );
  INV_X1 U10248 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8792) );
  MUX2_X1 U10249 ( .A(n8792), .B(n8791), .S(n9934), .Z(n8796) );
  AOI22_X1 U10250 ( .A1(n8794), .A2(n8807), .B1(n8806), .B2(n8793), .ZN(n8795)
         );
  NAND2_X1 U10251 ( .A1(n8796), .A2(n8795), .ZN(P2_U3441) );
  INV_X1 U10252 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8798) );
  MUX2_X1 U10253 ( .A(n8798), .B(n8797), .S(n9934), .Z(n8802) );
  AOI22_X1 U10254 ( .A1(n8800), .A2(n8807), .B1(n8806), .B2(n8799), .ZN(n8801)
         );
  NAND2_X1 U10255 ( .A1(n8802), .A2(n8801), .ZN(P2_U3438) );
  INV_X1 U10256 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8804) );
  MUX2_X1 U10257 ( .A(n8804), .B(n8803), .S(n9934), .Z(n8810) );
  AOI22_X1 U10258 ( .A1(n8808), .A2(n8807), .B1(n8806), .B2(n8805), .ZN(n8809)
         );
  NAND2_X1 U10259 ( .A1(n8810), .A2(n8809), .ZN(P2_U3435) );
  MUX2_X1 U10260 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8811), .S(n9934), .Z(
        P2_U3432) );
  MUX2_X1 U10261 ( .A(n8812), .B(P2_REG0_REG_0__SCAN_IN), .S(n9936), .Z(
        P2_U3390) );
  INV_X1 U10262 ( .A(n8813), .ZN(n9479) );
  NOR4_X1 U10263 ( .A1(n8814), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5090), .ZN(n8815) );
  AOI21_X1 U10264 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n8823), .A(n8815), .ZN(
        n8816) );
  OAI21_X1 U10265 ( .B1(n9479), .B2(n8825), .A(n8816), .ZN(P2_U3264) );
  AOI22_X1 U10266 ( .A1(n5094), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8823), .ZN(n8817) );
  OAI21_X1 U10267 ( .B1(n8818), .B2(n8825), .A(n8817), .ZN(P2_U3265) );
  AOI22_X1 U10268 ( .A1(n8819), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8823), .ZN(n8820) );
  OAI21_X1 U10269 ( .B1(n8821), .B2(n8825), .A(n8820), .ZN(P2_U3266) );
  AOI21_X1 U10270 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8823), .A(n8822), .ZN(
        n8824) );
  OAI21_X1 U10271 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(P2_U3267) );
  MUX2_X1 U10272 ( .A(n8827), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10273 ( .B1(n8830), .B2(n8829), .A(n8828), .ZN(n8831) );
  OAI21_X1 U10274 ( .B1(n8832), .B2(n8831), .A(n9531), .ZN(n8837) );
  AND2_X1 U10275 ( .A1(n8963), .A2(n9343), .ZN(n8833) );
  AOI21_X1 U10276 ( .B1(n8961), .B2(n9345), .A(n8833), .ZN(n9155) );
  AOI22_X1 U10277 ( .A1(n9163), .A2(n8955), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8834) );
  OAI21_X1 U10278 ( .B1(n9155), .B2(n8952), .A(n8834), .ZN(n8835) );
  AOI21_X1 U10279 ( .B1(n9162), .B2(n8943), .A(n8835), .ZN(n8836) );
  NAND2_X1 U10280 ( .A1(n8837), .A2(n8836), .ZN(P1_U3214) );
  AOI21_X1 U10281 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8846) );
  NAND2_X1 U10282 ( .A1(n9344), .A2(n9345), .ZN(n8842) );
  NAND2_X1 U10283 ( .A1(n8971), .A2(n9343), .ZN(n8841) );
  AND2_X1 U10284 ( .A1(n8842), .A2(n8841), .ZN(n9637) );
  NAND2_X1 U10285 ( .A1(n8955), .A2(n9640), .ZN(n8843) );
  NAND2_X1 U10286 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9604) );
  OAI211_X1 U10287 ( .C1(n9637), .C2(n8952), .A(n8843), .B(n9604), .ZN(n8844)
         );
  AOI21_X1 U10288 ( .B1(n9430), .B2(n8943), .A(n8844), .ZN(n8845) );
  OAI21_X1 U10289 ( .B1(n8846), .B2(n8945), .A(n8845), .ZN(P1_U3215) );
  INV_X1 U10290 ( .A(n9380), .ZN(n9227) );
  INV_X1 U10291 ( .A(n8847), .ZN(n8925) );
  INV_X1 U10292 ( .A(n8848), .ZN(n8850) );
  NOR3_X1 U10293 ( .A1(n8925), .A2(n8850), .A3(n8849), .ZN(n8853) );
  INV_X1 U10294 ( .A(n8851), .ZN(n8852) );
  OAI21_X1 U10295 ( .B1(n8853), .B2(n8852), .A(n9531), .ZN(n8857) );
  NOR2_X1 U10296 ( .A1(n9236), .A2(n9535), .ZN(n8855) );
  OAI22_X1 U10297 ( .A1(n4292), .A2(n8938), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10032), .ZN(n8854) );
  AOI211_X1 U10298 ( .C1(n8940), .C2(n8965), .A(n8855), .B(n8854), .ZN(n8856)
         );
  OAI211_X1 U10299 ( .C1(n9227), .C2(n9528), .A(n8857), .B(n8856), .ZN(
        P1_U3216) );
  XOR2_X1 U10300 ( .A(n8859), .B(n8858), .Z(n8860) );
  XNOR2_X1 U10301 ( .A(n8861), .B(n8860), .ZN(n8867) );
  NAND2_X1 U10302 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9106) );
  OAI21_X1 U10303 ( .B1(n8938), .B2(n8862), .A(n9106), .ZN(n8863) );
  AOI21_X1 U10304 ( .B1(n8940), .B2(n9296), .A(n8863), .ZN(n8864) );
  OAI21_X1 U10305 ( .B1(n9535), .B2(n9288), .A(n8864), .ZN(n8865) );
  AOI21_X1 U10306 ( .B1(n9399), .B2(n8943), .A(n8865), .ZN(n8866) );
  OAI21_X1 U10307 ( .B1(n8867), .B2(n8945), .A(n8866), .ZN(P1_U3219) );
  OAI21_X1 U10308 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8877) );
  NAND2_X1 U10309 ( .A1(n9265), .A2(n8943), .ZN(n8875) );
  OR2_X1 U10310 ( .A1(n4292), .A2(n9723), .ZN(n8873) );
  OR2_X1 U10311 ( .A1(n8871), .A2(n9721), .ZN(n8872) );
  NAND2_X1 U10312 ( .A1(n8873), .A2(n8872), .ZN(n9261) );
  AOI22_X1 U10313 ( .A1(n9261), .A2(n9526), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8874) );
  OAI211_X1 U10314 ( .C1(n9535), .C2(n9266), .A(n8875), .B(n8874), .ZN(n8876)
         );
  AOI21_X1 U10315 ( .B1(n8877), .B2(n9531), .A(n8876), .ZN(n8878) );
  INV_X1 U10316 ( .A(n8878), .ZN(P1_U3223) );
  OAI21_X1 U10317 ( .B1(n8880), .B2(n8879), .A(n6481), .ZN(n8881) );
  NAND2_X1 U10318 ( .A1(n8881), .A2(n9531), .ZN(n8887) );
  NAND2_X1 U10319 ( .A1(n8963), .A2(n9345), .ZN(n8883) );
  NAND2_X1 U10320 ( .A1(n8965), .A2(n9343), .ZN(n8882) );
  NAND2_X1 U10321 ( .A1(n8883), .A2(n8882), .ZN(n9187) );
  INV_X1 U10322 ( .A(n9195), .ZN(n8884) );
  OAI22_X1 U10323 ( .A1(n8884), .A2(n9535), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10031), .ZN(n8885) );
  AOI21_X1 U10324 ( .B1(n9187), .B2(n9526), .A(n8885), .ZN(n8886) );
  OAI211_X1 U10325 ( .C1(n4434), .C2(n9528), .A(n8887), .B(n8886), .ZN(
        P1_U3225) );
  OAI21_X1 U10326 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8891) );
  NAND2_X1 U10327 ( .A1(n8891), .A2(n9531), .ZN(n8897) );
  NOR2_X1 U10328 ( .A1(n9535), .A2(n9338), .ZN(n8894) );
  NAND2_X1 U10329 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9056) );
  OAI21_X1 U10330 ( .B1(n8892), .B2(n8937), .A(n9056), .ZN(n8893) );
  AOI211_X1 U10331 ( .C1(n8895), .C2(n9344), .A(n8894), .B(n8893), .ZN(n8896)
         );
  OAI211_X1 U10332 ( .C1(n4429), .C2(n9528), .A(n8897), .B(n8896), .ZN(
        P1_U3226) );
  INV_X1 U10333 ( .A(n8898), .ZN(n8903) );
  AOI21_X1 U10334 ( .B1(n8900), .B2(n8902), .A(n8899), .ZN(n8901) );
  AOI21_X1 U10335 ( .B1(n8903), .B2(n8902), .A(n8901), .ZN(n8908) );
  NOR2_X1 U10336 ( .A1(n9535), .A2(n9327), .ZN(n8906) );
  AND2_X1 U10337 ( .A1(n8969), .A2(n9343), .ZN(n8904) );
  AOI21_X1 U10338 ( .B1(n9295), .B2(n9345), .A(n8904), .ZN(n9318) );
  NAND2_X1 U10339 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9078) );
  OAI21_X1 U10340 ( .B1(n9318), .B2(n8952), .A(n9078), .ZN(n8905) );
  AOI211_X1 U10341 ( .C1(n9325), .C2(n8943), .A(n8906), .B(n8905), .ZN(n8907)
         );
  OAI21_X1 U10342 ( .B1(n8908), .B2(n8945), .A(n8907), .ZN(P1_U3228) );
  AND2_X1 U10343 ( .A1(n8966), .A2(n9343), .ZN(n8909) );
  AOI21_X1 U10344 ( .B1(n8964), .B2(n9345), .A(n8909), .ZN(n9206) );
  AOI22_X1 U10345 ( .A1(n9212), .A2(n8955), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8910) );
  OAI21_X1 U10346 ( .B1(n9206), .B2(n8952), .A(n8910), .ZN(n8914) );
  OAI21_X1 U10347 ( .B1(n8915), .B2(n8917), .A(n8916), .ZN(n8918) );
  NAND2_X1 U10348 ( .A1(n8918), .A2(n9531), .ZN(n8923) );
  AND2_X1 U10349 ( .A1(n9311), .A2(n9343), .ZN(n8919) );
  AOI21_X1 U10350 ( .B1(n8968), .B2(n9345), .A(n8919), .ZN(n9276) );
  OAI22_X1 U10351 ( .A1(n9276), .A2(n8952), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8920), .ZN(n8921) );
  AOI21_X1 U10352 ( .B1(n9280), .B2(n8955), .A(n8921), .ZN(n8922) );
  OAI211_X1 U10353 ( .C1(n6035), .C2(n9528), .A(n8923), .B(n8922), .ZN(
        P1_U3233) );
  AOI21_X1 U10354 ( .B1(n8926), .B2(n8924), .A(n8925), .ZN(n8931) );
  AND2_X1 U10355 ( .A1(n8968), .A2(n9343), .ZN(n8927) );
  AOI21_X1 U10356 ( .B1(n8966), .B2(n9345), .A(n8927), .ZN(n9243) );
  AOI22_X1 U10357 ( .A1(n9249), .A2(n8955), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8928) );
  OAI21_X1 U10358 ( .B1(n9243), .B2(n8952), .A(n8928), .ZN(n8929) );
  AOI21_X1 U10359 ( .B1(n9248), .B2(n8943), .A(n8929), .ZN(n8930) );
  OAI21_X1 U10360 ( .B1(n8931), .B2(n8945), .A(n8930), .ZN(P1_U3235) );
  XNOR2_X1 U10361 ( .A(n8933), .B(n8932), .ZN(n8934) );
  XNOR2_X1 U10362 ( .A(n8935), .B(n8934), .ZN(n8946) );
  OAI22_X1 U10363 ( .A1(n8938), .A2(n8937), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8936), .ZN(n8939) );
  AOI21_X1 U10364 ( .B1(n8940), .B2(n9311), .A(n8939), .ZN(n8941) );
  OAI21_X1 U10365 ( .B1(n9535), .B2(n9304), .A(n8941), .ZN(n8942) );
  AOI21_X1 U10366 ( .B1(n9405), .B2(n8943), .A(n8942), .ZN(n8944) );
  OAI21_X1 U10367 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(P1_U3238) );
  OAI21_X1 U10368 ( .B1(n8949), .B2(n8948), .A(n8947), .ZN(n8950) );
  NAND2_X1 U10369 ( .A1(n8950), .A2(n9531), .ZN(n8957) );
  NAND2_X1 U10370 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9617) );
  OAI21_X1 U10371 ( .B1(n8952), .B2(n8951), .A(n9617), .ZN(n8953) );
  AOI21_X1 U10372 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8956) );
  OAI211_X1 U10373 ( .C1(n8958), .C2(n9528), .A(n8957), .B(n8956), .ZN(
        P1_U3241) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8959), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8960), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8961), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8962), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8963), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8964), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8965), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8966), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8967), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n8968), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9296), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9311), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9295), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9346), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8969), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9344), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8970), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8971), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8972), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8973), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8974), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8975), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8976), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8977), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8978), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8979), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8980), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8981), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8982), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8983), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10404 ( .C1(n8986), .C2(n8985), .A(n9623), .B(n8984), .ZN(n8993)
         );
  AOI22_X1 U10405 ( .A1(n9076), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8992) );
  INV_X1 U10406 ( .A(n9629), .ZN(n9616) );
  NAND2_X1 U10407 ( .A1(n9616), .A2(n8987), .ZN(n8991) );
  OAI211_X1 U10408 ( .C1(n8998), .C2(n8989), .A(n9595), .B(n8988), .ZN(n8990)
         );
  NAND4_X1 U10409 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(
        P1_U3244) );
  NAND2_X1 U10410 ( .A1(n8995), .A2(n8994), .ZN(n9001) );
  AOI22_X1 U10411 ( .A1(n8999), .A2(n8998), .B1(n8997), .B2(n8996), .ZN(n9000)
         );
  OAI211_X1 U10412 ( .C1(n9002), .C2(n9001), .A(P1_U3973), .B(n9000), .ZN(
        n9044) );
  INV_X1 U10413 ( .A(n9003), .ZN(n9006) );
  INV_X1 U10414 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9004) );
  OAI22_X1 U10415 ( .A1(n9635), .A2(n9004), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5818), .ZN(n9005) );
  AOI21_X1 U10416 ( .B1(n9616), .B2(n9006), .A(n9005), .ZN(n9015) );
  OAI211_X1 U10417 ( .C1(n9009), .C2(n9008), .A(n9623), .B(n9007), .ZN(n9014)
         );
  OAI211_X1 U10418 ( .C1(n9012), .C2(n9011), .A(n9595), .B(n9010), .ZN(n9013)
         );
  NAND4_X1 U10419 ( .A1(n9044), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(
        P1_U3245) );
  OAI211_X1 U10420 ( .C1(n9018), .C2(n9017), .A(n9623), .B(n9016), .ZN(n9029)
         );
  INV_X1 U10421 ( .A(n9019), .ZN(n9023) );
  INV_X1 U10422 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10423 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9020) );
  OAI21_X1 U10424 ( .B1(n9635), .B2(n9021), .A(n9020), .ZN(n9022) );
  AOI21_X1 U10425 ( .B1(n9616), .B2(n9023), .A(n9022), .ZN(n9028) );
  OAI211_X1 U10426 ( .C1(n9026), .C2(n9025), .A(n9595), .B(n9024), .ZN(n9027)
         );
  NAND3_X1 U10427 ( .A1(n9029), .A2(n9028), .A3(n9027), .ZN(P1_U3246) );
  INV_X1 U10428 ( .A(n9030), .ZN(n9034) );
  INV_X1 U10429 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9032) );
  OAI21_X1 U10430 ( .B1(n9635), .B2(n9032), .A(n9031), .ZN(n9033) );
  AOI21_X1 U10431 ( .B1(n9616), .B2(n9034), .A(n9033), .ZN(n9043) );
  OAI211_X1 U10432 ( .C1(n9037), .C2(n9036), .A(n9595), .B(n9035), .ZN(n9042)
         );
  OAI211_X1 U10433 ( .C1(n9040), .C2(n9039), .A(n9623), .B(n9038), .ZN(n9041)
         );
  NAND4_X1 U10434 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(
        P1_U3247) );
  INV_X1 U10435 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9045) );
  MUX2_X1 U10436 ( .A(n9045), .B(P1_REG1_REG_13__SCAN_IN), .S(n9587), .Z(n9580) );
  OAI21_X1 U10437 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9060), .A(n9046), .ZN(
        n9581) );
  NOR2_X1 U10438 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  AOI21_X1 U10439 ( .B1(n9587), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9579), .ZN(
        n9598) );
  INV_X1 U10440 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10441 ( .A1(n9062), .A2(n9047), .ZN(n9049) );
  NAND2_X1 U10442 ( .A1(n9602), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9048) );
  AND2_X1 U10443 ( .A1(n9049), .A2(n9048), .ZN(n9597) );
  NOR2_X1 U10444 ( .A1(n9598), .A2(n9597), .ZN(n9596) );
  AOI21_X1 U10445 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9062), .A(n9596), .ZN(
        n9050) );
  NOR2_X1 U10446 ( .A1(n9050), .A2(n9064), .ZN(n9051) );
  INV_X1 U10447 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9610) );
  XNOR2_X1 U10448 ( .A(n9064), .B(n9050), .ZN(n9609) );
  NOR2_X1 U10449 ( .A1(n9610), .A2(n9609), .ZN(n9608) );
  NOR2_X1 U10450 ( .A1(n9051), .A2(n9608), .ZN(n9054) );
  INV_X1 U10451 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9052) );
  AOI22_X1 U10452 ( .A1(n9075), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9052), .B2(
        n9057), .ZN(n9053) );
  NAND2_X1 U10453 ( .A1(n9053), .A2(n9054), .ZN(n9074) );
  OAI21_X1 U10454 ( .B1(n9054), .B2(n9053), .A(n9074), .ZN(n9071) );
  NAND2_X1 U10455 ( .A1(n9076), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9055) );
  OAI211_X1 U10456 ( .C1(n9629), .C2(n9057), .A(n9056), .B(n9055), .ZN(n9070)
         );
  NAND2_X1 U10457 ( .A1(n9587), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9058) );
  OAI21_X1 U10458 ( .B1(n9587), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9058), .ZN(
        n9583) );
  OAI21_X1 U10459 ( .B1(n9060), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9059), .ZN(
        n9584) );
  NOR2_X1 U10460 ( .A1(n9583), .A2(n9584), .ZN(n9582) );
  NAND2_X1 U10461 ( .A1(n9062), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9061) );
  OAI21_X1 U10462 ( .B1(n9062), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9061), .ZN(
        n9593) );
  NOR2_X1 U10463 ( .A1(n9592), .A2(n9593), .ZN(n9591) );
  NOR2_X1 U10464 ( .A1(n9063), .A2(n9064), .ZN(n9065) );
  INV_X1 U10465 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10018) );
  XNOR2_X1 U10466 ( .A(n9064), .B(n9063), .ZN(n9612) );
  NOR2_X1 U10467 ( .A1(n10018), .A2(n9612), .ZN(n9611) );
  NAND2_X1 U10468 ( .A1(n9075), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9066) );
  OAI21_X1 U10469 ( .B1(n9075), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9066), .ZN(
        n9067) );
  NOR2_X1 U10470 ( .A1(n9068), .A2(n9067), .ZN(n9073) );
  AOI211_X1 U10471 ( .C1(n9068), .C2(n9067), .A(n9073), .B(n9620), .ZN(n9069)
         );
  AOI211_X1 U10472 ( .C1(n9623), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9072)
         );
  INV_X1 U10473 ( .A(n9072), .ZN(P1_U3259) );
  XNOR2_X1 U10474 ( .A(n9085), .B(n9328), .ZN(n9083) );
  XOR2_X1 U10475 ( .A(n9083), .B(n9084), .Z(n9082) );
  OAI21_X1 U10476 ( .B1(n9075), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9074), .ZN(
        n9093) );
  XOR2_X1 U10477 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9085), .Z(n9092) );
  XNOR2_X1 U10478 ( .A(n9093), .B(n9092), .ZN(n9080) );
  NAND2_X1 U10479 ( .A1(n9076), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9077) );
  OAI211_X1 U10480 ( .C1(n9629), .C2(n9091), .A(n9078), .B(n9077), .ZN(n9079)
         );
  AOI21_X1 U10481 ( .B1(n9080), .B2(n9623), .A(n9079), .ZN(n9081) );
  OAI21_X1 U10482 ( .B1(n9082), .B2(n9620), .A(n9081), .ZN(P1_U3260) );
  INV_X1 U10483 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U10484 ( .A1(n9084), .A2(n9083), .ZN(n9087) );
  OR2_X1 U10485 ( .A1(n9085), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U10486 ( .A1(n9087), .A2(n9086), .ZN(n9622) );
  NAND2_X1 U10487 ( .A1(n9094), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9088) );
  OAI21_X1 U10488 ( .B1(n9094), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9088), .ZN(
        n9621) );
  NAND2_X1 U10489 ( .A1(n9631), .A2(n9088), .ZN(n9090) );
  INV_X1 U10490 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U10491 ( .A(n9090), .B(n9089), .ZN(n9099) );
  INV_X1 U10492 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9412) );
  AOI22_X1 U10493 ( .A1(n9093), .A2(n9092), .B1(n9412), .B2(n9091), .ZN(n9626)
         );
  NAND2_X1 U10494 ( .A1(n9094), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9096) );
  OAI21_X1 U10495 ( .B1(n9094), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9096), .ZN(
        n9095) );
  INV_X1 U10496 ( .A(n9095), .ZN(n9625) );
  NAND2_X1 U10497 ( .A1(n9626), .A2(n9625), .ZN(n9624) );
  NAND2_X1 U10498 ( .A1(n9624), .A2(n9096), .ZN(n9098) );
  XNOR2_X1 U10499 ( .A(n9098), .B(n9097), .ZN(n9100) );
  AOI22_X1 U10500 ( .A1(n9099), .A2(n9595), .B1(n9623), .B2(n9100), .ZN(n9105)
         );
  INV_X1 U10501 ( .A(n9099), .ZN(n9102) );
  INV_X1 U10502 ( .A(n9623), .ZN(n9607) );
  OAI21_X1 U10503 ( .B1(n9100), .B2(n9607), .A(n9629), .ZN(n9101) );
  AOI21_X1 U10504 ( .B1(n9102), .B2(n9595), .A(n9101), .ZN(n9104) );
  OAI211_X1 U10505 ( .C1(n9108), .C2(n9635), .A(n9107), .B(n9106), .ZN(
        P1_U3262) );
  NOR2_X1 U10506 ( .A1(n9677), .A2(n6220), .ZN(n9117) );
  AOI21_X1 U10507 ( .B1(n9677), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9117), .ZN(
        n9111) );
  NAND2_X1 U10508 ( .A1(n9109), .A2(n9652), .ZN(n9110) );
  OAI211_X1 U10509 ( .C1(n9113), .C2(n9112), .A(n9111), .B(n9110), .ZN(
        P1_U3263) );
  AOI211_X1 U10510 ( .C1(n9115), .C2(n9132), .A(n9740), .B(n9114), .ZN(n9354)
         );
  NAND2_X1 U10511 ( .A1(n9354), .A2(n10148), .ZN(n9119) );
  AND2_X1 U10512 ( .A1(n9677), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9116) );
  NOR2_X1 U10513 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  OAI211_X1 U10514 ( .C1(n7761), .C2(n10140), .A(n9119), .B(n9118), .ZN(
        P1_U3264) );
  XNOR2_X1 U10515 ( .A(n9130), .B(n9129), .ZN(n9356) );
  AOI21_X1 U10516 ( .B1(n7742), .B2(n9131), .A(n9740), .ZN(n9133) );
  NAND2_X1 U10517 ( .A1(n9357), .A2(n10148), .ZN(n9139) );
  INV_X1 U10518 ( .A(n9134), .ZN(n9137) );
  INV_X1 U10519 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9135) );
  NOR2_X1 U10520 ( .A1(n9326), .A2(n9135), .ZN(n9136) );
  AOI22_X1 U10521 ( .A1(n9137), .A2(n9136), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9677), .ZN(n9138) );
  OAI211_X1 U10522 ( .C1(n6212), .C2(n10140), .A(n9139), .B(n9138), .ZN(n9140)
         );
  AOI21_X1 U10523 ( .B1(n9356), .B2(n10150), .A(n9140), .ZN(n9141) );
  OAI21_X1 U10524 ( .B1(n4361), .B2(n9677), .A(n9141), .ZN(P1_U3356) );
  AOI22_X1 U10525 ( .A1(n9143), .A2(n10146), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n9677), .ZN(n9144) );
  OAI21_X1 U10526 ( .B1(n9145), .B2(n10140), .A(n9144), .ZN(n9148) );
  NOR2_X1 U10527 ( .A1(n9146), .A2(n9677), .ZN(n9147) );
  AOI211_X1 U10528 ( .C1(n6152), .C2(n10148), .A(n9148), .B(n9147), .ZN(n9149)
         );
  OAI21_X1 U10529 ( .B1(n9150), .B2(n9352), .A(n9149), .ZN(P1_U3265) );
  NAND2_X1 U10530 ( .A1(n9151), .A2(n9157), .ZN(n9152) );
  NAND2_X1 U10531 ( .A1(n9152), .A2(n9665), .ZN(n9153) );
  OR2_X1 U10532 ( .A1(n9154), .A2(n9153), .ZN(n9156) );
  NAND2_X1 U10533 ( .A1(n9156), .A2(n9155), .ZN(n9358) );
  INV_X1 U10534 ( .A(n9358), .ZN(n9168) );
  XNOR2_X1 U10535 ( .A(n9158), .B(n9157), .ZN(n9360) );
  NAND2_X1 U10536 ( .A1(n9360), .A2(n10150), .ZN(n9167) );
  INV_X1 U10537 ( .A(n9176), .ZN(n9161) );
  INV_X1 U10538 ( .A(n9159), .ZN(n9160) );
  AOI211_X1 U10539 ( .C1(n9162), .C2(n9161), .A(n9740), .B(n9160), .ZN(n9359)
         );
  AOI22_X1 U10540 ( .A1(n9163), .A2(n10146), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9677), .ZN(n9164) );
  OAI21_X1 U10541 ( .B1(n9439), .B2(n10140), .A(n9164), .ZN(n9165) );
  AOI21_X1 U10542 ( .B1(n9359), .B2(n10148), .A(n9165), .ZN(n9166) );
  OAI211_X1 U10543 ( .C1(n9168), .C2(n9677), .A(n9167), .B(n9166), .ZN(
        P1_U3266) );
  XNOR2_X1 U10544 ( .A(n9169), .B(n9175), .ZN(n9170) );
  NAND2_X1 U10545 ( .A1(n9170), .A2(n9665), .ZN(n9173) );
  INV_X1 U10546 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U10547 ( .A1(n9173), .A2(n9172), .ZN(n9363) );
  INV_X1 U10548 ( .A(n9363), .ZN(n9184) );
  XOR2_X1 U10549 ( .A(n9175), .B(n9174), .Z(n9365) );
  NAND2_X1 U10550 ( .A1(n9365), .A2(n10150), .ZN(n9183) );
  AOI211_X1 U10551 ( .C1(n9177), .C2(n9192), .A(n9740), .B(n9176), .ZN(n9364)
         );
  INV_X1 U10552 ( .A(n9178), .ZN(n9179) );
  AOI22_X1 U10553 ( .A1(n9179), .A2(n10146), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9677), .ZN(n9180) );
  OAI21_X1 U10554 ( .B1(n9442), .B2(n10140), .A(n9180), .ZN(n9181) );
  AOI21_X1 U10555 ( .B1(n9364), .B2(n10148), .A(n9181), .ZN(n9182) );
  OAI211_X1 U10556 ( .C1(n9677), .C2(n9184), .A(n9183), .B(n9182), .ZN(
        P1_U3267) );
  OAI211_X1 U10557 ( .C1(n9186), .C2(n9190), .A(n9185), .B(n9665), .ZN(n9189)
         );
  INV_X1 U10558 ( .A(n9187), .ZN(n9188) );
  NAND2_X1 U10559 ( .A1(n9189), .A2(n9188), .ZN(n9368) );
  INV_X1 U10560 ( .A(n9368), .ZN(n9200) );
  XOR2_X1 U10561 ( .A(n9191), .B(n9190), .Z(n9370) );
  NAND2_X1 U10562 ( .A1(n9370), .A2(n10150), .ZN(n9199) );
  INV_X1 U10563 ( .A(n9192), .ZN(n9193) );
  AOI211_X1 U10564 ( .C1(n9194), .C2(n9209), .A(n9740), .B(n9193), .ZN(n9369)
         );
  AOI22_X1 U10565 ( .A1(n9195), .A2(n10146), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9677), .ZN(n9196) );
  OAI21_X1 U10566 ( .B1(n4434), .B2(n10140), .A(n9196), .ZN(n9197) );
  AOI21_X1 U10567 ( .B1(n9369), .B2(n10148), .A(n9197), .ZN(n9198) );
  OAI211_X1 U10568 ( .C1(n9677), .C2(n9200), .A(n9199), .B(n9198), .ZN(
        P1_U3268) );
  NAND2_X1 U10569 ( .A1(n9229), .A2(n9201), .ZN(n9203) );
  NAND2_X1 U10570 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  NAND3_X1 U10571 ( .A1(n9205), .A2(n9204), .A3(n9665), .ZN(n9207) );
  NAND2_X1 U10572 ( .A1(n9207), .A2(n9206), .ZN(n9373) );
  INV_X1 U10573 ( .A(n9373), .ZN(n9217) );
  XNOR2_X1 U10574 ( .A(n4316), .B(n9208), .ZN(n9375) );
  NAND2_X1 U10575 ( .A1(n9375), .A2(n10150), .ZN(n9216) );
  INV_X1 U10576 ( .A(n9209), .ZN(n9210) );
  AOI211_X1 U10577 ( .C1(n9211), .C2(n4438), .A(n9740), .B(n9210), .ZN(n9374)
         );
  AOI22_X1 U10578 ( .A1(n9212), .A2(n10146), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9677), .ZN(n9213) );
  OAI21_X1 U10579 ( .B1(n9448), .B2(n10140), .A(n9213), .ZN(n9214) );
  AOI21_X1 U10580 ( .B1(n9374), .B2(n10148), .A(n9214), .ZN(n9215) );
  OAI211_X1 U10581 ( .C1(n9677), .C2(n9217), .A(n9216), .B(n9215), .ZN(
        P1_U3269) );
  INV_X1 U10582 ( .A(n9218), .ZN(n9221) );
  AOI22_X1 U10583 ( .A1(n9222), .A2(n9221), .B1(n9220), .B2(n9219), .ZN(n9382)
         );
  NAND2_X1 U10584 ( .A1(n9380), .A2(n9245), .ZN(n9223) );
  NAND2_X1 U10585 ( .A1(n9223), .A2(n9711), .ZN(n9224) );
  NOR2_X1 U10586 ( .A1(n9225), .A2(n9224), .ZN(n9379) );
  INV_X1 U10587 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9226) );
  OAI22_X1 U10588 ( .A1(n9227), .A2(n10140), .B1(n9226), .B2(n10141), .ZN(
        n9228) );
  AOI21_X1 U10589 ( .B1(n9379), .B2(n10148), .A(n9228), .ZN(n9239) );
  INV_X1 U10590 ( .A(n9229), .ZN(n9230) );
  AOI21_X1 U10591 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9233) );
  OAI222_X1 U10592 ( .A1(n9723), .A2(n9235), .B1(n9721), .B2(n4292), .C1(n9719), .C2(n9233), .ZN(n9378) );
  NOR2_X1 U10593 ( .A1(n9236), .A2(n9326), .ZN(n9237) );
  OAI21_X1 U10594 ( .B1(n9378), .B2(n9237), .A(n10141), .ZN(n9238) );
  OAI211_X1 U10595 ( .C1(n9382), .C2(n9352), .A(n9239), .B(n9238), .ZN(
        P1_U3270) );
  XNOR2_X1 U10596 ( .A(n9240), .B(n9241), .ZN(n9385) );
  INV_X1 U10597 ( .A(n9385), .ZN(n9254) );
  XNOR2_X1 U10598 ( .A(n4317), .B(n4508), .ZN(n9242) );
  NAND2_X1 U10599 ( .A1(n9242), .A2(n9665), .ZN(n9244) );
  NAND2_X1 U10600 ( .A1(n9244), .A2(n9243), .ZN(n9383) );
  INV_X1 U10601 ( .A(n9264), .ZN(n9247) );
  INV_X1 U10602 ( .A(n9245), .ZN(n9246) );
  AOI211_X1 U10603 ( .C1(n9248), .C2(n9247), .A(n9740), .B(n9246), .ZN(n9384)
         );
  NAND2_X1 U10604 ( .A1(n9384), .A2(n10148), .ZN(n9251) );
  AOI22_X1 U10605 ( .A1(n9249), .A2(n10146), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9677), .ZN(n9250) );
  OAI211_X1 U10606 ( .C1(n9453), .C2(n10140), .A(n9251), .B(n9250), .ZN(n9252)
         );
  AOI21_X1 U10607 ( .B1(n10141), .B2(n9383), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10608 ( .B1(n9254), .B2(n9352), .A(n9253), .ZN(P1_U3271) );
  XOR2_X1 U10609 ( .A(n9260), .B(n9255), .Z(n9390) );
  INV_X1 U10610 ( .A(n9390), .ZN(n9272) );
  INV_X1 U10611 ( .A(n9256), .ZN(n9257) );
  AOI21_X1 U10612 ( .B1(n4312), .B2(n9258), .A(n9257), .ZN(n9259) );
  XNOR2_X1 U10613 ( .A(n9260), .B(n9259), .ZN(n9263) );
  INV_X1 U10614 ( .A(n9261), .ZN(n9262) );
  OAI21_X1 U10615 ( .B1(n9263), .B2(n9719), .A(n9262), .ZN(n9388) );
  AOI211_X1 U10616 ( .C1(n9265), .C2(n9279), .A(n9740), .B(n9264), .ZN(n9389)
         );
  NAND2_X1 U10617 ( .A1(n9389), .A2(n10148), .ZN(n9269) );
  INV_X1 U10618 ( .A(n9266), .ZN(n9267) );
  AOI22_X1 U10619 ( .A1(n9267), .A2(n10146), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n9677), .ZN(n9268) );
  OAI211_X1 U10620 ( .C1(n9457), .C2(n10140), .A(n9269), .B(n9268), .ZN(n9270)
         );
  AOI21_X1 U10621 ( .B1(n10141), .B2(n9388), .A(n9270), .ZN(n9271) );
  OAI21_X1 U10622 ( .B1(n9272), .B2(n9352), .A(n9271), .ZN(P1_U3272) );
  AOI21_X1 U10623 ( .B1(n7634), .B2(n9274), .A(n9273), .ZN(n9395) );
  XNOR2_X1 U10624 ( .A(n9275), .B(n4312), .ZN(n9278) );
  INV_X1 U10625 ( .A(n9276), .ZN(n9277) );
  AOI21_X1 U10626 ( .B1(n9278), .B2(n9665), .A(n9277), .ZN(n9394) );
  INV_X1 U10627 ( .A(n9394), .ZN(n9284) );
  OAI211_X1 U10628 ( .C1(n6035), .C2(n9287), .A(n9711), .B(n9279), .ZN(n9393)
         );
  NOR2_X1 U10629 ( .A1(n9393), .A2(n9655), .ZN(n9283) );
  AOI22_X1 U10630 ( .A1(n9280), .A2(n10146), .B1(n9677), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9281) );
  OAI21_X1 U10631 ( .B1(n6035), .B2(n10140), .A(n9281), .ZN(n9282) );
  AOI211_X1 U10632 ( .C1(n9284), .C2(n10141), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI21_X1 U10633 ( .B1(n9395), .B2(n9352), .A(n9285), .ZN(P1_U3273) );
  XOR2_X1 U10634 ( .A(n9286), .B(n9294), .Z(n9403) );
  AOI21_X1 U10635 ( .B1(n9399), .B2(n9302), .A(n9287), .ZN(n9400) );
  INV_X1 U10636 ( .A(n9288), .ZN(n9289) );
  AOI22_X1 U10637 ( .A1(n9677), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9289), .B2(
        n10146), .ZN(n9290) );
  OAI21_X1 U10638 ( .B1(n9291), .B2(n10140), .A(n9290), .ZN(n9299) );
  OAI21_X1 U10639 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9297) );
  AOI222_X1 U10640 ( .A1(n9665), .A2(n9297), .B1(n9296), .B2(n9345), .C1(n9295), .C2(n9343), .ZN(n9402) );
  NOR2_X1 U10641 ( .A1(n9402), .A2(n9677), .ZN(n9298) );
  AOI211_X1 U10642 ( .C1(n9400), .C2(n9350), .A(n9299), .B(n9298), .ZN(n9300)
         );
  OAI21_X1 U10643 ( .B1(n9403), .B2(n9352), .A(n9300), .ZN(P1_U3274) );
  XOR2_X1 U10644 ( .A(n9301), .B(n9310), .Z(n9408) );
  INV_X1 U10645 ( .A(n9302), .ZN(n9303) );
  AOI211_X1 U10646 ( .C1(n9405), .C2(n9322), .A(n9740), .B(n9303), .ZN(n9404)
         );
  INV_X1 U10647 ( .A(n9304), .ZN(n9305) );
  AOI22_X1 U10648 ( .A1(n9677), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9305), .B2(
        n10146), .ZN(n9306) );
  OAI21_X1 U10649 ( .B1(n9307), .B2(n10140), .A(n9306), .ZN(n9314) );
  OAI21_X1 U10650 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9312) );
  AOI222_X1 U10651 ( .A1(n9665), .A2(n9312), .B1(n9311), .B2(n9345), .C1(n9346), .C2(n9343), .ZN(n9407) );
  NOR2_X1 U10652 ( .A1(n9407), .A2(n9677), .ZN(n9313) );
  AOI211_X1 U10653 ( .C1(n9404), .C2(n10148), .A(n9314), .B(n9313), .ZN(n9315)
         );
  OAI21_X1 U10654 ( .B1(n9408), .B2(n9352), .A(n9315), .ZN(P1_U3275) );
  XNOR2_X1 U10655 ( .A(n9316), .B(n9320), .ZN(n9317) );
  OR2_X1 U10656 ( .A1(n9317), .A2(n9719), .ZN(n9319) );
  NAND2_X1 U10657 ( .A1(n9319), .A2(n9318), .ZN(n9409) );
  INV_X1 U10658 ( .A(n9409), .ZN(n9333) );
  XNOR2_X1 U10659 ( .A(n9321), .B(n9320), .ZN(n9411) );
  NAND2_X1 U10660 ( .A1(n9411), .A2(n10150), .ZN(n9332) );
  INV_X1 U10661 ( .A(n9336), .ZN(n9324) );
  INV_X1 U10662 ( .A(n9322), .ZN(n9323) );
  AOI211_X1 U10663 ( .C1(n9325), .C2(n9324), .A(n9740), .B(n9323), .ZN(n9410)
         );
  NOR2_X1 U10664 ( .A1(n9466), .A2(n10140), .ZN(n9330) );
  OAI22_X1 U10665 ( .A1(n10141), .A2(n9328), .B1(n9327), .B2(n9326), .ZN(n9329) );
  AOI211_X1 U10666 ( .C1(n9410), .C2(n10148), .A(n9330), .B(n9329), .ZN(n9331)
         );
  OAI211_X1 U10667 ( .C1(n9677), .C2(n9333), .A(n9332), .B(n9331), .ZN(
        P1_U3276) );
  XNOR2_X1 U10668 ( .A(n9335), .B(n9334), .ZN(n9420) );
  AOI21_X1 U10669 ( .B1(n9415), .B2(n9337), .A(n9336), .ZN(n9417) );
  INV_X1 U10670 ( .A(n9338), .ZN(n9339) );
  AOI22_X1 U10671 ( .A1(n9677), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9339), .B2(
        n10146), .ZN(n9340) );
  OAI21_X1 U10672 ( .B1(n4429), .B2(n10140), .A(n9340), .ZN(n9349) );
  XNOR2_X1 U10673 ( .A(n9342), .B(n9341), .ZN(n9347) );
  AOI222_X1 U10674 ( .A1(n9665), .A2(n9347), .B1(n9346), .B2(n9345), .C1(n9344), .C2(n9343), .ZN(n9419) );
  NOR2_X1 U10675 ( .A1(n9419), .A2(n9677), .ZN(n9348) );
  AOI211_X1 U10676 ( .C1(n9417), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9351)
         );
  OAI21_X1 U10677 ( .B1(n9420), .B2(n9352), .A(n9351), .ZN(P1_U3277) );
  INV_X1 U10678 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10078) );
  NOR2_X1 U10679 ( .A1(n9354), .A2(n9353), .ZN(n9432) );
  MUX2_X1 U10680 ( .A(n10078), .B(n9432), .S(n9770), .Z(n9355) );
  OAI21_X1 U10681 ( .B1(n7761), .B2(n9414), .A(n9355), .ZN(P1_U3552) );
  AOI211_X1 U10682 ( .C1(n9360), .C2(n9750), .A(n9359), .B(n9358), .ZN(n9436)
         );
  MUX2_X1 U10683 ( .A(n9361), .B(n9436), .S(n9770), .Z(n9362) );
  OAI21_X1 U10684 ( .B1(n9439), .B2(n9414), .A(n9362), .ZN(P1_U3549) );
  INV_X1 U10685 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9366) );
  AOI211_X1 U10686 ( .C1(n9365), .C2(n9750), .A(n9364), .B(n9363), .ZN(n9440)
         );
  MUX2_X1 U10687 ( .A(n9366), .B(n9440), .S(n9770), .Z(n9367) );
  OAI21_X1 U10688 ( .B1(n9442), .B2(n9414), .A(n9367), .ZN(P1_U3548) );
  AOI211_X1 U10689 ( .C1(n9370), .C2(n9750), .A(n9369), .B(n9368), .ZN(n9443)
         );
  MUX2_X1 U10690 ( .A(n9371), .B(n9443), .S(n9770), .Z(n9372) );
  OAI21_X1 U10691 ( .B1(n4434), .B2(n9414), .A(n9372), .ZN(P1_U3547) );
  INV_X1 U10692 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9376) );
  AOI211_X1 U10693 ( .C1(n9375), .C2(n9750), .A(n9374), .B(n9373), .ZN(n9446)
         );
  MUX2_X1 U10694 ( .A(n9376), .B(n9446), .S(n9770), .Z(n9377) );
  OAI21_X1 U10695 ( .B1(n9448), .B2(n9414), .A(n9377), .ZN(P1_U3546) );
  AOI211_X1 U10696 ( .C1(n9416), .C2(n9380), .A(n9379), .B(n9378), .ZN(n9381)
         );
  OAI21_X1 U10697 ( .B1(n9382), .B2(n9683), .A(n9381), .ZN(n9449) );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9449), .S(n9770), .Z(
        P1_U3545) );
  AOI211_X1 U10699 ( .C1(n9385), .C2(n9750), .A(n9384), .B(n9383), .ZN(n9450)
         );
  MUX2_X1 U10700 ( .A(n9386), .B(n9450), .S(n9770), .Z(n9387) );
  OAI21_X1 U10701 ( .B1(n9453), .B2(n9414), .A(n9387), .ZN(P1_U3544) );
  AOI211_X1 U10702 ( .C1(n9390), .C2(n9750), .A(n9389), .B(n9388), .ZN(n9454)
         );
  MUX2_X1 U10703 ( .A(n9391), .B(n9454), .S(n9770), .Z(n9392) );
  OAI21_X1 U10704 ( .B1(n9457), .B2(n9414), .A(n9392), .ZN(P1_U3543) );
  OAI211_X1 U10705 ( .C1(n9395), .C2(n9683), .A(n9394), .B(n9393), .ZN(n9396)
         );
  INV_X1 U10706 ( .A(n9396), .ZN(n9458) );
  MUX2_X1 U10707 ( .A(n9397), .B(n9458), .S(n9770), .Z(n9398) );
  OAI21_X1 U10708 ( .B1(n6035), .B2(n9414), .A(n9398), .ZN(P1_U3542) );
  AOI22_X1 U10709 ( .A1(n9400), .A2(n9711), .B1(n9416), .B2(n9399), .ZN(n9401)
         );
  OAI211_X1 U10710 ( .C1(n9403), .C2(n9683), .A(n9402), .B(n9401), .ZN(n9461)
         );
  MUX2_X1 U10711 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9461), .S(n9770), .Z(
        P1_U3541) );
  AOI21_X1 U10712 ( .B1(n9416), .B2(n9405), .A(n9404), .ZN(n9406) );
  OAI211_X1 U10713 ( .C1(n9408), .C2(n9683), .A(n9407), .B(n9406), .ZN(n9462)
         );
  MUX2_X1 U10714 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9462), .S(n9770), .Z(
        P1_U3540) );
  AOI211_X1 U10715 ( .C1(n9411), .C2(n9750), .A(n9410), .B(n9409), .ZN(n9463)
         );
  MUX2_X1 U10716 ( .A(n9412), .B(n9463), .S(n9770), .Z(n9413) );
  OAI21_X1 U10717 ( .B1(n9466), .B2(n9414), .A(n9413), .ZN(P1_U3539) );
  AOI22_X1 U10718 ( .A1(n9417), .A2(n9711), .B1(n9416), .B2(n9415), .ZN(n9418)
         );
  OAI211_X1 U10719 ( .C1(n9420), .C2(n9683), .A(n9419), .B(n9418), .ZN(n9467)
         );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9467), .S(n9770), .Z(
        P1_U3538) );
  XOR2_X1 U10721 ( .A(n9421), .B(n9422), .Z(n9639) );
  INV_X1 U10722 ( .A(n9639), .ZN(n9647) );
  AOI21_X1 U10723 ( .B1(n9423), .B2(n9422), .A(n9719), .ZN(n9425) );
  NAND2_X1 U10724 ( .A1(n9425), .A2(n9424), .ZN(n9636) );
  NAND2_X1 U10725 ( .A1(n9426), .A2(n9430), .ZN(n9427) );
  NAND3_X1 U10726 ( .A1(n4366), .A2(n9711), .A3(n9427), .ZN(n9645) );
  NAND3_X1 U10727 ( .A1(n9636), .A2(n9637), .A3(n9645), .ZN(n9428) );
  AOI21_X1 U10728 ( .B1(n9647), .B2(n9750), .A(n9428), .ZN(n9472) );
  AOI22_X1 U10729 ( .A1(n9430), .A2(n9429), .B1(n9768), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n9431) );
  OAI21_X1 U10730 ( .B1(n9472), .B2(n9768), .A(n9431), .ZN(P1_U3536) );
  INV_X1 U10731 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9433) );
  MUX2_X1 U10732 ( .A(n9433), .B(n9432), .S(n9753), .Z(n9434) );
  OAI21_X1 U10733 ( .B1(n7761), .B2(n9469), .A(n9434), .ZN(P1_U3520) );
  MUX2_X1 U10734 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9435), .S(n9753), .Z(
        P1_U3519) );
  INV_X1 U10735 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9437) );
  MUX2_X1 U10736 ( .A(n9437), .B(n9436), .S(n9753), .Z(n9438) );
  OAI21_X1 U10737 ( .B1(n9439), .B2(n9469), .A(n9438), .ZN(P1_U3517) );
  MUX2_X1 U10738 ( .A(n10014), .B(n9440), .S(n9753), .Z(n9441) );
  OAI21_X1 U10739 ( .B1(n9442), .B2(n9469), .A(n9441), .ZN(P1_U3516) );
  INV_X1 U10740 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9444) );
  MUX2_X1 U10741 ( .A(n9444), .B(n9443), .S(n9753), .Z(n9445) );
  OAI21_X1 U10742 ( .B1(n4434), .B2(n9469), .A(n9445), .ZN(P1_U3515) );
  MUX2_X1 U10743 ( .A(n10125), .B(n9446), .S(n9753), .Z(n9447) );
  OAI21_X1 U10744 ( .B1(n9448), .B2(n9469), .A(n9447), .ZN(P1_U3514) );
  MUX2_X1 U10745 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9449), .S(n9753), .Z(
        P1_U3513) );
  INV_X1 U10746 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9451) );
  MUX2_X1 U10747 ( .A(n9451), .B(n9450), .S(n9753), .Z(n9452) );
  OAI21_X1 U10748 ( .B1(n9453), .B2(n9469), .A(n9452), .ZN(P1_U3512) );
  INV_X1 U10749 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9455) );
  MUX2_X1 U10750 ( .A(n9455), .B(n9454), .S(n9753), .Z(n9456) );
  OAI21_X1 U10751 ( .B1(n9457), .B2(n9469), .A(n9456), .ZN(P1_U3511) );
  INV_X1 U10752 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U10753 ( .A(n9459), .B(n9458), .S(n9753), .Z(n9460) );
  OAI21_X1 U10754 ( .B1(n6035), .B2(n9469), .A(n9460), .ZN(P1_U3510) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9461), .S(n9753), .Z(
        P1_U3509) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9462), .S(n9753), .Z(
        P1_U3507) );
  INV_X1 U10757 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9464) );
  MUX2_X1 U10758 ( .A(n9464), .B(n9463), .S(n9753), .Z(n9465) );
  OAI21_X1 U10759 ( .B1(n9466), .B2(n9469), .A(n9465), .ZN(P1_U3504) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9467), .S(n9753), .Z(
        P1_U3501) );
  INV_X1 U10761 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9468) );
  OAI22_X1 U10762 ( .A1(n9642), .A2(n9469), .B1(n9753), .B2(n9468), .ZN(n9470)
         );
  INV_X1 U10763 ( .A(n9470), .ZN(n9471) );
  OAI21_X1 U10764 ( .B1(n9472), .B2(n9752), .A(n9471), .ZN(P1_U3495) );
  NOR4_X1 U10765 ( .A1(n9474), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9473), .ZN(n9475) );
  AOI21_X1 U10766 ( .B1(n9476), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9475), .ZN(
        n9477) );
  OAI21_X1 U10767 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(P1_U3324) );
  MUX2_X1 U10768 ( .A(n9480), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10769 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9491) );
  AOI211_X1 U10770 ( .C1(n9483), .C2(n9482), .A(n9607), .B(n9481), .ZN(n9488)
         );
  AOI211_X1 U10771 ( .C1(n9486), .C2(n9485), .A(n9620), .B(n9484), .ZN(n9487)
         );
  AOI211_X1 U10772 ( .C1(n9616), .C2(n9489), .A(n9488), .B(n9487), .ZN(n9490)
         );
  NAND2_X1 U10773 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9523) );
  OAI211_X1 U10774 ( .C1(n9635), .C2(n9491), .A(n9490), .B(n9523), .ZN(
        P1_U3253) );
  INV_X1 U10775 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10034) );
  AOI21_X1 U10776 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9495) );
  NAND2_X1 U10777 ( .A1(n9595), .A2(n9495), .ZN(n9501) );
  AOI21_X1 U10778 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9499) );
  NAND2_X1 U10779 ( .A1(n9623), .A2(n9499), .ZN(n9500) );
  OAI211_X1 U10780 ( .C1(n9629), .C2(n9502), .A(n9501), .B(n9500), .ZN(n9503)
         );
  INV_X1 U10781 ( .A(n9503), .ZN(n9505) );
  OAI211_X1 U10782 ( .C1(n9635), .C2(n10034), .A(n9505), .B(n9504), .ZN(
        P1_U3250) );
  INV_X1 U10783 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9520) );
  AOI21_X1 U10784 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9509) );
  NAND2_X1 U10785 ( .A1(n9595), .A2(n9509), .ZN(n9515) );
  AOI21_X1 U10786 ( .B1(n9512), .B2(n9511), .A(n9510), .ZN(n9513) );
  NAND2_X1 U10787 ( .A1(n9623), .A2(n9513), .ZN(n9514) );
  OAI211_X1 U10788 ( .C1(n9629), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9517)
         );
  INV_X1 U10789 ( .A(n9517), .ZN(n9519) );
  OAI211_X1 U10790 ( .C1(n9635), .C2(n9520), .A(n9519), .B(n9518), .ZN(
        P1_U3251) );
  OAI21_X1 U10791 ( .B1(n9522), .B2(n9521), .A(n7284), .ZN(n9532) );
  INV_X1 U10792 ( .A(n9523), .ZN(n9524) );
  AOI21_X1 U10793 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  OAI21_X1 U10794 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9530) );
  AOI21_X1 U10795 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9533) );
  OAI21_X1 U10796 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(P1_U3217) );
  INV_X1 U10797 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9536) );
  AOI22_X1 U10798 ( .A1(n9770), .A2(n9537), .B1(n9536), .B2(n9768), .ZN(
        P1_U3553) );
  INV_X1 U10799 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10047) );
  XOR2_X1 U10800 ( .A(n10047), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10801 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9551) );
  INV_X1 U10802 ( .A(n9538), .ZN(n9539) );
  OAI211_X1 U10803 ( .C1(n9541), .C2(n9540), .A(n9595), .B(n9539), .ZN(n9548)
         );
  NAND2_X1 U10804 ( .A1(n9616), .A2(n9542), .ZN(n9547) );
  OAI211_X1 U10805 ( .C1(n9545), .C2(n9544), .A(n9623), .B(n9543), .ZN(n9546)
         );
  AND3_X1 U10806 ( .A1(n9548), .A2(n9547), .A3(n9546), .ZN(n9550) );
  NAND2_X1 U10807 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9549) );
  OAI211_X1 U10808 ( .C1(n9635), .C2(n9551), .A(n9550), .B(n9549), .ZN(
        P1_U3248) );
  INV_X1 U10809 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9566) );
  AOI21_X1 U10810 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9555) );
  NAND2_X1 U10811 ( .A1(n9595), .A2(n9555), .ZN(n9561) );
  AOI21_X1 U10812 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9559) );
  NAND2_X1 U10813 ( .A1(n9623), .A2(n9559), .ZN(n9560) );
  OAI211_X1 U10814 ( .C1(n9629), .C2(n9562), .A(n9561), .B(n9560), .ZN(n9563)
         );
  INV_X1 U10815 ( .A(n9563), .ZN(n9565) );
  NAND2_X1 U10816 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9564) );
  OAI211_X1 U10817 ( .C1(n9635), .C2(n9566), .A(n9565), .B(n9564), .ZN(
        P1_U3249) );
  INV_X1 U10818 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9578) );
  AOI211_X1 U10819 ( .C1(n9569), .C2(n9568), .A(n9567), .B(n9620), .ZN(n9574)
         );
  AOI211_X1 U10820 ( .C1(n9572), .C2(n9571), .A(n9607), .B(n9570), .ZN(n9573)
         );
  AOI211_X1 U10821 ( .C1(n9616), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9577)
         );
  OAI211_X1 U10822 ( .C1(n9635), .C2(n9578), .A(n9577), .B(n9576), .ZN(
        P1_U3254) );
  INV_X1 U10823 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9590) );
  AOI211_X1 U10824 ( .C1(n9581), .C2(n9580), .A(n9579), .B(n9607), .ZN(n9586)
         );
  AOI211_X1 U10825 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9620), .ZN(n9585)
         );
  AOI211_X1 U10826 ( .C1(n9616), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9589)
         );
  OAI211_X1 U10827 ( .C1(n9635), .C2(n9590), .A(n9589), .B(n9588), .ZN(
        P1_U3256) );
  INV_X1 U10828 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9606) );
  AOI21_X1 U10829 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9594) );
  NAND2_X1 U10830 ( .A1(n9595), .A2(n9594), .ZN(n9601) );
  AOI21_X1 U10831 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  NAND2_X1 U10832 ( .A1(n9623), .A2(n9599), .ZN(n9600) );
  OAI211_X1 U10833 ( .C1(n9629), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9603)
         );
  INV_X1 U10834 ( .A(n9603), .ZN(n9605) );
  OAI211_X1 U10835 ( .C1(n9635), .C2(n9606), .A(n9605), .B(n9604), .ZN(
        P1_U3257) );
  INV_X1 U10836 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9619) );
  AOI211_X1 U10837 ( .C1(n9610), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9614)
         );
  AOI211_X1 U10838 ( .C1(n9612), .C2(n10018), .A(n9611), .B(n9620), .ZN(n9613)
         );
  AOI211_X1 U10839 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9618)
         );
  OAI211_X1 U10840 ( .C1(n9635), .C2(n9619), .A(n9618), .B(n9617), .ZN(
        P1_U3258) );
  AOI21_X1 U10841 ( .B1(n9622), .B2(n9621), .A(n9620), .ZN(n9632) );
  OAI211_X1 U10842 ( .C1(n9626), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9627)
         );
  OAI21_X1 U10843 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9630) );
  AOI21_X1 U10844 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9634) );
  NAND2_X1 U10845 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9633) );
  OAI211_X1 U10846 ( .C1(n9635), .C2(n9961), .A(n9634), .B(n9633), .ZN(
        P1_U3261) );
  OAI211_X1 U10847 ( .C1(n9639), .C2(n9638), .A(n9637), .B(n9636), .ZN(n9644)
         );
  AOI22_X1 U10848 ( .A1(n9677), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9640), .B2(
        n10146), .ZN(n9641) );
  OAI21_X1 U10849 ( .B1(n9642), .B2(n10140), .A(n9641), .ZN(n9643) );
  AOI21_X1 U10850 ( .B1(n9644), .B2(n10141), .A(n9643), .ZN(n9649) );
  INV_X1 U10851 ( .A(n9645), .ZN(n9646) );
  AOI22_X1 U10852 ( .A1(n9647), .A2(n9658), .B1(n10148), .B2(n9646), .ZN(n9648) );
  NAND2_X1 U10853 ( .A1(n9649), .A2(n9648), .ZN(P1_U3279) );
  AOI22_X1 U10854 ( .A1(n9677), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9650), .B2(
        n10146), .ZN(n9654) );
  NAND2_X1 U10855 ( .A1(n9652), .A2(n9651), .ZN(n9653) );
  OAI211_X1 U10856 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9657)
         );
  AOI21_X1 U10857 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(n9660) );
  OAI21_X1 U10858 ( .B1(n9677), .B2(n9661), .A(n9660), .ZN(P1_U3286) );
  XNOR2_X1 U10859 ( .A(n9669), .B(n9662), .ZN(n9666) );
  INV_X1 U10860 ( .A(n9663), .ZN(n9664) );
  AOI21_X1 U10861 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9697) );
  AOI22_X1 U10862 ( .A1(n9677), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10146), .ZN(n9667) );
  OAI21_X1 U10863 ( .B1(n10140), .B2(n5834), .A(n9667), .ZN(n9668) );
  INV_X1 U10864 ( .A(n9668), .ZN(n9676) );
  XNOR2_X1 U10865 ( .A(n9670), .B(n9669), .ZN(n9700) );
  OAI21_X1 U10866 ( .B1(n9671), .B2(n5834), .A(n9711), .ZN(n9673) );
  OR2_X1 U10867 ( .A1(n9673), .A2(n9672), .ZN(n9696) );
  INV_X1 U10868 ( .A(n9696), .ZN(n9674) );
  AOI22_X1 U10869 ( .A1(n9700), .A2(n10150), .B1(n9674), .B2(n10148), .ZN(
        n9675) );
  OAI211_X1 U10870 ( .C1(n9677), .C2(n9697), .A(n9676), .B(n9675), .ZN(
        P1_U3291) );
  AND2_X1 U10871 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9679), .ZN(P1_U3294) );
  AND2_X1 U10872 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9679), .ZN(P1_U3295) );
  AND2_X1 U10873 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9679), .ZN(P1_U3296) );
  AND2_X1 U10874 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9679), .ZN(P1_U3297) );
  AND2_X1 U10875 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9679), .ZN(P1_U3298) );
  AND2_X1 U10876 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9679), .ZN(P1_U3299) );
  AND2_X1 U10877 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9679), .ZN(P1_U3300) );
  AND2_X1 U10878 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9679), .ZN(P1_U3301) );
  AND2_X1 U10879 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9679), .ZN(P1_U3302) );
  AND2_X1 U10880 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9679), .ZN(P1_U3303) );
  AND2_X1 U10881 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9679), .ZN(P1_U3304) );
  AND2_X1 U10882 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9679), .ZN(P1_U3305) );
  AND2_X1 U10883 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9679), .ZN(P1_U3306) );
  AND2_X1 U10884 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9679), .ZN(P1_U3307) );
  AND2_X1 U10885 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9679), .ZN(P1_U3308) );
  INV_X1 U10886 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U10887 ( .A1(n9678), .A2(n10076), .ZN(P1_U3309) );
  AND2_X1 U10888 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9679), .ZN(P1_U3310) );
  AND2_X1 U10889 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9679), .ZN(P1_U3311) );
  AND2_X1 U10890 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9679), .ZN(P1_U3312) );
  AND2_X1 U10891 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9679), .ZN(P1_U3313) );
  AND2_X1 U10892 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9679), .ZN(P1_U3314) );
  AND2_X1 U10893 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9679), .ZN(P1_U3315) );
  AND2_X1 U10894 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9679), .ZN(P1_U3316) );
  AND2_X1 U10895 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9679), .ZN(P1_U3317) );
  AND2_X1 U10896 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9679), .ZN(P1_U3318) );
  AND2_X1 U10897 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9679), .ZN(P1_U3319) );
  AND2_X1 U10898 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9679), .ZN(P1_U3320) );
  AND2_X1 U10899 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9679), .ZN(P1_U3321) );
  AND2_X1 U10900 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9679), .ZN(P1_U3322) );
  AND2_X1 U10901 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9679), .ZN(P1_U3323) );
  INV_X1 U10902 ( .A(n9680), .ZN(n9685) );
  INV_X1 U10903 ( .A(n9681), .ZN(n9682) );
  AOI21_X1 U10904 ( .B1(n9683), .B2(n9719), .A(n9682), .ZN(n9684) );
  AOI211_X1 U10905 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9754)
         );
  INV_X1 U10906 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U10907 ( .A1(n9753), .A2(n9754), .B1(n9688), .B2(n9752), .ZN(
        P1_U3453) );
  INV_X1 U10908 ( .A(n9689), .ZN(n9731) );
  OAI21_X1 U10909 ( .B1(n9691), .B2(n9748), .A(n9690), .ZN(n9693) );
  AOI211_X1 U10910 ( .C1(n9731), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9756)
         );
  INV_X1 U10911 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10912 ( .A1(n9753), .A2(n9756), .B1(n9695), .B2(n9752), .ZN(
        P1_U3456) );
  OAI21_X1 U10913 ( .B1(n5834), .B2(n9748), .A(n9696), .ZN(n9699) );
  INV_X1 U10914 ( .A(n9697), .ZN(n9698) );
  AOI211_X1 U10915 ( .C1(n9750), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9757)
         );
  INV_X1 U10916 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9701) );
  AOI22_X1 U10917 ( .A1(n9753), .A2(n9757), .B1(n9701), .B2(n9752), .ZN(
        P1_U3459) );
  OAI21_X1 U10918 ( .B1(n9703), .B2(n9748), .A(n9702), .ZN(n9705) );
  AOI211_X1 U10919 ( .C1(n9750), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9759)
         );
  INV_X1 U10920 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U10921 ( .A1(n9753), .A2(n9759), .B1(n9707), .B2(n9752), .ZN(
        P1_U3462) );
  XNOR2_X1 U10922 ( .A(n9708), .B(n9714), .ZN(n10151) );
  INV_X1 U10923 ( .A(n9709), .ZN(n9712) );
  OAI211_X1 U10924 ( .C1(n9712), .C2(n10139), .A(n9711), .B(n9710), .ZN(n10147) );
  OAI21_X1 U10925 ( .B1(n10139), .B2(n9748), .A(n10147), .ZN(n9724) );
  NAND3_X1 U10926 ( .A1(n9715), .A2(n9714), .A3(n9713), .ZN(n9716) );
  AND2_X1 U10927 ( .A1(n9717), .A2(n9716), .ZN(n9718) );
  OAI222_X1 U10928 ( .A1(n9723), .A2(n9722), .B1(n9721), .B2(n9720), .C1(n9719), .C2(n9718), .ZN(n10142) );
  AOI211_X1 U10929 ( .C1(n9750), .C2(n10151), .A(n9724), .B(n10142), .ZN(n9761) );
  INV_X1 U10930 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10931 ( .A1(n9753), .A2(n9761), .B1(n9725), .B2(n9752), .ZN(
        P1_U3465) );
  OAI21_X1 U10932 ( .B1(n9727), .B2(n9748), .A(n9726), .ZN(n9729) );
  AOI211_X1 U10933 ( .C1(n9731), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9763)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U10935 ( .A1(n9753), .A2(n9763), .B1(n10083), .B2(n9752), .ZN(
        P1_U3477) );
  OAI21_X1 U10936 ( .B1(n9733), .B2(n9748), .A(n9732), .ZN(n9734) );
  AOI21_X1 U10937 ( .B1(n9735), .B2(n9750), .A(n9734), .ZN(n9736) );
  AND2_X1 U10938 ( .A1(n9737), .A2(n9736), .ZN(n9765) );
  INV_X1 U10939 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9738) );
  AOI22_X1 U10940 ( .A1(n9753), .A2(n9765), .B1(n9738), .B2(n9752), .ZN(
        P1_U3480) );
  OAI22_X1 U10941 ( .A1(n9741), .A2(n9740), .B1(n9739), .B2(n9748), .ZN(n9742)
         );
  AOI211_X1 U10942 ( .C1(n9744), .C2(n9750), .A(n9743), .B(n9742), .ZN(n9767)
         );
  INV_X1 U10943 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9745) );
  AOI22_X1 U10944 ( .A1(n9753), .A2(n9767), .B1(n9745), .B2(n9752), .ZN(
        P1_U3489) );
  OAI211_X1 U10945 ( .C1(n4772), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9749)
         );
  AOI21_X1 U10946 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9769) );
  INV_X1 U10947 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U10948 ( .A1(n9753), .A2(n9769), .B1(n10105), .B2(n9752), .ZN(
        P1_U3492) );
  AOI22_X1 U10949 ( .A1(n9770), .A2(n9754), .B1(n6554), .B2(n9768), .ZN(
        P1_U3522) );
  AOI22_X1 U10950 ( .A1(n9770), .A2(n9756), .B1(n9755), .B2(n9768), .ZN(
        P1_U3523) );
  AOI22_X1 U10951 ( .A1(n9770), .A2(n9757), .B1(n10096), .B2(n9768), .ZN(
        P1_U3524) );
  INV_X1 U10952 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U10953 ( .A1(n9770), .A2(n9759), .B1(n9758), .B2(n9768), .ZN(
        P1_U3525) );
  AOI22_X1 U10954 ( .A1(n9770), .A2(n9761), .B1(n9760), .B2(n9768), .ZN(
        P1_U3526) );
  INV_X1 U10955 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9762) );
  AOI22_X1 U10956 ( .A1(n9770), .A2(n9763), .B1(n9762), .B2(n9768), .ZN(
        P1_U3530) );
  AOI22_X1 U10957 ( .A1(n9770), .A2(n9765), .B1(n9764), .B2(n9768), .ZN(
        P1_U3531) );
  AOI22_X1 U10958 ( .A1(n9770), .A2(n9767), .B1(n9766), .B2(n9768), .ZN(
        P1_U3534) );
  AOI22_X1 U10959 ( .A1(n9770), .A2(n9769), .B1(n9045), .B2(n9768), .ZN(
        P1_U3535) );
  NAND2_X1 U10960 ( .A1(n9817), .A2(n9771), .ZN(n9786) );
  OAI21_X1 U10961 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9776) );
  NOR2_X1 U10962 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7620), .ZN(n9775) );
  AOI21_X1 U10963 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9785) );
  INV_X1 U10964 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9778) );
  OR2_X1 U10965 ( .A1(n9832), .A2(n9778), .ZN(n9784) );
  OAI21_X1 U10966 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9782) );
  NAND2_X1 U10967 ( .A1(n9821), .A2(n9782), .ZN(n9783) );
  AND4_X1 U10968 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(n9791)
         );
  XOR2_X1 U10969 ( .A(n9788), .B(n9787), .Z(n9789) );
  NAND2_X1 U10970 ( .A1(n9789), .A2(n9843), .ZN(n9790) );
  NAND2_X1 U10971 ( .A1(n9791), .A2(n9790), .ZN(P2_U3184) );
  AOI21_X1 U10972 ( .B1(n9794), .B2(n9793), .A(n9792), .ZN(n9795) );
  OAI22_X1 U10973 ( .A1(n9795), .A2(n9848), .B1(n4587), .B2(n9835), .ZN(n9796)
         );
  AOI21_X1 U10974 ( .B1(n9797), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9796), .ZN(
        n9808) );
  AOI21_X1 U10975 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  OR2_X1 U10976 ( .A1(n9801), .A2(n9826), .ZN(n9806) );
  OAI21_X1 U10977 ( .B1(n9803), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9802), .ZN(
        n9804) );
  NAND2_X1 U10978 ( .A1(n9804), .A2(n9821), .ZN(n9805) );
  NAND4_X1 U10979 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(
        P2_U3189) );
  INV_X1 U10980 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9830) );
  INV_X1 U10981 ( .A(n9809), .ZN(n9810) );
  OAI21_X1 U10982 ( .B1(n9811), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9810), .ZN(
        n9822) );
  AOI21_X1 U10983 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9819) );
  AOI21_X1 U10984 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9818) );
  OAI21_X1 U10985 ( .B1(n9819), .B2(n9848), .A(n9818), .ZN(n9820) );
  AOI21_X1 U10986 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9829) );
  AOI21_X1 U10987 ( .B1(n9825), .B2(n9824), .A(n9823), .ZN(n9827) );
  OR2_X1 U10988 ( .A1(n9827), .A2(n9826), .ZN(n9828) );
  OAI211_X1 U10989 ( .C1(n9830), .C2(n9832), .A(n9829), .B(n9828), .ZN(
        P2_U3191) );
  INV_X1 U10990 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9831) );
  OR2_X1 U10991 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  OAI21_X1 U10992 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  INV_X1 U10993 ( .A(n9836), .ZN(n9856) );
  AOI21_X1 U10994 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(n9853) );
  OAI21_X1 U10995 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9844) );
  NAND2_X1 U10996 ( .A1(n9844), .A2(n9843), .ZN(n9851) );
  AOI21_X1 U10997 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9849) );
  OR2_X1 U10998 ( .A1(n9849), .A2(n9848), .ZN(n9850) );
  OAI211_X1 U10999 ( .C1(n9853), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9854)
         );
  INV_X1 U11000 ( .A(n9854), .ZN(n9855) );
  OAI211_X1 U11001 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8294), .A(n9856), .B(
        n9855), .ZN(P2_U3199) );
  OAI21_X1 U11002 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9884) );
  INV_X1 U11003 ( .A(n9884), .ZN(n9875) );
  AOI22_X1 U11004 ( .A1(n9862), .A2(n7101), .B1(n9861), .B2(n9860), .ZN(n9869)
         );
  OAI21_X1 U11005 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9867) );
  NAND2_X1 U11006 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  OAI211_X1 U11007 ( .C1(n9875), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9882)
         );
  NOR2_X1 U11008 ( .A1(n9871), .A2(n9928), .ZN(n9883) );
  INV_X1 U11009 ( .A(n9883), .ZN(n9872) );
  OAI22_X1 U11010 ( .A1(n9875), .A2(n9874), .B1(n9873), .B2(n9872), .ZN(n9876)
         );
  AOI211_X1 U11011 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n9877), .A(n9882), .B(
        n9876), .ZN(n9879) );
  AOI22_X1 U11012 ( .A1(n9881), .A2(n9880), .B1(n9879), .B2(n9878), .ZN(
        P2_U3231) );
  AOI211_X1 U11013 ( .C1(n9926), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9938)
         );
  AOI22_X1 U11014 ( .A1(n9936), .A2(n5122), .B1(n9938), .B2(n9934), .ZN(
        P2_U3396) );
  INV_X1 U11015 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U11016 ( .A1(n9885), .A2(n9933), .ZN(n9888) );
  NAND2_X1 U11017 ( .A1(n9886), .A2(n9920), .ZN(n9887) );
  AND3_X1 U11018 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(n9940) );
  AOI22_X1 U11019 ( .A1(n9936), .A2(n9890), .B1(n9940), .B2(n9934), .ZN(
        P2_U3399) );
  AOI22_X1 U11020 ( .A1(n9892), .A2(n9933), .B1(n9920), .B2(n9891), .ZN(n9893)
         );
  AND2_X1 U11021 ( .A1(n9894), .A2(n9893), .ZN(n9942) );
  AOI22_X1 U11022 ( .A1(n9936), .A2(n5176), .B1(n9942), .B2(n9934), .ZN(
        P2_U3402) );
  INV_X1 U11023 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9899) );
  INV_X1 U11024 ( .A(n9926), .ZN(n9915) );
  OAI22_X1 U11025 ( .A1(n9896), .A2(n9915), .B1(n9895), .B2(n9928), .ZN(n9897)
         );
  NOR2_X1 U11026 ( .A1(n9898), .A2(n9897), .ZN(n9944) );
  AOI22_X1 U11027 ( .A1(n9936), .A2(n9899), .B1(n9944), .B2(n9934), .ZN(
        P2_U3405) );
  OR2_X1 U11028 ( .A1(n9900), .A2(n9911), .ZN(n9903) );
  NAND2_X1 U11029 ( .A1(n9901), .A2(n9920), .ZN(n9902) );
  AOI22_X1 U11030 ( .A1(n9936), .A2(n5220), .B1(n9945), .B2(n9934), .ZN(
        P2_U3408) );
  INV_X1 U11031 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9909) );
  OAI22_X1 U11032 ( .A1(n9906), .A2(n9915), .B1(n9905), .B2(n9928), .ZN(n9907)
         );
  NOR2_X1 U11033 ( .A1(n9908), .A2(n9907), .ZN(n9946) );
  AOI22_X1 U11034 ( .A1(n9936), .A2(n9909), .B1(n9946), .B2(n9934), .ZN(
        P2_U3411) );
  OAI22_X1 U11035 ( .A1(n9912), .A2(n9911), .B1(n9910), .B2(n9928), .ZN(n9913)
         );
  NOR2_X1 U11036 ( .A1(n9914), .A2(n9913), .ZN(n9947) );
  AOI22_X1 U11037 ( .A1(n9936), .A2(n5261), .B1(n9947), .B2(n9934), .ZN(
        P2_U3414) );
  INV_X1 U11038 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U11039 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  AOI211_X1 U11040 ( .C1(n9920), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9949)
         );
  AOI22_X1 U11041 ( .A1(n9936), .A2(n9921), .B1(n9949), .B2(n9934), .ZN(
        P2_U3417) );
  INV_X1 U11042 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U11043 ( .A1(n9922), .A2(n9928), .ZN(n9924) );
  AOI211_X1 U11044 ( .C1(n9926), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9951)
         );
  AOI22_X1 U11045 ( .A1(n9936), .A2(n9927), .B1(n9951), .B2(n9934), .ZN(
        P2_U3420) );
  INV_X1 U11046 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U11047 ( .A1(n9929), .A2(n9928), .ZN(n9931) );
  AOI211_X1 U11048 ( .C1(n9933), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9953)
         );
  AOI22_X1 U11049 ( .A1(n9936), .A2(n9935), .B1(n9953), .B2(n9934), .ZN(
        P2_U3423) );
  AOI22_X1 U11050 ( .A1(n9954), .A2(n9938), .B1(n9937), .B2(n5718), .ZN(
        P2_U3461) );
  AOI22_X1 U11051 ( .A1(n9954), .A2(n9940), .B1(n9939), .B2(n5718), .ZN(
        P2_U3462) );
  AOI22_X1 U11052 ( .A1(n9954), .A2(n9942), .B1(n9941), .B2(n5718), .ZN(
        P2_U3463) );
  AOI22_X1 U11053 ( .A1(n9954), .A2(n9944), .B1(n9943), .B2(n5718), .ZN(
        P2_U3464) );
  AOI22_X1 U11054 ( .A1(n9954), .A2(n9945), .B1(n5223), .B2(n5718), .ZN(
        P2_U3465) );
  AOI22_X1 U11055 ( .A1(n9954), .A2(n9946), .B1(n5240), .B2(n5718), .ZN(
        P2_U3466) );
  AOI22_X1 U11056 ( .A1(n9954), .A2(n9947), .B1(n5264), .B2(n5718), .ZN(
        P2_U3467) );
  AOI22_X1 U11057 ( .A1(n9954), .A2(n9949), .B1(n9948), .B2(n5718), .ZN(
        P2_U3468) );
  AOI22_X1 U11058 ( .A1(n9954), .A2(n9951), .B1(n9950), .B2(n5718), .ZN(
        P2_U3469) );
  AOI22_X1 U11059 ( .A1(n9954), .A2(n9953), .B1(n9952), .B2(n5718), .ZN(
        P2_U3470) );
  OAI222_X1 U11060 ( .A1(n9959), .A2(n9958), .B1(n9959), .B2(n9957), .C1(n9956), .C2(n9955), .ZN(ADD_1068_U5) );
  XOR2_X1 U11061 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11062 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9963) );
  INV_X1 U11063 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10057) );
  XOR2_X1 U11064 ( .A(n9963), .B(n10057), .Z(ADD_1068_U55) );
  OAI21_X1 U11065 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(ADD_1068_U56) );
  OAI21_X1 U11066 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(ADD_1068_U57) );
  OAI21_X1 U11067 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(ADD_1068_U58) );
  OAI21_X1 U11068 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(ADD_1068_U59) );
  OAI21_X1 U11069 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(ADD_1068_U60) );
  OAI21_X1 U11070 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(ADD_1068_U61) );
  OAI21_X1 U11071 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(ADD_1068_U62) );
  OAI21_X1 U11072 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(ADD_1068_U63) );
  NOR4_X1 U11073 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(n10092), .A4(n10108), .ZN(n10011) );
  NAND4_X1 U11074 ( .A1(SI_24_), .A2(P2_DATAO_REG_16__SCAN_IN), .A3(
        P2_DATAO_REG_9__SCAN_IN), .A4(P2_IR_REG_22__SCAN_IN), .ZN(n9990) );
  NAND4_X1 U11075 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P2_REG1_REG_27__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P2_ADDR_REG_11__SCAN_IN), .ZN(n9989)
         );
  NAND4_X1 U11076 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(
        P1_DATAO_REG_17__SCAN_IN), .A3(P2_D_REG_12__SCAN_IN), .A4(
        P2_REG0_REG_2__SCAN_IN), .ZN(n9988) );
  NOR3_X1 U11077 ( .A1(n9990), .A2(n9989), .A3(n9988), .ZN(n10010) );
  NAND4_X1 U11078 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(P2_REG1_REG_12__SCAN_IN), 
        .A3(P2_REG2_REG_8__SCAN_IN), .A4(P2_REG1_REG_13__SCAN_IN), .ZN(n9994)
         );
  NAND4_X1 U11079 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n9993)
         );
  NAND4_X1 U11080 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG2_REG_23__SCAN_IN), 
        .A3(P1_REG1_REG_6__SCAN_IN), .A4(P2_WR_REG_SCAN_IN), .ZN(n9992) );
  NAND4_X1 U11081 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(P2_REG2_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_19__SCAN_IN), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n9991)
         );
  NOR4_X1 U11082 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n10009)
         );
  NOR4_X1 U11083 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_29__SCAN_IN), .A4(P2_REG1_REG_25__SCAN_IN), .ZN(n9998)
         );
  NOR4_X1 U11084 ( .A1(SI_6_), .A2(SI_5_), .A3(P2_REG3_REG_9__SCAN_IN), .A4(
        P2_REG0_REG_4__SCAN_IN), .ZN(n9997) );
  NOR4_X1 U11085 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(P1_REG0_REG_13__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(P2_IR_REG_1__SCAN_IN), .ZN(n9996) );
  NOR4_X1 U11086 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(P1_REG2_REG_15__SCAN_IN), 
        .A3(P1_REG2_REG_11__SCAN_IN), .A4(P1_REG2_REG_18__SCAN_IN), .ZN(n9995)
         );
  NAND4_X1 U11087 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10007) );
  INV_X1 U11088 ( .A(n9999), .ZN(n10006) );
  INV_X1 U11089 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10114) );
  NAND4_X1 U11090 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10114), .A3(n5857), .A4(
        n10096), .ZN(n10005) );
  NAND4_X1 U11091 ( .A1(n10058), .A2(n10000), .A3(P1_IR_REG_28__SCAN_IN), .A4(
        P1_IR_REG_29__SCAN_IN), .ZN(n10003) );
  NAND4_X1 U11092 ( .A1(n10001), .A2(P1_DATAO_REG_2__SCAN_IN), .A3(
        P2_RD_REG_SCAN_IN), .A4(P1_IR_REG_12__SCAN_IN), .ZN(n10002) );
  OR4_X1 U11093 ( .A1(n10003), .A2(n10002), .A3(n10027), .A4(n10034), .ZN(
        n10004) );
  NOR4_X1 U11094 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n10008) );
  NAND4_X1 U11095 ( .A1(n10011), .A2(n10010), .A3(n10009), .A4(n10008), .ZN(
        n10157) );
  AOI22_X1 U11096 ( .A1(n10014), .A2(keyinput63), .B1(keyinput53), .B2(n10013), 
        .ZN(n10012) );
  OAI221_X1 U11097 ( .B1(n10014), .B2(keyinput63), .C1(n10013), .C2(keyinput53), .A(n10012), .ZN(n10025) );
  AOI22_X1 U11098 ( .A1(n10017), .A2(keyinput20), .B1(n10016), .B2(keyinput45), 
        .ZN(n10015) );
  OAI221_X1 U11099 ( .B1(n10017), .B2(keyinput20), .C1(n10016), .C2(keyinput45), .A(n10015), .ZN(n10024) );
  XOR2_X1 U11100 ( .A(n10018), .B(keyinput15), .Z(n10022) );
  XNOR2_X1 U11101 ( .A(SI_24_), .B(keyinput3), .ZN(n10021) );
  XNOR2_X1 U11102 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput40), .ZN(n10020)
         );
  XNOR2_X1 U11103 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput39), .ZN(n10019) );
  NAND4_X1 U11104 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10023) );
  NOR3_X1 U11105 ( .A1(n10025), .A2(n10024), .A3(n10023), .ZN(n10074) );
  AOI22_X1 U11106 ( .A1(n7318), .A2(keyinput34), .B1(keyinput42), .B2(n10027), 
        .ZN(n10026) );
  OAI221_X1 U11107 ( .B1(n7318), .B2(keyinput34), .C1(n10027), .C2(keyinput42), 
        .A(n10026), .ZN(n10039) );
  AOI22_X1 U11108 ( .A1(n5283), .A2(keyinput49), .B1(keyinput14), .B2(n10029), 
        .ZN(n10028) );
  OAI221_X1 U11109 ( .B1(n5283), .B2(keyinput49), .C1(n10029), .C2(keyinput14), 
        .A(n10028), .ZN(n10038) );
  AOI22_X1 U11110 ( .A1(n10032), .A2(keyinput43), .B1(n10031), .B2(keyinput6), 
        .ZN(n10030) );
  OAI221_X1 U11111 ( .B1(n10032), .B2(keyinput43), .C1(n10031), .C2(keyinput6), 
        .A(n10030), .ZN(n10037) );
  AOI22_X1 U11112 ( .A1(n10035), .A2(keyinput28), .B1(keyinput7), .B2(n10034), 
        .ZN(n10033) );
  OAI221_X1 U11113 ( .B1(n10035), .B2(keyinput28), .C1(n10034), .C2(keyinput7), 
        .A(n10033), .ZN(n10036) );
  NOR4_X1 U11114 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n10073) );
  XOR2_X1 U11115 ( .A(keyinput17), .B(n10040), .Z(n10044) );
  XNOR2_X1 U11116 ( .A(keyinput44), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10043) );
  XNOR2_X1 U11117 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput18), .ZN(n10042) );
  XNOR2_X1 U11118 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput2), .ZN(n10041) );
  NAND4_X1 U11119 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10053) );
  INV_X1 U11120 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11121 ( .A1(n10047), .A2(keyinput29), .B1(n10046), .B2(keyinput31), 
        .ZN(n10045) );
  OAI221_X1 U11122 ( .B1(n10047), .B2(keyinput29), .C1(n10046), .C2(keyinput31), .A(n10045), .ZN(n10052) );
  AOI22_X1 U11123 ( .A1(n10050), .A2(keyinput60), .B1(n10049), .B2(keyinput19), 
        .ZN(n10048) );
  OAI221_X1 U11124 ( .B1(n10050), .B2(keyinput60), .C1(n10049), .C2(keyinput19), .A(n10048), .ZN(n10051) );
  NOR3_X1 U11125 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10072) );
  INV_X1 U11126 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11127 ( .A1(n10056), .A2(keyinput38), .B1(keyinput22), .B2(n10055), 
        .ZN(n10054) );
  OAI221_X1 U11128 ( .B1(n10056), .B2(keyinput38), .C1(n10055), .C2(keyinput22), .A(n10054), .ZN(n10061) );
  XNOR2_X1 U11129 ( .A(n10057), .B(keyinput57), .ZN(n10060) );
  XNOR2_X1 U11130 ( .A(n10058), .B(keyinput0), .ZN(n10059) );
  OR3_X1 U11131 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10070) );
  INV_X1 U11132 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10064) );
  INV_X1 U11133 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11134 ( .A1(n10064), .A2(keyinput16), .B1(n10063), .B2(keyinput12), 
        .ZN(n10062) );
  OAI221_X1 U11135 ( .B1(n10064), .B2(keyinput16), .C1(n10063), .C2(keyinput12), .A(n10062), .ZN(n10069) );
  AOI22_X1 U11136 ( .A1(n10067), .A2(keyinput26), .B1(n10066), .B2(keyinput21), 
        .ZN(n10065) );
  OAI221_X1 U11137 ( .B1(n10067), .B2(keyinput26), .C1(n10066), .C2(keyinput21), .A(n10065), .ZN(n10068) );
  NOR3_X1 U11138 ( .A1(n10070), .A2(n10069), .A3(n10068), .ZN(n10071) );
  NAND4_X1 U11139 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10138) );
  AOI22_X1 U11140 ( .A1(n10076), .A2(keyinput48), .B1(keyinput8), .B2(n5176), 
        .ZN(n10075) );
  OAI221_X1 U11141 ( .B1(n10076), .B2(keyinput48), .C1(n5176), .C2(keyinput8), 
        .A(n10075), .ZN(n10089) );
  AOI22_X1 U11142 ( .A1(n10079), .A2(keyinput32), .B1(keyinput47), .B2(n10078), 
        .ZN(n10077) );
  OAI221_X1 U11143 ( .B1(n10079), .B2(keyinput32), .C1(n10078), .C2(keyinput47), .A(n10077), .ZN(n10088) );
  INV_X1 U11144 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11145 ( .A1(n10082), .A2(keyinput13), .B1(n10081), .B2(keyinput46), 
        .ZN(n10080) );
  OAI221_X1 U11146 ( .B1(n10082), .B2(keyinput13), .C1(n10081), .C2(keyinput46), .A(n10080), .ZN(n10087) );
  XOR2_X1 U11147 ( .A(n10083), .B(keyinput55), .Z(n10085) );
  XNOR2_X1 U11148 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput58), .ZN(n10084) );
  NAND2_X1 U11149 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  NOR4_X1 U11150 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10136) );
  AOI22_X1 U11151 ( .A1(n10092), .A2(keyinput4), .B1(n10091), .B2(keyinput41), 
        .ZN(n10090) );
  OAI221_X1 U11152 ( .B1(n10092), .B2(keyinput4), .C1(n10091), .C2(keyinput41), 
        .A(n10090), .ZN(n10103) );
  INV_X1 U11153 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11154 ( .A1(n9226), .A2(keyinput24), .B1(n10094), .B2(keyinput50), 
        .ZN(n10093) );
  OAI221_X1 U11155 ( .B1(n9226), .B2(keyinput24), .C1(n10094), .C2(keyinput50), 
        .A(n10093), .ZN(n10102) );
  AOI22_X1 U11156 ( .A1(n10097), .A2(keyinput36), .B1(n10096), .B2(keyinput35), 
        .ZN(n10095) );
  OAI221_X1 U11157 ( .B1(n10097), .B2(keyinput36), .C1(n10096), .C2(keyinput35), .A(n10095), .ZN(n10101) );
  XNOR2_X1 U11158 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput9), .ZN(n10099) );
  XNOR2_X1 U11159 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput62), .ZN(n10098) );
  NAND2_X1 U11160 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NOR4_X1 U11161 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10135) );
  INV_X1 U11162 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11163 ( .A1(n10106), .A2(keyinput25), .B1(n10105), .B2(keyinput54), 
        .ZN(n10104) );
  OAI221_X1 U11164 ( .B1(n10106), .B2(keyinput25), .C1(n10105), .C2(keyinput54), .A(n10104), .ZN(n10118) );
  AOI22_X1 U11165 ( .A1(n10109), .A2(keyinput23), .B1(n10108), .B2(keyinput52), 
        .ZN(n10107) );
  OAI221_X1 U11166 ( .B1(n10109), .B2(keyinput23), .C1(n10108), .C2(keyinput52), .A(n10107), .ZN(n10117) );
  INV_X1 U11167 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11168 ( .A1(n10112), .A2(keyinput37), .B1(n10111), .B2(keyinput51), 
        .ZN(n10110) );
  OAI221_X1 U11169 ( .B1(n10112), .B2(keyinput37), .C1(n10111), .C2(keyinput51), .A(n10110), .ZN(n10116) );
  AOI22_X1 U11170 ( .A1(n10114), .A2(keyinput5), .B1(n5857), .B2(keyinput1), 
        .ZN(n10113) );
  OAI221_X1 U11171 ( .B1(n10114), .B2(keyinput5), .C1(n5857), .C2(keyinput1), 
        .A(n10113), .ZN(n10115) );
  NOR4_X1 U11172 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10134) );
  AOI22_X1 U11173 ( .A1(n10121), .A2(keyinput10), .B1(keyinput33), .B2(n10120), 
        .ZN(n10119) );
  OAI221_X1 U11174 ( .B1(n10121), .B2(keyinput10), .C1(n10120), .C2(keyinput33), .A(n10119), .ZN(n10132) );
  AOI22_X1 U11175 ( .A1(n10123), .A2(keyinput59), .B1(keyinput27), .B2(n10001), 
        .ZN(n10122) );
  OAI221_X1 U11176 ( .B1(n10123), .B2(keyinput59), .C1(n10001), .C2(keyinput27), .A(n10122), .ZN(n10131) );
  AOI22_X1 U11177 ( .A1(n10125), .A2(keyinput56), .B1(keyinput11), .B2(n5122), 
        .ZN(n10124) );
  OAI221_X1 U11178 ( .B1(n10125), .B2(keyinput56), .C1(n5122), .C2(keyinput11), 
        .A(n10124), .ZN(n10130) );
  AOI22_X1 U11179 ( .A1(n10128), .A2(keyinput30), .B1(keyinput61), .B2(n10127), 
        .ZN(n10126) );
  OAI221_X1 U11180 ( .B1(n10128), .B2(keyinput30), .C1(n10127), .C2(keyinput61), .A(n10126), .ZN(n10129) );
  NOR4_X1 U11181 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10133) );
  NAND4_X1 U11182 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  NOR2_X1 U11183 ( .A1(n10138), .A2(n10137), .ZN(n10155) );
  NOR2_X1 U11184 ( .A1(n10140), .A2(n10139), .ZN(n10144) );
  MUX2_X1 U11185 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10142), .S(n10141), .Z(
        n10143) );
  AOI211_X1 U11186 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10153) );
  INV_X1 U11187 ( .A(n10147), .ZN(n10149) );
  AOI22_X1 U11188 ( .A1(n10151), .A2(n10150), .B1(n10149), .B2(n10148), .ZN(
        n10152) );
  NAND2_X1 U11189 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  XOR2_X1 U11190 ( .A(n10155), .B(n10154), .Z(n10156) );
  XNOR2_X1 U11191 ( .A(n10157), .B(n10156), .ZN(P1_U3289) );
  OAI21_X1 U11192 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(ADD_1068_U50) );
  OAI21_X1 U11193 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(ADD_1068_U51) );
  OAI21_X1 U11194 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(ADD_1068_U47) );
  OAI21_X1 U11195 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(ADD_1068_U49) );
  OAI21_X1 U11196 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(ADD_1068_U48) );
  AOI21_X1 U11197 ( .B1(n10175), .B2(n10174), .A(n10173), .ZN(ADD_1068_U54) );
  AOI21_X1 U11198 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(ADD_1068_U53) );
  OAI21_X1 U11199 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(ADD_1068_U52) );
  INV_X1 U4802 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9473) );
  INV_X2 U4871 ( .A(n8127), .ZN(n8128) );
  CLKBUF_X1 U4827 ( .A(n5325), .Z(n6513) );
  XNOR2_X1 U4852 ( .A(n5758), .B(n5757), .ZN(n8220) );
endmodule

