

module b14_C_SARLock_k_64_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621;

  INV_X2 U2266 ( .A(n2871), .ZN(n2854) );
  INV_X1 U2267 ( .A(n2837), .ZN(n2851) );
  INV_X1 U2269 ( .A(n2329), .ZN(n2507) );
  INV_X4 U2270 ( .A(n2350), .ZN(n2586) );
  XNOR2_X1 U2271 ( .A(n2640), .B(IR_REG_26__SCAN_IN), .ZN(n2652) );
  INV_X1 U2272 ( .A(n2655), .ZN(n3657) );
  INV_X1 U2273 ( .A(n2700), .ZN(n2022) );
  INV_X1 U2274 ( .A(n2700), .ZN(n2023) );
  INV_X1 U2275 ( .A(n2700), .ZN(n2871) );
  NAND2_X4 U2276 ( .A1(n4268), .A2(n2908), .ZN(n2328) );
  AND2_X1 U2278 ( .A1(n4134), .A2(n4135), .ZN(n2144) );
  OR2_X1 U2279 ( .A1(n4365), .A2(n4366), .ZN(n2166) );
  NAND2_X1 U2280 ( .A1(n2129), .A2(n2127), .ZN(n3862) );
  OR2_X1 U2281 ( .A1(n4026), .A2(n2130), .ZN(n2129) );
  OR2_X1 U2282 ( .A1(n4039), .A2(n4047), .ZN(n4037) );
  AOI21_X1 U2283 ( .B1(n4001), .B2(n2506), .A(n2276), .ZN(n3992) );
  NAND2_X1 U2284 ( .A1(n4019), .A2(n2491), .ZN(n4001) );
  NAND2_X1 U2285 ( .A1(n4021), .A2(n4020), .ZN(n4019) );
  OAI21_X1 U2286 ( .B1(n3260), .B2(n2204), .A(n2202), .ZN(n3312) );
  NAND2_X1 U2287 ( .A1(n2112), .A2(n2117), .ZN(n2113) );
  OAI22_X1 U2288 ( .A1(n3210), .A2(n2372), .B1(n3194), .B2(n3675), .ZN(n3184)
         );
  AOI21_X1 U2289 ( .B1(n3617), .B2(n2105), .A(n2104), .ZN(n2103) );
  AND2_X1 U2290 ( .A1(n3548), .A2(n3545), .ZN(n3617) );
  NOR2_X2 U2291 ( .A1(n2963), .A2(n2962), .ZN(n4461) );
  INV_X1 U2292 ( .A(n3678), .ZN(n3112) );
  AND4_X1 U2293 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(n3165)
         );
  AND4_X1 U2294 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), .ZN(n3212)
         );
  NAND3_X1 U2295 ( .A1(n2325), .A2(n2324), .A3(n2323), .ZN(n3678) );
  NAND2_X2 U2296 ( .A1(n2868), .A2(n3069), .ZN(n2837) );
  AND2_X2 U2297 ( .A1(n2682), .A2(n3069), .ZN(n2689) );
  AND2_X2 U2298 ( .A1(n2908), .A2(n2301), .ZN(n2350) );
  XNOR2_X1 U2300 ( .A(n2648), .B(IR_REG_24__SCAN_IN), .ZN(n2901) );
  NAND2_X1 U2301 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U2302 ( .A1(n2647), .A2(IR_REG_31__SCAN_IN), .ZN(n2648) );
  OR2_X1 U2303 ( .A1(n2523), .A2(n2641), .ZN(n2526) );
  AND2_X1 U2304 ( .A1(n2503), .A2(n2289), .ZN(n2523) );
  AND2_X1 U2305 ( .A1(n2036), .A2(n2266), .ZN(n2025) );
  AND4_X1 U2306 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(n2287)
         );
  AND2_X1 U2307 ( .A1(n2289), .A2(n2291), .ZN(n2266) );
  AND2_X1 U2308 ( .A1(n2277), .A2(n2243), .ZN(n2242) );
  NOR2_X1 U2309 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2285)
         );
  NOR2_X1 U2310 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2284)
         );
  NOR2_X1 U2311 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2283)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2286)
         );
  INV_X1 U2313 ( .A(IR_REG_18__SCAN_IN), .ZN(n2289) );
  NOR3_X1 U2314 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_15__SCAN_IN), .ZN(n2288) );
  NOR2_X1 U2315 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2277)
         );
  NOR2_X1 U2316 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2290)
         );
  NAND2_X1 U2317 ( .A1(n2676), .A2(n2675), .ZN(n4415) );
  AND2_X1 U2318 ( .A1(n3947), .A2(n3975), .ZN(n2528) );
  INV_X1 U2319 ( .A(n3385), .ZN(n2238) );
  NAND2_X1 U2320 ( .A1(n2911), .A2(IR_REG_28__SCAN_IN), .ZN(n2309) );
  AND2_X1 U2321 ( .A1(n2307), .A2(n2306), .ZN(n2310) );
  NAND2_X1 U2322 ( .A1(n2305), .A2(n2264), .ZN(n2307) );
  NOR2_X1 U2323 ( .A1(n2641), .A2(IR_REG_27__SCAN_IN), .ZN(n2264) );
  AND3_X1 U2324 ( .A1(n2081), .A2(n2080), .A3(n2061), .ZN(n3756) );
  NOR2_X1 U2325 ( .A1(n2422), .A2(n2211), .ZN(n2210) );
  INV_X1 U2326 ( .A(n2411), .ZN(n2211) );
  AND2_X1 U2327 ( .A1(n2025), .A2(n2141), .ZN(n2111) );
  CLKBUF_X1 U2328 ( .A(n2500), .Z(n2501) );
  OR2_X1 U2329 ( .A1(n2567), .A2(n3410), .ZN(n2576) );
  INV_X1 U2330 ( .A(n2328), .ZN(n2636) );
  NAND2_X1 U2331 ( .A1(n2063), .A2(n2944), .ZN(n2945) );
  NAND2_X1 U2332 ( .A1(n2064), .A2(n3707), .ZN(n2063) );
  INV_X1 U2333 ( .A(n3708), .ZN(n2064) );
  INV_X1 U2334 ( .A(IR_REG_9__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U2335 ( .A1(n2091), .A2(n2090), .ZN(n2218) );
  INV_X1 U2336 ( .A(n4294), .ZN(n2090) );
  NOR2_X1 U2337 ( .A1(n4304), .A2(n4305), .ZN(n4303) );
  INV_X1 U2338 ( .A(n2214), .ZN(n3752) );
  NAND2_X1 U2339 ( .A1(n3768), .A2(n2062), .ZN(n4365) );
  NAND2_X1 U2340 ( .A1(n2189), .A2(n2187), .ZN(n3781) );
  AOI21_X1 U2341 ( .B1(n2192), .B2(n2188), .A(n2051), .ZN(n2187) );
  INV_X1 U2342 ( .A(n2575), .ZN(n2196) );
  AND2_X1 U2343 ( .A1(n2565), .A2(n2055), .ZN(n2198) );
  NAND2_X1 U2344 ( .A1(n2031), .A2(n2046), .ZN(n2179) );
  NOR2_X1 U2345 ( .A1(n2185), .A2(n2184), .ZN(n2183) );
  NAND2_X1 U2346 ( .A1(n2046), .A2(n2181), .ZN(n2180) );
  INV_X1 U2347 ( .A(n2184), .ZN(n2181) );
  OR2_X1 U2348 ( .A1(n4101), .A2(n3400), .ZN(n2440) );
  OR2_X1 U2349 ( .A1(n3042), .A2(n2675), .ZN(n4099) );
  NAND2_X1 U2350 ( .A1(n3833), .A2(n3813), .ZN(n3812) );
  NAND2_X1 U2351 ( .A1(n2526), .A2(n2525), .ZN(n2604) );
  NAND2_X1 U2352 ( .A1(n3765), .A2(n2224), .ZN(n2223) );
  NAND2_X1 U2353 ( .A1(n3743), .A2(n4181), .ZN(n2224) );
  NAND2_X1 U2354 ( .A1(n2131), .A2(n3581), .ZN(n2130) );
  INV_X1 U2355 ( .A(n3638), .ZN(n2135) );
  AND2_X1 U2356 ( .A1(n2758), .A2(n2757), .ZN(n2761) );
  AOI21_X1 U2357 ( .B1(n2250), .B2(n2246), .A(n2780), .ZN(n2245) );
  NAND2_X1 U2358 ( .A1(n2054), .A2(n2250), .ZN(n2247) );
  INV_X1 U2359 ( .A(n2251), .ZN(n2250) );
  OAI21_X1 U2360 ( .B1(n2774), .B2(n2252), .A(n3418), .ZN(n2251) );
  OR2_X1 U2361 ( .A1(n2685), .A2(n4269), .ZN(n2868) );
  AND2_X1 U2362 ( .A1(n2226), .A2(n2225), .ZN(n3745) );
  NAND2_X1 U2363 ( .A1(n4270), .A2(REG1_REG_9__SCAN_IN), .ZN(n2225) );
  NOR2_X1 U2364 ( .A1(n3634), .A2(n2134), .ZN(n2133) );
  INV_X1 U2365 ( .A(n2045), .ZN(n2119) );
  NAND2_X1 U2366 ( .A1(n2106), .A2(n3539), .ZN(n3072) );
  NOR2_X1 U2367 ( .A1(n3538), .A2(n2107), .ZN(n2106) );
  INV_X1 U2368 ( .A(n2609), .ZN(n2107) );
  AND2_X1 U2369 ( .A1(n2786), .A2(n3975), .ZN(n2150) );
  OR2_X1 U2370 ( .A1(n4023), .A2(n4029), .ZN(n4009) );
  NAND2_X1 U2371 ( .A1(n3183), .A2(n2383), .ZN(n3201) );
  AND2_X1 U2372 ( .A1(n2036), .A2(n2289), .ZN(n2265) );
  AOI21_X1 U2373 ( .B1(n2241), .B2(n2236), .A(n2030), .ZN(n2235) );
  INV_X1 U2374 ( .A(n2703), .ZN(n2705) );
  XNOR2_X1 U2375 ( .A(n2701), .B(n2837), .ZN(n2704) );
  OAI22_X1 U2376 ( .A1(n3112), .A2(n2700), .B1(n2850), .B2(n2702), .ZN(n2701)
         );
  NAND2_X1 U2377 ( .A1(n3482), .A2(n2256), .ZN(n2254) );
  NAND2_X1 U2378 ( .A1(n2258), .A2(n2257), .ZN(n2256) );
  INV_X1 U2379 ( .A(n3483), .ZN(n2257) );
  INV_X1 U2380 ( .A(n3484), .ZN(n2258) );
  NAND2_X1 U2381 ( .A1(n2228), .A2(n2234), .ZN(n2227) );
  INV_X1 U2382 ( .A(n3188), .ZN(n2234) );
  INV_X1 U2383 ( .A(n3189), .ZN(n2228) );
  INV_X1 U2384 ( .A(n2232), .ZN(n2229) );
  OR2_X1 U2385 ( .A1(n2310), .A2(n2263), .ZN(n2260) );
  NAND2_X1 U2386 ( .A1(n2259), .A2(n2310), .ZN(n2261) );
  INV_X1 U2387 ( .A(DATAI_1_), .ZN(n2263) );
  AOI22_X1 U2388 ( .A1(n2691), .A2(n2022), .B1(n2689), .B2(n2690), .ZN(n2696)
         );
  NAND2_X1 U2389 ( .A1(n3444), .A2(n2240), .ZN(n2239) );
  NAND2_X1 U2390 ( .A1(n2310), .A2(n2309), .ZN(n2357) );
  AND2_X1 U2391 ( .A1(n2697), .A2(n2698), .ZN(n2699) );
  NAND2_X1 U2392 ( .A1(n2350), .A2(REG2_REG_0__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2393 ( .A1(n3693), .A2(n2943), .ZN(n3707) );
  NAND2_X1 U2394 ( .A1(n2947), .A2(n2946), .ZN(n2949) );
  XNOR2_X1 U2395 ( .A(n2949), .B(n4273), .ZN(n3721) );
  NOR2_X1 U2396 ( .A1(n2995), .A2(n2168), .ZN(n2975) );
  NOR2_X1 U2397 ( .A1(n2987), .A2(n3168), .ZN(n2168) );
  OR2_X1 U2398 ( .A1(n3006), .A2(n3007), .ZN(n2086) );
  NAND2_X1 U2399 ( .A1(n2996), .A2(n2152), .ZN(n2998) );
  NAND2_X1 U2400 ( .A1(n4271), .A2(REG2_REG_7__SCAN_IN), .ZN(n2152) );
  OR2_X1 U2401 ( .A1(n3011), .A2(n3010), .ZN(n2226) );
  XNOR2_X1 U2402 ( .A(n3745), .B(n4467), .ZN(n4457) );
  NOR2_X1 U2403 ( .A1(n4457), .A2(n4458), .ZN(n4456) );
  OR2_X1 U2404 ( .A1(n4303), .A2(n3750), .ZN(n2089) );
  NAND2_X1 U2405 ( .A1(n2089), .A2(n2088), .ZN(n2216) );
  INV_X1 U2406 ( .A(n4314), .ZN(n2088) );
  XNOR2_X1 U2407 ( .A(n2214), .B(n4332), .ZN(n4325) );
  OR2_X1 U2408 ( .A1(n4343), .A2(n4344), .ZN(n2171) );
  OR2_X1 U2409 ( .A1(n4325), .A2(n2083), .ZN(n2080) );
  OR2_X1 U2410 ( .A1(n4338), .A2(n4326), .ZN(n2083) );
  INV_X1 U2411 ( .A(n4338), .ZN(n2084) );
  OR2_X1 U2412 ( .A1(n4325), .A2(n4326), .ZN(n2085) );
  XNOR2_X1 U2413 ( .A(n3756), .B(n2490), .ZN(n4355) );
  NAND2_X1 U2414 ( .A1(n4355), .A2(n4354), .ZN(n4353) );
  INV_X1 U2415 ( .A(n3794), .ZN(n3797) );
  NAND2_X1 U2416 ( .A1(n3797), .A2(n3796), .ZN(n4127) );
  OR2_X1 U2417 ( .A1(n2576), .A2(n3496), .ZN(n2594) );
  AOI21_X1 U2418 ( .B1(n2195), .B2(n2193), .A(n2041), .ZN(n2192) );
  INV_X1 U2419 ( .A(n2198), .ZN(n2193) );
  NOR2_X1 U2420 ( .A1(n3805), .A2(n3810), .ZN(n3804) );
  OR2_X1 U2421 ( .A1(n2552), .A2(n2551), .ZN(n2560) );
  AND4_X1 U2422 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n3908)
         );
  INV_X1 U2423 ( .A(n2280), .ZN(n2186) );
  NOR2_X1 U2424 ( .A1(n2529), .A2(n2528), .ZN(n2184) );
  AOI22_X1 U2425 ( .A1(n4048), .A2(n2478), .B1(n4042), .B2(n4053), .ZN(n4021)
         );
  INV_X1 U2426 ( .A(n2206), .ZN(n2204) );
  AOI21_X1 U2427 ( .B1(n2206), .B2(n2203), .A(n2039), .ZN(n2202) );
  OAI22_X1 U2428 ( .A1(n2422), .A2(n2209), .B1(n3288), .B2(n3332), .ZN(n2208)
         );
  NAND2_X1 U2429 ( .A1(n2411), .A2(n2412), .ZN(n2209) );
  NOR2_X1 U2430 ( .A1(n2208), .A2(n4098), .ZN(n2206) );
  NAND2_X1 U2431 ( .A1(n3260), .A2(n2210), .ZN(n2207) );
  OR2_X1 U2432 ( .A1(n2423), .A2(n3331), .ZN(n2430) );
  NAND2_X1 U2433 ( .A1(n2095), .A2(n3536), .ZN(n3261) );
  NAND2_X1 U2434 ( .A1(n3197), .A2(n3557), .ZN(n2095) );
  OR2_X1 U2435 ( .A1(n2386), .A2(n2385), .ZN(n2399) );
  OR2_X1 U2436 ( .A1(n4278), .A2(n2848), .ZN(n4081) );
  INV_X1 U2437 ( .A(n4083), .ZN(n4109) );
  NAND2_X1 U2438 ( .A1(n2892), .A2(n4394), .ZN(n2957) );
  NAND2_X1 U2439 ( .A1(n2350), .A2(REG2_REG_1__SCAN_IN), .ZN(n2173) );
  NAND2_X1 U2440 ( .A1(n4278), .A2(n2959), .ZN(n4100) );
  INV_X1 U2441 ( .A(n2690), .ZN(n3043) );
  OR2_X1 U2442 ( .A1(n3812), .A2(n3779), .ZN(n3794) );
  AND2_X1 U2443 ( .A1(n4156), .A2(n2056), .ZN(n3833) );
  INV_X1 U2444 ( .A(n3970), .ZN(n3975) );
  INV_X1 U2445 ( .A(n3993), .ZN(n2786) );
  NAND2_X1 U2446 ( .A1(n4010), .A2(n2150), .ZN(n3978) );
  NAND3_X1 U2447 ( .A1(n2140), .A2(n2111), .A3(n2038), .ZN(n2298) );
  INV_X1 U2448 ( .A(n2293), .ZN(n2212) );
  AND2_X1 U2449 ( .A1(n2295), .A2(n2294), .ZN(n2213) );
  INV_X1 U2450 ( .A(IR_REG_29__SCAN_IN), .ZN(n2299) );
  XNOR2_X1 U2451 ( .A(n2297), .B(n3347), .ZN(n2302) );
  NAND2_X1 U2452 ( .A1(n3346), .A2(IR_REG_31__SCAN_IN), .ZN(n2297) );
  XNOR2_X1 U2453 ( .A(n2300), .B(n2299), .ZN(n2301) );
  NAND2_X1 U2454 ( .A1(n2298), .A2(IR_REG_31__SCAN_IN), .ZN(n2300) );
  NAND2_X1 U2455 ( .A1(n2305), .A2(IR_REG_31__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U2456 ( .A1(n2025), .A2(n2138), .ZN(n2137) );
  AND2_X1 U2457 ( .A1(n2139), .A2(n2294), .ZN(n2138) );
  INV_X1 U2458 ( .A(IR_REG_23__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U2459 ( .A1(n2646), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  XNOR2_X1 U2460 ( .A(n2654), .B(n2653), .ZN(n2958) );
  INV_X1 U2461 ( .A(IR_REG_20__SCAN_IN), .ZN(n2605) );
  AND2_X1 U2462 ( .A1(n2457), .A2(n2456), .ZN(n3751) );
  NOR2_X2 U2463 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2326)
         );
  AND2_X1 U2464 ( .A1(n4409), .A2(n2164), .ZN(n2163) );
  INV_X1 U2465 ( .A(n4012), .ZN(n4005) );
  INV_X1 U2466 ( .A(n4105), .ZN(n3332) );
  NAND2_X1 U2467 ( .A1(n2879), .A2(n4278), .ZN(n3513) );
  NAND2_X1 U2468 ( .A1(n2574), .A2(n2573), .ZN(n3867) );
  AOI21_X1 U2469 ( .B1(n4276), .B2(REG2_REG_1__SCAN_IN), .A(n2158), .ZN(n2157)
         );
  INV_X1 U2470 ( .A(n3704), .ZN(n2158) );
  XNOR2_X1 U2471 ( .A(n2975), .B(n2167), .ZN(n3047) );
  NAND2_X1 U2472 ( .A1(n4309), .A2(n3734), .ZN(n4320) );
  AND2_X1 U2473 ( .A1(n3687), .A2(n4278), .ZN(n4333) );
  INV_X1 U2474 ( .A(n2222), .ZN(n2221) );
  AOI21_X1 U2475 ( .B1(n2223), .B2(n4362), .A(n4455), .ZN(n2222) );
  AOI21_X1 U2476 ( .B1(n4461), .B2(ADDR_REG_18__SCAN_IN), .A(n4363), .ZN(n2220) );
  INV_X1 U2477 ( .A(n2166), .ZN(n4364) );
  AND2_X1 U2478 ( .A1(n2166), .A2(n2165), .ZN(n3772) );
  NAND2_X1 U2479 ( .A1(n3770), .A2(REG2_REG_18__SCAN_IN), .ZN(n2165) );
  AND2_X1 U2480 ( .A1(n3687), .A2(n3664), .ZN(n4463) );
  NOR2_X1 U2481 ( .A1(n2068), .A2(n2070), .ZN(n2067) );
  NOR2_X1 U2482 ( .A1(n3766), .A2(n2079), .ZN(n2070) );
  INV_X1 U2483 ( .A(n2071), .ZN(n2068) );
  INV_X1 U2484 ( .A(n3508), .ZN(n2252) );
  INV_X1 U2485 ( .A(IR_REG_28__SCAN_IN), .ZN(n2308) );
  INV_X1 U2486 ( .A(IR_REG_26__SCAN_IN), .ZN(n2304) );
  INV_X1 U2487 ( .A(IR_REG_21__SCAN_IN), .ZN(n2267) );
  AND2_X1 U2488 ( .A1(n2309), .A2(n2262), .ZN(n2259) );
  OAI21_X1 U2489 ( .B1(n3362), .B2(n3360), .A(n3359), .ZN(n2253) );
  NOR2_X1 U2490 ( .A1(n3863), .A2(n2108), .ZN(n3623) );
  NAND2_X1 U2491 ( .A1(n4027), .A2(n2109), .ZN(n2108) );
  INV_X1 U2492 ( .A(IR_REG_27__SCAN_IN), .ZN(n4535) );
  INV_X1 U2493 ( .A(IR_REG_6__SCAN_IN), .ZN(n4544) );
  AND2_X1 U2494 ( .A1(n2218), .A2(n2217), .ZN(n3749) );
  NAND2_X1 U2495 ( .A1(n3748), .A2(REG1_REG_11__SCAN_IN), .ZN(n2217) );
  NAND2_X1 U2496 ( .A1(n2216), .A2(n2215), .ZN(n2214) );
  NAND2_X1 U2497 ( .A1(n3751), .A2(REG1_REG_13__SCAN_IN), .ZN(n2215) );
  AND2_X1 U2498 ( .A1(n2171), .A2(n2170), .ZN(n3737) );
  NAND2_X1 U2499 ( .A1(n3755), .A2(REG2_REG_15__SCAN_IN), .ZN(n2170) );
  NOR2_X1 U2500 ( .A1(n2590), .A2(n2191), .ZN(n2190) );
  INV_X1 U2501 ( .A(n2192), .ZN(n2191) );
  NOR2_X1 U2502 ( .A1(n2195), .A2(n2590), .ZN(n2188) );
  INV_X1 U2503 ( .A(n2128), .ZN(n2127) );
  OAI21_X1 U2504 ( .B1(n2047), .B2(n2130), .A(n3641), .ZN(n2128) );
  NAND2_X1 U2505 ( .A1(n2135), .A2(n2132), .ZN(n2131) );
  NOR2_X1 U2506 ( .A1(n2467), .A2(n3512), .ZN(n2479) );
  INV_X1 U2507 ( .A(n2210), .ZN(n2203) );
  NOR2_X1 U2508 ( .A1(n2399), .A2(n3002), .ZN(n2413) );
  AOI21_X1 U2509 ( .B1(n2117), .B2(n2116), .A(n2115), .ZN(n2114) );
  INV_X1 U2510 ( .A(n3556), .ZN(n2116) );
  INV_X1 U2511 ( .A(n3553), .ZN(n2115) );
  NOR2_X1 U2512 ( .A1(n2348), .A2(n2986), .ZN(n2363) );
  INV_X1 U2513 ( .A(n3543), .ZN(n2105) );
  INV_X1 U2514 ( .A(n3548), .ZN(n2104) );
  NAND2_X1 U2515 ( .A1(n3680), .A2(n2683), .ZN(n3539) );
  NOR2_X1 U2516 ( .A1(n2814), .A2(n2147), .ZN(n2146) );
  AND2_X1 U2517 ( .A1(n2150), .A2(n3952), .ZN(n2149) );
  INV_X1 U2518 ( .A(n3115), .ZN(n3091) );
  NAND2_X1 U2519 ( .A1(n3092), .A2(n3091), .ZN(n3130) );
  NOR2_X1 U2520 ( .A1(n2293), .A2(IR_REG_17__SCAN_IN), .ZN(n2139) );
  NAND2_X1 U2521 ( .A1(n2254), .A2(n2052), .ZN(n3377) );
  NAND2_X1 U2522 ( .A1(n3484), .A2(n3483), .ZN(n2255) );
  OR2_X1 U2523 ( .A1(n2684), .A2(n2855), .ZN(n2688) );
  AND2_X1 U2524 ( .A1(n2762), .A2(n2761), .ZN(n3394) );
  NAND2_X1 U2525 ( .A1(n2250), .A2(n2249), .ZN(n2248) );
  AND2_X1 U2526 ( .A1(n2247), .A2(n2245), .ZN(n2244) );
  INV_X1 U2527 ( .A(n3360), .ZN(n2249) );
  INV_X1 U2528 ( .A(n2867), .ZN(n2882) );
  AND2_X1 U2529 ( .A1(n2600), .A2(n2599), .ZN(n3790) );
  OR2_X1 U2530 ( .A1(n2328), .A2(n3152), .ZN(n2342) );
  XNOR2_X1 U2531 ( .A(n2967), .B(n3029), .ZN(n3024) );
  INV_X1 U2532 ( .A(n2407), .ZN(n2409) );
  XNOR2_X1 U2533 ( .A(n3729), .B(n4467), .ZN(n4464) );
  NAND2_X1 U2534 ( .A1(n3727), .A2(n2151), .ZN(n3729) );
  NAND2_X1 U2535 ( .A1(n4270), .A2(REG2_REG_9__SCAN_IN), .ZN(n2151) );
  NAND2_X1 U2536 ( .A1(n4464), .A2(REG2_REG_10__SCAN_IN), .ZN(n4462) );
  OR2_X1 U2537 ( .A1(n4456), .A2(n3747), .ZN(n2091) );
  XNOR2_X1 U2538 ( .A(n3749), .B(n4405), .ZN(n4304) );
  NAND2_X1 U2539 ( .A1(n4298), .A2(n3731), .ZN(n3733) );
  XNOR2_X1 U2540 ( .A(n3737), .B(n2490), .ZN(n4352) );
  NAND2_X1 U2541 ( .A1(n3739), .A2(n3740), .ZN(n3768) );
  NAND2_X1 U2542 ( .A1(n4353), .A2(n3757), .ZN(n3758) );
  INV_X1 U2543 ( .A(n2079), .ZN(n2075) );
  NAND2_X1 U2544 ( .A1(n4362), .A2(n2075), .ZN(n2074) );
  NOR2_X1 U2545 ( .A1(n4127), .A2(n4130), .ZN(n4126) );
  AND3_X1 U2546 ( .A1(n2556), .A2(n2555), .A3(n2554), .ZN(n3865) );
  AOI21_X1 U2547 ( .B1(n2178), .B2(n2177), .A(n2176), .ZN(n3903) );
  NOR2_X1 U2548 ( .A1(n2180), .A2(n2029), .ZN(n2177) );
  OAI21_X1 U2549 ( .B1(n2179), .B2(n2029), .A(n2053), .ZN(n2176) );
  NAND2_X1 U2550 ( .A1(n2126), .A2(n2131), .ZN(n3922) );
  NAND2_X1 U2551 ( .A1(n4026), .A2(n2047), .ZN(n2126) );
  OR2_X1 U2552 ( .A1(n2516), .A2(n4598), .ZN(n2530) );
  NAND2_X1 U2553 ( .A1(n4026), .A2(n2133), .ZN(n3941) );
  OR2_X1 U2554 ( .A1(n2508), .A2(n3487), .ZN(n2516) );
  NAND2_X1 U2555 ( .A1(n4026), .A2(n3530), .ZN(n4003) );
  OR2_X1 U2556 ( .A1(n2459), .A2(n2458), .ZN(n2467) );
  AOI21_X1 U2557 ( .B1(n2024), .B2(n2028), .A(n2049), .ZN(n2200) );
  INV_X1 U2558 ( .A(n3518), .ZN(n4042) );
  OAI21_X1 U2559 ( .B1(n3261), .B2(n3565), .A(n3558), .ZN(n3283) );
  INV_X1 U2560 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3002) );
  INV_X1 U2561 ( .A(n4081), .ZN(n4106) );
  INV_X1 U2562 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2385) );
  INV_X1 U2563 ( .A(n3242), .ZN(n3179) );
  NAND2_X1 U2564 ( .A1(n2113), .A2(n2114), .ZN(n3175) );
  OAI21_X1 U2565 ( .B1(n3163), .B2(n2119), .A(n3556), .ZN(n3211) );
  INV_X1 U2566 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2986) );
  NAND2_X1 U2567 ( .A1(n3092), .A2(n2136), .ZN(n3169) );
  AND2_X1 U2568 ( .A1(n3131), .A2(n3091), .ZN(n2136) );
  NAND2_X1 U2569 ( .A1(n2102), .A2(n2103), .ZN(n3124) );
  NAND2_X1 U2570 ( .A1(n3086), .A2(n3617), .ZN(n3085) );
  NAND2_X1 U2571 ( .A1(n3074), .A2(n3543), .ZN(n3086) );
  NAND2_X1 U2572 ( .A1(n3539), .A2(n2609), .ZN(n2110) );
  INV_X1 U2573 ( .A(n4099), .ZN(n4129) );
  AOI21_X1 U2574 ( .B1(n2125), .B2(n4083), .A(n2124), .ZN(n3353) );
  OR2_X1 U2575 ( .A1(n2639), .A2(n2638), .ZN(n2124) );
  XNOR2_X1 U2576 ( .A(n2627), .B(n3780), .ZN(n2125) );
  NAND2_X1 U2577 ( .A1(n4156), .A2(n2032), .ZN(n3852) );
  NAND2_X1 U2578 ( .A1(n4156), .A2(n2146), .ZN(n3870) );
  NAND2_X1 U2579 ( .A1(n4156), .A2(n3893), .ZN(n3892) );
  AND2_X1 U2580 ( .A1(n3928), .A2(n3913), .ZN(n4156) );
  AND2_X1 U2581 ( .A1(n4010), .A2(n2148), .ZN(n3928) );
  AND2_X1 U2582 ( .A1(n2149), .A2(n3930), .ZN(n2148) );
  NAND2_X1 U2583 ( .A1(n4010), .A2(n2149), .ZN(n3951) );
  NOR2_X1 U2584 ( .A1(n4087), .A2(n4061), .ZN(n4062) );
  OR2_X1 U2585 ( .A1(n4086), .A2(n4077), .ZN(n4087) );
  OR2_X1 U2586 ( .A1(n4113), .A2(n3313), .ZN(n4086) );
  INV_X1 U2587 ( .A(n3400), .ZN(n3313) );
  NAND2_X1 U2588 ( .A1(n4111), .A2(n4110), .ZN(n4113) );
  INV_X1 U2589 ( .A(n3334), .ZN(n4110) );
  NOR2_X1 U2590 ( .A1(n3267), .A2(n3279), .ZN(n3289) );
  AND2_X1 U2591 ( .A1(n3289), .A2(n3288), .ZN(n4111) );
  OR2_X1 U2592 ( .A1(n3203), .A2(n3202), .ZN(n3267) );
  INV_X1 U2593 ( .A(n3194), .ZN(n3221) );
  NOR2_X1 U2594 ( .A1(n3169), .A2(n3170), .ZN(n3222) );
  AND2_X1 U2595 ( .A1(n3222), .A2(n3221), .ZN(n3219) );
  NOR2_X1 U2596 ( .A1(n3078), .A2(n3476), .ZN(n3092) );
  INV_X1 U2597 ( .A(n4415), .ZN(n4443) );
  AND3_X1 U2598 ( .A1(n2670), .A2(n2669), .A3(n2668), .ZN(n2677) );
  INV_X1 U2599 ( .A(n2957), .ZN(n3065) );
  XNOR2_X1 U2600 ( .A(n2607), .B(n2291), .ZN(n2685) );
  INV_X1 U2601 ( .A(IR_REG_7__SCAN_IN), .ZN(n2380) );
  INV_X1 U2602 ( .A(IR_REG_3__SCAN_IN), .ZN(n4545) );
  INV_X1 U2603 ( .A(n2282), .ZN(n2327) );
  NAND2_X1 U2604 ( .A1(n2233), .A2(n2232), .ZN(n3237) );
  INV_X1 U2605 ( .A(n2839), .ZN(n3813) );
  AND4_X1 U2606 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n3307)
         );
  NAND2_X1 U2607 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U2608 ( .A1(n2254), .A2(n2255), .ZN(n3376) );
  INV_X1 U2609 ( .A(n3236), .ZN(n2231) );
  AOI21_X1 U2610 ( .B1(n2229), .B2(n3236), .A(n2040), .ZN(n2230) );
  NAND2_X1 U2611 ( .A1(n3444), .A2(n3448), .ZN(n3389) );
  AND2_X1 U2612 ( .A1(n2576), .A2(n2568), .ZN(n3855) );
  AOI21_X1 U2613 ( .B1(n2779), .B2(n2778), .A(n2780), .ZN(n3418) );
  INV_X1 U2614 ( .A(n3675), .ZN(n3239) );
  INV_X1 U2615 ( .A(n2724), .ZN(n3170) );
  AND4_X1 U2616 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n3974)
         );
  INV_X1 U2617 ( .A(n2814), .ZN(n3871) );
  AND4_X1 U2618 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3276)
         );
  NAND2_X1 U2619 ( .A1(n2357), .A2(DATAI_0_), .ZN(n2316) );
  INV_X1 U2620 ( .A(n3517), .ZN(n3497) );
  NAND2_X1 U2621 ( .A1(n2239), .A2(n3385), .ZN(n3465) );
  AND4_X1 U2622 ( .A1(n2436), .A2(n2435), .A3(n2434), .A4(n2433), .ZN(n4101)
         );
  AND4_X1 U2623 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n3987)
         );
  AND4_X1 U2624 ( .A1(n2379), .A2(n2378), .A3(n2377), .A4(n2376), .ZN(n3213)
         );
  AND2_X1 U2625 ( .A1(n2594), .A2(n2577), .ZN(n3837) );
  AND2_X1 U2626 ( .A1(n2878), .A2(n3015), .ZN(n3521) );
  INV_X1 U2627 ( .A(n3499), .ZN(n3515) );
  AND2_X1 U2628 ( .A1(n2867), .A2(n2849), .ZN(n3510) );
  NAND2_X1 U2629 ( .A1(n2589), .A2(n2588), .ZN(n3830) );
  INV_X1 U2630 ( .A(n3803), .ZN(n3849) );
  INV_X1 U2631 ( .A(n3974), .ZN(n4006) );
  INV_X1 U2632 ( .A(n3987), .ZN(n4030) );
  INV_X1 U2633 ( .A(n4053), .ZN(n3419) );
  INV_X1 U2634 ( .A(n4101), .ZN(n3672) );
  INV_X1 U2635 ( .A(n3276), .ZN(n3264) );
  INV_X1 U2636 ( .A(n3213), .ZN(n3252) );
  INV_X1 U2637 ( .A(n2684), .ZN(n3680) );
  NAND2_X1 U2638 ( .A1(n2329), .A2(REG1_REG_0__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2639 ( .A1(n2892), .A2(n2891), .ZN(n3681) );
  AND2_X1 U2640 ( .A1(n2961), .A2(n2962), .ZN(n3687) );
  NAND2_X1 U2641 ( .A1(n3695), .A2(n3694), .ZN(n3693) );
  NAND2_X1 U2642 ( .A1(n3712), .A2(n3711), .ZN(n3710) );
  XNOR2_X1 U2643 ( .A(n2945), .B(n3029), .ZN(n3023) );
  OAI21_X1 U2644 ( .B1(n3721), .B2(n2948), .A(n2950), .ZN(n2990) );
  AND2_X1 U2645 ( .A1(n2984), .A2(n2169), .ZN(n2995) );
  INV_X1 U2646 ( .A(n2974), .ZN(n2169) );
  NAND2_X1 U2647 ( .A1(n2980), .A2(n2153), .ZN(n2996) );
  INV_X1 U2648 ( .A(n2978), .ZN(n2153) );
  XNOR2_X1 U2649 ( .A(n2998), .B(n4408), .ZN(n4290) );
  NAND2_X1 U2650 ( .A1(n2087), .A2(n2086), .ZN(n4285) );
  INV_X1 U2651 ( .A(n3008), .ZN(n2087) );
  NAND2_X1 U2652 ( .A1(n3001), .A2(n3000), .ZN(n3727) );
  NOR2_X1 U2653 ( .A1(n2033), .A2(n3008), .ZN(n3011) );
  INV_X1 U2654 ( .A(n2218), .ZN(n4293) );
  INV_X1 U2655 ( .A(n2091), .ZN(n4295) );
  XNOR2_X1 U2656 ( .A(n3733), .B(n4405), .ZN(n4310) );
  NAND2_X1 U2657 ( .A1(n4310), .A2(REG2_REG_12__SCAN_IN), .ZN(n4309) );
  INV_X1 U2658 ( .A(n2089), .ZN(n4315) );
  INV_X1 U2659 ( .A(n2216), .ZN(n4313) );
  NOR2_X1 U2660 ( .A1(n4328), .A2(n3736), .ZN(n4343) );
  INV_X1 U2661 ( .A(n2171), .ZN(n4342) );
  AND2_X1 U2662 ( .A1(n2082), .A2(n2085), .ZN(n4339) );
  NAND2_X1 U2663 ( .A1(n2081), .A2(n2080), .ZN(n4337) );
  INV_X1 U2664 ( .A(n3753), .ZN(n2082) );
  NAND2_X1 U2665 ( .A1(n2073), .A2(n2072), .ZN(n2071) );
  NAND2_X1 U2666 ( .A1(n3766), .A2(n2075), .ZN(n2072) );
  NAND2_X1 U2667 ( .A1(n2076), .A2(n2074), .ZN(n2073) );
  INV_X1 U2668 ( .A(n3766), .ZN(n2076) );
  NAND2_X1 U2669 ( .A1(n2078), .A2(n3766), .ZN(n2077) );
  INV_X1 U2670 ( .A(n4362), .ZN(n2078) );
  OAI21_X1 U2671 ( .B1(n2566), .B2(n2194), .A(n2192), .ZN(n3811) );
  NAND2_X1 U2672 ( .A1(n2197), .A2(n2575), .ZN(n3821) );
  NAND2_X1 U2673 ( .A1(n2566), .A2(n2198), .ZN(n2197) );
  NAND2_X1 U2674 ( .A1(n2566), .A2(n2565), .ZN(n3842) );
  OAI21_X1 U2675 ( .B1(n3990), .B2(n2180), .A(n2179), .ZN(n3920) );
  INV_X1 U2676 ( .A(n2182), .ZN(n3939) );
  AOI21_X1 U2677 ( .B1(n3990), .B2(n2185), .A(n2184), .ZN(n2182) );
  NAND2_X1 U2678 ( .A1(n2201), .A2(n2024), .ZN(n4058) );
  AND2_X1 U2679 ( .A1(n2201), .A2(n2048), .ZN(n4060) );
  OR2_X1 U2680 ( .A1(n4071), .A2(n2028), .ZN(n2201) );
  NAND2_X1 U2681 ( .A1(n2207), .A2(n2205), .ZN(n4096) );
  INV_X1 U2682 ( .A(n2208), .ZN(n2205) );
  INV_X1 U2683 ( .A(n4035), .ZN(n4068) );
  NAND2_X1 U2684 ( .A1(n3071), .A2(n2175), .ZN(n3076) );
  OR2_X1 U2685 ( .A1(n2684), .A2(n4081), .ZN(n2175) );
  OR2_X1 U2686 ( .A1(n2957), .A2(n2880), .ZN(n4370) );
  NAND2_X1 U2687 ( .A1(n3044), .A2(n2174), .ZN(n4383) );
  OR2_X1 U2688 ( .A1(n2684), .A2(n4100), .ZN(n2174) );
  INV_X1 U2689 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2120) );
  NAND2_X1 U2690 ( .A1(n2678), .A2(n4454), .ZN(n2121) );
  NAND2_X1 U2691 ( .A1(n2145), .A2(n2144), .ZN(n4214) );
  OR2_X1 U2692 ( .A1(n4133), .A2(n4415), .ZN(n2145) );
  NAND2_X1 U2693 ( .A1(n3353), .A2(n2122), .ZN(n2678) );
  NAND2_X1 U2694 ( .A1(n2123), .A2(n4432), .ZN(n2122) );
  INV_X1 U2695 ( .A(n3358), .ZN(n2123) );
  OAI21_X1 U2696 ( .B1(n2674), .B2(n2853), .A(n3794), .ZN(n3350) );
  AND2_X1 U2697 ( .A1(n4010), .A2(n2786), .ZN(n3976) );
  AND2_X2 U2698 ( .A1(n3067), .A2(n2677), .ZN(n4446) );
  NAND2_X1 U2699 ( .A1(n3065), .A2(n2914), .ZN(n4393) );
  INV_X1 U2700 ( .A(n2298), .ZN(n2296) );
  INV_X1 U2701 ( .A(IR_REG_30__SCAN_IN), .ZN(n3347) );
  XNOR2_X1 U2702 ( .A(n2631), .B(IR_REG_28__SCAN_IN), .ZN(n4278) );
  OR2_X1 U2703 ( .A1(n2303), .A2(n2641), .ZN(n2640) );
  AND2_X1 U2704 ( .A1(n2645), .A2(n2644), .ZN(n2905) );
  AOI21_X1 U2705 ( .B1(n2643), .B2(IR_REG_25__SCAN_IN), .A(n2642), .ZN(n2645)
         );
  AND2_X1 U2706 ( .A1(n2641), .A2(n2294), .ZN(n2642) );
  AND2_X1 U2707 ( .A1(n2958), .A2(STATE_REG_SCAN_IN), .ZN(n4394) );
  INV_X1 U2708 ( .A(n2685), .ZN(n3667) );
  AND2_X1 U2709 ( .A1(n2527), .A2(n2604), .ZN(n4269) );
  OAI21_X1 U2710 ( .B1(n2094), .B2(n2326), .A(n2093), .ZN(n2092) );
  NAND2_X1 U2711 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2094)
         );
  NAND2_X1 U2712 ( .A1(n2641), .A2(n2281), .ZN(n2093) );
  NAND2_X1 U2713 ( .A1(n2641), .A2(IR_REG_1__SCAN_IN), .ZN(n2154) );
  NAND2_X1 U2714 ( .A1(n2163), .A2(IR_REG_31__SCAN_IN), .ZN(n2162) );
  NAND2_X1 U2715 ( .A1(n2317), .A2(IR_REG_1__SCAN_IN), .ZN(n2155) );
  INV_X1 U2716 ( .A(n2219), .ZN(n4369) );
  OAI21_X1 U2717 ( .B1(n4361), .B2(n2221), .A(n2220), .ZN(n2219) );
  NAND2_X1 U2718 ( .A1(n2071), .A2(n2077), .ZN(n2069) );
  NAND2_X1 U2719 ( .A1(n2143), .A2(n2142), .ZN(U3547) );
  NAND2_X1 U2720 ( .A1(n4452), .A2(REG1_REG_29__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2721 ( .A1(n4214), .A2(n4454), .ZN(n2143) );
  OAI211_X1 U2722 ( .C1(n2309), .C2(n2263), .A(n2261), .B(n2260), .ZN(n2311)
         );
  AND2_X1 U2723 ( .A1(n4059), .A2(n2048), .ZN(n2024) );
  OR2_X1 U2724 ( .A1(n2253), .A2(n2774), .ZN(n3415) );
  AND2_X1 U2725 ( .A1(n2042), .A2(n2140), .ZN(n2026) );
  AOI21_X1 U2726 ( .B1(n2119), .B2(n3556), .A(n2118), .ZN(n2117) );
  AND2_X1 U2727 ( .A1(n2121), .A2(n2060), .ZN(n2027) );
  AND2_X1 U2728 ( .A1(n3613), .A2(n4088), .ZN(n2028) );
  AND2_X1 U2729 ( .A1(n3945), .A2(n2799), .ZN(n2029) );
  OR2_X1 U2730 ( .A1(n3368), .A2(n3369), .ZN(n2030) );
  OR2_X1 U2731 ( .A1(n2037), .A2(n2183), .ZN(n2031) );
  AND2_X1 U2732 ( .A1(n2146), .A2(n3853), .ZN(n2032) );
  AND2_X1 U2733 ( .A1(n2086), .A2(REG1_REG_8__SCAN_IN), .ZN(n2033) );
  INV_X1 U2734 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2161) );
  AND3_X1 U2735 ( .A1(n2173), .A2(n2172), .A3(n2096), .ZN(n2684) );
  OAI21_X1 U2736 ( .B1(n2357), .B2(n2317), .A(n2316), .ZN(n2690) );
  NAND2_X1 U2737 ( .A1(n2253), .A2(n2774), .ZN(n3416) );
  AND2_X1 U2738 ( .A1(n2239), .A2(n2236), .ZN(n2034) );
  NAND2_X1 U2739 ( .A1(n2503), .A2(n2265), .ZN(n2035) );
  NAND2_X1 U2740 ( .A1(n2140), .A2(n2111), .ZN(n2646) );
  AOI21_X1 U2741 ( .B1(n3405), .B2(n3406), .A(n3408), .ZN(n3491) );
  AND2_X1 U2742 ( .A1(n2290), .A2(n2267), .ZN(n2036) );
  AND2_X1 U2743 ( .A1(n3923), .A2(n3952), .ZN(n2037) );
  NAND2_X1 U2744 ( .A1(n2282), .A2(n2277), .ZN(n2355) );
  NAND2_X1 U2745 ( .A1(n2523), .A2(n2290), .ZN(n2601) );
  INV_X1 U2746 ( .A(n2195), .ZN(n2194) );
  NOR2_X1 U2747 ( .A1(n2583), .A2(n2196), .ZN(n2195) );
  NAND2_X1 U2748 ( .A1(n2684), .A2(n2311), .ZN(n2609) );
  AND2_X1 U2749 ( .A1(n2213), .A2(n2212), .ZN(n2038) );
  INV_X1 U2750 ( .A(IR_REG_2__SCAN_IN), .ZN(n2281) );
  AND2_X1 U2751 ( .A1(n3307), .A2(n4110), .ZN(n2039) );
  INV_X1 U2752 ( .A(IR_REG_17__SCAN_IN), .ZN(n2141) );
  AND2_X1 U2753 ( .A1(n2735), .A2(n2734), .ZN(n2040) );
  NOR2_X1 U2754 ( .A1(n3849), .A2(n2673), .ZN(n2041) );
  AND2_X1 U2755 ( .A1(n2025), .A2(n2139), .ZN(n2042) );
  AND2_X1 U2756 ( .A1(n2114), .A2(n2613), .ZN(n2043) );
  AND2_X1 U2757 ( .A1(n2242), .A2(n2282), .ZN(n2044) );
  NAND2_X1 U2758 ( .A1(n3165), .A2(n3149), .ZN(n3549) );
  INV_X1 U2759 ( .A(IR_REG_1__SCAN_IN), .ZN(n2164) );
  BUF_X1 U2760 ( .A(IR_REG_0__SCAN_IN), .Z(n4409) );
  AND3_X1 U2761 ( .A1(n2242), .A2(n2287), .A3(n2282), .ZN(n2455) );
  INV_X1 U2762 ( .A(n4272), .ZN(n2167) );
  INV_X1 U2763 ( .A(n3732), .ZN(n4405) );
  NAND2_X1 U2764 ( .A1(n3676), .A2(n2724), .ZN(n2045) );
  OR2_X1 U2765 ( .A1(n3923), .A2(n3952), .ZN(n2046) );
  AND2_X1 U2766 ( .A1(n2135), .A2(n2133), .ZN(n2047) );
  INV_X1 U2767 ( .A(IR_REG_5__SCAN_IN), .ZN(n2243) );
  OR2_X1 U2768 ( .A1(n3613), .A2(n4088), .ZN(n2048) );
  INV_X1 U2769 ( .A(n3554), .ZN(n2118) );
  OAI21_X1 U2770 ( .B1(n3260), .B2(n2412), .A(n2411), .ZN(n3287) );
  NAND2_X1 U2771 ( .A1(n3296), .A2(n2754), .ZN(n3326) );
  INV_X1 U2772 ( .A(n3530), .ZN(n2134) );
  AND2_X1 U2773 ( .A1(n3514), .A2(n4052), .ZN(n2049) );
  AND2_X1 U2774 ( .A1(n2207), .A2(n2206), .ZN(n2050) );
  AND2_X1 U2775 ( .A1(n3830), .A2(n2839), .ZN(n2051) );
  AND2_X1 U2776 ( .A1(n3940), .A2(n2623), .ZN(n3639) );
  INV_X1 U2777 ( .A(n3639), .ZN(n2132) );
  AND2_X1 U2778 ( .A1(n2791), .A2(n2255), .ZN(n2052) );
  NAND2_X1 U2779 ( .A1(n3908), .A2(n3930), .ZN(n2053) );
  INV_X1 U2780 ( .A(n2237), .ZN(n2236) );
  OR2_X1 U2781 ( .A1(n3466), .A2(n2238), .ZN(n2237) );
  INV_X1 U2782 ( .A(n2241), .ZN(n2240) );
  NAND2_X1 U2783 ( .A1(n3448), .A2(n2058), .ZN(n2241) );
  AND2_X1 U2784 ( .A1(n2774), .A2(n2252), .ZN(n2054) );
  OR2_X1 U2785 ( .A1(n3867), .A2(n2825), .ZN(n2055) );
  OR2_X1 U2786 ( .A1(n3184), .A2(n3607), .ZN(n3183) );
  INV_X1 U2787 ( .A(n3359), .ZN(n2246) );
  INV_X1 U2788 ( .A(n3835), .ZN(n2673) );
  AND2_X1 U2789 ( .A1(n2032), .A2(n3835), .ZN(n2056) );
  AND2_X1 U2790 ( .A1(n3528), .A2(DATAI_25_), .ZN(n2825) );
  AND2_X1 U2791 ( .A1(n2033), .A2(n2087), .ZN(n2057) );
  NAND2_X1 U2792 ( .A1(n2803), .A2(n2802), .ZN(n2058) );
  AND2_X1 U2793 ( .A1(n3528), .A2(DATAI_21_), .ZN(n2799) );
  NAND2_X1 U2794 ( .A1(n3062), .A2(n3118), .ZN(n2059) );
  INV_X1 U2795 ( .A(n3893), .ZN(n2147) );
  AND2_X2 U2796 ( .A1(n2677), .A2(n2847), .ZN(n4454) );
  INV_X1 U2797 ( .A(n4454), .ZN(n4452) );
  INV_X1 U2798 ( .A(n4438), .ZN(n4432) );
  OR2_X1 U2799 ( .A1(n4454), .A2(n2120), .ZN(n2060) );
  INV_X1 U2800 ( .A(n4357), .ZN(n4455) );
  AND2_X1 U2801 ( .A1(n3687), .A2(n3703), .ZN(n4357) );
  NAND2_X1 U2802 ( .A1(n3755), .A2(REG1_REG_15__SCAN_IN), .ZN(n2061) );
  NAND3_X1 U2803 ( .A1(n2162), .A2(n2155), .A3(n2154), .ZN(n4276) );
  INV_X1 U2804 ( .A(n2160), .ZN(n2262) );
  OR2_X1 U2805 ( .A1(n3769), .A2(REG2_REG_17__SCAN_IN), .ZN(n2062) );
  NAND2_X1 U2806 ( .A1(n2693), .A2(n2691), .ZN(n2694) );
  NAND2_X1 U2807 ( .A1(n2765), .A2(n2764), .ZN(n3362) );
  AOI21_X1 U2808 ( .B1(n3426), .B2(n3427), .A(n3429), .ZN(n3482) );
  NOR2_X1 U2809 ( .A1(n3053), .A2(n3055), .ZN(n3054) );
  AOI21_X1 U2810 ( .B1(n3273), .B2(n3274), .A(n2278), .ZN(n3298) );
  NAND2_X2 U2811 ( .A1(n2689), .A2(n4415), .ZN(n2855) );
  AOI21_X1 U2812 ( .B1(n3491), .B2(n3493), .A(n3492), .ZN(n3339) );
  NAND2_X2 U2813 ( .A1(n3445), .A2(n3446), .ZN(n3444) );
  NAND2_X1 U2814 ( .A1(n2223), .A2(n2067), .ZN(n2066) );
  NOR2_X1 U2815 ( .A1(n2223), .A2(n4362), .ZN(n4361) );
  NAND2_X1 U2816 ( .A1(n3778), .A2(n2065), .ZN(U3259) );
  OAI211_X1 U2817 ( .C1(n2223), .C2(n2069), .A(n2066), .B(n4357), .ZN(n2065)
         );
  AND2_X1 U2818 ( .A1(n3770), .A2(REG1_REG_18__SCAN_IN), .ZN(n2079) );
  NAND2_X1 U2819 ( .A1(n3753), .A2(n2084), .ZN(n2081) );
  INV_X1 U2820 ( .A(n2085), .ZN(n4324) );
  NAND2_X1 U2822 ( .A1(n2908), .A2(REG3_REG_1__SCAN_IN), .ZN(n2099) );
  NAND2_X1 U2823 ( .A1(n2097), .A2(n4268), .ZN(n2096) );
  NAND2_X1 U2824 ( .A1(n2099), .A2(n2098), .ZN(n2097) );
  AND2_X1 U2825 ( .A1(n4268), .A2(n2302), .ZN(n2329) );
  NAND2_X1 U2826 ( .A1(n2302), .A2(REG1_REG_1__SCAN_IN), .ZN(n2098) );
  INV_X1 U2827 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2100) );
  INV_X1 U2828 ( .A(n3074), .ZN(n2101) );
  NAND2_X1 U2829 ( .A1(n2101), .A2(n3617), .ZN(n2102) );
  NAND3_X1 U2830 ( .A1(n2102), .A2(n2103), .A3(n3549), .ZN(n2612) );
  NAND2_X1 U2831 ( .A1(n2110), .A2(n3538), .ZN(n3030) );
  AOI21_X1 U2832 ( .B1(n2110), .B2(n3035), .A(n2272), .ZN(n3063) );
  XNOR2_X1 U2833 ( .A(n2110), .B(n3036), .ZN(n3141) );
  NOR2_X1 U2834 ( .A1(n4387), .A2(n2110), .ZN(n2109) );
  INV_X1 U2835 ( .A(n3163), .ZN(n2112) );
  NAND2_X1 U2836 ( .A1(n2113), .A2(n2043), .ZN(n2614) );
  INV_X1 U2837 ( .A(n2500), .ZN(n2140) );
  NOR2_X1 U2838 ( .A1(n2137), .A2(n2501), .ZN(n2303) );
  NOR2_X2 U2839 ( .A1(n2500), .A2(IR_REG_17__SCAN_IN), .ZN(n2503) );
  OAI21_X1 U2840 ( .B1(n2161), .B2(n2262), .A(n2156), .ZN(n3692) );
  NAND2_X1 U2841 ( .A1(n2262), .A2(n2161), .ZN(n2156) );
  NAND2_X1 U2842 ( .A1(n2159), .A2(n2157), .ZN(n3691) );
  NAND2_X1 U2843 ( .A1(n2160), .A2(n2161), .ZN(n2159) );
  INV_X1 U2844 ( .A(n4276), .ZN(n2160) );
  OAI22_X1 U2845 ( .A1(n4318), .A2(n4320), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3751), .ZN(n3735) );
  OAI22_X1 U2846 ( .A1(n3716), .A2(n2973), .B1(n2972), .B2(n2971), .ZN(n2984)
         );
  XOR2_X1 U2847 ( .A(n4332), .B(n3735), .Z(n4329) );
  NAND2_X1 U2848 ( .A1(n2318), .A2(REG0_REG_1__SCAN_IN), .ZN(n2172) );
  AND2_X1 U2849 ( .A1(n2302), .A2(n2301), .ZN(n2318) );
  NAND4_X1 U2850 ( .A1(n2287), .A2(n2288), .A3(n2282), .A4(n2242), .ZN(n2500)
         );
  AND2_X2 U2851 ( .A1(n2326), .A2(n2281), .ZN(n2282) );
  INV_X1 U2852 ( .A(n3990), .ZN(n2178) );
  NAND2_X1 U2853 ( .A1(n3990), .A2(n2280), .ZN(n3960) );
  NOR2_X1 U2854 ( .A1(n2528), .A2(n2186), .ZN(n2185) );
  NAND2_X1 U2855 ( .A1(n2566), .A2(n2190), .ZN(n2189) );
  NAND2_X1 U2856 ( .A1(n4071), .A2(n2024), .ZN(n2199) );
  NAND2_X1 U2857 ( .A1(n2199), .A2(n2200), .ZN(n4048) );
  INV_X1 U2858 ( .A(n2226), .ZN(n3744) );
  NAND2_X1 U2859 ( .A1(n3187), .A2(n2227), .ZN(n2233) );
  NAND2_X1 U2860 ( .A1(n3189), .A2(n3188), .ZN(n2232) );
  OAI21_X2 U2861 ( .B1(n2233), .B2(n2231), .A(n2230), .ZN(n3246) );
  OAI21_X2 U2862 ( .B1(n3444), .B2(n2237), .A(n2235), .ZN(n3370) );
  OAI21_X1 U2863 ( .B1(n3362), .B2(n2248), .A(n2244), .ZN(n3426) );
  AND2_X2 U2864 ( .A1(n2269), .A2(n2268), .ZN(n3398) );
  NAND2_X1 U2865 ( .A1(n3326), .A2(n3327), .ZN(n2268) );
  OAI21_X1 U2866 ( .B1(n3326), .B2(n3327), .A(n3328), .ZN(n2269) );
  NAND2_X1 U2867 ( .A1(n3298), .A2(n3297), .ZN(n3296) );
  XNOR2_X1 U2868 ( .A(n3781), .B(n3780), .ZN(n3358) );
  XNOR2_X1 U2869 ( .A(n2704), .B(n2705), .ZN(n3474) );
  AND2_X1 U2870 ( .A1(n3123), .A2(n3122), .ZN(n4424) );
  AOI21_X2 U2871 ( .B1(n3398), .B2(n3395), .A(n3394), .ZN(n3456) );
  AND2_X1 U2872 ( .A1(n2715), .A2(n2714), .ZN(n2270) );
  OR2_X1 U2873 ( .A1(n3672), .A2(n3313), .ZN(n2271) );
  AND2_X1 U2874 ( .A1(n3680), .A2(n2311), .ZN(n2272) );
  NAND2_X2 U2875 ( .A1(n3068), .A2(n4370), .ZN(n4372) );
  INV_X1 U2876 ( .A(n4372), .ZN(n4391) );
  AND2_X1 U2877 ( .A1(n2862), .A2(n3510), .ZN(n2273) );
  OR2_X1 U2878 ( .A1(n3350), .A2(n4266), .ZN(n2274) );
  OR2_X1 U2879 ( .A1(n3350), .A2(n4208), .ZN(n2275) );
  AND2_X1 U2880 ( .A1(n4030), .A2(n4005), .ZN(n2276) );
  AND2_X1 U2881 ( .A1(n2747), .A2(n2746), .ZN(n2278) );
  INV_X1 U2882 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2429) );
  INV_X1 U2883 ( .A(IR_REG_22__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U2884 ( .A1(n3370), .A2(n2279), .ZN(n3436) );
  AND2_X1 U2885 ( .A1(n2817), .A2(n2818), .ZN(n2279) );
  INV_X1 U2886 ( .A(n2610), .ZN(n3061) );
  NAND2_X1 U2887 ( .A1(n3546), .A2(n3543), .ZN(n2610) );
  INV_X1 U2888 ( .A(n3913), .ZN(n2548) );
  AND4_X1 U2889 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3514)
         );
  INV_X1 U2890 ( .A(n3923), .ZN(n3971) );
  AND4_X1 U2891 ( .A1(n2535), .A2(n2534), .A3(n2533), .A4(n2532), .ZN(n3923)
         );
  INV_X1 U2892 ( .A(n3925), .ZN(n3891) );
  NAND2_X1 U2893 ( .A1(n2547), .A2(n2546), .ZN(n3925) );
  AND4_X1 U2894 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n4036)
         );
  OR2_X1 U2895 ( .A1(n4006), .A2(n3993), .ZN(n2280) );
  INV_X1 U2896 ( .A(n3613), .ZN(n4055) );
  AND4_X1 U2897 ( .A1(n2448), .A2(n2447), .A3(n2446), .A4(n2445), .ZN(n3613)
         );
  INV_X1 U2898 ( .A(n4409), .ZN(n2317) );
  NAND2_X1 U2899 ( .A1(n3153), .A2(n2728), .ZN(n3187) );
  INV_X1 U2900 ( .A(n3952), .ZN(n3944) );
  NAND2_X1 U2901 ( .A1(n2726), .A2(n2727), .ZN(n2728) );
  AND2_X1 U2902 ( .A1(n2625), .A2(n3822), .ZN(n3582) );
  AND2_X1 U2903 ( .A1(n4072), .A2(n2617), .ZN(n3566) );
  INV_X1 U2904 ( .A(n3476), .ZN(n2702) );
  INV_X1 U2905 ( .A(IR_REG_25__SCAN_IN), .ZN(n2294) );
  INV_X1 U2906 ( .A(n3379), .ZN(n2791) );
  INV_X1 U2907 ( .A(n3582), .ZN(n3647) );
  INV_X1 U2908 ( .A(n2560), .ZN(n2559) );
  NAND2_X1 U2909 ( .A1(n3677), .A2(n3131), .ZN(n3551) );
  AND3_X1 U2910 ( .A1(n4535), .A2(n2308), .A3(n2304), .ZN(n2295) );
  AND2_X1 U2911 ( .A1(n2768), .A2(n2767), .ZN(n2769) );
  INV_X1 U2912 ( .A(n2855), .ZN(n2841) );
  AOI22_X1 U2913 ( .A1(n2690), .A2(n2023), .B1(n2692), .B2(n4409), .ZN(n2695)
         );
  OR3_X1 U2914 ( .A1(n2405), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2407) );
  OR2_X1 U2915 ( .A1(n3830), .A2(n3813), .ZN(n3522) );
  NAND2_X1 U2916 ( .A1(n2559), .A2(REG3_REG_24__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U2917 ( .A1(n3671), .A2(n4029), .ZN(n2491) );
  INV_X1 U2918 ( .A(n3254), .ZN(n3202) );
  OR2_X1 U2919 ( .A1(n2656), .A2(n2848), .ZN(n3064) );
  INV_X1 U2920 ( .A(n3119), .ZN(n2345) );
  INV_X1 U2921 ( .A(n3337), .ZN(n3338) );
  NOR2_X1 U2922 ( .A1(n2530), .A2(n3450), .ZN(n2536) );
  AND2_X1 U2923 ( .A1(n2479), .A2(REG3_REG_16__SCAN_IN), .ZN(n2492) );
  NOR2_X1 U2924 ( .A1(n2430), .A2(n2429), .ZN(n2442) );
  AND2_X1 U2925 ( .A1(n3066), .A2(n2847), .ZN(n2867) );
  OR2_X1 U2926 ( .A1(n3352), .A2(n2328), .ZN(n2600) );
  AND4_X1 U2927 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n3947)
         );
  INV_X1 U2928 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4484) );
  INV_X1 U2929 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3331) );
  INV_X1 U2930 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3512) );
  INV_X1 U2931 ( .A(n4269), .ZN(n3775) );
  AND4_X1 U2932 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n4053)
         );
  AND2_X1 U2933 ( .A1(n2613), .A2(n3537), .ZN(n3607) );
  OR2_X1 U2934 ( .A1(n3995), .A2(n4415), .ZN(n4066) );
  INV_X1 U2935 ( .A(n2914), .ZN(n2846) );
  INV_X1 U2936 ( .A(n3301), .ZN(n3288) );
  INV_X1 U2937 ( .A(n2905), .ZN(n2651) );
  OR2_X1 U2938 ( .A1(n2374), .A2(n4484), .ZN(n2386) );
  NAND2_X1 U2939 ( .A1(n2413), .A2(REG3_REG_10__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U2940 ( .A1(n2536), .A2(REG3_REG_21__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U2941 ( .A1(n2492), .A2(REG3_REG_17__SCAN_IN), .ZN(n2508) );
  INV_X1 U2942 ( .A(n4088), .ZN(n4077) );
  NOR2_X1 U2943 ( .A1(n2872), .A2(n4278), .ZN(n3499) );
  INV_X1 U2944 ( .A(n3521), .ZN(n3503) );
  AND2_X1 U2945 ( .A1(n2582), .A2(n2581), .ZN(n3803) );
  INV_X1 U2946 ( .A(n3947), .ZN(n3985) );
  NAND2_X1 U2947 ( .A1(n2409), .A2(n2408), .ZN(n2453) );
  INV_X1 U2948 ( .A(n4100), .ZN(n4078) );
  INV_X1 U2949 ( .A(n3514), .ZN(n4079) );
  AND2_X1 U2950 ( .A1(n3572), .A2(n3535), .ZN(n4098) );
  NAND2_X1 U2951 ( .A1(n2629), .A2(n2628), .ZN(n4083) );
  INV_X1 U2952 ( .A(n4066), .ZN(n4377) );
  AOI21_X1 U2953 ( .B1(n2846), .B2(n4596), .A(n2915), .ZN(n2847) );
  INV_X1 U2954 ( .A(n2799), .ZN(n3930) );
  AND2_X1 U2955 ( .A1(n4102), .A2(n4416), .ZN(n4438) );
  AND2_X1 U2956 ( .A1(n4382), .A2(n2685), .ZN(n4423) );
  NAND2_X1 U2957 ( .A1(n2652), .A2(n2650), .ZN(n2914) );
  AND2_X1 U2958 ( .A1(n2487), .A2(n2477), .ZN(n3755) );
  AND2_X1 U2959 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  INV_X1 U2960 ( .A(n3510), .ZN(n3505) );
  INV_X1 U2961 ( .A(n3790), .ZN(n3809) );
  OAI211_X1 U2962 ( .C1(n2586), .C2(n3874), .A(n2563), .B(n2562), .ZN(n3888)
         );
  INV_X1 U2963 ( .A(n3681), .ZN(n3679) );
  INV_X1 U2964 ( .A(n4333), .ZN(n4468) );
  NAND2_X1 U2965 ( .A1(n4372), .A2(n3161), .ZN(n4035) );
  NAND2_X1 U2966 ( .A1(n4454), .A2(n4443), .ZN(n4208) );
  NAND2_X1 U2967 ( .A1(n4446), .A2(n4443), .ZN(n4266) );
  INV_X1 U2968 ( .A(n4446), .ZN(n4444) );
  INV_X1 U2969 ( .A(n4393), .ZN(n4392) );
  AND2_X1 U2970 ( .A1(n2672), .A2(n2671), .ZN(n2915) );
  INV_X1 U2971 ( .A(n2301), .ZN(n4268) );
  INV_X1 U2972 ( .A(n3751), .ZN(n4403) );
  AND2_X1 U2973 ( .A1(n2392), .A2(n2382), .ZN(n4271) );
  INV_X1 U2974 ( .A(n3681), .ZN(U4043) );
  INV_X1 U2975 ( .A(IR_REG_24__SCAN_IN), .ZN(n2292) );
  NAND2_X1 U2976 ( .A1(n2653), .A2(n2292), .ZN(n2293) );
  NAND2_X1 U2977 ( .A1(n2296), .A2(n2299), .ZN(n3346) );
  NAND2_X1 U2978 ( .A1(n2303), .A2(n2304), .ZN(n2305) );
  NAND2_X1 U2979 ( .A1(n2308), .A2(IR_REG_27__SCAN_IN), .ZN(n2306) );
  INV_X1 U2980 ( .A(n2311), .ZN(n2683) );
  INV_X1 U2981 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3022) );
  OR2_X1 U2982 ( .A1(n2328), .A2(n3022), .ZN(n2314) );
  NAND2_X1 U2983 ( .A1(n2318), .A2(REG0_REG_0__SCAN_IN), .ZN(n2313) );
  NAND4_X1 U2984 ( .A1(n2315), .A2(n2314), .A3(n2313), .A4(n2312), .ZN(n2691)
         );
  AND2_X1 U2985 ( .A1(n2691), .A2(n2690), .ZN(n3035) );
  NAND2_X1 U2986 ( .A1(n2350), .A2(REG2_REG_2__SCAN_IN), .ZN(n2325) );
  INV_X1 U2987 ( .A(n2318), .ZN(n2331) );
  INV_X1 U2988 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2319) );
  OR2_X1 U2989 ( .A1(n2331), .A2(n2319), .ZN(n2324) );
  INV_X1 U2990 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2320) );
  OR2_X1 U2991 ( .A1(n2328), .A2(n2320), .ZN(n2322) );
  NAND2_X1 U2992 ( .A1(n2329), .A2(REG1_REG_2__SCAN_IN), .ZN(n2321) );
  AND2_X1 U2993 ( .A1(n2322), .A2(n2321), .ZN(n2323) );
  MUX2_X1 U2994 ( .A(n4275), .B(DATAI_2_), .S(n2357), .Z(n3476) );
  NAND2_X1 U2995 ( .A1(n3678), .A2(n2702), .ZN(n3546) );
  NAND2_X1 U2996 ( .A1(n3112), .A2(n3476), .ZN(n3543) );
  NAND2_X1 U2997 ( .A1(n3063), .A2(n2610), .ZN(n3062) );
  NAND2_X1 U2998 ( .A1(n3112), .A2(n2702), .ZN(n3083) );
  OR2_X1 U2999 ( .A1(n2328), .A2(REG3_REG_3__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U3000 ( .A1(n2329), .A2(REG1_REG_3__SCAN_IN), .ZN(n2335) );
  INV_X1 U3001 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2330) );
  OR2_X1 U3002 ( .A1(n2586), .A2(n2330), .ZN(n2334) );
  INV_X1 U3003 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2332) );
  OR2_X1 U3004 ( .A1(n2331), .A2(n2332), .ZN(n2333) );
  NAND4_X1 U3005 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n2708)
         );
  NAND2_X1 U3006 ( .A1(n2327), .A2(IR_REG_31__SCAN_IN), .ZN(n2338) );
  XNOR2_X1 U3007 ( .A(n2338), .B(IR_REG_3__SCAN_IN), .ZN(n4274) );
  MUX2_X1 U3008 ( .A(n4274), .B(DATAI_3_), .S(n2357), .Z(n3115) );
  OR2_X1 U3009 ( .A1(n2708), .A2(n3115), .ZN(n2337) );
  AND2_X1 U3010 ( .A1(n3083), .A2(n2337), .ZN(n3118) );
  NAND2_X1 U3011 ( .A1(n2318), .A2(REG0_REG_4__SCAN_IN), .ZN(n2344) );
  INV_X1 U3012 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2948) );
  OR2_X1 U3013 ( .A1(n2507), .A2(n2948), .ZN(n2343) );
  NAND2_X1 U3014 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2348) );
  OAI21_X1 U3015 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2348), .ZN(n3152) );
  INV_X1 U3016 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2973) );
  OR2_X1 U3017 ( .A1(n2586), .A2(n2973), .ZN(n2341) );
  NAND2_X1 U3018 ( .A1(n2338), .A2(n4545), .ZN(n2339) );
  NAND2_X1 U3019 ( .A1(n2339), .A2(IR_REG_31__SCAN_IN), .ZN(n2340) );
  XNOR2_X1 U3020 ( .A(n2340), .B(IR_REG_4__SCAN_IN), .ZN(n4273) );
  MUX2_X1 U3021 ( .A(n4273), .B(DATAI_4_), .S(n2357), .Z(n3149) );
  NAND4_X1 U3022 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(n3677)
         );
  INV_X1 U3023 ( .A(n3149), .ZN(n3131) );
  NAND2_X1 U3024 ( .A1(n3549), .A2(n3551), .ZN(n3120) );
  AND2_X1 U3025 ( .A1(n3118), .A2(n3120), .ZN(n2346) );
  INV_X1 U3026 ( .A(n2708), .ZN(n3146) );
  NAND2_X1 U3027 ( .A1(n2708), .A2(n3115), .ZN(n3119) );
  AOI22_X1 U3028 ( .A1(n3062), .A2(n2346), .B1(n2345), .B2(n3120), .ZN(n3123)
         );
  NAND2_X1 U3029 ( .A1(n3677), .A2(n3149), .ZN(n2347) );
  NAND2_X1 U3030 ( .A1(n3123), .A2(n2347), .ZN(n3162) );
  NAND2_X1 U3031 ( .A1(n2918), .A2(REG0_REG_5__SCAN_IN), .ZN(n2354) );
  INV_X1 U3032 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2951) );
  OR2_X1 U3033 ( .A1(n2507), .A2(n2951), .ZN(n2353) );
  INV_X1 U3034 ( .A(n2363), .ZN(n2365) );
  NAND2_X1 U3035 ( .A1(n2348), .A2(n2986), .ZN(n2349) );
  NAND2_X1 U3036 ( .A1(n2365), .A2(n2349), .ZN(n3171) );
  OR2_X1 U3037 ( .A1(n2328), .A2(n3171), .ZN(n2352) );
  INV_X1 U3038 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3168) );
  OR2_X1 U3039 ( .A1(n2586), .A2(n3168), .ZN(n2351) );
  NAND2_X1 U3040 ( .A1(n2355), .A2(IR_REG_31__SCAN_IN), .ZN(n2356) );
  XNOR2_X1 U3041 ( .A(n2356), .B(n2243), .ZN(n2987) );
  INV_X1 U3042 ( .A(DATAI_5_), .ZN(n2358) );
  CLKBUF_X3 U3043 ( .A(n2357), .Z(n3528) );
  MUX2_X1 U3044 ( .A(n2987), .B(n2358), .S(n3528), .Z(n2724) );
  NAND2_X1 U3045 ( .A1(n3212), .A2(n2724), .ZN(n2359) );
  NAND2_X1 U3046 ( .A1(n3162), .A2(n2359), .ZN(n2361) );
  INV_X1 U3047 ( .A(n3212), .ZN(n3676) );
  NAND2_X1 U3048 ( .A1(n3676), .A2(n3170), .ZN(n2360) );
  NAND2_X1 U3049 ( .A1(n2361), .A2(n2360), .ZN(n3210) );
  NAND2_X1 U3050 ( .A1(n2918), .A2(REG0_REG_6__SCAN_IN), .ZN(n2370) );
  INV_X1 U3051 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2362) );
  OR2_X1 U3052 ( .A1(n2507), .A2(n2362), .ZN(n2369) );
  NAND2_X1 U3053 ( .A1(n2363), .A2(REG3_REG_6__SCAN_IN), .ZN(n2374) );
  INV_X1 U3054 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2364) );
  NAND2_X1 U3055 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  NAND2_X1 U3056 ( .A1(n2374), .A2(n2366), .ZN(n4371) );
  OR2_X1 U3057 ( .A1(n2328), .A2(n4371), .ZN(n2368) );
  INV_X1 U3058 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2976) );
  OR2_X1 U3059 ( .A1(n2586), .A2(n2976), .ZN(n2367) );
  NAND4_X1 U3060 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .ZN(n3675)
         );
  OR2_X1 U3061 ( .A1(n2044), .A2(n2641), .ZN(n2371) );
  XNOR2_X1 U3062 ( .A(n2371), .B(IR_REG_6__SCAN_IN), .ZN(n4272) );
  MUX2_X1 U3063 ( .A(n4272), .B(DATAI_6_), .S(n3528), .Z(n3194) );
  AND2_X1 U3064 ( .A1(n3675), .A2(n3194), .ZN(n2372) );
  NAND2_X1 U3065 ( .A1(n2918), .A2(REG0_REG_7__SCAN_IN), .ZN(n2379) );
  INV_X1 U3066 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2373) );
  OR2_X1 U3067 ( .A1(n2507), .A2(n2373), .ZN(n2378) );
  NAND2_X1 U3068 ( .A1(n2374), .A2(n4484), .ZN(n2375) );
  NAND2_X1 U3069 ( .A1(n2386), .A2(n2375), .ZN(n3245) );
  OR2_X1 U3070 ( .A1(n2328), .A2(n3245), .ZN(n2377) );
  INV_X1 U3071 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2977) );
  OR2_X1 U3072 ( .A1(n2586), .A2(n2977), .ZN(n2376) );
  NAND2_X1 U3073 ( .A1(n2044), .A2(n4544), .ZN(n2405) );
  NAND2_X1 U3074 ( .A1(n2405), .A2(IR_REG_31__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3075 ( .A1(n2381), .A2(n2380), .ZN(n2392) );
  OR2_X1 U3076 ( .A1(n2381), .A2(n2380), .ZN(n2382) );
  MUX2_X1 U3077 ( .A(n4271), .B(DATAI_7_), .S(n3528), .Z(n3242) );
  NAND2_X1 U3078 ( .A1(n3213), .A2(n3242), .ZN(n2613) );
  NAND2_X1 U3079 ( .A1(n3252), .A2(n3179), .ZN(n3537) );
  NAND2_X1 U3080 ( .A1(n3252), .A2(n3242), .ZN(n2383) );
  NAND2_X1 U3081 ( .A1(n2918), .A2(REG0_REG_8__SCAN_IN), .ZN(n2391) );
  INV_X1 U3082 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2384) );
  OR2_X1 U3083 ( .A1(n2507), .A2(n2384), .ZN(n2390) );
  NAND2_X1 U3084 ( .A1(n2386), .A2(n2385), .ZN(n2387) );
  NAND2_X1 U3085 ( .A1(n2399), .A2(n2387), .ZN(n3251) );
  OR2_X1 U3086 ( .A1(n2328), .A2(n3251), .ZN(n2389) );
  INV_X1 U3087 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3205) );
  OR2_X1 U3088 ( .A1(n2586), .A2(n3205), .ZN(n2388) );
  NAND2_X1 U3089 ( .A1(n2392), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  INV_X1 U3090 ( .A(IR_REG_8__SCAN_IN), .ZN(n2393) );
  XNOR2_X1 U3091 ( .A(n2394), .B(n2393), .ZN(n4408) );
  INV_X1 U3092 ( .A(DATAI_8_), .ZN(n2395) );
  MUX2_X1 U3093 ( .A(n4408), .B(n2395), .S(n3528), .Z(n3254) );
  NAND2_X1 U3094 ( .A1(n3276), .A2(n3254), .ZN(n2396) );
  NAND2_X1 U3095 ( .A1(n3201), .A2(n2396), .ZN(n2398) );
  NAND2_X1 U3096 ( .A1(n3264), .A2(n3202), .ZN(n2397) );
  NAND2_X1 U3097 ( .A1(n2398), .A2(n2397), .ZN(n3260) );
  NAND2_X1 U3098 ( .A1(n2918), .A2(REG0_REG_9__SCAN_IN), .ZN(n2404) );
  INV_X1 U3099 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3009) );
  OR2_X1 U3100 ( .A1(n2507), .A2(n3009), .ZN(n2403) );
  INV_X1 U3101 ( .A(n2413), .ZN(n2415) );
  NAND2_X1 U3102 ( .A1(n2399), .A2(n3002), .ZN(n2400) );
  NAND2_X1 U3103 ( .A1(n2415), .A2(n2400), .ZN(n3282) );
  OR2_X1 U3104 ( .A1(n2328), .A2(n3282), .ZN(n2402) );
  INV_X1 U3105 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3269) );
  OR2_X1 U3106 ( .A1(n2586), .A2(n3269), .ZN(n2401) );
  NAND4_X1 U3107 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n3674)
         );
  NAND2_X1 U3108 ( .A1(n2407), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  MUX2_X1 U3109 ( .A(n2406), .B(IR_REG_31__SCAN_IN), .S(n2408), .Z(n2410) );
  NAND2_X1 U3110 ( .A1(n2410), .A2(n2453), .ZN(n3728) );
  INV_X1 U3111 ( .A(n3728), .ZN(n4270) );
  MUX2_X1 U3112 ( .A(n4270), .B(DATAI_9_), .S(n3528), .Z(n3279) );
  AND2_X1 U3113 ( .A1(n3674), .A2(n3279), .ZN(n2412) );
  INV_X1 U3114 ( .A(n3674), .ZN(n3299) );
  INV_X1 U3115 ( .A(n3279), .ZN(n3262) );
  NAND2_X1 U3116 ( .A1(n3299), .A2(n3262), .ZN(n2411) );
  NAND2_X1 U3117 ( .A1(n2918), .A2(REG0_REG_10__SCAN_IN), .ZN(n2420) );
  INV_X1 U3118 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4458) );
  OR2_X1 U3119 ( .A1(n2507), .A2(n4458), .ZN(n2419) );
  INV_X1 U3120 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3121 ( .A1(n2415), .A2(n2414), .ZN(n2416) );
  NAND2_X1 U3122 ( .A1(n2423), .A2(n2416), .ZN(n3304) );
  OR2_X1 U3123 ( .A1(n2328), .A2(n3304), .ZN(n2418) );
  INV_X1 U3124 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3291) );
  OR2_X1 U3125 ( .A1(n2586), .A2(n3291), .ZN(n2417) );
  NAND4_X1 U3126 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n4105)
         );
  NAND2_X1 U3127 ( .A1(n2453), .A2(IR_REG_31__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U3128 ( .A(n2421), .B(IR_REG_10__SCAN_IN), .ZN(n3746) );
  MUX2_X1 U3129 ( .A(n3746), .B(DATAI_10_), .S(n3528), .Z(n3301) );
  NOR2_X1 U3130 ( .A1(n4105), .A2(n3301), .ZN(n2422) );
  NAND2_X1 U3131 ( .A1(n2918), .A2(REG0_REG_11__SCAN_IN), .ZN(n2428) );
  INV_X1 U3132 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4206) );
  OR2_X1 U3133 ( .A1(n2507), .A2(n4206), .ZN(n2427) );
  NAND2_X1 U3134 ( .A1(n2423), .A2(n3331), .ZN(n2424) );
  NAND2_X1 U3135 ( .A1(n2430), .A2(n2424), .ZN(n4114) );
  OR2_X1 U3136 ( .A1(n2328), .A2(n4114), .ZN(n2426) );
  INV_X1 U3137 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4115) );
  OR2_X1 U3138 ( .A1(n2586), .A2(n4115), .ZN(n2425) );
  OAI21_X1 U3139 ( .B1(n2453), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2437) );
  XNOR2_X1 U3140 ( .A(n2437), .B(IR_REG_11__SCAN_IN), .ZN(n3748) );
  MUX2_X1 U3141 ( .A(n3748), .B(DATAI_11_), .S(n3528), .Z(n3334) );
  NAND2_X1 U3142 ( .A1(n3307), .A2(n3334), .ZN(n3572) );
  INV_X1 U3143 ( .A(n3307), .ZN(n3673) );
  NAND2_X1 U3144 ( .A1(n3673), .A2(n4110), .ZN(n3535) );
  NAND2_X1 U3145 ( .A1(n2918), .A2(REG0_REG_12__SCAN_IN), .ZN(n2436) );
  INV_X1 U3146 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4305) );
  OR2_X1 U3147 ( .A1(n2507), .A2(n4305), .ZN(n2435) );
  INV_X1 U31480 ( .A(n2442), .ZN(n2443) );
  NAND2_X1 U31490 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  NAND2_X1 U3150 ( .A1(n2443), .A2(n2431), .ZN(n3315) );
  OR2_X1 U3151 ( .A1(n2328), .A2(n3315), .ZN(n2434) );
  INV_X1 U3152 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2432) );
  OR2_X1 U3153 ( .A1(n2586), .A2(n2432), .ZN(n2433) );
  INV_X1 U3154 ( .A(IR_REG_11__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U3155 ( .A1(n2437), .A2(n2451), .ZN(n2438) );
  NAND2_X1 U3156 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  XNOR2_X1 U3157 ( .A(n2439), .B(IR_REG_12__SCAN_IN), .ZN(n3732) );
  INV_X1 U3158 ( .A(DATAI_12_), .ZN(n4404) );
  MUX2_X1 U3159 ( .A(n4405), .B(n4404), .S(n3528), .Z(n3400) );
  NAND2_X1 U3160 ( .A1(n3312), .A2(n2440), .ZN(n2441) );
  NAND2_X1 U3161 ( .A1(n2441), .A2(n2271), .ZN(n4071) );
  NAND2_X1 U3162 ( .A1(n2918), .A2(REG0_REG_13__SCAN_IN), .ZN(n2448) );
  INV_X1 U3163 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4197) );
  OR2_X1 U3164 ( .A1(n2507), .A2(n4197), .ZN(n2447) );
  NAND2_X1 U3165 ( .A1(n2442), .A2(REG3_REG_13__SCAN_IN), .ZN(n2459) );
  INV_X1 U3166 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U3167 ( .A1(n2443), .A2(n3461), .ZN(n2444) );
  NAND2_X1 U3168 ( .A1(n2459), .A2(n2444), .ZN(n4090) );
  OR2_X1 U3169 ( .A1(n2328), .A2(n4090), .ZN(n2446) );
  INV_X1 U3170 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4091) );
  OR2_X1 U3171 ( .A1(n2586), .A2(n4091), .ZN(n2445) );
  INV_X1 U3172 ( .A(IR_REG_10__SCAN_IN), .ZN(n2450) );
  INV_X1 U3173 ( .A(IR_REG_12__SCAN_IN), .ZN(n2449) );
  NAND3_X1 U3174 ( .A1(n2451), .A2(n2450), .A3(n2449), .ZN(n2452) );
  OAI21_X1 U3175 ( .B1(n2453), .B2(n2452), .A(IR_REG_31__SCAN_IN), .ZN(n2454)
         );
  MUX2_X1 U3176 ( .A(IR_REG_31__SCAN_IN), .B(n2454), .S(IR_REG_13__SCAN_IN), 
        .Z(n2457) );
  INV_X1 U3177 ( .A(n2455), .ZN(n2456) );
  INV_X1 U3178 ( .A(DATAI_13_), .ZN(n4402) );
  MUX2_X1 U3179 ( .A(n4403), .B(n4402), .S(n3528), .Z(n4088) );
  NAND2_X1 U3180 ( .A1(n2918), .A2(REG0_REG_14__SCAN_IN), .ZN(n2465) );
  INV_X1 U3181 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4326) );
  OR2_X1 U3182 ( .A1(n2507), .A2(n4326), .ZN(n2464) );
  INV_X1 U3183 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3184 ( .A1(n2459), .A2(n2458), .ZN(n2460) );
  NAND2_X1 U3185 ( .A1(n2467), .A2(n2460), .ZN(n3363) );
  OR2_X1 U3186 ( .A1(n2328), .A2(n3363), .ZN(n2463) );
  INV_X1 U3187 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2461) );
  OR2_X1 U3188 ( .A1(n2586), .A2(n2461), .ZN(n2462) );
  OR2_X1 U3189 ( .A1(n2455), .A2(n2641), .ZN(n2466) );
  XNOR2_X1 U3190 ( .A(n2466), .B(IR_REG_14__SCAN_IN), .ZN(n4332) );
  MUX2_X1 U3191 ( .A(n4332), .B(DATAI_14_), .S(n3528), .Z(n4061) );
  NAND2_X1 U3192 ( .A1(n3514), .A2(n4061), .ZN(n3568) );
  INV_X1 U3193 ( .A(n4061), .ZN(n4052) );
  NAND2_X1 U3194 ( .A1(n4079), .A2(n4052), .ZN(n3531) );
  NAND2_X1 U3195 ( .A1(n3568), .A2(n3531), .ZN(n4059) );
  NAND2_X1 U3196 ( .A1(n2918), .A2(REG0_REG_15__SCAN_IN), .ZN(n2472) );
  INV_X1 U3197 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3754) );
  OR2_X1 U3198 ( .A1(n2507), .A2(n3754), .ZN(n2471) );
  INV_X1 U3199 ( .A(n2479), .ZN(n2481) );
  NAND2_X1 U3200 ( .A1(n2467), .A2(n3512), .ZN(n2468) );
  NAND2_X1 U3201 ( .A1(n2481), .A2(n2468), .ZN(n4043) );
  OR2_X1 U3202 ( .A1(n2328), .A2(n4043), .ZN(n2470) );
  INV_X1 U3203 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4044) );
  OR2_X1 U3204 ( .A1(n2586), .A2(n4044), .ZN(n2469) );
  INV_X1 U3205 ( .A(IR_REG_14__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3206 ( .A1(n2455), .A2(n2473), .ZN(n2474) );
  NAND2_X1 U3207 ( .A1(n2474), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  INV_X1 U3208 ( .A(IR_REG_15__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3209 ( .A1(n2476), .A2(n2475), .ZN(n2487) );
  OR2_X1 U32100 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  MUX2_X1 U32110 ( .A(n3755), .B(DATAI_15_), .S(n3528), .Z(n3518) );
  NAND2_X1 U32120 ( .A1(n3419), .A2(n3518), .ZN(n2478) );
  NAND2_X1 U32130 ( .A1(n2350), .A2(REG2_REG_16__SCAN_IN), .ZN(n2486) );
  INV_X1 U32140 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4527) );
  OR2_X1 U32150 ( .A1(n2331), .A2(n4527), .ZN(n2485) );
  INV_X1 U32160 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4354) );
  OR2_X1 U32170 ( .A1(n2507), .A2(n4354), .ZN(n2484) );
  INV_X1 U32180 ( .A(n2492), .ZN(n2494) );
  INV_X1 U32190 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U32200 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  NAND2_X1 U32210 ( .A1(n2494), .A2(n2482), .ZN(n4024) );
  OR2_X1 U32220 ( .A1(n2328), .A2(n4024), .ZN(n2483) );
  NAND2_X1 U32230 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2489) );
  INV_X1 U32240 ( .A(IR_REG_16__SCAN_IN), .ZN(n2488) );
  XNOR2_X1 U32250 ( .A(n2489), .B(n2488), .ZN(n4398) );
  INV_X1 U32260 ( .A(n4398), .ZN(n2490) );
  MUX2_X1 U32270 ( .A(n2490), .B(DATAI_16_), .S(n3528), .Z(n4029) );
  NAND2_X1 U32280 ( .A1(n4036), .A2(n4029), .ZN(n3635) );
  INV_X1 U32290 ( .A(n4036), .ZN(n3671) );
  INV_X1 U32300 ( .A(n4029), .ZN(n3421) );
  NAND2_X1 U32310 ( .A1(n3671), .A2(n3421), .ZN(n3530) );
  NAND2_X1 U32320 ( .A1(n3635), .A2(n3530), .ZN(n4020) );
  NAND2_X1 U32330 ( .A1(n2918), .A2(REG0_REG_17__SCAN_IN), .ZN(n2499) );
  INV_X1 U32340 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4181) );
  OR2_X1 U32350 ( .A1(n2507), .A2(n4181), .ZN(n2498) );
  INV_X1 U32360 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U32370 ( .A1(n2494), .A2(n2493), .ZN(n2495) );
  NAND2_X1 U32380 ( .A1(n2508), .A2(n2495), .ZN(n4013) );
  OR2_X1 U32390 ( .A1(n2328), .A2(n4013), .ZN(n2497) );
  INV_X1 U32400 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4014) );
  OR2_X1 U32410 ( .A1(n2586), .A2(n4014), .ZN(n2496) );
  NAND2_X1 U32420 ( .A1(n2501), .A2(IR_REG_31__SCAN_IN), .ZN(n2502) );
  MUX2_X1 U32430 ( .A(IR_REG_31__SCAN_IN), .B(n2502), .S(IR_REG_17__SCAN_IN), 
        .Z(n2504) );
  INV_X1 U32440 ( .A(n2503), .ZN(n2514) );
  NAND2_X1 U32450 ( .A1(n2504), .A2(n2514), .ZN(n3743) );
  INV_X1 U32460 ( .A(DATAI_17_), .ZN(n2505) );
  MUX2_X1 U32470 ( .A(n3743), .B(n2505), .S(n3528), .Z(n4012) );
  NAND2_X1 U32480 ( .A1(n3987), .A2(n4012), .ZN(n2506) );
  NAND2_X1 U32490 ( .A1(n2918), .A2(REG0_REG_18__SCAN_IN), .ZN(n2513) );
  INV_X1 U32500 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3764) );
  OR2_X1 U32510 ( .A1(n2507), .A2(n3764), .ZN(n2512) );
  INV_X1 U32520 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U32530 ( .A1(n2508), .A2(n3487), .ZN(n2509) );
  NAND2_X1 U32540 ( .A1(n2516), .A2(n2509), .ZN(n3996) );
  OR2_X1 U32550 ( .A1(n2328), .A2(n3996), .ZN(n2511) );
  INV_X1 U32560 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3997) );
  OR2_X1 U32570 ( .A1(n2586), .A2(n3997), .ZN(n2510) );
  NAND2_X1 U32580 ( .A1(n2514), .A2(IR_REG_31__SCAN_IN), .ZN(n2515) );
  XNOR2_X1 U32590 ( .A(n2515), .B(IR_REG_18__SCAN_IN), .ZN(n3770) );
  MUX2_X1 U32600 ( .A(n3770), .B(DATAI_18_), .S(n3528), .Z(n3993) );
  NAND2_X1 U32610 ( .A1(n3974), .A2(n3993), .ZN(n3964) );
  NAND2_X1 U32620 ( .A1(n4006), .A2(n2786), .ZN(n3965) );
  NAND2_X1 U32630 ( .A1(n3964), .A2(n3965), .ZN(n3991) );
  NAND2_X1 U32640 ( .A1(n3992), .A2(n3991), .ZN(n3990) );
  NAND2_X1 U32650 ( .A1(n2918), .A2(REG0_REG_19__SCAN_IN), .ZN(n2522) );
  INV_X1 U32660 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4173) );
  OR2_X1 U32670 ( .A1(n2507), .A2(n4173), .ZN(n2521) );
  INV_X1 U32680 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U32690 ( .A1(n2516), .A2(n4598), .ZN(n2517) );
  NAND2_X1 U32700 ( .A1(n2530), .A2(n2517), .ZN(n3381) );
  OR2_X1 U32710 ( .A1(n2328), .A2(n3381), .ZN(n2520) );
  INV_X1 U32720 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2518) );
  OR2_X1 U32730 ( .A1(n2586), .A2(n2518), .ZN(n2519) );
  INV_X1 U32740 ( .A(n2526), .ZN(n2524) );
  NAND2_X1 U32750 ( .A1(n2524), .A2(IR_REG_19__SCAN_IN), .ZN(n2527) );
  INV_X1 U32760 ( .A(IR_REG_19__SCAN_IN), .ZN(n2525) );
  MUX2_X1 U32770 ( .A(n4269), .B(DATAI_19_), .S(n3528), .Z(n3970) );
  NAND2_X1 U32780 ( .A1(n3985), .A2(n3970), .ZN(n2529) );
  NAND2_X1 U32790 ( .A1(n2918), .A2(REG0_REG_20__SCAN_IN), .ZN(n2535) );
  INV_X1 U32800 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4169) );
  OR2_X1 U32810 ( .A1(n2507), .A2(n4169), .ZN(n2534) );
  INV_X1 U32820 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3450) );
  INV_X1 U32830 ( .A(n2536), .ZN(n2537) );
  NAND2_X1 U32840 ( .A1(n2530), .A2(n3450), .ZN(n2531) );
  NAND2_X1 U32850 ( .A1(n2537), .A2(n2531), .ZN(n3954) );
  OR2_X1 U32860 ( .A1(n2328), .A2(n3954), .ZN(n2533) );
  INV_X1 U32870 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3955) );
  OR2_X1 U32880 ( .A1(n2586), .A2(n3955), .ZN(n2532) );
  NAND2_X1 U32890 ( .A1(n3528), .A2(DATAI_20_), .ZN(n3952) );
  INV_X1 U32900 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U32910 ( .A1(n2537), .A2(n4587), .ZN(n2538) );
  NAND2_X1 U32920 ( .A1(n2552), .A2(n2538), .ZN(n3932) );
  OR2_X1 U32930 ( .A1(n3932), .A2(n2328), .ZN(n2542) );
  NAND2_X1 U32940 ( .A1(n2918), .A2(REG0_REG_21__SCAN_IN), .ZN(n2541) );
  INV_X1 U32950 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4164) );
  OR2_X1 U32960 ( .A1(n2507), .A2(n4164), .ZN(n2540) );
  INV_X1 U32970 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3933) );
  OR2_X1 U32980 ( .A1(n2586), .A2(n3933), .ZN(n2539) );
  INV_X1 U32990 ( .A(n3908), .ZN(n3945) );
  INV_X1 U33000 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U33010 ( .A1(n2918), .A2(REG0_REG_22__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U33020 ( .A1(n2350), .A2(REG2_REG_22__SCAN_IN), .ZN(n2543) );
  OAI211_X1 U33030 ( .C1(n2507), .C2(n4531), .A(n2544), .B(n2543), .ZN(n2545)
         );
  INV_X1 U33040 ( .A(n2545), .ZN(n2547) );
  XNOR2_X1 U33050 ( .A(n2552), .B(REG3_REG_22__SCAN_IN), .ZN(n3914) );
  NAND2_X1 U33060 ( .A1(n3914), .A2(n2636), .ZN(n2546) );
  NAND2_X1 U33070 ( .A1(n3528), .A2(DATAI_22_), .ZN(n3913) );
  OR2_X1 U33080 ( .A1(n3925), .A2(n3913), .ZN(n3884) );
  NAND2_X1 U33090 ( .A1(n3925), .A2(n3913), .ZN(n2624) );
  NAND2_X1 U33100 ( .A1(n3884), .A2(n2624), .ZN(n3902) );
  NAND2_X1 U33110 ( .A1(n3903), .A2(n3902), .ZN(n3901) );
  NAND2_X1 U33120 ( .A1(n3925), .A2(n2548), .ZN(n2549) );
  NAND2_X1 U33130 ( .A1(n3901), .A2(n2549), .ZN(n3879) );
  INV_X1 U33140 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3467) );
  INV_X1 U33150 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2550) );
  OAI21_X1 U33160 ( .B1(n2552), .B2(n3467), .A(n2550), .ZN(n2553) );
  NAND2_X1 U33170 ( .A1(REG3_REG_22__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .ZN(
        n2551) );
  AND2_X1 U33180 ( .A1(n2553), .A2(n2560), .ZN(n3894) );
  NAND2_X1 U33190 ( .A1(n3894), .A2(n2636), .ZN(n2556) );
  AOI22_X1 U33200 ( .A1(n2329), .A2(REG1_REG_23__SCAN_IN), .B1(n2918), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U33210 ( .A1(n2350), .A2(REG2_REG_23__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U33220 ( .A1(n3528), .A2(DATAI_23_), .ZN(n3893) );
  NAND2_X1 U33230 ( .A1(n3865), .A2(n3893), .ZN(n2558) );
  NOR2_X1 U33240 ( .A1(n3865), .A2(n3893), .ZN(n2557) );
  AOI21_X2 U33250 ( .B1(n3879), .B2(n2558), .A(n2557), .ZN(n3860) );
  INV_X1 U33260 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3874) );
  INV_X1 U33270 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U33280 ( .A1(n2560), .A2(n4511), .ZN(n2561) );
  NAND2_X1 U33290 ( .A1(n2567), .A2(n2561), .ZN(n3873) );
  OR2_X1 U33300 ( .A1(n3873), .A2(n2328), .ZN(n2563) );
  AOI22_X1 U33310 ( .A1(n2329), .A2(REG1_REG_24__SCAN_IN), .B1(n2918), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2562) );
  AND2_X1 U33320 ( .A1(n3528), .A2(DATAI_24_), .ZN(n2814) );
  NAND2_X1 U33330 ( .A1(n3888), .A2(n2814), .ZN(n2564) );
  NAND2_X1 U33340 ( .A1(n3860), .A2(n2564), .ZN(n2566) );
  INV_X1 U33350 ( .A(n3888), .ZN(n3847) );
  NAND2_X1 U33360 ( .A1(n3847), .A2(n3871), .ZN(n2565) );
  INV_X1 U33370 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U33380 ( .A1(n2567), .A2(n3410), .ZN(n2568) );
  NAND2_X1 U33390 ( .A1(n3855), .A2(n2636), .ZN(n2574) );
  INV_X1 U33400 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U33410 ( .A1(n2329), .A2(REG1_REG_25__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U33420 ( .A1(n2918), .A2(REG0_REG_25__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U33430 ( .C1(n2571), .C2(n2586), .A(n2570), .B(n2569), .ZN(n2572)
         );
  INV_X1 U33440 ( .A(n2572), .ZN(n2573) );
  NAND2_X1 U33450 ( .A1(n3867), .A2(n2825), .ZN(n2575) );
  INV_X1 U33460 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U33470 ( .A1(n2576), .A2(n3496), .ZN(n2577) );
  NAND2_X1 U33480 ( .A1(n3837), .A2(n2636), .ZN(n2582) );
  INV_X1 U33490 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U33500 ( .A1(n2329), .A2(REG1_REG_26__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33510 ( .A1(n2350), .A2(REG2_REG_26__SCAN_IN), .ZN(n2578) );
  OAI211_X1 U33520 ( .C1(n2331), .C2(n4533), .A(n2579), .B(n2578), .ZN(n2580)
         );
  INV_X1 U3353 ( .A(n2580), .ZN(n2581) );
  NAND2_X1 U33540 ( .A1(n3528), .A2(DATAI_26_), .ZN(n3835) );
  NOR2_X1 U3355 ( .A1(n3803), .A2(n3835), .ZN(n2583) );
  XNOR2_X1 U3356 ( .A(n2594), .B(REG3_REG_27__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U3357 ( .A1(n3814), .A2(n2636), .ZN(n2589) );
  INV_X1 U3358 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U3359 ( .A1(n2329), .A2(REG1_REG_27__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U3360 ( .A1(n2918), .A2(REG0_REG_27__SCAN_IN), .ZN(n2584) );
  OAI211_X1 U3361 ( .C1(n3815), .C2(n2586), .A(n2585), .B(n2584), .ZN(n2587)
         );
  INV_X1 U3362 ( .A(n2587), .ZN(n2588) );
  AND2_X1 U3363 ( .A1(n3528), .A2(DATAI_27_), .ZN(n2839) );
  NOR2_X1 U3364 ( .A1(n3830), .A2(n2839), .ZN(n2590) );
  INV_X1 U3365 ( .A(n2594), .ZN(n2592) );
  AND2_X1 U3366 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2591) );
  NAND2_X1 U3367 ( .A1(n2592), .A2(n2591), .ZN(n3793) );
  INV_X1 U3368 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3341) );
  INV_X1 U3369 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2593) );
  OAI21_X1 U3370 ( .B1(n2594), .B2(n3341), .A(n2593), .ZN(n2595) );
  NAND2_X1 U3371 ( .A1(n3793), .A2(n2595), .ZN(n3352) );
  INV_X1 U3372 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U3373 ( .A1(n2329), .A2(REG1_REG_28__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U3374 ( .A1(n2918), .A2(REG0_REG_28__SCAN_IN), .ZN(n2596) );
  OAI211_X1 U3375 ( .C1(n3351), .C2(n2586), .A(n2597), .B(n2596), .ZN(n2598)
         );
  INV_X1 U3376 ( .A(n2598), .ZN(n2599) );
  AND2_X1 U3377 ( .A1(n3528), .A2(DATAI_28_), .ZN(n3779) );
  NAND2_X1 U3378 ( .A1(n3790), .A2(n3779), .ZN(n3523) );
  INV_X1 U3379 ( .A(n3779), .ZN(n2853) );
  NAND2_X1 U3380 ( .A1(n3809), .A2(n2853), .ZN(n3783) );
  NAND2_X1 U3381 ( .A1(n3523), .A2(n3783), .ZN(n3780) );
  NAND2_X1 U3382 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2602) );
  MUX2_X1 U3383 ( .A(IR_REG_31__SCAN_IN), .B(n2602), .S(IR_REG_21__SCAN_IN), 
        .Z(n2603) );
  NAND2_X1 U3384 ( .A1(n2603), .A2(n2035), .ZN(n2655) );
  XNOR2_X2 U3385 ( .A(n2606), .B(n2605), .ZN(n2675) );
  NAND2_X2 U3386 ( .A1(n3657), .A2(n2675), .ZN(n3069) );
  NAND2_X1 U3387 ( .A1(n2035), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  XNOR2_X1 U3388 ( .A(n3069), .B(n3667), .ZN(n2608) );
  NAND2_X1 U3389 ( .A1(n2608), .A2(n3775), .ZN(n4102) );
  AND2_X1 U3390 ( .A1(n2675), .A2(n4269), .ZN(n4382) );
  INV_X1 U3391 ( .A(n4423), .ZN(n4416) );
  INV_X1 U3392 ( .A(n2691), .ZN(n3056) );
  NAND2_X1 U3393 ( .A1(n3056), .A2(n2690), .ZN(n3538) );
  NAND2_X1 U3394 ( .A1(n3072), .A2(n2609), .ZN(n2611) );
  NAND2_X1 U3395 ( .A1(n2611), .A2(n3061), .ZN(n3074) );
  NAND2_X1 U3396 ( .A1(n3146), .A2(n3115), .ZN(n3548) );
  NAND2_X1 U3397 ( .A1(n2708), .A2(n3091), .ZN(n3545) );
  NAND2_X1 U3398 ( .A1(n2612), .A2(n3551), .ZN(n3163) );
  NAND2_X1 U3399 ( .A1(n3212), .A2(n3170), .ZN(n3556) );
  NAND2_X1 U3400 ( .A1(n3675), .A2(n3221), .ZN(n3554) );
  NAND2_X1 U3401 ( .A1(n3239), .A2(n3194), .ZN(n3553) );
  NAND2_X1 U3402 ( .A1(n2614), .A2(n3537), .ZN(n3197) );
  NAND2_X1 U3403 ( .A1(n3276), .A2(n3202), .ZN(n3557) );
  NAND2_X1 U3404 ( .A1(n3264), .A2(n3254), .ZN(n3536) );
  AND2_X1 U3405 ( .A1(n3674), .A2(n3262), .ZN(n3565) );
  NAND2_X1 U3406 ( .A1(n3299), .A2(n3279), .ZN(n3558) );
  NAND2_X1 U3407 ( .A1(n4105), .A2(n3288), .ZN(n3534) );
  NAND2_X1 U3408 ( .A1(n3283), .A2(n3534), .ZN(n2615) );
  NAND2_X1 U3409 ( .A1(n3332), .A2(n3301), .ZN(n3563) );
  NAND2_X1 U3410 ( .A1(n2615), .A2(n3563), .ZN(n4097) );
  NAND2_X1 U3411 ( .A1(n4097), .A2(n3535), .ZN(n2616) );
  NAND2_X1 U3412 ( .A1(n2616), .A2(n3572), .ZN(n4074) );
  NAND2_X1 U3413 ( .A1(n3672), .A2(n3400), .ZN(n4072) );
  NAND2_X1 U3414 ( .A1(n4055), .A2(n4088), .ZN(n2617) );
  NAND2_X1 U3415 ( .A1(n4074), .A2(n3566), .ZN(n2619) );
  NOR2_X1 U3416 ( .A1(n3672), .A2(n3400), .ZN(n4073) );
  NOR2_X1 U3417 ( .A1(n4055), .A2(n4088), .ZN(n2618) );
  AOI21_X1 U3418 ( .B1(n3566), .B2(n4073), .A(n2618), .ZN(n3570) );
  NAND2_X1 U3419 ( .A1(n2619), .A2(n3570), .ZN(n4051) );
  INV_X1 U3420 ( .A(n4059), .ZN(n3608) );
  NAND2_X1 U3421 ( .A1(n4051), .A2(n3608), .ZN(n2620) );
  NAND2_X1 U3422 ( .A1(n2620), .A2(n3568), .ZN(n4039) );
  NAND2_X1 U3423 ( .A1(n4053), .A2(n3518), .ZN(n3567) );
  NAND2_X1 U3424 ( .A1(n3419), .A2(n4042), .ZN(n3532) );
  NAND2_X1 U3425 ( .A1(n3567), .A2(n3532), .ZN(n4047) );
  NAND2_X1 U3426 ( .A1(n4037), .A2(n3532), .ZN(n4028) );
  INV_X1 U3427 ( .A(n4020), .ZN(n4027) );
  NAND2_X1 U3428 ( .A1(n4028), .A2(n4027), .ZN(n4026) );
  NAND2_X1 U3429 ( .A1(n3985), .A2(n3975), .ZN(n3593) );
  AND2_X1 U3430 ( .A1(n3965), .A2(n3593), .ZN(n2621) );
  NAND2_X1 U3431 ( .A1(n4030), .A2(n4012), .ZN(n3961) );
  NAND2_X1 U3432 ( .A1(n2621), .A2(n3961), .ZN(n3634) );
  NAND2_X1 U3433 ( .A1(n3987), .A2(n4005), .ZN(n3962) );
  NAND2_X1 U3434 ( .A1(n3964), .A2(n3962), .ZN(n2622) );
  NOR2_X1 U3435 ( .A1(n3985), .A2(n3975), .ZN(n3594) );
  AOI21_X1 U3436 ( .B1(n2622), .B2(n2621), .A(n3594), .ZN(n3940) );
  NAND2_X1 U3437 ( .A1(n3923), .A2(n3944), .ZN(n2623) );
  AND2_X1 U3438 ( .A1(n3971), .A2(n3952), .ZN(n3638) );
  NAND2_X1 U3439 ( .A1(n3908), .A2(n2799), .ZN(n3882) );
  AND2_X1 U3440 ( .A1(n3884), .A2(n3882), .ZN(n3581) );
  INV_X1 U3441 ( .A(n3581), .ZN(n3642) );
  NOR2_X1 U3442 ( .A1(n3908), .A2(n2799), .ZN(n3880) );
  INV_X1 U3443 ( .A(n3865), .ZN(n3910) );
  NAND2_X1 U3444 ( .A1(n3910), .A2(n3893), .ZN(n3598) );
  NAND2_X1 U3445 ( .A1(n3598), .A2(n2624), .ZN(n3584) );
  AOI21_X1 U3446 ( .B1(n3880), .B2(n3884), .A(n3584), .ZN(n3641) );
  NOR2_X1 U3447 ( .A1(n3888), .A2(n3871), .ZN(n3621) );
  NOR2_X1 U3448 ( .A1(n3910), .A2(n3893), .ZN(n3597) );
  NOR2_X1 U3449 ( .A1(n3621), .A2(n3597), .ZN(n3644) );
  NAND2_X1 U3450 ( .A1(n3862), .A2(n3644), .ZN(n3844) );
  NAND2_X1 U3451 ( .A1(n3803), .A2(n2673), .ZN(n2625) );
  INV_X1 U3452 ( .A(n3867), .ZN(n3828) );
  NAND2_X1 U3453 ( .A1(n3828), .A2(n2825), .ZN(n3822) );
  INV_X1 U3454 ( .A(n2825), .ZN(n3853) );
  NAND2_X1 U3455 ( .A1(n3867), .A2(n3853), .ZN(n3592) );
  NAND2_X1 U3456 ( .A1(n3888), .A2(n3871), .ZN(n3843) );
  NAND2_X1 U3457 ( .A1(n3592), .A2(n3843), .ZN(n3823) );
  NOR2_X1 U34580 ( .A1(n3803), .A2(n2673), .ZN(n3630) );
  AOI21_X1 U34590 ( .B1(n3582), .B2(n3823), .A(n3630), .ZN(n3587) );
  OAI21_X1 U3460 ( .B1(n3844), .B2(n3647), .A(n3587), .ZN(n3805) );
  NAND2_X1 U3461 ( .A1(n3830), .A2(n3813), .ZN(n3585) );
  NAND2_X1 U3462 ( .A1(n3522), .A2(n3585), .ZN(n3810) );
  INV_X1 U3463 ( .A(n3522), .ZN(n2626) );
  NOR2_X1 U3464 ( .A1(n3804), .A2(n2626), .ZN(n2627) );
  NAND2_X1 U3465 ( .A1(n3667), .A2(n4269), .ZN(n2629) );
  INV_X1 U3466 ( .A(n2675), .ZN(n3660) );
  NAND2_X1 U34670 ( .A1(n3657), .A2(n3660), .ZN(n2628) );
  INV_X1 U3468 ( .A(n3830), .ZN(n3501) );
  NAND2_X1 U34690 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(
        n2630) );
  NAND2_X1 U3470 ( .A1(n2911), .A2(n2630), .ZN(n2631) );
  NAND2_X1 U34710 ( .A1(n3667), .A2(n3657), .ZN(n2848) );
  NOR2_X1 U3472 ( .A1(n3501), .A2(n4081), .ZN(n2639) );
  INV_X1 U34730 ( .A(n3793), .ZN(n2637) );
  INV_X1 U3474 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U34750 ( .A1(n2918), .A2(REG0_REG_29__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3476 ( .A1(n2350), .A2(REG2_REG_29__SCAN_IN), .ZN(n2632) );
  OAI211_X1 U34770 ( .C1(n2507), .C2(n2634), .A(n2633), .B(n2632), .ZN(n2635)
         );
  AOI21_X1 U3478 ( .B1(n2637), .B2(n2636), .A(n2635), .ZN(n3524) );
  INV_X1 U34790 ( .A(n2848), .ZN(n2959) );
  NAND2_X1 U3480 ( .A1(n2685), .A2(n2655), .ZN(n3042) );
  OAI22_X1 U34810 ( .A1(n3524), .A2(n4100), .B1(n4099), .B2(n2853), .ZN(n2638)
         );
  NOR2_X1 U3482 ( .A1(n2026), .A2(n2641), .ZN(n2643) );
  INV_X1 U34830 ( .A(n2303), .ZN(n2644) );
  NAND2_X1 U3484 ( .A1(n2651), .A2(B_REG_SCAN_IN), .ZN(n2649) );
  NAND2_X1 U34850 ( .A1(n2654), .A2(n2653), .ZN(n2647) );
  MUX2_X1 U3486 ( .A(n2649), .B(B_REG_SCAN_IN), .S(n2901), .Z(n2650) );
  INV_X1 U34870 ( .A(n2652), .ZN(n2672) );
  NAND2_X1 U3488 ( .A1(n2672), .A2(n2651), .ZN(n2844) );
  OAI21_X1 U34890 ( .B1(n2914), .B2(D_REG_1__SCAN_IN), .A(n2844), .ZN(n2670)
         );
  NAND3_X1 U3490 ( .A1(n2652), .A2(n2901), .A3(n2905), .ZN(n2682) );
  NAND2_X1 U34910 ( .A1(n4423), .A2(n2655), .ZN(n2880) );
  AND2_X1 U3492 ( .A1(n2675), .A2(n3775), .ZN(n2656) );
  NAND2_X1 U34930 ( .A1(n2880), .A2(n3064), .ZN(n2657) );
  NOR2_X1 U3494 ( .A1(n2957), .A2(n2657), .ZN(n2669) );
  NOR4_X1 U34950 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2661) );
  NOR4_X1 U3496 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2660) );
  NOR4_X1 U34970 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2659) );
  NOR4_X1 U3498 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2658) );
  AND4_X1 U34990 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n2667)
         );
  NOR2_X1 U3500 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_7__SCAN_IN), .ZN(n2665) );
  NOR4_X1 U35010 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2664) );
  NOR4_X1 U3502 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2663) );
  NOR4_X1 U35030 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2662) );
  AND4_X1 U3504 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n2666)
         );
  NAND2_X1 U35050 ( .A1(n2667), .A2(n2666), .ZN(n2842) );
  NAND2_X1 U35060 ( .A1(n2846), .A2(n2842), .ZN(n2668) );
  INV_X1 U35070 ( .A(D_REG_0__SCAN_IN), .ZN(n4596) );
  INV_X1 U35080 ( .A(n2901), .ZN(n2671) );
  NAND2_X1 U35090 ( .A1(n2683), .A2(n3043), .ZN(n3078) );
  NAND2_X1 U35100 ( .A1(n3219), .A2(n3179), .ZN(n3203) );
  NAND2_X1 U35110 ( .A1(n4062), .A2(n4042), .ZN(n4023) );
  NOR2_X4 U35120 ( .A1(n4009), .A2(n4005), .ZN(n4010) );
  INV_X1 U35130 ( .A(n3812), .ZN(n2674) );
  INV_X1 U35140 ( .A(n3042), .ZN(n2676) );
  NAND2_X1 U35150 ( .A1(n2027), .A2(n2275), .ZN(U3546) );
  INV_X1 U35160 ( .A(n2847), .ZN(n3067) );
  MUX2_X1 U35170 ( .A(REG0_REG_28__SCAN_IN), .B(n2678), .S(n4446), .Z(n2679)
         );
  INV_X1 U35180 ( .A(n2679), .ZN(n2680) );
  NAND2_X1 U35190 ( .A1(n2680), .A2(n2274), .ZN(U3514) );
  INV_X2 U35200 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U35210 ( .A(n3069), .ZN(n2681) );
  NAND2_X2 U35220 ( .A1(n2892), .A2(n2681), .ZN(n2700) );
  INV_X4 U35230 ( .A(n2689), .ZN(n2850) );
  OAI22_X1 U35240 ( .A1(n2684), .A2(n2700), .B1(n2683), .B2(n2850), .ZN(n2686)
         );
  XNOR2_X1 U35250 ( .A(n2686), .B(n2837), .ZN(n2697) );
  NAND2_X1 U35260 ( .A1(n2311), .A2(n2871), .ZN(n2687) );
  NAND2_X1 U35270 ( .A1(n2688), .A2(n2687), .ZN(n2698) );
  XNOR2_X1 U35280 ( .A(n2697), .B(n2698), .ZN(n3053) );
  INV_X1 U35290 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3682) );
  OAI21_X1 U35300 ( .B1(n2892), .B2(n3682), .A(n2696), .ZN(n3019) );
  INV_X1 U35310 ( .A(n2892), .ZN(n2692) );
  INV_X1 U35320 ( .A(n2855), .ZN(n2693) );
  NAND2_X1 U35330 ( .A1(n2695), .A2(n2694), .ZN(n3018) );
  AOI22_X1 U35340 ( .A1(n3019), .A2(n3018), .B1(n2851), .B2(n2696), .ZN(n3055)
         );
  NOR2_X1 U35350 ( .A1(n3054), .A2(n2699), .ZN(n3473) );
  OAI22_X1 U35360 ( .A1(n3112), .A2(n2855), .B1(n2700), .B2(n2702), .ZN(n2703)
         );
  NAND2_X1 U35370 ( .A1(n3473), .A2(n3474), .ZN(n3472) );
  INV_X1 U35380 ( .A(n2704), .ZN(n2706) );
  NAND2_X1 U35390 ( .A1(n3472), .A2(n2707), .ZN(n3110) );
  OAI22_X1 U35400 ( .A1(n3146), .A2(n2855), .B1(n2700), .B2(n3091), .ZN(n2713)
         );
  NAND2_X1 U35410 ( .A1(n2708), .A2(n2871), .ZN(n2710) );
  NAND2_X1 U35420 ( .A1(n3115), .A2(n2689), .ZN(n2709) );
  NAND2_X1 U35430 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  XNOR2_X1 U35440 ( .A(n2711), .B(n2837), .ZN(n2712) );
  XOR2_X1 U35450 ( .A(n2713), .B(n2712), .Z(n3109) );
  INV_X1 U35460 ( .A(n2712), .ZN(n2715) );
  INV_X1 U35470 ( .A(n2713), .ZN(n2714) );
  AOI21_X2 U35480 ( .B1(n3110), .B2(n3109), .A(n2270), .ZN(n3145) );
  OR2_X1 U35490 ( .A1(n3165), .A2(n2855), .ZN(n2717) );
  NAND2_X1 U35500 ( .A1(n3149), .A2(n2023), .ZN(n2716) );
  NAND2_X1 U35510 ( .A1(n2717), .A2(n2716), .ZN(n2720) );
  OAI22_X1 U35520 ( .A1(n3165), .A2(n2700), .B1(n2850), .B2(n3131), .ZN(n2718)
         );
  XNOR2_X1 U35530 ( .A(n2718), .B(n2837), .ZN(n2719) );
  XOR2_X1 U35540 ( .A(n2720), .B(n2719), .Z(n3144) );
  NAND2_X1 U35550 ( .A1(n3145), .A2(n3144), .ZN(n3143) );
  NAND2_X1 U35560 ( .A1(n2719), .A2(n2720), .ZN(n2721) );
  NAND2_X1 U35570 ( .A1(n3143), .A2(n2721), .ZN(n3155) );
  OR2_X1 U35580 ( .A1(n3212), .A2(n2855), .ZN(n2723) );
  NAND2_X1 U35590 ( .A1(n3170), .A2(n2023), .ZN(n2722) );
  NAND2_X1 U35600 ( .A1(n2723), .A2(n2722), .ZN(n2727) );
  OAI22_X1 U35610 ( .A1(n3212), .A2(n2854), .B1(n2850), .B2(n2724), .ZN(n2725)
         );
  XNOR2_X1 U35620 ( .A(n2725), .B(n2837), .ZN(n2726) );
  XOR2_X1 U35630 ( .A(n2727), .B(n2726), .Z(n3154) );
  NAND2_X1 U35640 ( .A1(n3155), .A2(n3154), .ZN(n3153) );
  OAI22_X1 U35650 ( .A1(n3239), .A2(n2855), .B1(n2854), .B2(n3221), .ZN(n3188)
         );
  OAI22_X1 U35660 ( .A1(n3239), .A2(n2854), .B1(n2850), .B2(n3221), .ZN(n2729)
         );
  XNOR2_X1 U35670 ( .A(n2729), .B(n2837), .ZN(n3189) );
  OAI22_X1 U35680 ( .A1(n3213), .A2(n2854), .B1(n2850), .B2(n3179), .ZN(n2730)
         );
  XNOR2_X1 U35690 ( .A(n2730), .B(n2851), .ZN(n2733) );
  OR2_X1 U35700 ( .A1(n3213), .A2(n2855), .ZN(n2732) );
  NAND2_X1 U35710 ( .A1(n3242), .A2(n2023), .ZN(n2731) );
  NAND2_X1 U35720 ( .A1(n2732), .A2(n2731), .ZN(n2734) );
  XNOR2_X1 U35730 ( .A(n2733), .B(n2734), .ZN(n3236) );
  INV_X1 U35740 ( .A(n2733), .ZN(n2735) );
  OAI22_X1 U35750 ( .A1(n3276), .A2(n2854), .B1(n2850), .B2(n3254), .ZN(n2736)
         );
  XNOR2_X1 U35760 ( .A(n2736), .B(n2851), .ZN(n2740) );
  OR2_X1 U35770 ( .A1(n3276), .A2(n2855), .ZN(n2738) );
  NAND2_X1 U35780 ( .A1(n3202), .A2(n2871), .ZN(n2737) );
  AND2_X1 U35790 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NOR2_X1 U35800 ( .A1(n2740), .A2(n2739), .ZN(n3249) );
  NAND2_X1 U35810 ( .A1(n2740), .A2(n2739), .ZN(n3247) );
  OAI21_X1 U3582 ( .B1(n3246), .B2(n3249), .A(n3247), .ZN(n3273) );
  OAI22_X1 U3583 ( .A1(n3299), .A2(n2855), .B1(n2854), .B2(n3262), .ZN(n2745)
         );
  NAND2_X1 U3584 ( .A1(n3674), .A2(n2023), .ZN(n2742) );
  NAND2_X1 U3585 ( .A1(n3279), .A2(n2689), .ZN(n2741) );
  NAND2_X1 U3586 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  XNOR2_X1 U3587 ( .A(n2743), .B(n2837), .ZN(n2744) );
  XOR2_X1 U3588 ( .A(n2745), .B(n2744), .Z(n3274) );
  INV_X1 U3589 ( .A(n2744), .ZN(n2747) );
  INV_X1 U3590 ( .A(n2745), .ZN(n2746) );
  NAND2_X1 U3591 ( .A1(n4105), .A2(n2023), .ZN(n2749) );
  NAND2_X1 U3592 ( .A1(n3301), .A2(n2689), .ZN(n2748) );
  NAND2_X1 U3593 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  XNOR2_X1 U3594 ( .A(n2750), .B(n2837), .ZN(n2751) );
  AOI22_X1 U3595 ( .A1(n4105), .A2(n2841), .B1(n2023), .B2(n3301), .ZN(n2752)
         );
  XNOR2_X1 U3596 ( .A(n2751), .B(n2752), .ZN(n3297) );
  INV_X1 U3597 ( .A(n2751), .ZN(n2753) );
  OR2_X1 U3598 ( .A1(n2753), .A2(n2752), .ZN(n2754) );
  OAI22_X1 U3599 ( .A1(n3307), .A2(n2855), .B1(n2854), .B2(n4110), .ZN(n3327)
         );
  OAI22_X1 U3600 ( .A1(n3307), .A2(n2854), .B1(n2850), .B2(n4110), .ZN(n2755)
         );
  XNOR2_X1 U3601 ( .A(n2755), .B(n2837), .ZN(n3328) );
  OAI22_X1 U3602 ( .A1(n4101), .A2(n2854), .B1(n2850), .B2(n3400), .ZN(n2756)
         );
  XNOR2_X1 U3603 ( .A(n2756), .B(n2851), .ZN(n2762) );
  INV_X1 U3604 ( .A(n2762), .ZN(n2760) );
  OR2_X1 U3605 ( .A1(n4101), .A2(n2855), .ZN(n2758) );
  NAND2_X1 U3606 ( .A1(n3313), .A2(n2023), .ZN(n2757) );
  INV_X1 U3607 ( .A(n2761), .ZN(n2759) );
  NAND2_X1 U3608 ( .A1(n2760), .A2(n2759), .ZN(n3395) );
  OAI22_X1 U3609 ( .A1(n3613), .A2(n2854), .B1(n2850), .B2(n4088), .ZN(n2763)
         );
  XNOR2_X1 U3610 ( .A(n2763), .B(n2837), .ZN(n3458) );
  OAI22_X1 U3611 ( .A1(n3613), .A2(n2855), .B1(n2854), .B2(n4088), .ZN(n3457)
         );
  OAI21_X2 U3612 ( .B1(n3456), .B2(n3458), .A(n3457), .ZN(n2765) );
  NAND2_X1 U3613 ( .A1(n3456), .A2(n3458), .ZN(n2764) );
  OAI22_X1 U3614 ( .A1(n3514), .A2(n2854), .B1(n2850), .B2(n4052), .ZN(n2766)
         );
  XNOR2_X1 U3615 ( .A(n2766), .B(n2851), .ZN(n2770) );
  OR2_X1 U3616 ( .A1(n3514), .A2(n2855), .ZN(n2768) );
  NAND2_X1 U3617 ( .A1(n4061), .A2(n2022), .ZN(n2767) );
  NOR2_X1 U3618 ( .A1(n2770), .A2(n2769), .ZN(n3360) );
  NAND2_X1 U3619 ( .A1(n2770), .A2(n2769), .ZN(n3359) );
  OAI22_X1 U3620 ( .A1(n4053), .A2(n2854), .B1(n2850), .B2(n4042), .ZN(n2771)
         );
  XOR2_X1 U3621 ( .A(n2837), .B(n2771), .Z(n2774) );
  OR2_X1 U3622 ( .A1(n4053), .A2(n2855), .ZN(n2773) );
  NAND2_X1 U3623 ( .A1(n3518), .A2(n2022), .ZN(n2772) );
  NAND2_X1 U3624 ( .A1(n2773), .A2(n2772), .ZN(n3508) );
  OAI22_X1 U3625 ( .A1(n4036), .A2(n2854), .B1(n2850), .B2(n3421), .ZN(n2775)
         );
  XNOR2_X1 U3626 ( .A(n2775), .B(n2837), .ZN(n2779) );
  OR2_X1 U3627 ( .A1(n4036), .A2(n2855), .ZN(n2777) );
  NAND2_X1 U3628 ( .A1(n4029), .A2(n2871), .ZN(n2776) );
  NAND2_X1 U3629 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  NOR2_X1 U3630 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  OAI22_X1 U3631 ( .A1(n3987), .A2(n2854), .B1(n2850), .B2(n4012), .ZN(n2781)
         );
  XNOR2_X1 U3632 ( .A(n2781), .B(n2837), .ZN(n2785) );
  OR2_X1 U3633 ( .A1(n3987), .A2(n2855), .ZN(n2783) );
  NAND2_X1 U3634 ( .A1(n4005), .A2(n2022), .ZN(n2782) );
  NAND2_X1 U3635 ( .A1(n2783), .A2(n2782), .ZN(n2784) );
  NAND2_X1 U3636 ( .A1(n2785), .A2(n2784), .ZN(n3427) );
  NOR2_X1 U3637 ( .A1(n2785), .A2(n2784), .ZN(n3429) );
  OAI22_X1 U3638 ( .A1(n3974), .A2(n2855), .B1(n2854), .B2(n2786), .ZN(n3483)
         );
  OAI22_X1 U3639 ( .A1(n3974), .A2(n2854), .B1(n2850), .B2(n2786), .ZN(n2787)
         );
  XNOR2_X1 U3640 ( .A(n2787), .B(n2837), .ZN(n3484) );
  OAI22_X1 U3641 ( .A1(n3947), .A2(n2854), .B1(n2850), .B2(n3975), .ZN(n2788)
         );
  XOR2_X1 U3642 ( .A(n2837), .B(n2788), .Z(n2790) );
  AOI22_X1 U3643 ( .A1(n3985), .A2(n2841), .B1(n2023), .B2(n3970), .ZN(n2789)
         );
  NAND2_X1 U3644 ( .A1(n2790), .A2(n2789), .ZN(n2792) );
  OAI21_X1 U3645 ( .B1(n2790), .B2(n2789), .A(n2792), .ZN(n3379) );
  NAND2_X1 U3646 ( .A1(n3377), .A2(n2792), .ZN(n3445) );
  OAI22_X1 U3647 ( .A1(n3923), .A2(n2854), .B1(n2850), .B2(n3952), .ZN(n2793)
         );
  XNOR2_X1 U3648 ( .A(n2793), .B(n2837), .ZN(n2794) );
  OAI22_X1 U3649 ( .A1(n3923), .A2(n2855), .B1(n2854), .B2(n3952), .ZN(n2795)
         );
  NAND2_X1 U3650 ( .A1(n2794), .A2(n2795), .ZN(n3446) );
  INV_X1 U3651 ( .A(n2794), .ZN(n2797) );
  INV_X1 U3652 ( .A(n2795), .ZN(n2796) );
  NAND2_X1 U3653 ( .A1(n2797), .A2(n2796), .ZN(n3448) );
  OAI22_X1 U3654 ( .A1(n3908), .A2(n2854), .B1(n2850), .B2(n3930), .ZN(n2798)
         );
  XNOR2_X1 U3655 ( .A(n2798), .B(n2851), .ZN(n2803) );
  OR2_X1 U3656 ( .A1(n3908), .A2(n2855), .ZN(n2801) );
  NAND2_X1 U3657 ( .A1(n2799), .A2(n2022), .ZN(n2800) );
  NAND2_X1 U3658 ( .A1(n2801), .A2(n2800), .ZN(n2804) );
  INV_X1 U3659 ( .A(n2804), .ZN(n2802) );
  INV_X1 U3660 ( .A(n2803), .ZN(n2805) );
  NAND2_X1 U3661 ( .A1(n2805), .A2(n2804), .ZN(n3385) );
  NAND2_X1 U3662 ( .A1(n3925), .A2(n2871), .ZN(n2807) );
  NAND2_X1 U3663 ( .A1(n2548), .A2(n2689), .ZN(n2806) );
  NAND2_X1 U3664 ( .A1(n2807), .A2(n2806), .ZN(n2808) );
  XNOR2_X1 U3665 ( .A(n2808), .B(n2837), .ZN(n2811) );
  OAI22_X1 U3666 ( .A1(n3891), .A2(n2855), .B1(n2854), .B2(n3913), .ZN(n2810)
         );
  XNOR2_X1 U3667 ( .A(n2811), .B(n2810), .ZN(n3466) );
  OAI22_X1 U3668 ( .A1(n3865), .A2(n2854), .B1(n2850), .B2(n3893), .ZN(n2809)
         );
  XNOR2_X1 U3669 ( .A(n2809), .B(n2837), .ZN(n2813) );
  OAI22_X1 U3670 ( .A1(n3865), .A2(n2855), .B1(n2854), .B2(n3893), .ZN(n2812)
         );
  XNOR2_X1 U3671 ( .A(n2813), .B(n2812), .ZN(n3368) );
  NOR2_X1 U3672 ( .A1(n2811), .A2(n2810), .ZN(n3369) );
  NAND2_X1 U3673 ( .A1(n2813), .A2(n2812), .ZN(n2817) );
  AND2_X1 U3674 ( .A1(n2814), .A2(n2871), .ZN(n2815) );
  AOI21_X1 U3675 ( .B1(n3888), .B2(n2841), .A(n2815), .ZN(n2818) );
  OAI22_X1 U3676 ( .A1(n3847), .A2(n2854), .B1(n2850), .B2(n3871), .ZN(n2816)
         );
  XNOR2_X1 U3677 ( .A(n2816), .B(n2837), .ZN(n3438) );
  NAND2_X1 U3678 ( .A1(n3436), .A2(n3438), .ZN(n2821) );
  NAND2_X1 U3679 ( .A1(n3370), .A2(n2817), .ZN(n2820) );
  INV_X1 U3680 ( .A(n2818), .ZN(n2819) );
  NAND2_X1 U3681 ( .A1(n2820), .A2(n2819), .ZN(n3435) );
  NAND2_X1 U3682 ( .A1(n2821), .A2(n3435), .ZN(n3405) );
  NAND2_X1 U3683 ( .A1(n3867), .A2(n2022), .ZN(n2823) );
  NAND2_X1 U3684 ( .A1(n2825), .A2(n2689), .ZN(n2822) );
  NAND2_X1 U3685 ( .A1(n2823), .A2(n2822), .ZN(n2824) );
  XNOR2_X1 U3686 ( .A(n2824), .B(n2851), .ZN(n2828) );
  AND2_X1 U3687 ( .A1(n2825), .A2(n2871), .ZN(n2826) );
  AOI21_X1 U3688 ( .B1(n3867), .B2(n2841), .A(n2826), .ZN(n2827) );
  NAND2_X1 U3689 ( .A1(n2828), .A2(n2827), .ZN(n3406) );
  NOR2_X1 U3690 ( .A1(n2828), .A2(n2827), .ZN(n3408) );
  OAI22_X1 U3691 ( .A1(n3803), .A2(n2854), .B1(n2850), .B2(n3835), .ZN(n2829)
         );
  XNOR2_X1 U3692 ( .A(n2829), .B(n2851), .ZN(n2834) );
  INV_X1 U3693 ( .A(n2834), .ZN(n2832) );
  NOR2_X1 U3694 ( .A1(n3835), .A2(n2854), .ZN(n2830) );
  AOI21_X1 U3695 ( .B1(n3849), .B2(n2841), .A(n2830), .ZN(n2833) );
  INV_X1 U3696 ( .A(n2833), .ZN(n2831) );
  NAND2_X1 U3697 ( .A1(n2832), .A2(n2831), .ZN(n3493) );
  AND2_X1 U3698 ( .A1(n2834), .A2(n2833), .ZN(n3492) );
  NAND2_X1 U3699 ( .A1(n3830), .A2(n2871), .ZN(n2836) );
  NAND2_X1 U3700 ( .A1(n2839), .A2(n2689), .ZN(n2835) );
  NAND2_X1 U3701 ( .A1(n2836), .A2(n2835), .ZN(n2838) );
  XNOR2_X1 U3702 ( .A(n2838), .B(n2837), .ZN(n2860) );
  AND2_X1 U3703 ( .A1(n2839), .A2(n2871), .ZN(n2840) );
  AOI21_X1 U3704 ( .B1(n3830), .B2(n2841), .A(n2840), .ZN(n2858) );
  XNOR2_X1 U3705 ( .A(n2860), .B(n2858), .ZN(n3337) );
  NAND2_X1 U3706 ( .A1(n3339), .A2(n3337), .ZN(n2861) );
  INV_X1 U3707 ( .A(n2842), .ZN(n2843) );
  NAND2_X1 U3708 ( .A1(n2843), .A2(D_REG_1__SCAN_IN), .ZN(n2845) );
  INV_X1 U3709 ( .A(n2844), .ZN(n2916) );
  AOI21_X1 U3710 ( .B1(n2846), .B2(n2845), .A(n2916), .ZN(n3066) );
  OAI211_X1 U3711 ( .C1(n3042), .C2(n3775), .A(n4099), .B(n2848), .ZN(n2873)
         );
  NOR2_X1 U3712 ( .A1(n2957), .A2(n2873), .ZN(n2849) );
  OAI22_X1 U3713 ( .A1(n3790), .A2(n2854), .B1(n2850), .B2(n2853), .ZN(n2852)
         );
  XNOR2_X1 U3714 ( .A(n2852), .B(n2851), .ZN(n2857) );
  OAI22_X1 U3715 ( .A1(n3790), .A2(n2855), .B1(n2854), .B2(n2853), .ZN(n2856)
         );
  XNOR2_X1 U3716 ( .A(n2857), .B(n2856), .ZN(n2864) );
  INV_X1 U3717 ( .A(n2858), .ZN(n2859) );
  NAND2_X1 U3718 ( .A1(n2860), .A2(n2859), .ZN(n2865) );
  NAND4_X1 U3719 ( .A1(n2861), .A2(n3510), .A3(n2864), .A4(n2865), .ZN(n2890)
         );
  INV_X1 U3720 ( .A(n2861), .ZN(n2863) );
  INV_X1 U3721 ( .A(n2864), .ZN(n2862) );
  NAND2_X1 U3722 ( .A1(n2863), .A2(n2273), .ZN(n2889) );
  INV_X1 U3723 ( .A(n2865), .ZN(n2866) );
  NAND3_X1 U3724 ( .A1(n2862), .A2(n3510), .A3(n2866), .ZN(n2887) );
  INV_X1 U3725 ( .A(n2868), .ZN(n2869) );
  AND2_X1 U3726 ( .A1(n4394), .A2(n2869), .ZN(n2870) );
  NAND2_X1 U3727 ( .A1(n2023), .A2(n2870), .ZN(n2877) );
  NOR2_X1 U3728 ( .A1(n2882), .A2(n2877), .ZN(n2879) );
  INV_X1 U3729 ( .A(n2879), .ZN(n2872) );
  NAND2_X1 U3730 ( .A1(n2873), .A2(n4099), .ZN(n2874) );
  NAND2_X1 U3731 ( .A1(n2882), .A2(n2874), .ZN(n2875) );
  NAND2_X1 U3732 ( .A1(n2875), .A2(n3064), .ZN(n3017) );
  NAND2_X1 U3733 ( .A1(n2892), .A2(n2958), .ZN(n2876) );
  OAI21_X1 U3734 ( .B1(n3017), .B2(n2876), .A(STATE_REG_SCAN_IN), .ZN(n2878)
         );
  INV_X1 U3735 ( .A(n2877), .ZN(n3665) );
  NAND2_X1 U3736 ( .A1(n2882), .A2(n3665), .ZN(n3015) );
  NOR2_X1 U3737 ( .A1(n3521), .A2(n3352), .ZN(n2885) );
  NAND2_X1 U3738 ( .A1(n3065), .A2(n4129), .ZN(n2881) );
  OAI21_X2 U3739 ( .B1(n2882), .B2(n2881), .A(n4370), .ZN(n3517) );
  AOI22_X1 U3740 ( .A1(n3517), .A2(n3779), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2883) );
  OAI21_X1 U3741 ( .B1(n3524), .B2(n3513), .A(n2883), .ZN(n2884) );
  AOI211_X1 U3742 ( .C1(n3499), .C2(n3830), .A(n2885), .B(n2884), .ZN(n2886)
         );
  NAND3_X1 U3743 ( .A1(n2890), .A2(n2889), .A3(n2888), .ZN(U3217) );
  INV_X1 U3744 ( .A(n4394), .ZN(n2891) );
  MUX2_X1 U3745 ( .A(n2987), .B(n2358), .S(U3149), .Z(n2893) );
  INV_X1 U3746 ( .A(n2893), .ZN(U3347) );
  INV_X1 U3747 ( .A(n3743), .ZN(n3769) );
  NAND2_X1 U3748 ( .A1(n3769), .A2(STATE_REG_SCAN_IN), .ZN(n2894) );
  OAI21_X1 U3749 ( .B1(STATE_REG_SCAN_IN), .B2(n2505), .A(n2894), .ZN(U3335)
         );
  INV_X1 U3750 ( .A(DATAI_21_), .ZN(n2896) );
  NAND2_X1 U3751 ( .A1(n3657), .A2(STATE_REG_SCAN_IN), .ZN(n2895) );
  OAI21_X1 U3752 ( .B1(STATE_REG_SCAN_IN), .B2(n2896), .A(n2895), .ZN(U3331)
         );
  INV_X1 U3753 ( .A(DATAI_20_), .ZN(n2898) );
  NAND2_X1 U3754 ( .A1(n3660), .A2(STATE_REG_SCAN_IN), .ZN(n2897) );
  OAI21_X1 U3755 ( .B1(STATE_REG_SCAN_IN), .B2(n2898), .A(n2897), .ZN(U3332)
         );
  INV_X1 U3756 ( .A(DATAI_22_), .ZN(n2900) );
  NAND2_X1 U3757 ( .A1(n3667), .A2(STATE_REG_SCAN_IN), .ZN(n2899) );
  OAI21_X1 U3758 ( .B1(STATE_REG_SCAN_IN), .B2(n2900), .A(n2899), .ZN(U3330)
         );
  INV_X1 U3759 ( .A(DATAI_24_), .ZN(n2903) );
  NAND2_X1 U3760 ( .A1(n2901), .A2(STATE_REG_SCAN_IN), .ZN(n2902) );
  OAI21_X1 U3761 ( .B1(STATE_REG_SCAN_IN), .B2(n2903), .A(n2902), .ZN(U3328)
         );
  INV_X1 U3762 ( .A(DATAI_26_), .ZN(n4583) );
  NAND2_X1 U3763 ( .A1(n2652), .A2(STATE_REG_SCAN_IN), .ZN(n2904) );
  OAI21_X1 U3764 ( .B1(STATE_REG_SCAN_IN), .B2(n4583), .A(n2904), .ZN(U3326)
         );
  INV_X1 U3765 ( .A(DATAI_25_), .ZN(n2907) );
  NAND2_X1 U3766 ( .A1(n2905), .A2(STATE_REG_SCAN_IN), .ZN(n2906) );
  OAI21_X1 U3767 ( .B1(STATE_REG_SCAN_IN), .B2(n2907), .A(n2906), .ZN(U3327)
         );
  INV_X1 U3768 ( .A(DATAI_30_), .ZN(n2910) );
  NAND2_X1 U3769 ( .A1(n2908), .A2(STATE_REG_SCAN_IN), .ZN(n2909) );
  OAI21_X1 U3770 ( .B1(STATE_REG_SCAN_IN), .B2(n2910), .A(n2909), .ZN(U3322)
         );
  INV_X1 U3771 ( .A(DATAI_27_), .ZN(n2913) );
  XNOR2_X1 U3772 ( .A(n2911), .B(IR_REG_27__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U3773 ( .A1(n3787), .A2(STATE_REG_SCAN_IN), .ZN(n2912) );
  OAI21_X1 U3774 ( .B1(STATE_REG_SCAN_IN), .B2(n2913), .A(n2912), .ZN(U3325)
         );
  AOI22_X1 U3775 ( .A1(n4393), .A2(n4596), .B1(n2915), .B2(n4394), .ZN(U3458)
         );
  INV_X1 U3776 ( .A(D_REG_1__SCAN_IN), .ZN(n2917) );
  AOI22_X1 U3777 ( .A1(n4393), .A2(n2917), .B1(n2916), .B2(n4394), .ZN(U3459)
         );
  INV_X1 U3778 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n2923) );
  INV_X1 U3779 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2921) );
  NAND2_X1 U3780 ( .A1(n2350), .A2(REG2_REG_30__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3781 ( .A1(n2918), .A2(REG0_REG_30__SCAN_IN), .ZN(n2919) );
  OAI211_X1 U3782 ( .C1(n2507), .C2(n2921), .A(n2920), .B(n2919), .ZN(n3788)
         );
  NAND2_X1 U3783 ( .A1(n3788), .A2(n3679), .ZN(n2922) );
  OAI21_X1 U3784 ( .B1(n3679), .B2(n2923), .A(n2922), .ZN(U3580) );
  INV_X1 U3785 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n2925) );
  NAND2_X1 U3786 ( .A1(n2708), .A2(n3679), .ZN(n2924) );
  OAI21_X1 U3787 ( .B1(U4043), .B2(n2925), .A(n2924), .ZN(U3553) );
  INV_X1 U3788 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U3789 ( .A1(n3264), .A2(n3679), .ZN(n2926) );
  OAI21_X1 U3790 ( .B1(U4043), .B2(n2927), .A(n2926), .ZN(U3558) );
  INV_X1 U3791 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U3792 ( .A1(n3419), .A2(U4043), .ZN(n2928) );
  OAI21_X1 U3793 ( .B1(U4043), .B2(n2929), .A(n2928), .ZN(U3565) );
  INV_X1 U3794 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3795 ( .A1(n4079), .A2(n3679), .ZN(n2930) );
  OAI21_X1 U3796 ( .B1(U4043), .B2(n2931), .A(n2930), .ZN(U3564) );
  INV_X1 U3797 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n2933) );
  NAND2_X1 U3798 ( .A1(n3252), .A2(U4043), .ZN(n2932) );
  OAI21_X1 U3799 ( .B1(U4043), .B2(n2933), .A(n2932), .ZN(U3557) );
  INV_X1 U3800 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n2935) );
  NAND2_X1 U3801 ( .A1(n3971), .A2(n3679), .ZN(n2934) );
  OAI21_X1 U3802 ( .B1(U4043), .B2(n2935), .A(n2934), .ZN(U3570) );
  INV_X1 U3803 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n2937) );
  NAND2_X1 U3804 ( .A1(n4006), .A2(n3679), .ZN(n2936) );
  OAI21_X1 U3805 ( .B1(n3679), .B2(n2937), .A(n2936), .ZN(U3568) );
  INV_X1 U3806 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n2939) );
  NAND2_X1 U3807 ( .A1(n3985), .A2(n3679), .ZN(n2938) );
  OAI21_X1 U3808 ( .B1(n3679), .B2(n2939), .A(n2938), .ZN(U3569) );
  INV_X1 U3809 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U3810 ( .A1(n4055), .A2(n3679), .ZN(n2940) );
  OAI21_X1 U3811 ( .B1(U4043), .B2(n2941), .A(n2940), .ZN(U3563) );
  NAND2_X1 U3812 ( .A1(n3681), .A2(DATAO_REG_29__SCAN_IN), .ZN(n2942) );
  OAI21_X1 U3813 ( .B1(n3524), .B2(n3681), .A(n2942), .ZN(U3579) );
  XNOR2_X1 U3814 ( .A(n4275), .B(REG1_REG_2__SCAN_IN), .ZN(n3708) );
  INV_X1 U3815 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4534) );
  XNOR2_X1 U3816 ( .A(n4276), .B(n4534), .ZN(n3695) );
  AND2_X1 U3817 ( .A1(n4409), .A2(REG1_REG_0__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U3818 ( .A1(n4276), .A2(REG1_REG_1__SCAN_IN), .ZN(n2943) );
  NAND2_X1 U3819 ( .A1(n4275), .A2(REG1_REG_2__SCAN_IN), .ZN(n2944) );
  INV_X1 U3820 ( .A(n4274), .ZN(n3029) );
  NAND2_X1 U3821 ( .A1(n3023), .A2(REG1_REG_3__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U3822 ( .A1(n2945), .A2(n4274), .ZN(n2946) );
  NAND2_X1 U3823 ( .A1(n2949), .A2(n4273), .ZN(n2950) );
  MUX2_X1 U3824 ( .A(n2951), .B(REG1_REG_5__SCAN_IN), .S(n2987), .Z(n2991) );
  NAND2_X1 U3825 ( .A1(n2990), .A2(n2991), .ZN(n2989) );
  OR2_X1 U3826 ( .A1(n2987), .A2(n2951), .ZN(n2952) );
  NAND2_X1 U3827 ( .A1(n2989), .A2(n2952), .ZN(n2953) );
  XNOR2_X1 U3828 ( .A(n2953), .B(n2167), .ZN(n3046) );
  AND2_X1 U3829 ( .A1(n2953), .A2(n4272), .ZN(n2954) );
  AOI21_X1 U3830 ( .B1(n3046), .B2(REG1_REG_6__SCAN_IN), .A(n2954), .ZN(n3005)
         );
  XOR2_X1 U3831 ( .A(n2373), .B(n4271), .Z(n2955) );
  XNOR2_X1 U3832 ( .A(n3005), .B(n2955), .ZN(n2983) );
  INV_X1 U3833 ( .A(n2958), .ZN(n2956) );
  NAND2_X1 U3834 ( .A1(n2956), .A2(STATE_REG_SCAN_IN), .ZN(n3669) );
  NAND2_X1 U3835 ( .A1(n2957), .A2(n3669), .ZN(n2961) );
  NAND2_X1 U3836 ( .A1(n2959), .A2(n2958), .ZN(n2960) );
  AND2_X1 U3837 ( .A1(n3528), .A2(n2960), .ZN(n2962) );
  INV_X1 U3838 ( .A(n3787), .ZN(n3703) );
  INV_X1 U3839 ( .A(n2961), .ZN(n2963) );
  NOR2_X1 U3840 ( .A1(STATE_REG_SCAN_IN), .A2(n4484), .ZN(n3241) );
  INV_X1 U3841 ( .A(n4271), .ZN(n2997) );
  NOR2_X1 U3842 ( .A1(n4468), .A2(n2997), .ZN(n2964) );
  AOI211_X1 U3843 ( .C1(n4461), .C2(ADDR_REG_7__SCAN_IN), .A(n3241), .B(n2964), 
        .ZN(n2982) );
  INV_X1 U3844 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3077) );
  MUX2_X1 U3845 ( .A(REG2_REG_2__SCAN_IN), .B(n3077), .S(n4275), .Z(n3712) );
  AND2_X1 U3846 ( .A1(n4409), .A2(REG2_REG_0__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U3847 ( .A1(n4276), .A2(REG2_REG_1__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U3848 ( .A1(n3691), .A2(n2965), .ZN(n3711) );
  NAND2_X1 U3849 ( .A1(n4275), .A2(REG2_REG_2__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3850 ( .A1(n3710), .A2(n2966), .ZN(n2967) );
  NAND2_X1 U3851 ( .A1(n3024), .A2(REG2_REG_3__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3852 ( .A1(n2967), .A2(n4274), .ZN(n2968) );
  NAND2_X1 U3853 ( .A1(n2969), .A2(n2968), .ZN(n2970) );
  XNOR2_X1 U3854 ( .A(n2970), .B(n4273), .ZN(n3716) );
  INV_X1 U3855 ( .A(n2970), .ZN(n2972) );
  INV_X1 U3856 ( .A(n4273), .ZN(n2971) );
  MUX2_X1 U3857 ( .A(REG2_REG_5__SCAN_IN), .B(n3168), .S(n2987), .Z(n2974) );
  OAI22_X1 U3858 ( .A1(n3047), .A2(n2976), .B1(n2975), .B2(n2167), .ZN(n2980)
         );
  MUX2_X1 U3859 ( .A(REG2_REG_7__SCAN_IN), .B(n2977), .S(n4271), .Z(n2979) );
  NOR2_X1 U3860 ( .A1(n4278), .A2(n3703), .ZN(n3664) );
  MUX2_X1 U3861 ( .A(n2977), .B(REG2_REG_7__SCAN_IN), .S(n4271), .Z(n2978) );
  OAI211_X1 U3862 ( .C1(n2980), .C2(n2979), .A(n4463), .B(n2996), .ZN(n2981)
         );
  OAI211_X1 U3863 ( .C1(n2983), .C2(n4455), .A(n2982), .B(n2981), .ZN(U3247)
         );
  MUX2_X1 U3864 ( .A(n3168), .B(REG2_REG_5__SCAN_IN), .S(n2987), .Z(n2985) );
  OAI21_X1 U3865 ( .B1(n2985), .B2(n2984), .A(n4463), .ZN(n2994) );
  NOR2_X1 U3866 ( .A1(n2986), .A2(STATE_REG_SCAN_IN), .ZN(n3157) );
  NOR2_X1 U3867 ( .A1(n4468), .A2(n2987), .ZN(n2988) );
  AOI211_X1 U3868 ( .C1(n4461), .C2(ADDR_REG_5__SCAN_IN), .A(n3157), .B(n2988), 
        .ZN(n2993) );
  OAI211_X1 U3869 ( .C1(n2991), .C2(n2990), .A(n4357), .B(n2989), .ZN(n2992)
         );
  OAI211_X1 U3870 ( .C1(n2995), .C2(n2994), .A(n2993), .B(n2992), .ZN(U3245)
         );
  NOR2_X1 U3871 ( .A1(n4461), .A2(U4043), .ZN(U3148) );
  INV_X1 U3872 ( .A(n4408), .ZN(n3007) );
  NAND2_X1 U3873 ( .A1(n2998), .A2(n3007), .ZN(n2999) );
  NAND2_X1 U3874 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4290), .ZN(n4289) );
  NAND2_X1 U3875 ( .A1(n2999), .A2(n4289), .ZN(n3001) );
  MUX2_X1 U3876 ( .A(n3269), .B(REG2_REG_9__SCAN_IN), .S(n3728), .Z(n3000) );
  OAI211_X1 U3877 ( .C1(n3001), .C2(n3000), .A(n3727), .B(n4463), .ZN(n3014)
         );
  NOR2_X1 U3878 ( .A1(STATE_REG_SCAN_IN), .A2(n3002), .ZN(n3278) );
  NAND2_X1 U3879 ( .A1(n4271), .A2(REG1_REG_7__SCAN_IN), .ZN(n3004) );
  NOR2_X1 U3880 ( .A1(n4271), .A2(REG1_REG_7__SCAN_IN), .ZN(n3003) );
  AOI21_X1 U3881 ( .B1(n3005), .B2(n3004), .A(n3003), .ZN(n3006) );
  AND2_X1 U3882 ( .A1(n3006), .A2(n3007), .ZN(n3008) );
  MUX2_X1 U3883 ( .A(REG1_REG_9__SCAN_IN), .B(n3009), .S(n3728), .Z(n3010) );
  AOI211_X1 U3884 ( .C1(n3011), .C2(n3010), .A(n3744), .B(n4455), .ZN(n3012)
         );
  AOI211_X1 U3885 ( .C1(n4461), .C2(ADDR_REG_9__SCAN_IN), .A(n3278), .B(n3012), 
        .ZN(n3013) );
  OAI211_X1 U3886 ( .C1(n4468), .C2(n3728), .A(n3014), .B(n3013), .ZN(U3249)
         );
  NAND2_X1 U3887 ( .A1(n3015), .A2(n3065), .ZN(n3016) );
  OR2_X1 U3888 ( .A1(n3017), .A2(n3016), .ZN(n3477) );
  INV_X1 U3889 ( .A(n3477), .ZN(n3057) );
  XOR2_X1 U3890 ( .A(n3019), .B(n3018), .Z(n3700) );
  NAND2_X1 U3891 ( .A1(n3700), .A2(n3510), .ZN(n3021) );
  INV_X1 U3892 ( .A(n3513), .ZN(n3478) );
  AOI22_X1 U3893 ( .A1(n3478), .A2(n3680), .B1(n2690), .B2(n3517), .ZN(n3020)
         );
  OAI211_X1 U3894 ( .C1(n3057), .C2(n3022), .A(n3021), .B(n3020), .ZN(U3229)
         );
  XOR2_X1 U3895 ( .A(REG1_REG_3__SCAN_IN), .B(n3023), .Z(n3026) );
  XOR2_X1 U3896 ( .A(REG2_REG_3__SCAN_IN), .B(n3024), .Z(n3025) );
  AOI22_X1 U3897 ( .A1(n4357), .A2(n3026), .B1(n4463), .B2(n3025), .ZN(n3028)
         );
  INV_X1 U3898 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3093) );
  NOR2_X1 U3899 ( .A1(STATE_REG_SCAN_IN), .A2(n3093), .ZN(n3114) );
  AOI21_X1 U3900 ( .B1(n4461), .B2(ADDR_REG_3__SCAN_IN), .A(n3114), .ZN(n3027)
         );
  OAI211_X1 U3901 ( .C1(n3029), .C2(n4468), .A(n3028), .B(n3027), .ZN(U3243)
         );
  NAND2_X1 U3902 ( .A1(n3072), .A2(n3030), .ZN(n3034) );
  NAND2_X1 U3903 ( .A1(n2311), .A2(n4129), .ZN(n3032) );
  NAND2_X1 U3904 ( .A1(n2691), .A2(n4106), .ZN(n3031) );
  OAI211_X1 U3905 ( .C1(n3112), .C2(n4100), .A(n3032), .B(n3031), .ZN(n3033)
         );
  AOI21_X1 U3906 ( .B1(n3034), .B2(n4083), .A(n3033), .ZN(n3038) );
  INV_X1 U3907 ( .A(n3035), .ZN(n3036) );
  INV_X1 U3908 ( .A(n4102), .ZN(n3127) );
  NAND2_X1 U3909 ( .A1(n3141), .A2(n3127), .ZN(n3037) );
  NAND2_X1 U3910 ( .A1(n3038), .A2(n3037), .ZN(n3138) );
  INV_X1 U3911 ( .A(n3141), .ZN(n3039) );
  OAI21_X1 U3912 ( .B1(n3043), .B2(n2683), .A(n3078), .ZN(n3137) );
  OAI22_X1 U3913 ( .A1(n3039), .A2(n4416), .B1(n4415), .B2(n3137), .ZN(n3040)
         );
  NOR2_X1 U3914 ( .A1(n3138), .A2(n3040), .ZN(n4413) );
  NAND2_X1 U3915 ( .A1(n4452), .A2(REG1_REG_1__SCAN_IN), .ZN(n3041) );
  OAI21_X1 U3916 ( .B1(n4413), .B2(n4452), .A(n3041), .ZN(U3519) );
  NAND2_X1 U3917 ( .A1(n2691), .A2(n3043), .ZN(n3540) );
  NAND2_X1 U3918 ( .A1(n3538), .A2(n3540), .ZN(n4387) );
  NOR2_X1 U3919 ( .A1(n3043), .A2(n3042), .ZN(n4385) );
  OAI21_X1 U3920 ( .B1(n3127), .B2(n4083), .A(n4387), .ZN(n3044) );
  AOI211_X1 U3921 ( .C1(n4423), .C2(n4387), .A(n4385), .B(n4383), .ZN(n4412)
         );
  NAND2_X1 U3922 ( .A1(n4452), .A2(REG1_REG_0__SCAN_IN), .ZN(n3045) );
  OAI21_X1 U3923 ( .B1(n4412), .B2(n4452), .A(n3045), .ZN(U3518) );
  XNOR2_X1 U3924 ( .A(n3046), .B(REG1_REG_6__SCAN_IN), .ZN(n3052) );
  XNOR2_X1 U3925 ( .A(n3047), .B(REG2_REG_6__SCAN_IN), .ZN(n3050) );
  AND2_X1 U3926 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3193) );
  AOI21_X1 U3927 ( .B1(n4461), .B2(ADDR_REG_6__SCAN_IN), .A(n3193), .ZN(n3048)
         );
  OAI21_X1 U3928 ( .B1(n4468), .B2(n2167), .A(n3048), .ZN(n3049) );
  AOI21_X1 U3929 ( .B1(n3050), .B2(n4463), .A(n3049), .ZN(n3051) );
  OAI21_X1 U3930 ( .B1(n3052), .B2(n4455), .A(n3051), .ZN(U3246) );
  AOI211_X1 U3931 ( .C1(n3055), .C2(n3053), .A(n3505), .B(n3054), .ZN(n3060)
         );
  OAI22_X1 U3932 ( .A1(n3515), .A2(n3056), .B1(n3497), .B2(n2683), .ZN(n3059)
         );
  OAI22_X1 U3933 ( .A1(n3057), .A2(n2100), .B1(n3513), .B2(n3112), .ZN(n3058)
         );
  OR3_X1 U3934 ( .A1(n3060), .A2(n3059), .A3(n3058), .ZN(U3219) );
  OAI21_X1 U3935 ( .B1(n3063), .B2(n2610), .A(n3062), .ZN(n3101) );
  INV_X1 U3936 ( .A(n3101), .ZN(n3082) );
  NAND4_X1 U3937 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(n3068)
         );
  OR2_X1 U3938 ( .A1(n3069), .A2(n3775), .ZN(n3160) );
  INV_X1 U3939 ( .A(n3160), .ZN(n3070) );
  NAND2_X1 U3940 ( .A1(n4372), .A2(n3070), .ZN(n4120) );
  AOI22_X1 U3941 ( .A1(n2708), .A2(n4078), .B1(n4129), .B2(n3476), .ZN(n3071)
         );
  NAND3_X1 U3942 ( .A1(n2610), .A2(n2609), .A3(n3072), .ZN(n3073) );
  AOI21_X1 U3943 ( .B1(n3074), .B2(n3073), .A(n4109), .ZN(n3075) );
  AOI211_X1 U3944 ( .C1(n3127), .C2(n3101), .A(n3076), .B(n3075), .ZN(n3099)
         );
  MUX2_X1 U3945 ( .A(n3077), .B(n3099), .S(n4372), .Z(n3081) );
  NAND2_X1 U3946 ( .A1(n4372), .A2(n3775), .ZN(n3995) );
  AND2_X1 U3947 ( .A1(n3078), .A2(n3476), .ZN(n3079) );
  NOR2_X1 U3948 ( .A1(n3092), .A2(n3079), .ZN(n3106) );
  INV_X1 U3949 ( .A(n4370), .ZN(n4386) );
  AOI22_X1 U3950 ( .A1(n4377), .A2(n3106), .B1(REG3_REG_2__SCAN_IN), .B2(n4386), .ZN(n3080) );
  OAI211_X1 U3951 ( .C1(n3082), .C2(n4120), .A(n3081), .B(n3080), .ZN(U3288)
         );
  NAND2_X1 U3952 ( .A1(n3062), .A2(n3083), .ZN(n3084) );
  XNOR2_X1 U3953 ( .A(n3084), .B(n3617), .ZN(n4417) );
  OAI21_X1 U3954 ( .B1(n3617), .B2(n3086), .A(n3085), .ZN(n3089) );
  AOI22_X1 U3955 ( .A1(n3677), .A2(n4078), .B1(n4129), .B2(n3115), .ZN(n3087)
         );
  OAI21_X1 U3956 ( .B1(n3112), .B2(n4081), .A(n3087), .ZN(n3088) );
  AOI21_X1 U3957 ( .B1(n3089), .B2(n4083), .A(n3088), .ZN(n3090) );
  OAI21_X1 U3958 ( .B1(n4417), .B2(n4102), .A(n3090), .ZN(n4419) );
  INV_X1 U3959 ( .A(n4419), .ZN(n3098) );
  INV_X1 U3960 ( .A(n4417), .ZN(n3096) );
  INV_X1 U3961 ( .A(n4120), .ZN(n4388) );
  OAI21_X1 U3962 ( .B1(n3092), .B2(n3091), .A(n3130), .ZN(n4414) );
  AOI22_X1 U3963 ( .A1(n4391), .A2(REG2_REG_3__SCAN_IN), .B1(n4386), .B2(n3093), .ZN(n3094) );
  OAI21_X1 U3964 ( .B1(n4066), .B2(n4414), .A(n3094), .ZN(n3095) );
  AOI21_X1 U3965 ( .B1(n3096), .B2(n4388), .A(n3095), .ZN(n3097) );
  OAI21_X1 U3966 ( .B1(n3098), .B2(n4391), .A(n3097), .ZN(U3287) );
  INV_X1 U3967 ( .A(n3099), .ZN(n3100) );
  AOI21_X1 U3968 ( .B1(n4423), .B2(n3101), .A(n3100), .ZN(n3108) );
  INV_X1 U3969 ( .A(n4266), .ZN(n3103) );
  NOR2_X1 U3970 ( .A1(n4446), .A2(n2319), .ZN(n3102) );
  AOI21_X1 U3971 ( .B1(n3103), .B2(n3106), .A(n3102), .ZN(n3104) );
  OAI21_X1 U3972 ( .B1(n3108), .B2(n4444), .A(n3104), .ZN(U3471) );
  INV_X1 U3973 ( .A(n4208), .ZN(n3105) );
  AOI22_X1 U3974 ( .A1(n3106), .A2(n3105), .B1(REG1_REG_2__SCAN_IN), .B2(n4452), .ZN(n3107) );
  OAI21_X1 U3975 ( .B1(n3108), .B2(n4452), .A(n3107), .ZN(U3520) );
  XNOR2_X1 U3976 ( .A(n3110), .B(n3109), .ZN(n3111) );
  NAND2_X1 U3977 ( .A1(n3111), .A2(n3510), .ZN(n3117) );
  OAI22_X1 U3978 ( .A1(n3515), .A2(n3112), .B1(n3165), .B2(n3513), .ZN(n3113)
         );
  AOI211_X1 U3979 ( .C1(n3115), .C2(n3517), .A(n3114), .B(n3113), .ZN(n3116)
         );
  OAI211_X1 U3980 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3521), .A(n3117), .B(n3116), 
        .ZN(U3215) );
  AND2_X1 U3981 ( .A1(n2059), .A2(n3119), .ZN(n3121) );
  INV_X1 U3982 ( .A(n3120), .ZN(n3606) );
  NAND2_X1 U3983 ( .A1(n3121), .A2(n3606), .ZN(n3122) );
  INV_X1 U3984 ( .A(n4424), .ZN(n3136) );
  XOR2_X1 U3985 ( .A(n3606), .B(n3124), .Z(n3129) );
  AOI22_X1 U3986 ( .A1(n2708), .A2(n4106), .B1(n4129), .B2(n3149), .ZN(n3125)
         );
  OAI21_X1 U3987 ( .B1(n3212), .B2(n4100), .A(n3125), .ZN(n3126) );
  AOI21_X1 U3988 ( .B1(n4424), .B2(n3127), .A(n3126), .ZN(n3128) );
  OAI21_X1 U3989 ( .B1(n3129), .B2(n4109), .A(n3128), .ZN(n4421) );
  INV_X1 U3990 ( .A(n3130), .ZN(n3132) );
  OAI211_X1 U3991 ( .C1(n3132), .C2(n3131), .A(n4443), .B(n3169), .ZN(n4420)
         );
  OAI22_X1 U3992 ( .A1(n4420), .A2(n4269), .B1(n4370), .B2(n3152), .ZN(n3133)
         );
  OAI21_X1 U3993 ( .B1(n4421), .B2(n3133), .A(n4372), .ZN(n3135) );
  NAND2_X1 U3994 ( .A1(n4391), .A2(REG2_REG_4__SCAN_IN), .ZN(n3134) );
  OAI211_X1 U3995 ( .C1(n3136), .C2(n4120), .A(n3135), .B(n3134), .ZN(U3286)
         );
  OAI22_X1 U3996 ( .A1(n4066), .A2(n3137), .B1(n2100), .B2(n4370), .ZN(n3140)
         );
  MUX2_X1 U3997 ( .A(REG2_REG_1__SCAN_IN), .B(n3138), .S(n4372), .Z(n3139) );
  AOI211_X1 U3998 ( .C1(n4388), .C2(n3141), .A(n3140), .B(n3139), .ZN(n3142)
         );
  INV_X1 U3999 ( .A(n3142), .ZN(U3289) );
  OAI211_X1 U4000 ( .C1(n3145), .C2(n3144), .A(n3143), .B(n3510), .ZN(n3151)
         );
  NAND2_X1 U4001 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3718) );
  INV_X1 U4002 ( .A(n3718), .ZN(n3148) );
  OAI22_X1 U4003 ( .A1(n3515), .A2(n3146), .B1(n3212), .B2(n3513), .ZN(n3147)
         );
  AOI211_X1 U4004 ( .C1(n3149), .C2(n3517), .A(n3148), .B(n3147), .ZN(n3150)
         );
  OAI211_X1 U4005 ( .C1(n3521), .C2(n3152), .A(n3151), .B(n3150), .ZN(U3227)
         );
  OAI211_X1 U4006 ( .C1(n3155), .C2(n3154), .A(n3153), .B(n3510), .ZN(n3159)
         );
  OAI22_X1 U4007 ( .A1(n3515), .A2(n3165), .B1(n3239), .B2(n3513), .ZN(n3156)
         );
  AOI211_X1 U4008 ( .C1(n3170), .C2(n3517), .A(n3157), .B(n3156), .ZN(n3158)
         );
  OAI211_X1 U4009 ( .C1(n3521), .C2(n3171), .A(n3159), .B(n3158), .ZN(U3224)
         );
  NAND2_X1 U4010 ( .A1(n4102), .A2(n3160), .ZN(n3161) );
  NAND2_X1 U4011 ( .A1(n2045), .A2(n3556), .ZN(n3604) );
  XNOR2_X1 U4012 ( .A(n3162), .B(n3604), .ZN(n4426) );
  XNOR2_X1 U4013 ( .A(n3163), .B(n3604), .ZN(n3167) );
  AOI22_X1 U4014 ( .A1(n4078), .A2(n3675), .B1(n3170), .B2(n4129), .ZN(n3164)
         );
  OAI21_X1 U4015 ( .B1(n3165), .B2(n4081), .A(n3164), .ZN(n3166) );
  AOI21_X1 U4016 ( .B1(n3167), .B2(n4083), .A(n3166), .ZN(n4427) );
  MUX2_X1 U4017 ( .A(n4427), .B(n3168), .S(n4391), .Z(n3174) );
  AOI21_X1 U4018 ( .B1(n3170), .B2(n3169), .A(n3222), .ZN(n4430) );
  INV_X1 U4019 ( .A(n3171), .ZN(n3172) );
  AOI22_X1 U4020 ( .A1(n4430), .A2(n4377), .B1(n3172), .B2(n4386), .ZN(n3173)
         );
  OAI211_X1 U4021 ( .C1(n4035), .C2(n4426), .A(n3174), .B(n3173), .ZN(U3285)
         );
  XNOR2_X1 U4022 ( .A(n3175), .B(n3607), .ZN(n3178) );
  AOI22_X1 U4023 ( .A1(n3264), .A2(n4078), .B1(n4129), .B2(n3242), .ZN(n3176)
         );
  OAI21_X1 U4024 ( .B1(n3239), .B2(n4081), .A(n3176), .ZN(n3177) );
  AOI21_X1 U4025 ( .B1(n3178), .B2(n4083), .A(n3177), .ZN(n4436) );
  OAI211_X1 U4026 ( .C1(n3219), .C2(n3179), .A(n4443), .B(n3203), .ZN(n4435)
         );
  INV_X1 U4027 ( .A(n4435), .ZN(n3182) );
  INV_X1 U4028 ( .A(n3995), .ZN(n3181) );
  OAI22_X1 U4029 ( .A1(n4372), .A2(n2977), .B1(n3245), .B2(n4370), .ZN(n3180)
         );
  AOI21_X1 U4030 ( .B1(n3182), .B2(n3181), .A(n3180), .ZN(n3186) );
  NAND2_X1 U4031 ( .A1(n3184), .A2(n3607), .ZN(n4433) );
  NAND3_X1 U4032 ( .A1(n3183), .A2(n4433), .A3(n4068), .ZN(n3185) );
  OAI211_X1 U4033 ( .C1(n4436), .C2(n4391), .A(n3186), .B(n3185), .ZN(U3283)
         );
  XNOR2_X1 U4034 ( .A(n3189), .B(n3188), .ZN(n3190) );
  XNOR2_X1 U4035 ( .A(n3187), .B(n3190), .ZN(n3191) );
  NAND2_X1 U4036 ( .A1(n3191), .A2(n3510), .ZN(n3196) );
  OAI22_X1 U4037 ( .A1(n3515), .A2(n3212), .B1(n3213), .B2(n3513), .ZN(n3192)
         );
  AOI211_X1 U4038 ( .C1(n3194), .C2(n3517), .A(n3193), .B(n3192), .ZN(n3195)
         );
  OAI211_X1 U4039 ( .C1(n3521), .C2(n4371), .A(n3196), .B(n3195), .ZN(U3236)
         );
  NAND2_X1 U4040 ( .A1(n3557), .A2(n3536), .ZN(n3603) );
  XNOR2_X1 U4041 ( .A(n3197), .B(n3603), .ZN(n3200) );
  AOI22_X1 U4042 ( .A1(n4078), .A2(n3674), .B1(n3202), .B2(n4129), .ZN(n3198)
         );
  OAI21_X1 U40430 ( .B1(n3213), .B2(n4081), .A(n3198), .ZN(n3199) );
  AOI21_X1 U4044 ( .B1(n3200), .B2(n4083), .A(n3199), .ZN(n3228) );
  XNOR2_X1 U4045 ( .A(n3201), .B(n3603), .ZN(n3229) );
  INV_X1 U4046 ( .A(n3229), .ZN(n3208) );
  NAND2_X1 U4047 ( .A1(n3203), .A2(n3202), .ZN(n3204) );
  NAND2_X1 U4048 ( .A1(n3267), .A2(n3204), .ZN(n3232) );
  NOR2_X1 U4049 ( .A1(n3232), .A2(n4066), .ZN(n3207) );
  OAI22_X1 U4050 ( .A1(n4372), .A2(n3205), .B1(n3251), .B2(n4370), .ZN(n3206)
         );
  AOI211_X1 U4051 ( .C1(n3208), .C2(n4068), .A(n3207), .B(n3206), .ZN(n3209)
         );
  OAI21_X1 U4052 ( .B1(n4391), .B2(n3228), .A(n3209), .ZN(U3282) );
  NAND2_X1 U4053 ( .A1(n3553), .A2(n3554), .ZN(n3620) );
  XNOR2_X1 U4054 ( .A(n3210), .B(n3620), .ZN(n4374) );
  XOR2_X1 U4055 ( .A(n3620), .B(n3211), .Z(n3216) );
  NOR2_X1 U4056 ( .A1(n3212), .A2(n4081), .ZN(n3215) );
  OAI22_X1 U4057 ( .A1(n3213), .A2(n4100), .B1(n4099), .B2(n3221), .ZN(n3214)
         );
  AOI211_X1 U4058 ( .C1(n3216), .C2(n4083), .A(n3215), .B(n3214), .ZN(n3217)
         );
  OAI21_X1 U4059 ( .B1(n4102), .B2(n4374), .A(n3217), .ZN(n3218) );
  INV_X1 U4060 ( .A(n3218), .ZN(n4381) );
  OAI21_X1 U4061 ( .B1(n4416), .B2(n4374), .A(n4381), .ZN(n3226) );
  INV_X1 U4062 ( .A(n3219), .ZN(n3220) );
  OAI21_X1 U4063 ( .B1(n3222), .B2(n3221), .A(n3220), .ZN(n4375) );
  OAI22_X1 U4064 ( .A1(n4375), .A2(n4208), .B1(n4454), .B2(n2362), .ZN(n3223)
         );
  AOI21_X1 U4065 ( .B1(n3226), .B2(n4454), .A(n3223), .ZN(n3224) );
  INV_X1 U4066 ( .A(n3224), .ZN(U3524) );
  INV_X1 U4067 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4476) );
  OAI22_X1 U4068 ( .A1(n4375), .A2(n4266), .B1(n4446), .B2(n4476), .ZN(n3225)
         );
  AOI21_X1 U4069 ( .B1(n3226), .B2(n4446), .A(n3225), .ZN(n3227) );
  INV_X1 U4070 ( .A(n3227), .ZN(U3479) );
  OAI21_X1 U4071 ( .B1(n4438), .B2(n3229), .A(n3228), .ZN(n3234) );
  OAI22_X1 U4072 ( .A1(n3232), .A2(n4208), .B1(n4454), .B2(n2384), .ZN(n3230)
         );
  AOI21_X1 U4073 ( .B1(n3234), .B2(n4454), .A(n3230), .ZN(n3231) );
  INV_X1 U4074 ( .A(n3231), .ZN(U3526) );
  INV_X1 U4075 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4483) );
  OAI22_X1 U4076 ( .A1(n3232), .A2(n4266), .B1(n4446), .B2(n4483), .ZN(n3233)
         );
  AOI21_X1 U4077 ( .B1(n3234), .B2(n4446), .A(n3233), .ZN(n3235) );
  INV_X1 U4078 ( .A(n3235), .ZN(U3483) );
  XOR2_X1 U4079 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND2_X1 U4080 ( .A1(n3238), .A2(n3510), .ZN(n3244) );
  OAI22_X1 U4081 ( .A1(n3515), .A2(n3239), .B1(n3276), .B2(n3513), .ZN(n3240)
         );
  AOI211_X1 U4082 ( .C1(n3242), .C2(n3517), .A(n3241), .B(n3240), .ZN(n3243)
         );
  OAI211_X1 U4083 ( .C1(n3521), .C2(n3245), .A(n3244), .B(n3243), .ZN(U3210)
         );
  INV_X1 U4084 ( .A(n3247), .ZN(n3248) );
  NOR2_X1 U4085 ( .A1(n3249), .A2(n3248), .ZN(n3250) );
  XNOR2_X1 U4086 ( .A(n3246), .B(n3250), .ZN(n3258) );
  INV_X1 U4087 ( .A(n3251), .ZN(n3256) );
  AOI22_X1 U4088 ( .A1(n3478), .A2(n3674), .B1(n3499), .B2(n3252), .ZN(n3253)
         );
  NAND2_X1 U4089 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4286) );
  OAI211_X1 U4090 ( .C1(n3497), .C2(n3254), .A(n3253), .B(n4286), .ZN(n3255)
         );
  AOI21_X1 U4091 ( .B1(n3256), .B2(n3503), .A(n3255), .ZN(n3257) );
  OAI21_X1 U4092 ( .B1(n3258), .B2(n3505), .A(n3257), .ZN(U3218) );
  INV_X1 U4093 ( .A(n3565), .ZN(n3259) );
  NAND2_X1 U4094 ( .A1(n3259), .A2(n3558), .ZN(n3605) );
  XNOR2_X1 U4095 ( .A(n3260), .B(n3605), .ZN(n4439) );
  XOR2_X1 U4096 ( .A(n3605), .B(n3261), .Z(n3266) );
  OAI22_X1 U4097 ( .A1(n3332), .A2(n4100), .B1(n4099), .B2(n3262), .ZN(n3263)
         );
  AOI21_X1 U4098 ( .B1(n4106), .B2(n3264), .A(n3263), .ZN(n3265) );
  OAI21_X1 U4099 ( .B1(n3266), .B2(n4109), .A(n3265), .ZN(n4440) );
  NAND2_X1 U4100 ( .A1(n4440), .A2(n4372), .ZN(n3272) );
  AND2_X1 U4101 ( .A1(n3267), .A2(n3279), .ZN(n3268) );
  NOR2_X1 U4102 ( .A1(n3289), .A2(n3268), .ZN(n4442) );
  OAI22_X1 U4103 ( .A1(n4372), .A2(n3269), .B1(n3282), .B2(n4370), .ZN(n3270)
         );
  AOI21_X1 U4104 ( .B1(n4442), .B2(n4377), .A(n3270), .ZN(n3271) );
  OAI211_X1 U4105 ( .C1(n4439), .C2(n4035), .A(n3272), .B(n3271), .ZN(U3281)
         );
  XNOR2_X1 U4106 ( .A(n3273), .B(n3274), .ZN(n3275) );
  NAND2_X1 U4107 ( .A1(n3275), .A2(n3510), .ZN(n3281) );
  OAI22_X1 U4108 ( .A1(n3515), .A2(n3276), .B1(n3332), .B2(n3513), .ZN(n3277)
         );
  AOI211_X1 U4109 ( .C1(n3279), .C2(n3517), .A(n3278), .B(n3277), .ZN(n3280)
         );
  OAI211_X1 U4110 ( .C1(n3521), .C2(n3282), .A(n3281), .B(n3280), .ZN(U3228)
         );
  NAND2_X1 U4111 ( .A1(n3563), .A2(n3534), .ZN(n3600) );
  XNOR2_X1 U4112 ( .A(n3283), .B(n3600), .ZN(n3286) );
  OAI22_X1 U4113 ( .A1(n3307), .A2(n4100), .B1(n4099), .B2(n3288), .ZN(n3284)
         );
  AOI21_X1 U4114 ( .B1(n4106), .B2(n3674), .A(n3284), .ZN(n3285) );
  OAI21_X1 U4115 ( .B1(n3286), .B2(n4109), .A(n3285), .ZN(n3319) );
  INV_X1 U4116 ( .A(n3319), .ZN(n3295) );
  XNOR2_X1 U4117 ( .A(n3287), .B(n3600), .ZN(n3320) );
  NOR2_X1 U4118 ( .A1(n3289), .A2(n3288), .ZN(n3290) );
  OR2_X1 U4119 ( .A1(n4111), .A2(n3290), .ZN(n3325) );
  NOR2_X1 U4120 ( .A1(n3325), .A2(n4066), .ZN(n3293) );
  OAI22_X1 U4121 ( .A1(n4372), .A2(n3291), .B1(n3304), .B2(n4370), .ZN(n3292)
         );
  AOI211_X1 U4122 ( .C1(n3320), .C2(n4068), .A(n3293), .B(n3292), .ZN(n3294)
         );
  OAI21_X1 U4123 ( .B1(n3295), .B2(n4391), .A(n3294), .ZN(U3280) );
  OAI211_X1 U4124 ( .C1(n3298), .C2(n3297), .A(n3296), .B(n3510), .ZN(n3303)
         );
  AND2_X1 U4125 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4459) );
  OAI22_X1 U4126 ( .A1(n3515), .A2(n3299), .B1(n3307), .B2(n3513), .ZN(n3300)
         );
  AOI211_X1 U4127 ( .C1(n3301), .C2(n3517), .A(n4459), .B(n3300), .ZN(n3302)
         );
  OAI211_X1 U4128 ( .C1(n3521), .C2(n3304), .A(n3303), .B(n3302), .ZN(U3214)
         );
  INV_X1 U4129 ( .A(n4072), .ZN(n3305) );
  OR2_X1 U4130 ( .A1(n3305), .A2(n4073), .ZN(n3601) );
  INV_X1 U4131 ( .A(n3601), .ZN(n3306) );
  XNOR2_X1 U4132 ( .A(n4074), .B(n3306), .ZN(n3311) );
  OR2_X1 U4133 ( .A1(n3307), .A2(n4081), .ZN(n3309) );
  NAND2_X1 U4134 ( .A1(n3313), .A2(n4129), .ZN(n3308) );
  OAI211_X1 U4135 ( .C1(n3613), .C2(n4100), .A(n3309), .B(n3308), .ZN(n3310)
         );
  AOI21_X1 U4136 ( .B1(n3311), .B2(n4083), .A(n3310), .ZN(n4200) );
  XNOR2_X1 U4137 ( .A(n3312), .B(n3601), .ZN(n4199) );
  NAND2_X1 U4138 ( .A1(n4113), .A2(n3313), .ZN(n3314) );
  NAND2_X1 U4139 ( .A1(n4086), .A2(n3314), .ZN(n4262) );
  INV_X1 U4140 ( .A(n3315), .ZN(n3402) );
  AOI22_X1 U4141 ( .A1(n4391), .A2(REG2_REG_12__SCAN_IN), .B1(n3402), .B2(
        n4386), .ZN(n3316) );
  OAI21_X1 U4142 ( .B1(n4262), .B2(n4066), .A(n3316), .ZN(n3317) );
  AOI21_X1 U4143 ( .B1(n4199), .B2(n4068), .A(n3317), .ZN(n3318) );
  OAI21_X1 U4144 ( .B1(n4391), .B2(n4200), .A(n3318), .ZN(U3278) );
  INV_X1 U4145 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3321) );
  AOI21_X1 U4146 ( .B1(n4432), .B2(n3320), .A(n3319), .ZN(n3323) );
  MUX2_X1 U4147 ( .A(n3321), .B(n3323), .S(n4446), .Z(n3322) );
  OAI21_X1 U4148 ( .B1(n3325), .B2(n4266), .A(n3322), .ZN(U3487) );
  MUX2_X1 U4149 ( .A(n4458), .B(n3323), .S(n4454), .Z(n3324) );
  OAI21_X1 U4150 ( .B1(n4208), .B2(n3325), .A(n3324), .ZN(U3528) );
  XNOR2_X1 U4151 ( .A(n3328), .B(n3327), .ZN(n3329) );
  XNOR2_X1 U4152 ( .A(n3326), .B(n3329), .ZN(n3330) );
  NAND2_X1 U4153 ( .A1(n3330), .A2(n3510), .ZN(n3336) );
  NOR2_X1 U4154 ( .A1(STATE_REG_SCAN_IN), .A2(n3331), .ZN(n4296) );
  OAI22_X1 U4155 ( .A1(n3515), .A2(n3332), .B1(n4101), .B2(n3513), .ZN(n3333)
         );
  AOI211_X1 U4156 ( .C1(n3334), .C2(n3517), .A(n4296), .B(n3333), .ZN(n3335)
         );
  OAI211_X1 U4157 ( .C1(n3521), .C2(n4114), .A(n3336), .B(n3335), .ZN(U3233)
         );
  XNOR2_X1 U4158 ( .A(n3339), .B(n3338), .ZN(n3340) );
  NAND2_X1 U4159 ( .A1(n3340), .A2(n3510), .ZN(n3345) );
  OAI22_X1 U4160 ( .A1(n3497), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n3341), 
        .ZN(n3343) );
  OAI22_X1 U4161 ( .A1(n3790), .A2(n3513), .B1(n3803), .B2(n3515), .ZN(n3342)
         );
  AOI211_X1 U4162 ( .C1(n3814), .C2(n3503), .A(n3343), .B(n3342), .ZN(n3344)
         );
  NAND2_X1 U4163 ( .A1(n3345), .A2(n3344), .ZN(U3211) );
  NAND3_X1 U4164 ( .A1(n3347), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3349) );
  INV_X1 U4165 ( .A(DATAI_31_), .ZN(n3348) );
  OAI22_X1 U4166 ( .A1(n3346), .A2(n3349), .B1(STATE_REG_SCAN_IN), .B2(n3348), 
        .ZN(U3321) );
  INV_X1 U4167 ( .A(n3350), .ZN(n3356) );
  OAI22_X1 U4168 ( .A1(n3352), .A2(n4370), .B1(n3351), .B2(n4372), .ZN(n3355)
         );
  NOR2_X1 U4169 ( .A1(n3353), .A2(n4391), .ZN(n3354) );
  AOI211_X1 U4170 ( .C1(n4377), .C2(n3356), .A(n3355), .B(n3354), .ZN(n3357)
         );
  OAI21_X1 U4171 ( .B1(n3358), .B2(n4035), .A(n3357), .ZN(U3262) );
  NOR2_X1 U4172 ( .A1(n3360), .A2(n2246), .ZN(n3361) );
  XNOR2_X1 U4173 ( .A(n3362), .B(n3361), .ZN(n3367) );
  INV_X1 U4174 ( .A(n3363), .ZN(n4064) );
  AOI22_X1 U4175 ( .A1(n3478), .A2(n3419), .B1(n3499), .B2(n4055), .ZN(n3364)
         );
  NAND2_X1 U4176 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4334) );
  OAI211_X1 U4177 ( .C1(n3497), .C2(n4052), .A(n3364), .B(n4334), .ZN(n3365)
         );
  AOI21_X1 U4178 ( .B1(n4064), .B2(n3503), .A(n3365), .ZN(n3366) );
  OAI21_X1 U4179 ( .B1(n3367), .B2(n3505), .A(n3366), .ZN(U3212) );
  OAI21_X1 U4180 ( .B1(n2034), .B2(n3369), .A(n3368), .ZN(n3371) );
  NAND3_X1 U4181 ( .A1(n3371), .A2(n3510), .A3(n3370), .ZN(n3375) );
  AOI22_X1 U4182 ( .A1(n3517), .A2(n2147), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3374) );
  AOI22_X1 U4183 ( .A1(n3478), .A2(n3888), .B1(n3499), .B2(n3925), .ZN(n3373)
         );
  NAND2_X1 U4184 ( .A1(n3503), .A2(n3894), .ZN(n3372) );
  NAND4_X1 U4185 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(U3213)
         );
  INV_X1 U4186 ( .A(n3377), .ZN(n3378) );
  AOI21_X1 U4187 ( .B1(n3379), .B2(n3376), .A(n3378), .ZN(n3384) );
  NOR2_X1 U4188 ( .A1(n4598), .A2(STATE_REG_SCAN_IN), .ZN(n3773) );
  OAI22_X1 U4189 ( .A1(n3515), .A2(n3974), .B1(n3923), .B2(n3513), .ZN(n3380)
         );
  AOI211_X1 U4190 ( .C1(n3970), .C2(n3517), .A(n3773), .B(n3380), .ZN(n3383)
         );
  INV_X1 U4191 ( .A(n3381), .ZN(n3979) );
  NAND2_X1 U4192 ( .A1(n3503), .A2(n3979), .ZN(n3382) );
  OAI211_X1 U4193 ( .C1(n3384), .C2(n3505), .A(n3383), .B(n3382), .ZN(U3216)
         );
  NAND2_X1 U4194 ( .A1(n2058), .A2(n3385), .ZN(n3388) );
  INV_X1 U4195 ( .A(n3448), .ZN(n3386) );
  OAI211_X1 U4196 ( .C1(n3445), .C2(n3386), .A(n3446), .B(n3388), .ZN(n3387)
         );
  OAI211_X1 U4197 ( .C1(n3389), .C2(n3388), .A(n3510), .B(n3387), .ZN(n3393)
         );
  OAI22_X1 U4198 ( .A1(n3515), .A2(n3923), .B1(n3891), .B2(n3513), .ZN(n3391)
         );
  OAI22_X1 U4199 ( .A1(n3497), .A2(n3930), .B1(STATE_REG_SCAN_IN), .B2(n4587), 
        .ZN(n3390) );
  NOR2_X1 U4200 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  OAI211_X1 U4201 ( .C1(n3521), .C2(n3932), .A(n3393), .B(n3392), .ZN(U3220)
         );
  INV_X1 U4202 ( .A(n3394), .ZN(n3396) );
  NAND2_X1 U4203 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  XNOR2_X1 U4204 ( .A(n3398), .B(n3397), .ZN(n3404) );
  AOI22_X1 U4205 ( .A1(n3478), .A2(n4055), .B1(n3499), .B2(n3673), .ZN(n3399)
         );
  NAND2_X1 U4206 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4306) );
  OAI211_X1 U4207 ( .C1(n3497), .C2(n3400), .A(n3399), .B(n4306), .ZN(n3401)
         );
  AOI21_X1 U4208 ( .B1(n3402), .B2(n3503), .A(n3401), .ZN(n3403) );
  OAI21_X1 U4209 ( .B1(n3404), .B2(n3505), .A(n3403), .ZN(U3221) );
  INV_X1 U4210 ( .A(n3406), .ZN(n3407) );
  NOR2_X1 U4211 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  XNOR2_X1 U4212 ( .A(n3405), .B(n3409), .ZN(n3414) );
  OAI22_X1 U4213 ( .A1(n3497), .A2(n3853), .B1(STATE_REG_SCAN_IN), .B2(n3410), 
        .ZN(n3412) );
  OAI22_X1 U4214 ( .A1(n3803), .A2(n3513), .B1(n3515), .B2(n3847), .ZN(n3411)
         );
  AOI211_X1 U4215 ( .C1(n3855), .C2(n3503), .A(n3412), .B(n3411), .ZN(n3413)
         );
  OAI21_X1 U4216 ( .B1(n3414), .B2(n3505), .A(n3413), .ZN(U3222) );
  INV_X1 U4217 ( .A(n3415), .ZN(n3507) );
  OAI21_X1 U4218 ( .B1(n3507), .B2(n3508), .A(n3416), .ZN(n3417) );
  XOR2_X1 U4219 ( .A(n3418), .B(n3417), .Z(n3425) );
  INV_X1 U4220 ( .A(n4024), .ZN(n3423) );
  AOI22_X1 U4221 ( .A1(n3478), .A2(n4030), .B1(n3499), .B2(n3419), .ZN(n3420)
         );
  NAND2_X1 U4222 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4348) );
  OAI211_X1 U4223 ( .C1(n3497), .C2(n3421), .A(n3420), .B(n4348), .ZN(n3422)
         );
  AOI21_X1 U4224 ( .B1(n3423), .B2(n3503), .A(n3422), .ZN(n3424) );
  OAI21_X1 U4225 ( .B1(n3425), .B2(n3505), .A(n3424), .ZN(U3223) );
  INV_X1 U4226 ( .A(n3427), .ZN(n3428) );
  NOR2_X1 U4227 ( .A1(n3429), .A2(n3428), .ZN(n3430) );
  XNOR2_X1 U4228 ( .A(n3426), .B(n3430), .ZN(n3431) );
  NAND2_X1 U4229 ( .A1(n3431), .A2(n3510), .ZN(n3434) );
  AND2_X1 U4230 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3742) );
  OAI22_X1 U4231 ( .A1(n3515), .A2(n4036), .B1(n3974), .B2(n3513), .ZN(n3432)
         );
  AOI211_X1 U4232 ( .C1(n4005), .C2(n3517), .A(n3742), .B(n3432), .ZN(n3433)
         );
  OAI211_X1 U4233 ( .C1(n3521), .C2(n4013), .A(n3434), .B(n3433), .ZN(U3225)
         );
  NAND2_X1 U4234 ( .A1(n3435), .A2(n3436), .ZN(n3437) );
  XOR2_X1 U4235 ( .A(n3438), .B(n3437), .Z(n3443) );
  INV_X1 U4236 ( .A(n3873), .ZN(n3441) );
  OAI22_X1 U4237 ( .A1(n3497), .A2(n3871), .B1(STATE_REG_SCAN_IN), .B2(n4511), 
        .ZN(n3440) );
  OAI22_X1 U4238 ( .A1(n3515), .A2(n3865), .B1(n3828), .B2(n3513), .ZN(n3439)
         );
  AOI211_X1 U4239 ( .C1(n3441), .C2(n3503), .A(n3440), .B(n3439), .ZN(n3442)
         );
  OAI21_X1 U4240 ( .B1(n3443), .B2(n3505), .A(n3442), .ZN(U3226) );
  INV_X1 U4241 ( .A(n3444), .ZN(n3449) );
  AOI21_X1 U4242 ( .B1(n3446), .B2(n3448), .A(n3445), .ZN(n3447) );
  AOI21_X1 U4243 ( .B1(n3449), .B2(n3448), .A(n3447), .ZN(n3455) );
  INV_X1 U4244 ( .A(n3954), .ZN(n3453) );
  OAI22_X1 U4245 ( .A1(n3497), .A2(n3952), .B1(STATE_REG_SCAN_IN), .B2(n3450), 
        .ZN(n3452) );
  OAI22_X1 U4246 ( .A1(n3515), .A2(n3947), .B1(n3908), .B2(n3513), .ZN(n3451)
         );
  AOI211_X1 U4247 ( .C1(n3453), .C2(n3503), .A(n3452), .B(n3451), .ZN(n3454)
         );
  OAI21_X1 U4248 ( .B1(n3455), .B2(n3505), .A(n3454), .ZN(U3230) );
  XNOR2_X1 U4249 ( .A(n3458), .B(n3457), .ZN(n3459) );
  XNOR2_X1 U4250 ( .A(n3456), .B(n3459), .ZN(n3460) );
  NAND2_X1 U4251 ( .A1(n3460), .A2(n3510), .ZN(n3464) );
  NOR2_X1 U4252 ( .A1(STATE_REG_SCAN_IN), .A2(n3461), .ZN(n4316) );
  OAI22_X1 U4253 ( .A1(n3515), .A2(n4101), .B1(n3514), .B2(n3513), .ZN(n3462)
         );
  AOI211_X1 U4254 ( .C1(n4077), .C2(n3517), .A(n4316), .B(n3462), .ZN(n3463)
         );
  OAI211_X1 U4255 ( .C1(n3521), .C2(n4090), .A(n3464), .B(n3463), .ZN(U3231)
         );
  AOI21_X1 U4256 ( .B1(n3466), .B2(n3465), .A(n2034), .ZN(n3471) );
  OAI22_X1 U4257 ( .A1(n3497), .A2(n3913), .B1(STATE_REG_SCAN_IN), .B2(n3467), 
        .ZN(n3469) );
  OAI22_X1 U4258 ( .A1(n3515), .A2(n3908), .B1(n3865), .B2(n3513), .ZN(n3468)
         );
  AOI211_X1 U4259 ( .C1(n3914), .C2(n3503), .A(n3469), .B(n3468), .ZN(n3470)
         );
  OAI21_X1 U4260 ( .B1(n3471), .B2(n3505), .A(n3470), .ZN(U3232) );
  OAI21_X1 U4261 ( .B1(n3474), .B2(n3473), .A(n3472), .ZN(n3475) );
  NAND2_X1 U4262 ( .A1(n3475), .A2(n3510), .ZN(n3481) );
  AOI22_X1 U4263 ( .A1(n3499), .A2(n3680), .B1(n3476), .B2(n3517), .ZN(n3480)
         );
  AOI22_X1 U4264 ( .A1(n3478), .A2(n2708), .B1(REG3_REG_2__SCAN_IN), .B2(n3477), .ZN(n3479) );
  NAND3_X1 U4265 ( .A1(n3481), .A2(n3480), .A3(n3479), .ZN(U3234) );
  XNOR2_X1 U4266 ( .A(n3484), .B(n3483), .ZN(n3485) );
  XNOR2_X1 U4267 ( .A(n3482), .B(n3485), .ZN(n3486) );
  NAND2_X1 U4268 ( .A1(n3486), .A2(n3510), .ZN(n3490) );
  NOR2_X1 U4269 ( .A1(n3487), .A2(STATE_REG_SCAN_IN), .ZN(n4363) );
  OAI22_X1 U4270 ( .A1(n3515), .A2(n3987), .B1(n3947), .B2(n3513), .ZN(n3488)
         );
  AOI211_X1 U4271 ( .C1(n3993), .C2(n3517), .A(n4363), .B(n3488), .ZN(n3489)
         );
  OAI211_X1 U4272 ( .C1(n3521), .C2(n3996), .A(n3490), .B(n3489), .ZN(U3235)
         );
  INV_X1 U4273 ( .A(n3492), .ZN(n3494) );
  NAND2_X1 U4274 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  XNOR2_X1 U4275 ( .A(n3491), .B(n3495), .ZN(n3506) );
  OAI22_X1 U4276 ( .A1(n3497), .A2(n3835), .B1(STATE_REG_SCAN_IN), .B2(n3496), 
        .ZN(n3498) );
  AOI21_X1 U4277 ( .B1(n3499), .B2(n3867), .A(n3498), .ZN(n3500) );
  OAI21_X1 U4278 ( .B1(n3501), .B2(n3513), .A(n3500), .ZN(n3502) );
  AOI21_X1 U4279 ( .B1(n3837), .B2(n3503), .A(n3502), .ZN(n3504) );
  OAI21_X1 U4280 ( .B1(n3506), .B2(n3505), .A(n3504), .ZN(U3237) );
  NAND2_X1 U4281 ( .A1(n3415), .A2(n3416), .ZN(n3509) );
  XNOR2_X1 U4282 ( .A(n3509), .B(n3508), .ZN(n3511) );
  NAND2_X1 U4283 ( .A1(n3511), .A2(n3510), .ZN(n3520) );
  NOR2_X1 U4284 ( .A1(STATE_REG_SCAN_IN), .A2(n3512), .ZN(n4341) );
  OAI22_X1 U4285 ( .A1(n3515), .A2(n3514), .B1(n4036), .B2(n3513), .ZN(n3516)
         );
  AOI211_X1 U4286 ( .C1(n3518), .C2(n3517), .A(n4341), .B(n3516), .ZN(n3519)
         );
  OAI211_X1 U4287 ( .C1(n3521), .C2(n4043), .A(n3520), .B(n3519), .ZN(U3238)
         );
  AND2_X1 U4288 ( .A1(n3528), .A2(DATAI_29_), .ZN(n3795) );
  OR2_X1 U4289 ( .A1(n3524), .A2(n3795), .ZN(n3616) );
  AND2_X1 U4290 ( .A1(n3783), .A2(n3616), .ZN(n3629) );
  NAND2_X1 U4291 ( .A1(n3523), .A2(n3522), .ZN(n3784) );
  NAND2_X1 U4292 ( .A1(n3524), .A2(n3795), .ZN(n3615) );
  INV_X1 U4293 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U4294 ( .A1(n2350), .A2(REG2_REG_31__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4295 ( .A1(n2918), .A2(REG0_REG_31__SCAN_IN), .ZN(n3525) );
  OAI211_X1 U4296 ( .C1(n2507), .C2(n3527), .A(n3526), .B(n3525), .ZN(n4123)
         );
  NAND2_X1 U4297 ( .A1(n3528), .A2(DATAI_31_), .ZN(n4121) );
  NAND2_X1 U4298 ( .A1(n4123), .A2(n4121), .ZN(n3590) );
  AND2_X1 U4299 ( .A1(n3528), .A2(DATAI_30_), .ZN(n4130) );
  INV_X1 U4300 ( .A(n4130), .ZN(n3588) );
  OR2_X1 U4301 ( .A1(n3788), .A2(n3588), .ZN(n3529) );
  AND2_X1 U4302 ( .A1(n3590), .A2(n3529), .ZN(n3599) );
  NAND2_X1 U4303 ( .A1(n3615), .A2(n3599), .ZN(n3646) );
  AOI21_X1 U4304 ( .B1(n3629), .B2(n3784), .A(n3646), .ZN(n3651) );
  INV_X1 U4305 ( .A(n3634), .ZN(n3578) );
  NAND2_X1 U4306 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  NAND2_X1 U4307 ( .A1(n3567), .A2(n3533), .ZN(n3632) );
  AND4_X1 U4308 ( .A1(n3566), .A2(n3535), .A3(n3534), .A4(n3632), .ZN(n3575)
         );
  NAND2_X1 U4309 ( .A1(n3537), .A2(n3536), .ZN(n3555) );
  INV_X1 U4310 ( .A(n3555), .ZN(n3562) );
  INV_X1 U4311 ( .A(n3538), .ZN(n3541) );
  OAI211_X1 U4312 ( .C1(n3657), .C2(n3541), .A(n3540), .B(n3539), .ZN(n3542)
         );
  NAND3_X1 U4313 ( .A1(n3543), .A2(n2609), .A3(n3542), .ZN(n3544) );
  NAND3_X1 U4314 ( .A1(n3546), .A2(n3545), .A3(n3544), .ZN(n3547) );
  NAND3_X1 U4315 ( .A1(n3549), .A2(n3548), .A3(n3547), .ZN(n3550) );
  NAND4_X1 U4316 ( .A1(n3551), .A2(n2045), .A3(n3554), .A4(n3550), .ZN(n3552)
         );
  NAND3_X1 U4317 ( .A1(n3607), .A2(n3553), .A3(n3552), .ZN(n3561) );
  NOR3_X1 U4318 ( .A1(n2118), .A2(n3556), .A3(n3555), .ZN(n3560) );
  NAND2_X1 U4319 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  AOI211_X1 U4320 ( .C1(n3562), .C2(n3561), .A(n3560), .B(n3559), .ZN(n3564)
         );
  OAI21_X1 U4321 ( .B1(n3565), .B2(n3564), .A(n3563), .ZN(n3574) );
  INV_X1 U4322 ( .A(n3566), .ZN(n3571) );
  NAND2_X1 U4323 ( .A1(n3568), .A2(n3567), .ZN(n3633) );
  INV_X1 U4324 ( .A(n3633), .ZN(n3569) );
  OAI211_X1 U4325 ( .C1(n3572), .C2(n3571), .A(n3570), .B(n3569), .ZN(n3573)
         );
  AOI22_X1 U4326 ( .A1(n3575), .A2(n3574), .B1(n3632), .B2(n3573), .ZN(n3576)
         );
  OAI21_X1 U4327 ( .B1(n2134), .B2(n3576), .A(n3635), .ZN(n3577) );
  AOI21_X1 U4328 ( .B1(n3578), .B2(n3577), .A(n2132), .ZN(n3579) );
  OR3_X1 U4329 ( .A1(n3638), .A2(n3880), .A3(n3579), .ZN(n3580) );
  AND2_X1 U4330 ( .A1(n3581), .A2(n3580), .ZN(n3583) );
  OAI211_X1 U4331 ( .C1(n3584), .C2(n3583), .A(n3582), .B(n3644), .ZN(n3586)
         );
  NAND4_X1 U4332 ( .A1(n3587), .A2(n3629), .A3(n3586), .A4(n3585), .ZN(n3591)
         );
  NAND2_X1 U4333 ( .A1(n3788), .A2(n3588), .ZN(n3654) );
  OR2_X1 U4334 ( .A1(n4123), .A2(n4121), .ZN(n3589) );
  NAND2_X1 U4335 ( .A1(n3654), .A2(n3589), .ZN(n3596) );
  AOI22_X1 U4336 ( .A1(n3651), .A2(n3591), .B1(n3590), .B2(n3596), .ZN(n3662)
         );
  NAND2_X1 U4337 ( .A1(n3822), .A2(n3592), .ZN(n3846) );
  INV_X1 U4338 ( .A(n3593), .ZN(n3595) );
  OR2_X1 U4339 ( .A1(n3595), .A2(n3594), .ZN(n3967) );
  NOR3_X1 U4340 ( .A1(n3846), .A2(n3596), .A3(n3967), .ZN(n3612) );
  INV_X1 U4341 ( .A(n3597), .ZN(n3861) );
  NAND2_X1 U4342 ( .A1(n3861), .A2(n3598), .ZN(n3886) );
  INV_X1 U4343 ( .A(n3599), .ZN(n3602) );
  NOR4_X1 U4344 ( .A1(n3886), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3611)
         );
  NOR4_X1 U4345 ( .A1(n3605), .A2(n3604), .A3(n3991), .A4(n3603), .ZN(n3610)
         );
  AND4_X1 U4346 ( .A1(n3608), .A2(n4098), .A3(n3607), .A4(n3606), .ZN(n3609)
         );
  AND4_X1 U4347 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3614)
         );
  XNOR2_X1 U4348 ( .A(n3803), .B(n3835), .ZN(n3825) );
  XNOR2_X1 U4349 ( .A(n3923), .B(n3944), .ZN(n3938) );
  INV_X1 U4350 ( .A(n3938), .ZN(n3942) );
  XNOR2_X1 U4351 ( .A(n3613), .B(n4088), .ZN(n4076) );
  NAND4_X1 U4352 ( .A1(n3614), .A2(n3825), .A3(n3942), .A4(n4076), .ZN(n3628)
         );
  NAND2_X1 U4353 ( .A1(n3616), .A2(n3615), .ZN(n3785) );
  INV_X1 U4354 ( .A(n3785), .ZN(n3626) );
  INV_X1 U4355 ( .A(n3617), .ZN(n3619) );
  INV_X1 U4356 ( .A(n3882), .ZN(n3618) );
  OR2_X1 U4357 ( .A1(n3880), .A2(n3618), .ZN(n3921) );
  NOR4_X1 U4358 ( .A1(n2610), .A2(n3619), .A3(n3921), .A4(n4047), .ZN(n3625)
         );
  NAND2_X1 U4359 ( .A1(n3962), .A2(n3961), .ZN(n4002) );
  NOR3_X1 U4360 ( .A1(n3902), .A2(n4002), .A3(n3620), .ZN(n3624) );
  INV_X1 U4361 ( .A(n3843), .ZN(n3622) );
  OR2_X1 U4362 ( .A1(n3622), .A2(n3621), .ZN(n3863) );
  NAND4_X1 U4363 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  NOR4_X1 U4364 ( .A1(n3628), .A2(n3627), .A3(n3780), .A4(n3810), .ZN(n3659)
         );
  INV_X1 U4365 ( .A(n4123), .ZN(n3653) );
  INV_X1 U4366 ( .A(n3629), .ZN(n3631) );
  OR3_X1 U4367 ( .A1(n3810), .A2(n3631), .A3(n3630), .ZN(n3650) );
  OAI21_X1 U4368 ( .B1(n4051), .B2(n3633), .A(n3632), .ZN(n3636) );
  AOI211_X1 U4369 ( .C1(n3636), .C2(n3635), .A(n2134), .B(n3634), .ZN(n3637)
         );
  INV_X1 U4370 ( .A(n3637), .ZN(n3640) );
  AOI21_X1 U4371 ( .B1(n3640), .B2(n3639), .A(n3638), .ZN(n3643) );
  OAI21_X1 U4372 ( .B1(n3643), .B2(n3642), .A(n3641), .ZN(n3645) );
  AOI21_X1 U4373 ( .B1(n3645), .B2(n3644), .A(n3823), .ZN(n3648) );
  NOR4_X1 U4374 ( .A1(n3648), .A2(n3784), .A3(n3647), .A4(n3646), .ZN(n3649)
         );
  AOI21_X1 U4375 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(n3652) );
  AOI21_X1 U4376 ( .B1(n4130), .B2(n3653), .A(n3652), .ZN(n3656) );
  AOI21_X1 U4377 ( .B1(n3654), .B2(n4123), .A(n4121), .ZN(n3655) );
  NOR2_X1 U4378 ( .A1(n3656), .A2(n3655), .ZN(n3658) );
  MUX2_X1 U4379 ( .A(n3659), .B(n3658), .S(n3657), .Z(n3661) );
  MUX2_X1 U4380 ( .A(n3662), .B(n3661), .S(n3660), .Z(n3663) );
  XNOR2_X1 U4381 ( .A(n3663), .B(n4269), .ZN(n3670) );
  NAND2_X1 U4382 ( .A1(n3665), .A2(n3664), .ZN(n3666) );
  OAI211_X1 U4383 ( .C1(n3667), .C2(n3669), .A(n3666), .B(B_REG_SCAN_IN), .ZN(
        n3668) );
  OAI21_X1 U4384 ( .B1(n3670), .B2(n3669), .A(n3668), .ZN(U3239) );
  MUX2_X1 U4385 ( .A(DATAO_REG_31__SCAN_IN), .B(n4123), .S(n3679), .Z(U3581)
         );
  MUX2_X1 U4386 ( .A(DATAO_REG_28__SCAN_IN), .B(n3809), .S(n3679), .Z(U3578)
         );
  MUX2_X1 U4387 ( .A(DATAO_REG_27__SCAN_IN), .B(n3830), .S(n3679), .Z(U3577)
         );
  MUX2_X1 U4388 ( .A(n3849), .B(DATAO_REG_26__SCAN_IN), .S(n3681), .Z(U3576)
         );
  MUX2_X1 U4389 ( .A(n3867), .B(DATAO_REG_25__SCAN_IN), .S(n3681), .Z(U3575)
         );
  MUX2_X1 U4390 ( .A(n3888), .B(DATAO_REG_24__SCAN_IN), .S(n3681), .Z(U3574)
         );
  MUX2_X1 U4391 ( .A(n3910), .B(DATAO_REG_23__SCAN_IN), .S(n3681), .Z(U3573)
         );
  MUX2_X1 U4392 ( .A(n3925), .B(DATAO_REG_22__SCAN_IN), .S(n3681), .Z(U3572)
         );
  MUX2_X1 U4393 ( .A(n3945), .B(DATAO_REG_21__SCAN_IN), .S(n3681), .Z(U3571)
         );
  MUX2_X1 U4394 ( .A(DATAO_REG_17__SCAN_IN), .B(n4030), .S(n3679), .Z(U3567)
         );
  MUX2_X1 U4395 ( .A(DATAO_REG_16__SCAN_IN), .B(n3671), .S(n3679), .Z(U3566)
         );
  MUX2_X1 U4396 ( .A(DATAO_REG_12__SCAN_IN), .B(n3672), .S(n3679), .Z(U3562)
         );
  MUX2_X1 U4397 ( .A(DATAO_REG_11__SCAN_IN), .B(n3673), .S(n3679), .Z(U3561)
         );
  MUX2_X1 U4398 ( .A(n4105), .B(DATAO_REG_10__SCAN_IN), .S(n3681), .Z(U3560)
         );
  MUX2_X1 U4399 ( .A(n3674), .B(DATAO_REG_9__SCAN_IN), .S(n3681), .Z(U3559) );
  MUX2_X1 U4400 ( .A(n3675), .B(DATAO_REG_6__SCAN_IN), .S(n3681), .Z(U3556) );
  MUX2_X1 U4401 ( .A(DATAO_REG_5__SCAN_IN), .B(n3676), .S(n3679), .Z(U3555) );
  MUX2_X1 U4402 ( .A(DATAO_REG_4__SCAN_IN), .B(n3677), .S(n3679), .Z(U3554) );
  MUX2_X1 U4403 ( .A(DATAO_REG_2__SCAN_IN), .B(n3678), .S(n3679), .Z(U3552) );
  MUX2_X1 U4404 ( .A(DATAO_REG_1__SCAN_IN), .B(n3680), .S(n3679), .Z(U3551) );
  MUX2_X1 U4405 ( .A(n2691), .B(DATAO_REG_0__SCAN_IN), .S(n3681), .Z(U3550) );
  AOI22_X1 U4406 ( .A1(n4461), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3690) );
  NAND3_X1 U4407 ( .A1(n4357), .A2(n3682), .A3(n4409), .ZN(n3689) );
  INV_X1 U4408 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3683) );
  AND2_X1 U4409 ( .A1(n3787), .A2(n3683), .ZN(n3684) );
  NOR2_X1 U4410 ( .A1(n3684), .A2(n4278), .ZN(n3706) );
  NOR2_X1 U4411 ( .A1(n3787), .A2(REG1_REG_0__SCAN_IN), .ZN(n3685) );
  OAI21_X1 U4412 ( .B1(n4409), .B2(n3685), .A(n3706), .ZN(n3686) );
  OAI211_X1 U4413 ( .C1(n3706), .C2(n4409), .A(n3687), .B(n3686), .ZN(n3688)
         );
  NAND3_X1 U4414 ( .A1(n3690), .A2(n3689), .A3(n3688), .ZN(U3240) );
  AOI22_X1 U4415 ( .A1(n4461), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3699) );
  NAND2_X1 U4416 ( .A1(n4333), .A2(n4276), .ZN(n3698) );
  OAI211_X1 U4417 ( .C1(n3704), .C2(n3692), .A(n4463), .B(n3691), .ZN(n3697)
         );
  OAI211_X1 U4418 ( .C1(n3695), .C2(n3694), .A(n4357), .B(n3693), .ZN(n3696)
         );
  NAND4_X1 U4419 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(U3241)
         );
  NAND2_X1 U4420 ( .A1(n3700), .A2(n3703), .ZN(n3702) );
  INV_X1 U4421 ( .A(n4278), .ZN(n3701) );
  OAI211_X1 U4422 ( .C1(n3704), .C2(n3703), .A(n3702), .B(n3701), .ZN(n3705)
         );
  OAI211_X1 U4423 ( .C1(n4409), .C2(n3706), .A(n3705), .B(U4043), .ZN(n3726)
         );
  AOI22_X1 U4424 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4461), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3715) );
  XNOR2_X1 U4425 ( .A(n3708), .B(n3707), .ZN(n3709) );
  AOI22_X1 U4426 ( .A1(n4275), .A2(n4333), .B1(n4357), .B2(n3709), .ZN(n3714)
         );
  OAI211_X1 U4427 ( .C1(n3712), .C2(n3711), .A(n4463), .B(n3710), .ZN(n3713)
         );
  NAND4_X1 U4428 ( .A1(n3726), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(U3242)
         );
  NAND2_X1 U4429 ( .A1(n4461), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3725) );
  XNOR2_X1 U4430 ( .A(n3716), .B(REG2_REG_4__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U4431 ( .A1(n4463), .A2(n3717), .ZN(n3720) );
  NAND2_X1 U4432 ( .A1(n4333), .A2(n4273), .ZN(n3719) );
  AND3_X1 U4433 ( .A1(n3720), .A2(n3719), .A3(n3718), .ZN(n3724) );
  XNOR2_X1 U4434 ( .A(n3721), .B(REG1_REG_4__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4435 ( .A1(n4357), .A2(n3722), .ZN(n3723) );
  NAND4_X1 U4436 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(U3244)
         );
  XNOR2_X1 U4437 ( .A(n3743), .B(REG2_REG_17__SCAN_IN), .ZN(n3740) );
  INV_X1 U4438 ( .A(n4332), .ZN(n4401) );
  NOR2_X1 U4439 ( .A1(n4091), .A2(n4403), .ZN(n4318) );
  NAND2_X1 U4440 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3748), .ZN(n3731) );
  INV_X1 U4441 ( .A(n3748), .ZN(n4406) );
  AOI22_X1 U4442 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3748), .B1(n4406), .B2(
        n4115), .ZN(n4300) );
  NAND2_X1 U4443 ( .A1(n3746), .A2(n3729), .ZN(n3730) );
  INV_X1 U4444 ( .A(n3746), .ZN(n4467) );
  NAND2_X1 U4445 ( .A1(n3730), .A2(n4462), .ZN(n4299) );
  NAND2_X1 U4446 ( .A1(n4300), .A2(n4299), .ZN(n4298) );
  NAND2_X1 U4447 ( .A1(n3732), .A2(n3733), .ZN(n3734) );
  NOR2_X1 U4448 ( .A1(n4401), .A2(n3735), .ZN(n3736) );
  NOR2_X1 U4449 ( .A1(n2461), .A2(n4329), .ZN(n4328) );
  INV_X1 U4450 ( .A(n3755), .ZN(n4400) );
  AOI22_X1 U4451 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4400), .B1(n3755), .B2(
        n4044), .ZN(n4344) );
  NAND2_X1 U4452 ( .A1(n3737), .A2(n4398), .ZN(n3738) );
  INV_X1 U4453 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U4454 ( .A1(n4352), .A2(n4351), .ZN(n4350) );
  NAND2_X1 U4455 ( .A1(n3738), .A2(n4350), .ZN(n3739) );
  OAI21_X1 U4456 ( .B1(n3740), .B2(n3739), .A(n3768), .ZN(n3741) );
  AOI22_X1 U4457 ( .A1(n3769), .A2(n4333), .B1(n4463), .B2(n3741), .ZN(n3763)
         );
  AOI21_X1 U4458 ( .B1(n4461), .B2(ADDR_REG_17__SCAN_IN), .A(n3742), .ZN(n3762) );
  XNOR2_X1 U4459 ( .A(n3743), .B(REG1_REG_17__SCAN_IN), .ZN(n3759) );
  NOR2_X1 U4460 ( .A1(n3745), .A2(n4467), .ZN(n3747) );
  AOI22_X1 U4461 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4406), .B1(n3748), .B2(
        n4206), .ZN(n4294) );
  NOR2_X1 U4462 ( .A1(n3749), .A2(n4405), .ZN(n3750) );
  AOI22_X1 U4463 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4403), .B1(n3751), .B2(
        n4197), .ZN(n4314) );
  NOR2_X1 U4464 ( .A1(n3752), .A2(n4401), .ZN(n3753) );
  AOI22_X1 U4465 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4400), .B1(n3755), .B2(
        n3754), .ZN(n4338) );
  NAND2_X1 U4466 ( .A1(n3756), .A2(n4398), .ZN(n3757) );
  NAND2_X1 U4467 ( .A1(n3758), .A2(n3759), .ZN(n3765) );
  OAI21_X1 U4468 ( .B1(n3759), .B2(n3758), .A(n3765), .ZN(n3760) );
  NAND2_X1 U4469 ( .A1(n4357), .A2(n3760), .ZN(n3761) );
  NAND3_X1 U4470 ( .A1(n3763), .A2(n3762), .A3(n3761), .ZN(U3257) );
  INV_X1 U4471 ( .A(n3770), .ZN(n4396) );
  AOI22_X1 U4472 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4396), .B1(n3770), .B2(
        n3764), .ZN(n4362) );
  XNOR2_X1 U4473 ( .A(n4269), .B(REG1_REG_19__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4474 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3770), .ZN(n3767) );
  OAI21_X1 U4475 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3770), .A(n3767), .ZN(n4366) );
  MUX2_X1 U4476 ( .A(REG2_REG_19__SCAN_IN), .B(n2518), .S(n4269), .Z(n3771) );
  XNOR2_X1 U4477 ( .A(n3772), .B(n3771), .ZN(n3777) );
  AOI21_X1 U4478 ( .B1(n4461), .B2(ADDR_REG_19__SCAN_IN), .A(n3773), .ZN(n3774) );
  OAI21_X1 U4479 ( .B1(n4468), .B2(n3775), .A(n3774), .ZN(n3776) );
  AOI21_X1 U4480 ( .B1(n3777), .B2(n4463), .A(n3776), .ZN(n3778) );
  AOI22_X1 U4481 ( .A1(n3781), .A2(n3780), .B1(n3779), .B2(n3809), .ZN(n3782)
         );
  XNOR2_X1 U4482 ( .A(n3782), .B(n3785), .ZN(n4132) );
  INV_X1 U4483 ( .A(n4132), .ZN(n3802) );
  OAI21_X1 U4484 ( .B1(n3804), .B2(n3784), .A(n3783), .ZN(n3786) );
  XNOR2_X1 U4485 ( .A(n3786), .B(n3785), .ZN(n3792) );
  AOI21_X1 U4486 ( .B1(B_REG_SCAN_IN), .B2(n3787), .A(n4100), .ZN(n4122) );
  AOI22_X1 U4487 ( .A1(n3788), .A2(n4122), .B1(n4129), .B2(n3795), .ZN(n3789)
         );
  OAI21_X1 U4488 ( .B1(n3790), .B2(n4081), .A(n3789), .ZN(n3791) );
  AOI21_X1 U4489 ( .B1(n3792), .B2(n4083), .A(n3791), .ZN(n4134) );
  OAI21_X1 U4490 ( .B1(n4370), .B2(n3793), .A(n4134), .ZN(n3800) );
  INV_X1 U4491 ( .A(n3795), .ZN(n3796) );
  OAI21_X1 U4492 ( .B1(n3797), .B2(n3796), .A(n4127), .ZN(n4133) );
  INV_X1 U4493 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3798) );
  OAI22_X1 U4494 ( .A1(n4133), .A2(n4066), .B1(n3798), .B2(n4372), .ZN(n3799)
         );
  AOI21_X1 U4495 ( .B1(n3800), .B2(n4372), .A(n3799), .ZN(n3801) );
  OAI21_X1 U4496 ( .B1(n3802), .B2(n4035), .A(n3801), .ZN(U3354) );
  OAI22_X1 U4497 ( .A1(n3803), .A2(n4081), .B1(n4099), .B2(n3813), .ZN(n3808)
         );
  AOI21_X1 U4498 ( .B1(n3805), .B2(n3810), .A(n3804), .ZN(n3806) );
  NOR2_X1 U4499 ( .A1(n3806), .A2(n4109), .ZN(n3807) );
  AOI211_X1 U4500 ( .C1(n4078), .C2(n3809), .A(n3808), .B(n3807), .ZN(n4137)
         );
  XNOR2_X1 U4501 ( .A(n3811), .B(n3810), .ZN(n4136) );
  NAND2_X1 U4502 ( .A1(n4136), .A2(n4068), .ZN(n3820) );
  OAI21_X1 U4503 ( .B1(n3833), .B2(n3813), .A(n3812), .ZN(n4139) );
  INV_X1 U4504 ( .A(n4139), .ZN(n3818) );
  INV_X1 U4505 ( .A(n3814), .ZN(n3816) );
  OAI22_X1 U4506 ( .A1(n3816), .A2(n4370), .B1(n3815), .B2(n4372), .ZN(n3817)
         );
  AOI21_X1 U4507 ( .B1(n3818), .B2(n4377), .A(n3817), .ZN(n3819) );
  OAI211_X1 U4508 ( .C1(n4137), .C2(n4391), .A(n3820), .B(n3819), .ZN(U3263)
         );
  XNOR2_X1 U4509 ( .A(n3821), .B(n3825), .ZN(n4141) );
  INV_X1 U4510 ( .A(n4141), .ZN(n3841) );
  INV_X1 U4511 ( .A(n3844), .ZN(n3824) );
  OAI21_X1 U4512 ( .B1(n3824), .B2(n3823), .A(n3822), .ZN(n3827) );
  INV_X1 U4513 ( .A(n3825), .ZN(n3826) );
  XNOR2_X1 U4514 ( .A(n3827), .B(n3826), .ZN(n3832) );
  OAI22_X1 U4515 ( .A1(n3828), .A2(n4081), .B1(n4099), .B2(n3835), .ZN(n3829)
         );
  AOI21_X1 U4516 ( .B1(n4078), .B2(n3830), .A(n3829), .ZN(n3831) );
  OAI21_X1 U4517 ( .B1(n3832), .B2(n4109), .A(n3831), .ZN(n4140) );
  INV_X1 U4518 ( .A(n3852), .ZN(n3836) );
  INV_X1 U4519 ( .A(n3833), .ZN(n3834) );
  OAI21_X1 U4520 ( .B1(n3836), .B2(n3835), .A(n3834), .ZN(n4218) );
  AOI22_X1 U4521 ( .A1(REG2_REG_26__SCAN_IN), .A2(n4391), .B1(n3837), .B2(
        n4386), .ZN(n3838) );
  OAI21_X1 U4522 ( .B1(n4218), .B2(n4066), .A(n3838), .ZN(n3839) );
  AOI21_X1 U4523 ( .B1(n4140), .B2(n4372), .A(n3839), .ZN(n3840) );
  OAI21_X1 U4524 ( .B1(n3841), .B2(n4035), .A(n3840), .ZN(U3264) );
  XNOR2_X1 U4525 ( .A(n3842), .B(n3846), .ZN(n4145) );
  INV_X1 U4526 ( .A(n4145), .ZN(n3859) );
  NAND2_X1 U4527 ( .A1(n3844), .A2(n3843), .ZN(n3845) );
  XOR2_X1 U4528 ( .A(n3846), .B(n3845), .Z(n3851) );
  OAI22_X1 U4529 ( .A1(n3847), .A2(n4081), .B1(n4099), .B2(n3853), .ZN(n3848)
         );
  AOI21_X1 U4530 ( .B1(n3849), .B2(n4078), .A(n3848), .ZN(n3850) );
  OAI21_X1 U4531 ( .B1(n3851), .B2(n4109), .A(n3850), .ZN(n4144) );
  INV_X1 U4532 ( .A(n3870), .ZN(n3854) );
  OAI21_X1 U4533 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n4222) );
  AOI22_X1 U4534 ( .A1(n4391), .A2(REG2_REG_25__SCAN_IN), .B1(n3855), .B2(
        n4386), .ZN(n3856) );
  OAI21_X1 U4535 ( .B1(n4222), .B2(n4066), .A(n3856), .ZN(n3857) );
  AOI21_X1 U4536 ( .B1(n4144), .B2(n4372), .A(n3857), .ZN(n3858) );
  OAI21_X1 U4537 ( .B1(n3859), .B2(n4035), .A(n3858), .ZN(U3265) );
  XNOR2_X1 U4538 ( .A(n3860), .B(n3863), .ZN(n4149) );
  INV_X1 U4539 ( .A(n4149), .ZN(n3878) );
  NAND2_X1 U4540 ( .A1(n3862), .A2(n3861), .ZN(n3864) );
  XNOR2_X1 U4541 ( .A(n3864), .B(n3863), .ZN(n3869) );
  OAI22_X1 U4542 ( .A1(n3865), .A2(n4081), .B1(n4099), .B2(n3871), .ZN(n3866)
         );
  AOI21_X1 U4543 ( .B1(n4078), .B2(n3867), .A(n3866), .ZN(n3868) );
  OAI21_X1 U4544 ( .B1(n3869), .B2(n4109), .A(n3868), .ZN(n4148) );
  INV_X1 U4545 ( .A(n3892), .ZN(n3872) );
  OAI21_X1 U4546 ( .B1(n3872), .B2(n3871), .A(n3870), .ZN(n4226) );
  NOR2_X1 U4547 ( .A1(n4226), .A2(n4066), .ZN(n3876) );
  OAI22_X1 U4548 ( .A1(n4372), .A2(n3874), .B1(n3873), .B2(n4370), .ZN(n3875)
         );
  AOI211_X1 U4549 ( .C1(n4148), .C2(n4372), .A(n3876), .B(n3875), .ZN(n3877)
         );
  OAI21_X1 U4550 ( .B1(n3878), .B2(n4035), .A(n3877), .ZN(U3266) );
  XOR2_X1 U4551 ( .A(n3886), .B(n3879), .Z(n4153) );
  INV_X1 U4552 ( .A(n4153), .ZN(n3900) );
  INV_X1 U4553 ( .A(n3880), .ZN(n3881) );
  NAND2_X1 U4554 ( .A1(n3922), .A2(n3881), .ZN(n3883) );
  NAND2_X1 U4555 ( .A1(n3883), .A2(n3882), .ZN(n3905) );
  INV_X1 U4556 ( .A(n3902), .ZN(n3906) );
  NAND2_X1 U4557 ( .A1(n3905), .A2(n3906), .ZN(n3904) );
  NAND2_X1 U4558 ( .A1(n3904), .A2(n3884), .ZN(n3885) );
  XOR2_X1 U4559 ( .A(n3886), .B(n3885), .Z(n3887) );
  NAND2_X1 U4560 ( .A1(n3887), .A2(n4083), .ZN(n3890) );
  AOI22_X1 U4561 ( .A1(n3888), .A2(n4078), .B1(n4129), .B2(n2147), .ZN(n3889)
         );
  OAI211_X1 U4562 ( .C1(n3891), .C2(n4081), .A(n3890), .B(n3889), .ZN(n4152)
         );
  OAI21_X1 U4563 ( .B1(n4156), .B2(n3893), .A(n3892), .ZN(n4230) );
  NOR2_X1 U4564 ( .A1(n4230), .A2(n4066), .ZN(n3898) );
  INV_X1 U4565 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3896) );
  INV_X1 U4566 ( .A(n3894), .ZN(n3895) );
  OAI22_X1 U4567 ( .A1(n4372), .A2(n3896), .B1(n3895), .B2(n4370), .ZN(n3897)
         );
  AOI211_X1 U4568 ( .C1(n4152), .C2(n4372), .A(n3898), .B(n3897), .ZN(n3899)
         );
  OAI21_X1 U4569 ( .B1(n3900), .B2(n4035), .A(n3899), .ZN(U3267) );
  OAI21_X1 U4570 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(n4161) );
  OAI21_X1 U4571 ( .B1(n3906), .B2(n3905), .A(n3904), .ZN(n3907) );
  NAND2_X1 U4572 ( .A1(n3907), .A2(n4083), .ZN(n3912) );
  OAI22_X1 U4573 ( .A1(n3908), .A2(n4081), .B1(n4099), .B2(n3913), .ZN(n3909)
         );
  AOI21_X1 U4574 ( .B1(n3910), .B2(n4078), .A(n3909), .ZN(n3911) );
  NAND2_X1 U4575 ( .A1(n3912), .A2(n3911), .ZN(n4159) );
  INV_X1 U4576 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3917) );
  NOR2_X1 U4577 ( .A1(n3928), .A2(n3913), .ZN(n4157) );
  OR3_X1 U4578 ( .A1(n4156), .A2(n4157), .A3(n4066), .ZN(n3916) );
  NAND2_X1 U4579 ( .A1(n3914), .A2(n4386), .ZN(n3915) );
  OAI211_X1 U4580 ( .C1(n4372), .C2(n3917), .A(n3916), .B(n3915), .ZN(n3918)
         );
  AOI21_X1 U4581 ( .B1(n4159), .B2(n4372), .A(n3918), .ZN(n3919) );
  OAI21_X1 U4582 ( .B1(n4161), .B2(n4035), .A(n3919), .ZN(U3268) );
  XNOR2_X1 U4583 ( .A(n3920), .B(n3921), .ZN(n4163) );
  INV_X1 U4584 ( .A(n4163), .ZN(n3937) );
  XNOR2_X1 U4585 ( .A(n3922), .B(n3921), .ZN(n3927) );
  OAI22_X1 U4586 ( .A1(n3923), .A2(n4081), .B1(n4099), .B2(n3930), .ZN(n3924)
         );
  AOI21_X1 U4587 ( .B1(n4078), .B2(n3925), .A(n3924), .ZN(n3926) );
  OAI21_X1 U4588 ( .B1(n3927), .B2(n4109), .A(n3926), .ZN(n4162) );
  INV_X1 U4589 ( .A(n3951), .ZN(n3931) );
  INV_X1 U4590 ( .A(n3928), .ZN(n3929) );
  OAI21_X1 U4591 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n4235) );
  NOR2_X1 U4592 ( .A1(n4235), .A2(n4066), .ZN(n3935) );
  OAI22_X1 U4593 ( .A1(n4372), .A2(n3933), .B1(n3932), .B2(n4370), .ZN(n3934)
         );
  AOI211_X1 U4594 ( .C1(n4162), .C2(n4372), .A(n3935), .B(n3934), .ZN(n3936)
         );
  OAI21_X1 U4595 ( .B1(n3937), .B2(n4035), .A(n3936), .ZN(U3269) );
  XNOR2_X1 U4596 ( .A(n3939), .B(n3938), .ZN(n4166) );
  NAND2_X1 U4597 ( .A1(n3941), .A2(n3940), .ZN(n3943) );
  XNOR2_X1 U4598 ( .A(n3943), .B(n3942), .ZN(n3949) );
  AOI22_X1 U4599 ( .A1(n3945), .A2(n4078), .B1(n4129), .B2(n3944), .ZN(n3946)
         );
  OAI21_X1 U4600 ( .B1(n3947), .B2(n4081), .A(n3946), .ZN(n3948) );
  AOI21_X1 U4601 ( .B1(n3949), .B2(n4083), .A(n3948), .ZN(n3950) );
  OAI21_X1 U4602 ( .B1(n4166), .B2(n4102), .A(n3950), .ZN(n4167) );
  NAND2_X1 U4603 ( .A1(n4167), .A2(n4372), .ZN(n3959) );
  INV_X1 U4604 ( .A(n3978), .ZN(n3953) );
  OAI21_X1 U4605 ( .B1(n3953), .B2(n3952), .A(n3951), .ZN(n4239) );
  INV_X1 U4606 ( .A(n4239), .ZN(n3957) );
  OAI22_X1 U4607 ( .A1(n4372), .A2(n3955), .B1(n3954), .B2(n4370), .ZN(n3956)
         );
  AOI21_X1 U4608 ( .B1(n3957), .B2(n4377), .A(n3956), .ZN(n3958) );
  OAI211_X1 U4609 ( .C1(n4166), .C2(n4120), .A(n3959), .B(n3958), .ZN(U3270)
         );
  XNOR2_X1 U4610 ( .A(n3960), .B(n3967), .ZN(n4172) );
  INV_X1 U4611 ( .A(n4172), .ZN(n3983) );
  INV_X1 U4612 ( .A(n3961), .ZN(n3963) );
  OAI21_X1 U4613 ( .B1(n4003), .B2(n3963), .A(n3962), .ZN(n3984) );
  INV_X1 U4614 ( .A(n3964), .ZN(n3966) );
  OAI21_X1 U4615 ( .B1(n3984), .B2(n3966), .A(n3965), .ZN(n3968) );
  XNOR2_X1 U4616 ( .A(n3968), .B(n3967), .ZN(n3969) );
  NAND2_X1 U4617 ( .A1(n3969), .A2(n4083), .ZN(n3973) );
  AOI22_X1 U4618 ( .A1(n3971), .A2(n4078), .B1(n4129), .B2(n3970), .ZN(n3972)
         );
  OAI211_X1 U4619 ( .C1(n3974), .C2(n4081), .A(n3973), .B(n3972), .ZN(n4171)
         );
  OR2_X1 U4620 ( .A1(n3976), .A2(n3975), .ZN(n3977) );
  NAND2_X1 U4621 ( .A1(n3978), .A2(n3977), .ZN(n4243) );
  AOI22_X1 U4622 ( .A1(n4391), .A2(REG2_REG_19__SCAN_IN), .B1(n3979), .B2(
        n4386), .ZN(n3980) );
  OAI21_X1 U4623 ( .B1(n4243), .B2(n4066), .A(n3980), .ZN(n3981) );
  AOI21_X1 U4624 ( .B1(n4171), .B2(n4372), .A(n3981), .ZN(n3982) );
  OAI21_X1 U4625 ( .B1(n3983), .B2(n4035), .A(n3982), .ZN(U3271) );
  XOR2_X1 U4626 ( .A(n3991), .B(n3984), .Z(n3989) );
  AOI22_X1 U4627 ( .A1(n3985), .A2(n4078), .B1(n4129), .B2(n3993), .ZN(n3986)
         );
  OAI21_X1 U4628 ( .B1(n3987), .B2(n4081), .A(n3986), .ZN(n3988) );
  AOI21_X1 U4629 ( .B1(n3989), .B2(n4083), .A(n3988), .ZN(n4177) );
  OAI21_X1 U4630 ( .B1(n3992), .B2(n3991), .A(n3990), .ZN(n4175) );
  XNOR2_X1 U4631 ( .A(n4010), .B(n3993), .ZN(n3994) );
  NAND2_X1 U4632 ( .A1(n3994), .A2(n4443), .ZN(n4176) );
  NOR2_X1 U4633 ( .A1(n4176), .A2(n3995), .ZN(n3999) );
  OAI22_X1 U4634 ( .A1(n4372), .A2(n3997), .B1(n3996), .B2(n4370), .ZN(n3998)
         );
  AOI211_X1 U4635 ( .C1(n4175), .C2(n4068), .A(n3999), .B(n3998), .ZN(n4000)
         );
  OAI21_X1 U4636 ( .B1(n4391), .B2(n4177), .A(n4000), .ZN(U3272) );
  XOR2_X1 U4637 ( .A(n4002), .B(n4001), .Z(n4180) );
  INV_X1 U4638 ( .A(n4180), .ZN(n4018) );
  XNOR2_X1 U4639 ( .A(n4003), .B(n4002), .ZN(n4004) );
  NAND2_X1 U4640 ( .A1(n4004), .A2(n4083), .ZN(n4008) );
  AOI22_X1 U4641 ( .A1(n4006), .A2(n4078), .B1(n4129), .B2(n4005), .ZN(n4007)
         );
  OAI211_X1 U4642 ( .C1(n4036), .C2(n4081), .A(n4008), .B(n4007), .ZN(n4179)
         );
  INV_X1 U4643 ( .A(n4009), .ZN(n4022) );
  INV_X1 U4644 ( .A(n4010), .ZN(n4011) );
  OAI21_X1 U4645 ( .B1(n4022), .B2(n4012), .A(n4011), .ZN(n4248) );
  NOR2_X1 U4646 ( .A1(n4248), .A2(n4066), .ZN(n4016) );
  OAI22_X1 U4647 ( .A1(n4372), .A2(n4014), .B1(n4013), .B2(n4370), .ZN(n4015)
         );
  AOI211_X1 U4648 ( .C1(n4179), .C2(n4372), .A(n4016), .B(n4015), .ZN(n4017)
         );
  OAI21_X1 U4649 ( .B1(n4018), .B2(n4035), .A(n4017), .ZN(U3273) );
  OAI21_X1 U4650 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4186) );
  AOI21_X1 U4651 ( .B1(n4029), .B2(n4023), .A(n4022), .ZN(n4184) );
  OAI22_X1 U4652 ( .A1(n4372), .A2(n4351), .B1(n4024), .B2(n4370), .ZN(n4025)
         );
  AOI21_X1 U4653 ( .B1(n4184), .B2(n4377), .A(n4025), .ZN(n4034) );
  OAI211_X1 U4654 ( .C1(n4028), .C2(n4027), .A(n4026), .B(n4083), .ZN(n4032)
         );
  AOI22_X1 U4655 ( .A1(n4030), .A2(n4078), .B1(n4129), .B2(n4029), .ZN(n4031)
         );
  OAI211_X1 U4656 ( .C1(n4053), .C2(n4081), .A(n4032), .B(n4031), .ZN(n4183)
         );
  NAND2_X1 U4657 ( .A1(n4183), .A2(n4372), .ZN(n4033) );
  OAI211_X1 U4658 ( .C1(n4186), .C2(n4035), .A(n4034), .B(n4033), .ZN(U3274)
         );
  OAI22_X1 U4659 ( .A1(n4036), .A2(n4100), .B1(n4099), .B2(n4042), .ZN(n4041)
         );
  INV_X1 U4660 ( .A(n4037), .ZN(n4038) );
  AOI211_X1 U4661 ( .C1(n4039), .C2(n4047), .A(n4109), .B(n4038), .ZN(n4040)
         );
  AOI211_X1 U4662 ( .C1(n4106), .C2(n4079), .A(n4041), .B(n4040), .ZN(n4189)
         );
  XNOR2_X1 U4663 ( .A(n4062), .B(n4042), .ZN(n4190) );
  INV_X1 U4664 ( .A(n4190), .ZN(n4046) );
  OAI22_X1 U4665 ( .A1(n4372), .A2(n4044), .B1(n4043), .B2(n4370), .ZN(n4045)
         );
  AOI21_X1 U4666 ( .B1(n4046), .B2(n4377), .A(n4045), .ZN(n4050) );
  XNOR2_X1 U4667 ( .A(n4048), .B(n4047), .ZN(n4187) );
  NAND2_X1 U4668 ( .A1(n4187), .A2(n4068), .ZN(n4049) );
  OAI211_X1 U4669 ( .C1(n4189), .C2(n4391), .A(n4050), .B(n4049), .ZN(U3275)
         );
  XNOR2_X1 U4670 ( .A(n4051), .B(n4059), .ZN(n4057) );
  OAI22_X1 U4671 ( .A1(n4053), .A2(n4100), .B1(n4099), .B2(n4052), .ZN(n4054)
         );
  AOI21_X1 U4672 ( .B1(n4106), .B2(n4055), .A(n4054), .ZN(n4056) );
  OAI21_X1 U4673 ( .B1(n4057), .B2(n4109), .A(n4056), .ZN(n4191) );
  INV_X1 U4674 ( .A(n4191), .ZN(n4070) );
  OAI21_X1 U4675 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(n4192) );
  AND2_X1 U4676 ( .A1(n4087), .A2(n4061), .ZN(n4063) );
  OR2_X1 U4677 ( .A1(n4063), .A2(n4062), .ZN(n4254) );
  AOI22_X1 U4678 ( .A1(n4391), .A2(REG2_REG_14__SCAN_IN), .B1(n4064), .B2(
        n4386), .ZN(n4065) );
  OAI21_X1 U4679 ( .B1(n4254), .B2(n4066), .A(n4065), .ZN(n4067) );
  AOI21_X1 U4680 ( .B1(n4192), .B2(n4068), .A(n4067), .ZN(n4069) );
  OAI21_X1 U4681 ( .B1(n4391), .B2(n4070), .A(n4069), .ZN(U3276) );
  XNOR2_X1 U4682 ( .A(n4071), .B(n4076), .ZN(n4194) );
  OAI21_X1 U4683 ( .B1(n4074), .B2(n4073), .A(n4072), .ZN(n4075) );
  XOR2_X1 U4684 ( .A(n4076), .B(n4075), .Z(n4084) );
  AOI22_X1 U4685 ( .A1(n4079), .A2(n4078), .B1(n4129), .B2(n4077), .ZN(n4080)
         );
  OAI21_X1 U4686 ( .B1(n4101), .B2(n4081), .A(n4080), .ZN(n4082) );
  AOI21_X1 U4687 ( .B1(n4084), .B2(n4083), .A(n4082), .ZN(n4085) );
  OAI21_X1 U4688 ( .B1(n4194), .B2(n4102), .A(n4085), .ZN(n4195) );
  NAND2_X1 U4689 ( .A1(n4195), .A2(n4372), .ZN(n4095) );
  INV_X1 U4690 ( .A(n4086), .ZN(n4089) );
  OAI21_X1 U4691 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4258) );
  INV_X1 U4692 ( .A(n4258), .ZN(n4093) );
  OAI22_X1 U4693 ( .A1(n4372), .A2(n4091), .B1(n4090), .B2(n4370), .ZN(n4092)
         );
  AOI21_X1 U4694 ( .B1(n4093), .B2(n4377), .A(n4092), .ZN(n4094) );
  OAI211_X1 U4695 ( .C1(n4194), .C2(n4120), .A(n4095), .B(n4094), .ZN(U3277)
         );
  AOI21_X1 U4696 ( .B1(n4098), .B2(n4096), .A(n2050), .ZN(n4203) );
  XOR2_X1 U4697 ( .A(n4098), .B(n4097), .Z(n4108) );
  OAI22_X1 U4698 ( .A1(n4101), .A2(n4100), .B1(n4099), .B2(n4110), .ZN(n4104)
         );
  NOR2_X1 U4699 ( .A1(n4203), .A2(n4102), .ZN(n4103) );
  AOI211_X1 U4700 ( .C1(n4106), .C2(n4105), .A(n4104), .B(n4103), .ZN(n4107)
         );
  OAI21_X1 U4701 ( .B1(n4109), .B2(n4108), .A(n4107), .ZN(n4204) );
  NAND2_X1 U4702 ( .A1(n4204), .A2(n4372), .ZN(n4119) );
  OR2_X1 U4703 ( .A1(n4111), .A2(n4110), .ZN(n4112) );
  NAND2_X1 U4704 ( .A1(n4113), .A2(n4112), .ZN(n4267) );
  INV_X1 U4705 ( .A(n4267), .ZN(n4117) );
  OAI22_X1 U4706 ( .A1(n4372), .A2(n4115), .B1(n4114), .B2(n4370), .ZN(n4116)
         );
  AOI21_X1 U4707 ( .B1(n4117), .B2(n4377), .A(n4116), .ZN(n4118) );
  OAI211_X1 U4708 ( .C1(n4203), .C2(n4120), .A(n4119), .B(n4118), .ZN(U3279)
         );
  XOR2_X1 U4709 ( .A(n4121), .B(n4126), .Z(n4279) );
  INV_X1 U4710 ( .A(n4279), .ZN(n4210) );
  INV_X1 U4711 ( .A(n4121), .ZN(n4124) );
  AND2_X1 U4712 ( .A1(n4123), .A2(n4122), .ZN(n4128) );
  AOI21_X1 U4713 ( .B1(n4124), .B2(n4129), .A(n4128), .ZN(n4281) );
  MUX2_X1 U4714 ( .A(n3527), .B(n4281), .S(n4454), .Z(n4125) );
  OAI21_X1 U4715 ( .B1(n4210), .B2(n4208), .A(n4125), .ZN(U3549) );
  AOI21_X1 U4716 ( .B1(n4130), .B2(n4127), .A(n4126), .ZN(n4282) );
  INV_X1 U4717 ( .A(n4282), .ZN(n4213) );
  AOI21_X1 U4718 ( .B1(n4130), .B2(n4129), .A(n4128), .ZN(n4284) );
  MUX2_X1 U4719 ( .A(n2921), .B(n4284), .S(n4454), .Z(n4131) );
  OAI21_X1 U4720 ( .B1(n4213), .B2(n4208), .A(n4131), .ZN(U3548) );
  NAND2_X1 U4721 ( .A1(n4132), .A2(n4432), .ZN(n4135) );
  NAND2_X1 U4722 ( .A1(n4136), .A2(n4432), .ZN(n4138) );
  OAI211_X1 U4723 ( .C1(n4415), .C2(n4139), .A(n4138), .B(n4137), .ZN(n4215)
         );
  MUX2_X1 U4724 ( .A(REG1_REG_27__SCAN_IN), .B(n4215), .S(n4454), .Z(U3545) );
  INV_X1 U4725 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4142) );
  AOI21_X1 U4726 ( .B1(n4141), .B2(n4432), .A(n4140), .ZN(n4216) );
  MUX2_X1 U4727 ( .A(n4142), .B(n4216), .S(n4454), .Z(n4143) );
  OAI21_X1 U4728 ( .B1(n4208), .B2(n4218), .A(n4143), .ZN(U3544) );
  INV_X1 U4729 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4146) );
  AOI21_X1 U4730 ( .B1(n4145), .B2(n4432), .A(n4144), .ZN(n4219) );
  MUX2_X1 U4731 ( .A(n4146), .B(n4219), .S(n4454), .Z(n4147) );
  OAI21_X1 U4732 ( .B1(n4208), .B2(n4222), .A(n4147), .ZN(U3543) );
  INV_X1 U4733 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4150) );
  AOI21_X1 U4734 ( .B1(n4149), .B2(n4432), .A(n4148), .ZN(n4223) );
  MUX2_X1 U4735 ( .A(n4150), .B(n4223), .S(n4454), .Z(n4151) );
  OAI21_X1 U4736 ( .B1(n4208), .B2(n4226), .A(n4151), .ZN(U3542) );
  INV_X1 U4737 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4154) );
  AOI21_X1 U4738 ( .B1(n4153), .B2(n4432), .A(n4152), .ZN(n4227) );
  MUX2_X1 U4739 ( .A(n4154), .B(n4227), .S(n4454), .Z(n4155) );
  OAI21_X1 U4740 ( .B1(n4208), .B2(n4230), .A(n4155), .ZN(U3541) );
  NOR3_X1 U4741 ( .A1(n4157), .A2(n4156), .A3(n4415), .ZN(n4158) );
  NOR2_X1 U4742 ( .A1(n4159), .A2(n4158), .ZN(n4160) );
  OAI21_X1 U4743 ( .B1(n4161), .B2(n4438), .A(n4160), .ZN(n4231) );
  MUX2_X1 U4744 ( .A(REG1_REG_22__SCAN_IN), .B(n4231), .S(n4454), .Z(U3540) );
  AOI21_X1 U4745 ( .B1(n4163), .B2(n4432), .A(n4162), .ZN(n4232) );
  MUX2_X1 U4746 ( .A(n4164), .B(n4232), .S(n4454), .Z(n4165) );
  OAI21_X1 U4747 ( .B1(n4208), .B2(n4235), .A(n4165), .ZN(U3539) );
  INV_X1 U4748 ( .A(n4166), .ZN(n4168) );
  AOI21_X1 U4749 ( .B1(n4423), .B2(n4168), .A(n4167), .ZN(n4236) );
  MUX2_X1 U4750 ( .A(n4169), .B(n4236), .S(n4454), .Z(n4170) );
  OAI21_X1 U4751 ( .B1(n4208), .B2(n4239), .A(n4170), .ZN(U3538) );
  AOI21_X1 U4752 ( .B1(n4172), .B2(n4432), .A(n4171), .ZN(n4240) );
  MUX2_X1 U4753 ( .A(n4173), .B(n4240), .S(n4454), .Z(n4174) );
  OAI21_X1 U4754 ( .B1(n4208), .B2(n4243), .A(n4174), .ZN(U3537) );
  INV_X1 U4755 ( .A(n4175), .ZN(n4178) );
  OAI211_X1 U4756 ( .C1(n4178), .C2(n4438), .A(n4177), .B(n4176), .ZN(n4244)
         );
  MUX2_X1 U4757 ( .A(REG1_REG_18__SCAN_IN), .B(n4244), .S(n4454), .Z(U3536) );
  AOI21_X1 U4758 ( .B1(n4180), .B2(n4432), .A(n4179), .ZN(n4245) );
  MUX2_X1 U4759 ( .A(n4181), .B(n4245), .S(n4454), .Z(n4182) );
  OAI21_X1 U4760 ( .B1(n4208), .B2(n4248), .A(n4182), .ZN(U3535) );
  AOI21_X1 U4761 ( .B1(n4443), .B2(n4184), .A(n4183), .ZN(n4185) );
  OAI21_X1 U4762 ( .B1(n4186), .B2(n4438), .A(n4185), .ZN(n4249) );
  MUX2_X1 U4763 ( .A(REG1_REG_16__SCAN_IN), .B(n4249), .S(n4454), .Z(U3534) );
  NAND2_X1 U4764 ( .A1(n4187), .A2(n4432), .ZN(n4188) );
  OAI211_X1 U4765 ( .C1(n4190), .C2(n4415), .A(n4189), .B(n4188), .ZN(n4250)
         );
  MUX2_X1 U4766 ( .A(REG1_REG_15__SCAN_IN), .B(n4250), .S(n4454), .Z(U3533) );
  AOI21_X1 U4767 ( .B1(n4192), .B2(n4432), .A(n4191), .ZN(n4251) );
  MUX2_X1 U4768 ( .A(n4326), .B(n4251), .S(n4454), .Z(n4193) );
  OAI21_X1 U4769 ( .B1(n4208), .B2(n4254), .A(n4193), .ZN(U3532) );
  INV_X1 U4770 ( .A(n4194), .ZN(n4196) );
  AOI21_X1 U4771 ( .B1(n4423), .B2(n4196), .A(n4195), .ZN(n4255) );
  MUX2_X1 U4772 ( .A(n4197), .B(n4255), .S(n4454), .Z(n4198) );
  OAI21_X1 U4773 ( .B1(n4208), .B2(n4258), .A(n4198), .ZN(U3531) );
  NAND2_X1 U4774 ( .A1(n4199), .A2(n4432), .ZN(n4201) );
  AND2_X1 U4775 ( .A1(n4201), .A2(n4200), .ZN(n4259) );
  MUX2_X1 U4776 ( .A(n4259), .B(n4305), .S(n4452), .Z(n4202) );
  OAI21_X1 U4777 ( .B1(n4208), .B2(n4262), .A(n4202), .ZN(U3530) );
  INV_X1 U4778 ( .A(n4203), .ZN(n4205) );
  AOI21_X1 U4779 ( .B1(n4423), .B2(n4205), .A(n4204), .ZN(n4263) );
  MUX2_X1 U4780 ( .A(n4206), .B(n4263), .S(n4454), .Z(n4207) );
  OAI21_X1 U4781 ( .B1(n4208), .B2(n4267), .A(n4207), .ZN(U3529) );
  INV_X1 U4782 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4600) );
  MUX2_X1 U4783 ( .A(n4600), .B(n4281), .S(n4446), .Z(n4209) );
  OAI21_X1 U4784 ( .B1(n4210), .B2(n4266), .A(n4209), .ZN(U3517) );
  INV_X1 U4785 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4211) );
  MUX2_X1 U4786 ( .A(n4211), .B(n4284), .S(n4446), .Z(n4212) );
  OAI21_X1 U4787 ( .B1(n4213), .B2(n4266), .A(n4212), .ZN(U3516) );
  MUX2_X1 U4788 ( .A(REG0_REG_29__SCAN_IN), .B(n4214), .S(n4446), .Z(U3515) );
  MUX2_X1 U4789 ( .A(REG0_REG_27__SCAN_IN), .B(n4215), .S(n4446), .Z(U3513) );
  MUX2_X1 U4790 ( .A(n4533), .B(n4216), .S(n4446), .Z(n4217) );
  OAI21_X1 U4791 ( .B1(n4218), .B2(n4266), .A(n4217), .ZN(U3512) );
  INV_X1 U4792 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4220) );
  MUX2_X1 U4793 ( .A(n4220), .B(n4219), .S(n4446), .Z(n4221) );
  OAI21_X1 U4794 ( .B1(n4222), .B2(n4266), .A(n4221), .ZN(U3511) );
  INV_X1 U4795 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4224) );
  MUX2_X1 U4796 ( .A(n4224), .B(n4223), .S(n4446), .Z(n4225) );
  OAI21_X1 U4797 ( .B1(n4226), .B2(n4266), .A(n4225), .ZN(U3510) );
  INV_X1 U4798 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4228) );
  MUX2_X1 U4799 ( .A(n4228), .B(n4227), .S(n4446), .Z(n4229) );
  OAI21_X1 U4800 ( .B1(n4230), .B2(n4266), .A(n4229), .ZN(U3509) );
  MUX2_X1 U4801 ( .A(REG0_REG_22__SCAN_IN), .B(n4231), .S(n4446), .Z(U3508) );
  INV_X1 U4802 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4233) );
  MUX2_X1 U4803 ( .A(n4233), .B(n4232), .S(n4446), .Z(n4234) );
  OAI21_X1 U4804 ( .B1(n4235), .B2(n4266), .A(n4234), .ZN(U3507) );
  INV_X1 U4805 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4237) );
  MUX2_X1 U4806 ( .A(n4237), .B(n4236), .S(n4446), .Z(n4238) );
  OAI21_X1 U4807 ( .B1(n4239), .B2(n4266), .A(n4238), .ZN(U3506) );
  INV_X1 U4808 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4241) );
  MUX2_X1 U4809 ( .A(n4241), .B(n4240), .S(n4446), .Z(n4242) );
  OAI21_X1 U4810 ( .B1(n4243), .B2(n4266), .A(n4242), .ZN(U3505) );
  MUX2_X1 U4811 ( .A(REG0_REG_18__SCAN_IN), .B(n4244), .S(n4446), .Z(U3503) );
  INV_X1 U4812 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4246) );
  MUX2_X1 U4813 ( .A(n4246), .B(n4245), .S(n4446), .Z(n4247) );
  OAI21_X1 U4814 ( .B1(n4248), .B2(n4266), .A(n4247), .ZN(U3501) );
  MUX2_X1 U4815 ( .A(REG0_REG_16__SCAN_IN), .B(n4249), .S(n4446), .Z(U3499) );
  MUX2_X1 U4816 ( .A(REG0_REG_15__SCAN_IN), .B(n4250), .S(n4446), .Z(U3497) );
  INV_X1 U4817 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4252) );
  MUX2_X1 U4818 ( .A(n4252), .B(n4251), .S(n4446), .Z(n4253) );
  OAI21_X1 U4819 ( .B1(n4254), .B2(n4266), .A(n4253), .ZN(U3495) );
  INV_X1 U4820 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4256) );
  MUX2_X1 U4821 ( .A(n4256), .B(n4255), .S(n4446), .Z(n4257) );
  OAI21_X1 U4822 ( .B1(n4258), .B2(n4266), .A(n4257), .ZN(U3493) );
  INV_X1 U4823 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4260) );
  MUX2_X1 U4824 ( .A(n4260), .B(n4259), .S(n4446), .Z(n4261) );
  OAI21_X1 U4825 ( .B1(n4262), .B2(n4266), .A(n4261), .ZN(U3491) );
  INV_X1 U4826 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4264) );
  MUX2_X1 U4827 ( .A(n4264), .B(n4263), .S(n4446), .Z(n4265) );
  OAI21_X1 U4828 ( .B1(n4267), .B2(n4266), .A(n4265), .ZN(U3489) );
  MUX2_X1 U4829 ( .A(n4268), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4830 ( .A(n4269), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4831 ( .A(n4270), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4832 ( .A(n4271), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4833 ( .A(n4272), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4834 ( .A(DATAI_4_), .B(n4273), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4835 ( .A(DATAI_3_), .B(n4274), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4836 ( .A(DATAI_2_), .B(n4275), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U4837 ( .A(n4276), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4838 ( .A(DATAI_28_), .ZN(n4277) );
  AOI22_X1 U4839 ( .A1(STATE_REG_SCAN_IN), .A2(n4278), .B1(n4277), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4840 ( .A1(n4279), .A2(n4377), .B1(n4391), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4280) );
  OAI21_X1 U4841 ( .B1(n4391), .B2(n4281), .A(n4280), .ZN(U3260) );
  AOI22_X1 U4842 ( .A1(n4282), .A2(n4377), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4391), .ZN(n4283) );
  OAI21_X1 U4843 ( .B1(n4391), .B2(n4284), .A(n4283), .ZN(U3261) );
  AOI211_X1 U4844 ( .C1(n2384), .C2(n4285), .A(n2057), .B(n4455), .ZN(n4288)
         );
  INV_X1 U4845 ( .A(n4286), .ZN(n4287) );
  AOI211_X1 U4846 ( .C1(n4461), .C2(ADDR_REG_8__SCAN_IN), .A(n4288), .B(n4287), 
        .ZN(n4292) );
  OAI211_X1 U4847 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4290), .A(n4463), .B(n4289), 
        .ZN(n4291) );
  OAI211_X1 U4848 ( .C1(n4468), .C2(n4408), .A(n4292), .B(n4291), .ZN(U3248)
         );
  AOI211_X1 U4849 ( .C1(n4295), .C2(n4294), .A(n4293), .B(n4455), .ZN(n4297)
         );
  AOI211_X1 U4850 ( .C1(n4461), .C2(ADDR_REG_11__SCAN_IN), .A(n4297), .B(n4296), .ZN(n4302) );
  OAI211_X1 U4851 ( .C1(n4300), .C2(n4299), .A(n4463), .B(n4298), .ZN(n4301)
         );
  OAI211_X1 U4852 ( .C1(n4468), .C2(n4406), .A(n4302), .B(n4301), .ZN(U3251)
         );
  AOI211_X1 U4853 ( .C1(n4305), .C2(n4304), .A(n4303), .B(n4455), .ZN(n4308)
         );
  INV_X1 U4854 ( .A(n4306), .ZN(n4307) );
  AOI211_X1 U4855 ( .C1(n4461), .C2(ADDR_REG_12__SCAN_IN), .A(n4308), .B(n4307), .ZN(n4312) );
  OAI211_X1 U4856 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4310), .A(n4463), .B(n4309), .ZN(n4311) );
  OAI211_X1 U4857 ( .C1(n4468), .C2(n4405), .A(n4312), .B(n4311), .ZN(U3252)
         );
  AOI211_X1 U4858 ( .C1(n4315), .C2(n4314), .A(n4313), .B(n4455), .ZN(n4317)
         );
  AOI211_X1 U4859 ( .C1(n4461), .C2(ADDR_REG_13__SCAN_IN), .A(n4317), .B(n4316), .ZN(n4323) );
  AOI21_X1 U4860 ( .B1(n4091), .B2(n4403), .A(n4318), .ZN(n4321) );
  INV_X1 U4861 ( .A(n4463), .ZN(n4327) );
  AOI21_X1 U4862 ( .B1(n4321), .B2(n4320), .A(n4327), .ZN(n4319) );
  OAI21_X1 U4863 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4322) );
  OAI211_X1 U4864 ( .C1(n4468), .C2(n4403), .A(n4323), .B(n4322), .ZN(U3253)
         );
  NAND2_X1 U4865 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4461), .ZN(n4336) );
  AOI211_X1 U4866 ( .C1(n4326), .C2(n4325), .A(n4324), .B(n4455), .ZN(n4331)
         );
  AOI211_X1 U4867 ( .C1(n2461), .C2(n4329), .A(n4328), .B(n4327), .ZN(n4330)
         );
  AOI211_X1 U4868 ( .C1(n4333), .C2(n4332), .A(n4331), .B(n4330), .ZN(n4335)
         );
  NAND3_X1 U4869 ( .A1(n4336), .A2(n4335), .A3(n4334), .ZN(U3254) );
  AOI211_X1 U4870 ( .C1(n4339), .C2(n4338), .A(n4337), .B(n4455), .ZN(n4340)
         );
  AOI211_X1 U4871 ( .C1(n4461), .C2(ADDR_REG_15__SCAN_IN), .A(n4341), .B(n4340), .ZN(n4347) );
  AOI21_X1 U4872 ( .B1(n4344), .B2(n4343), .A(n4342), .ZN(n4345) );
  NAND2_X1 U4873 ( .A1(n4463), .A2(n4345), .ZN(n4346) );
  OAI211_X1 U4874 ( .C1(n4468), .C2(n4400), .A(n4347), .B(n4346), .ZN(U3255)
         );
  INV_X1 U4875 ( .A(n4348), .ZN(n4349) );
  AOI21_X1 U4876 ( .B1(n4461), .B2(ADDR_REG_16__SCAN_IN), .A(n4349), .ZN(n4360) );
  OAI21_X1 U4877 ( .B1(n4352), .B2(n4351), .A(n4350), .ZN(n4358) );
  OAI21_X1 U4878 ( .B1(n4355), .B2(n4354), .A(n4353), .ZN(n4356) );
  AOI22_X1 U4879 ( .A1(n4463), .A2(n4358), .B1(n4357), .B2(n4356), .ZN(n4359)
         );
  OAI211_X1 U4880 ( .C1(n4398), .C2(n4468), .A(n4360), .B(n4359), .ZN(U3256)
         );
  AOI21_X1 U4881 ( .B1(n4366), .B2(n4365), .A(n4364), .ZN(n4367) );
  NAND2_X1 U4882 ( .A1(n4463), .A2(n4367), .ZN(n4368) );
  OAI211_X1 U4883 ( .C1(n4468), .C2(n4396), .A(n4369), .B(n4368), .ZN(U3258)
         );
  OAI22_X1 U4884 ( .A1(n4372), .A2(n2976), .B1(n4371), .B2(n4370), .ZN(n4373)
         );
  INV_X1 U4885 ( .A(n4373), .ZN(n4380) );
  INV_X1 U4886 ( .A(n4374), .ZN(n4378) );
  INV_X1 U4887 ( .A(n4375), .ZN(n4376) );
  AOI22_X1 U4888 ( .A1(n4378), .A2(n4388), .B1(n4377), .B2(n4376), .ZN(n4379)
         );
  OAI211_X1 U4889 ( .C1(n4391), .C2(n4381), .A(n4380), .B(n4379), .ZN(U3284)
         );
  INV_X1 U4890 ( .A(n4382), .ZN(n4384) );
  AOI21_X1 U4891 ( .B1(n4385), .B2(n4384), .A(n4383), .ZN(n4390) );
  AOI22_X1 U4892 ( .A1(n4388), .A2(n4387), .B1(REG3_REG_0__SCAN_IN), .B2(n4386), .ZN(n4389) );
  OAI221_X1 U4893 ( .B1(n4391), .B2(n4390), .C1(n4372), .C2(n3683), .A(n4389), 
        .ZN(U3290) );
  INV_X1 U4894 ( .A(D_REG_31__SCAN_IN), .ZN(n4488) );
  NOR2_X1 U4895 ( .A1(n4392), .A2(n4488), .ZN(U3291) );
  AND2_X1 U4896 ( .A1(D_REG_30__SCAN_IN), .A2(n4393), .ZN(U3292) );
  AND2_X1 U4897 ( .A1(D_REG_29__SCAN_IN), .A2(n4393), .ZN(U3293) );
  AND2_X1 U4898 ( .A1(D_REG_28__SCAN_IN), .A2(n4393), .ZN(U3294) );
  AND2_X1 U4899 ( .A1(D_REG_27__SCAN_IN), .A2(n4393), .ZN(U3295) );
  AND2_X1 U4900 ( .A1(D_REG_26__SCAN_IN), .A2(n4393), .ZN(U3296) );
  AND2_X1 U4901 ( .A1(D_REG_25__SCAN_IN), .A2(n4393), .ZN(U3297) );
  AND2_X1 U4902 ( .A1(D_REG_24__SCAN_IN), .A2(n4393), .ZN(U3298) );
  AND2_X1 U4903 ( .A1(D_REG_23__SCAN_IN), .A2(n4393), .ZN(U3299) );
  INV_X1 U4904 ( .A(D_REG_22__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U4905 ( .A1(n4392), .A2(n4486), .ZN(U3300) );
  INV_X1 U4906 ( .A(D_REG_21__SCAN_IN), .ZN(n4492) );
  NOR2_X1 U4907 ( .A1(n4392), .A2(n4492), .ZN(U3301) );
  AND2_X1 U4908 ( .A1(D_REG_20__SCAN_IN), .A2(n4393), .ZN(U3302) );
  AND2_X1 U4909 ( .A1(D_REG_19__SCAN_IN), .A2(n4393), .ZN(U3303) );
  AND2_X1 U4910 ( .A1(D_REG_18__SCAN_IN), .A2(n4393), .ZN(U3304) );
  AND2_X1 U4911 ( .A1(D_REG_17__SCAN_IN), .A2(n4393), .ZN(U3305) );
  AND2_X1 U4912 ( .A1(D_REG_16__SCAN_IN), .A2(n4393), .ZN(U3306) );
  AND2_X1 U4913 ( .A1(D_REG_15__SCAN_IN), .A2(n4393), .ZN(U3307) );
  AND2_X1 U4914 ( .A1(D_REG_14__SCAN_IN), .A2(n4393), .ZN(U3308) );
  INV_X1 U4915 ( .A(D_REG_13__SCAN_IN), .ZN(n4528) );
  NOR2_X1 U4916 ( .A1(n4392), .A2(n4528), .ZN(U3309) );
  AND2_X1 U4917 ( .A1(D_REG_12__SCAN_IN), .A2(n4393), .ZN(U3310) );
  AND2_X1 U4918 ( .A1(D_REG_11__SCAN_IN), .A2(n4393), .ZN(U3311) );
  INV_X1 U4919 ( .A(D_REG_10__SCAN_IN), .ZN(n4491) );
  NOR2_X1 U4920 ( .A1(n4392), .A2(n4491), .ZN(U3312) );
  AND2_X1 U4921 ( .A1(D_REG_9__SCAN_IN), .A2(n4393), .ZN(U3313) );
  AND2_X1 U4922 ( .A1(D_REG_8__SCAN_IN), .A2(n4393), .ZN(U3314) );
  INV_X1 U4923 ( .A(D_REG_7__SCAN_IN), .ZN(n4489) );
  NOR2_X1 U4924 ( .A1(n4392), .A2(n4489), .ZN(U3315) );
  AND2_X1 U4925 ( .A1(D_REG_6__SCAN_IN), .A2(n4393), .ZN(U3316) );
  AND2_X1 U4926 ( .A1(D_REG_5__SCAN_IN), .A2(n4393), .ZN(U3317) );
  AND2_X1 U4927 ( .A1(D_REG_4__SCAN_IN), .A2(n4393), .ZN(U3318) );
  AND2_X1 U4928 ( .A1(D_REG_3__SCAN_IN), .A2(n4393), .ZN(U3319) );
  AND2_X1 U4929 ( .A1(D_REG_2__SCAN_IN), .A2(n4393), .ZN(U3320) );
  INV_X1 U4930 ( .A(DATAI_23_), .ZN(n4395) );
  AOI21_X1 U4931 ( .B1(U3149), .B2(n4395), .A(n4394), .ZN(U3329) );
  INV_X1 U4932 ( .A(DATAI_18_), .ZN(n4584) );
  AOI22_X1 U4933 ( .A1(STATE_REG_SCAN_IN), .A2(n4396), .B1(n4584), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U4934 ( .A(DATAI_16_), .ZN(n4397) );
  AOI22_X1 U4935 ( .A1(STATE_REG_SCAN_IN), .A2(n4398), .B1(n4397), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4936 ( .A(DATAI_15_), .ZN(n4399) );
  AOI22_X1 U4937 ( .A1(STATE_REG_SCAN_IN), .A2(n4400), .B1(n4399), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U4938 ( .A(DATAI_14_), .ZN(n4604) );
  AOI22_X1 U4939 ( .A1(STATE_REG_SCAN_IN), .A2(n4401), .B1(n4604), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U4940 ( .A1(STATE_REG_SCAN_IN), .A2(n4403), .B1(n4402), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U4941 ( .A1(STATE_REG_SCAN_IN), .A2(n4405), .B1(n4404), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U4942 ( .A(DATAI_11_), .ZN(n4603) );
  AOI22_X1 U4943 ( .A1(STATE_REG_SCAN_IN), .A2(n4406), .B1(n4603), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U4944 ( .A(DATAI_10_), .ZN(n4407) );
  AOI22_X1 U4945 ( .A1(STATE_REG_SCAN_IN), .A2(n4467), .B1(n4407), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U4946 ( .A1(STATE_REG_SCAN_IN), .A2(n4408), .B1(n2395), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U4947 ( .A(DATAI_0_), .ZN(n4410) );
  AOI22_X1 U4948 ( .A1(STATE_REG_SCAN_IN), .A2(n2317), .B1(n4410), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U4949 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4950 ( .A1(n4446), .A2(n4412), .B1(n4411), .B2(n4444), .ZN(U3467)
         );
  INV_X1 U4951 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U4952 ( .A1(n4446), .A2(n4413), .B1(n4477), .B2(n4444), .ZN(U3469)
         );
  OAI22_X1 U4953 ( .A1(n4417), .A2(n4416), .B1(n4415), .B2(n4414), .ZN(n4418)
         );
  NOR2_X1 U4954 ( .A1(n4419), .A2(n4418), .ZN(n4448) );
  AOI22_X1 U4955 ( .A1(n4446), .A2(n4448), .B1(n2332), .B2(n4444), .ZN(U3473)
         );
  INV_X1 U4956 ( .A(n4420), .ZN(n4422) );
  AOI211_X1 U4957 ( .C1(n4424), .C2(n4423), .A(n4422), .B(n4421), .ZN(n4449)
         );
  INV_X1 U4958 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U4959 ( .A1(n4446), .A2(n4449), .B1(n4425), .B2(n4444), .ZN(U3475)
         );
  NOR2_X1 U4960 ( .A1(n4426), .A2(n4438), .ZN(n4429) );
  INV_X1 U4961 ( .A(n4427), .ZN(n4428) );
  AOI211_X1 U4962 ( .C1(n4443), .C2(n4430), .A(n4429), .B(n4428), .ZN(n4450)
         );
  INV_X1 U4963 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U4964 ( .A1(n4446), .A2(n4450), .B1(n4431), .B2(n4444), .ZN(U3477)
         );
  NAND3_X1 U4965 ( .A1(n3183), .A2(n4433), .A3(n4432), .ZN(n4434) );
  AND3_X1 U4966 ( .A1(n4436), .A2(n4435), .A3(n4434), .ZN(n4451) );
  INV_X1 U4967 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U4968 ( .A1(n4446), .A2(n4451), .B1(n4437), .B2(n4444), .ZN(U3481)
         );
  NOR2_X1 U4969 ( .A1(n4439), .A2(n4438), .ZN(n4441) );
  AOI211_X1 U4970 ( .C1(n4443), .C2(n4442), .A(n4441), .B(n4440), .ZN(n4453)
         );
  INV_X1 U4971 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4972 ( .A1(n4446), .A2(n4453), .B1(n4445), .B2(n4444), .ZN(U3485)
         );
  INV_X1 U4973 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U4974 ( .A1(n4454), .A2(n4448), .B1(n4447), .B2(n4452), .ZN(U3521)
         );
  AOI22_X1 U4975 ( .A1(n4454), .A2(n4449), .B1(n2948), .B2(n4452), .ZN(U3522)
         );
  AOI22_X1 U4976 ( .A1(n4454), .A2(n4450), .B1(n2951), .B2(n4452), .ZN(U3523)
         );
  AOI22_X1 U4977 ( .A1(n4454), .A2(n4451), .B1(n2373), .B2(n4452), .ZN(U3525)
         );
  AOI22_X1 U4978 ( .A1(n4454), .A2(n4453), .B1(n3009), .B2(n4452), .ZN(U3527)
         );
  AOI211_X1 U4979 ( .C1(n4458), .C2(n4457), .A(n4456), .B(n4455), .ZN(n4460)
         );
  AOI211_X1 U4980 ( .C1(n4461), .C2(ADDR_REG_10__SCAN_IN), .A(n4460), .B(n4459), .ZN(n4466) );
  OAI211_X1 U4981 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4464), .A(n4463), .B(n4462), .ZN(n4465) );
  OAI211_X1 U4982 ( .C1(n4468), .C2(n4467), .A(n4466), .B(n4465), .ZN(n4621)
         );
  INV_X1 U4983 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4471) );
  INV_X1 U4984 ( .A(keyinput43), .ZN(n4470) );
  AOI22_X1 U4985 ( .A1(n4471), .A2(keyinput30), .B1(ADDR_REG_13__SCAN_IN), 
        .B2(n4470), .ZN(n4469) );
  OAI221_X1 U4986 ( .B1(n4471), .B2(keyinput30), .C1(n4470), .C2(
        ADDR_REG_13__SCAN_IN), .A(n4469), .ZN(n4481) );
  INV_X1 U4987 ( .A(keyinput23), .ZN(n4473) );
  AOI22_X1 U4988 ( .A1(n4091), .A2(keyinput32), .B1(ADDR_REG_17__SCAN_IN), 
        .B2(n4473), .ZN(n4472) );
  OAI221_X1 U4989 ( .B1(n4091), .B2(keyinput32), .C1(n4473), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4472), .ZN(n4480) );
  AOI22_X1 U4990 ( .A1(n4115), .A2(keyinput63), .B1(keyinput60), .B2(n3291), 
        .ZN(n4474) );
  OAI221_X1 U4991 ( .B1(n4115), .B2(keyinput63), .C1(n3291), .C2(keyinput60), 
        .A(n4474), .ZN(n4479) );
  AOI22_X1 U4992 ( .A1(n4477), .A2(keyinput25), .B1(n4476), .B2(keyinput52), 
        .ZN(n4475) );
  OAI221_X1 U4993 ( .B1(n4477), .B2(keyinput25), .C1(n4476), .C2(keyinput52), 
        .A(n4475), .ZN(n4478) );
  NOR4_X1 U4994 ( .A1(n4481), .A2(n4480), .A3(n4479), .A4(n4478), .ZN(n4619)
         );
  AOI22_X1 U4995 ( .A1(n4484), .A2(keyinput22), .B1(keyinput50), .B2(n4483), 
        .ZN(n4482) );
  OAI221_X1 U4996 ( .B1(n4484), .B2(keyinput22), .C1(n4483), .C2(keyinput50), 
        .A(n4482), .ZN(n4496) );
  AOI22_X1 U4997 ( .A1(n3269), .A2(keyinput37), .B1(n4486), .B2(keyinput24), 
        .ZN(n4485) );
  OAI221_X1 U4998 ( .B1(n3269), .B2(keyinput37), .C1(n4486), .C2(keyinput24), 
        .A(n4485), .ZN(n4495) );
  AOI22_X1 U4999 ( .A1(n4489), .A2(keyinput28), .B1(keyinput11), .B2(n4488), 
        .ZN(n4487) );
  OAI221_X1 U5000 ( .B1(n4489), .B2(keyinput28), .C1(n4488), .C2(keyinput11), 
        .A(n4487), .ZN(n4494) );
  AOI22_X1 U5001 ( .A1(n4492), .A2(keyinput46), .B1(keyinput0), .B2(n4491), 
        .ZN(n4490) );
  OAI221_X1 U5002 ( .B1(n4492), .B2(keyinput46), .C1(n4491), .C2(keyinput0), 
        .A(n4490), .ZN(n4493) );
  NOR4_X1 U5003 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), .ZN(n4618)
         );
  INV_X1 U5004 ( .A(keyinput55), .ZN(n4564) );
  AOI22_X1 U5005 ( .A1(n3022), .A2(keyinput40), .B1(ADDR_REG_19__SCAN_IN), 
        .B2(n4564), .ZN(n4497) );
  OAI221_X1 U5006 ( .B1(n3022), .B2(keyinput40), .C1(n4564), .C2(
        ADDR_REG_19__SCAN_IN), .A(n4497), .ZN(n4522) );
  INV_X1 U5007 ( .A(keyinput42), .ZN(n4500) );
  INV_X1 U5008 ( .A(keyinput51), .ZN(n4499) );
  AOI22_X1 U5009 ( .A1(n4500), .A2(DATAO_REG_8__SCAN_IN), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n4499), .ZN(n4498) );
  OAI221_X1 U5010 ( .B1(n4500), .B2(DATAO_REG_8__SCAN_IN), .C1(n4499), .C2(
        DATAO_REG_3__SCAN_IN), .A(n4498), .ZN(n4521) );
  INV_X1 U5011 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4506) );
  INV_X1 U5012 ( .A(keyinput14), .ZN(n4503) );
  INV_X1 U5013 ( .A(keyinput62), .ZN(n4502) );
  OAI22_X1 U5014 ( .A1(n4503), .A2(DATAO_REG_13__SCAN_IN), .B1(n4502), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n4501) );
  AOI221_X1 U5015 ( .B1(n4503), .B2(DATAO_REG_13__SCAN_IN), .C1(
        DATAO_REG_15__SCAN_IN), .C2(n4502), .A(n4501), .ZN(n4505) );
  XNOR2_X1 U5016 ( .A(REG2_REG_17__SCAN_IN), .B(keyinput20), .ZN(n4504) );
  OAI211_X1 U5017 ( .C1(keyinput35), .C2(n4506), .A(n4505), .B(n4504), .ZN(
        n4520) );
  INV_X1 U5018 ( .A(keyinput58), .ZN(n4509) );
  INV_X1 U5019 ( .A(keyinput5), .ZN(n4508) );
  OAI22_X1 U5020 ( .A1(n4509), .A2(DATAO_REG_14__SCAN_IN), .B1(n4508), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n4507) );
  AOI221_X1 U5021 ( .B1(n4509), .B2(DATAO_REG_14__SCAN_IN), .C1(
        DATAO_REG_7__SCAN_IN), .C2(n4508), .A(n4507), .ZN(n4518) );
  OAI22_X1 U5022 ( .A1(n4511), .A2(keyinput36), .B1(n3815), .B2(keyinput12), 
        .ZN(n4510) );
  AOI221_X1 U5023 ( .B1(n4511), .B2(keyinput36), .C1(keyinput12), .C2(n3815), 
        .A(n4510), .ZN(n4517) );
  OAI22_X1 U5024 ( .A1(n2317), .A2(keyinput44), .B1(n2976), .B2(keyinput4), 
        .ZN(n4512) );
  AOI221_X1 U5025 ( .B1(n2317), .B2(keyinput44), .C1(keyinput4), .C2(n2976), 
        .A(n4512), .ZN(n4516) );
  INV_X1 U5026 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4514) );
  INV_X1 U5027 ( .A(keyinput3), .ZN(n4559) );
  OAI22_X1 U5028 ( .A1(n4514), .A2(keyinput19), .B1(n4559), .B2(
        ADDR_REG_7__SCAN_IN), .ZN(n4513) );
  AOI221_X1 U5029 ( .B1(n4514), .B2(keyinput19), .C1(ADDR_REG_7__SCAN_IN), 
        .C2(n4559), .A(n4513), .ZN(n4515) );
  NAND4_X1 U5030 ( .A1(n4518), .A2(n4517), .A3(n4516), .A4(n4515), .ZN(n4519)
         );
  NOR4_X1 U5031 ( .A1(n4522), .A2(n4521), .A3(n4520), .A4(n4519), .ZN(n4617)
         );
  INV_X1 U5032 ( .A(keyinput18), .ZN(n4525) );
  INV_X1 U5033 ( .A(keyinput38), .ZN(n4524) );
  AOI22_X1 U5034 ( .A1(n4525), .A2(DATAO_REG_18__SCAN_IN), .B1(
        DATAO_REG_19__SCAN_IN), .B2(n4524), .ZN(n4523) );
  OAI221_X1 U5035 ( .B1(n4525), .B2(DATAO_REG_18__SCAN_IN), .C1(n4524), .C2(
        DATAO_REG_19__SCAN_IN), .A(n4523), .ZN(n4615) );
  AOI22_X1 U5036 ( .A1(n4528), .A2(keyinput29), .B1(keyinput48), .B2(n4527), 
        .ZN(n4526) );
  OAI221_X1 U5037 ( .B1(n4528), .B2(keyinput29), .C1(n4527), .C2(keyinput48), 
        .A(n4526), .ZN(n4614) );
  INV_X1 U5038 ( .A(keyinput34), .ZN(n4530) );
  AOI22_X1 U5039 ( .A1(n4531), .A2(keyinput9), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n4530), .ZN(n4529) );
  OAI221_X1 U5040 ( .B1(n4531), .B2(keyinput9), .C1(n4530), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4529), .ZN(n4539) );
  AOI22_X1 U5041 ( .A1(n3896), .A2(keyinput53), .B1(n4533), .B2(keyinput1), 
        .ZN(n4532) );
  OAI221_X1 U5042 ( .B1(n3896), .B2(keyinput53), .C1(n4533), .C2(keyinput1), 
        .A(n4532), .ZN(n4538) );
  XNOR2_X1 U5043 ( .A(n4534), .B(keyinput17), .ZN(n4537) );
  XNOR2_X1 U5044 ( .A(n4535), .B(keyinput31), .ZN(n4536) );
  NOR4_X1 U5045 ( .A1(n4539), .A2(n4538), .A3(n4537), .A4(n4536), .ZN(n4552)
         );
  INV_X1 U5046 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4542) );
  INV_X1 U5047 ( .A(keyinput39), .ZN(n4541) );
  OAI22_X1 U5048 ( .A1(n4542), .A2(keyinput49), .B1(n4541), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4540) );
  AOI221_X1 U5049 ( .B1(n4542), .B2(keyinput49), .C1(DATAO_REG_30__SCAN_IN), 
        .C2(n4541), .A(n4540), .ZN(n4551) );
  XOR2_X1 U5050 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput26), .Z(n4549) );
  INV_X1 U5051 ( .A(keyinput27), .ZN(n4543) );
  XNOR2_X1 U5052 ( .A(n4543), .B(ADDR_REG_10__SCAN_IN), .ZN(n4548) );
  XNOR2_X1 U5053 ( .A(n4544), .B(keyinput59), .ZN(n4547) );
  XNOR2_X1 U5054 ( .A(n4545), .B(keyinput16), .ZN(n4546) );
  NOR4_X1 U5055 ( .A1(n4549), .A2(n4548), .A3(n4547), .A4(n4546), .ZN(n4550)
         );
  NAND3_X1 U5056 ( .A1(n4552), .A2(n4551), .A3(n4550), .ZN(n4613) );
  NAND2_X1 U5057 ( .A1(keyinput1), .A2(keyinput27), .ZN(n4558) );
  NOR2_X1 U5058 ( .A1(keyinput17), .A2(keyinput59), .ZN(n4556) );
  NAND3_X1 U5059 ( .A1(keyinput0), .A2(keyinput29), .A3(keyinput18), .ZN(n4554) );
  NAND3_X1 U5060 ( .A1(keyinput38), .A2(keyinput34), .A3(keyinput53), .ZN(
        n4553) );
  NOR4_X1 U5061 ( .A1(keyinput48), .A2(keyinput9), .A3(n4554), .A4(n4553), 
        .ZN(n4555) );
  NAND4_X1 U5062 ( .A1(keyinput26), .A2(keyinput16), .A3(n4556), .A4(n4555), 
        .ZN(n4557) );
  NOR4_X1 U5063 ( .A1(keyinput49), .A2(keyinput39), .A3(n4558), .A4(n4557), 
        .ZN(n4581) );
  NAND2_X1 U5064 ( .A1(keyinput51), .A2(keyinput14), .ZN(n4563) );
  NOR2_X1 U5065 ( .A1(keyinput58), .A2(keyinput5), .ZN(n4561) );
  NOR4_X1 U5066 ( .A1(keyinput12), .A2(keyinput44), .A3(keyinput4), .A4(n4559), 
        .ZN(n4560) );
  NAND4_X1 U5067 ( .A1(keyinput62), .A2(keyinput36), .A3(n4561), .A4(n4560), 
        .ZN(n4562) );
  NOR4_X1 U5068 ( .A1(keyinput40), .A2(keyinput42), .A3(n4563), .A4(n4562), 
        .ZN(n4565) );
  NAND4_X1 U5069 ( .A1(keyinput20), .A2(keyinput13), .A3(n4565), .A4(n4564), 
        .ZN(n4579) );
  NAND4_X1 U5070 ( .A1(keyinput52), .A2(keyinput22), .A3(keyinput50), .A4(
        keyinput37), .ZN(n4578) );
  NOR2_X1 U5071 ( .A1(keyinput63), .A2(keyinput60), .ZN(n4569) );
  NAND3_X1 U5072 ( .A1(keyinput43), .A2(keyinput30), .A3(keyinput23), .ZN(
        n4567) );
  NAND3_X1 U5073 ( .A1(keyinput28), .A2(keyinput11), .A3(keyinput46), .ZN(
        n4566) );
  NOR4_X1 U5074 ( .A1(keyinput19), .A2(keyinput24), .A3(n4567), .A4(n4566), 
        .ZN(n4568) );
  NAND4_X1 U5075 ( .A1(keyinput32), .A2(keyinput25), .A3(n4569), .A4(n4568), 
        .ZN(n4577) );
  NOR3_X1 U5076 ( .A1(keyinput31), .A2(keyinput7), .A3(keyinput2), .ZN(n4575)
         );
  NAND2_X1 U5077 ( .A1(keyinput54), .A2(keyinput10), .ZN(n4570) );
  NOR3_X1 U5078 ( .A1(keyinput15), .A2(keyinput47), .A3(n4570), .ZN(n4574) );
  NAND4_X1 U5079 ( .A1(keyinput56), .A2(keyinput8), .A3(keyinput57), .A4(
        keyinput61), .ZN(n4572) );
  NAND2_X1 U5080 ( .A1(keyinput41), .A2(keyinput45), .ZN(n4571) );
  NOR4_X1 U5081 ( .A1(keyinput21), .A2(keyinput33), .A3(n4572), .A4(n4571), 
        .ZN(n4573) );
  NAND4_X1 U5082 ( .A1(keyinput6), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(
        n4576) );
  NOR4_X1 U5083 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4580)
         );
  AOI21_X1 U5084 ( .B1(n4581), .B2(n4580), .A(keyinput35), .ZN(n4611) );
  AOI22_X1 U5085 ( .A1(n4584), .A2(keyinput45), .B1(n4583), .B2(keyinput33), 
        .ZN(n4582) );
  OAI221_X1 U5086 ( .B1(n4584), .B2(keyinput45), .C1(n4583), .C2(keyinput33), 
        .A(n4582), .ZN(n4594) );
  INV_X1 U5087 ( .A(DATAI_2_), .ZN(n4586) );
  AOI22_X1 U5088 ( .A1(n4587), .A2(keyinput13), .B1(keyinput21), .B2(n4586), 
        .ZN(n4585) );
  OAI221_X1 U5089 ( .B1(n4587), .B2(keyinput13), .C1(n4586), .C2(keyinput21), 
        .A(n4585), .ZN(n4593) );
  AOI22_X1 U5090 ( .A1(n2429), .A2(keyinput8), .B1(n2243), .B2(keyinput57), 
        .ZN(n4588) );
  OAI221_X1 U5091 ( .B1(n2429), .B2(keyinput8), .C1(n2243), .C2(keyinput57), 
        .A(n4588), .ZN(n4592) );
  XNOR2_X1 U5092 ( .A(IR_REG_14__SCAN_IN), .B(keyinput41), .ZN(n4590) );
  XNOR2_X1 U5093 ( .A(IR_REG_4__SCAN_IN), .B(keyinput61), .ZN(n4589) );
  NAND2_X1 U5094 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  NOR4_X1 U5095 ( .A1(n4594), .A2(n4593), .A3(n4592), .A4(n4591), .ZN(n4610)
         );
  AOI22_X1 U5096 ( .A1(n2281), .A2(keyinput2), .B1(keyinput15), .B2(n4596), 
        .ZN(n4595) );
  OAI221_X1 U5097 ( .B1(n2281), .B2(keyinput2), .C1(n4596), .C2(keyinput15), 
        .A(n4595), .ZN(n4608) );
  AOI22_X1 U5098 ( .A1(n2505), .A2(keyinput6), .B1(n4598), .B2(keyinput7), 
        .ZN(n4597) );
  OAI221_X1 U5099 ( .B1(n2505), .B2(keyinput6), .C1(n4598), .C2(keyinput7), 
        .A(n4597), .ZN(n4607) );
  INV_X1 U5100 ( .A(DATAI_7_), .ZN(n4601) );
  AOI22_X1 U5101 ( .A1(n4601), .A2(keyinput47), .B1(keyinput56), .B2(n4600), 
        .ZN(n4599) );
  OAI221_X1 U5102 ( .B1(n4601), .B2(keyinput47), .C1(n4600), .C2(keyinput56), 
        .A(n4599), .ZN(n4606) );
  AOI22_X1 U5103 ( .A1(n4604), .A2(keyinput10), .B1(keyinput54), .B2(n4603), 
        .ZN(n4602) );
  OAI221_X1 U5104 ( .B1(n4604), .B2(keyinput10), .C1(n4603), .C2(keyinput54), 
        .A(n4602), .ZN(n4605) );
  NOR4_X1 U5105 ( .A1(n4608), .A2(n4607), .A3(n4606), .A4(n4605), .ZN(n4609)
         );
  OAI211_X1 U5106 ( .C1(ADDR_REG_5__SCAN_IN), .C2(n4611), .A(n4610), .B(n4609), 
        .ZN(n4612) );
  NOR4_X1 U5107 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4616)
         );
  NAND4_X1 U5108 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4620)
         );
  XNOR2_X1 U5109 ( .A(n4621), .B(n4620), .ZN(U3250) );
  INV_X2 U2265 ( .A(IR_REG_31__SCAN_IN), .ZN(n2641) );
  NOR2_X1 U2821 ( .A1(n2282), .A2(n2092), .ZN(n4275) );
  CLKBUF_X1 U2268 ( .A(n2318), .Z(n2918) );
  CLKBUF_X1 U2277 ( .A(n2682), .Z(n2892) );
  INV_X1 U2299 ( .A(n2302), .ZN(n2908) );
endmodule

