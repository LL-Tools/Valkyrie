

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2002, n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741;

  INV_X1 U2244 ( .A(n3267), .ZN(n4576) );
  INV_X1 U2245 ( .A(n3061), .ZN(n3723) );
  CLKBUF_X2 U2246 ( .A(n2416), .Z(n2805) );
  INV_X1 U2248 ( .A(n2858), .ZN(n2794) );
  INV_X1 U2249 ( .A(n3717), .ZN(n3061) );
  NAND2_X1 U2250 ( .A1(n2997), .A2(n2339), .ZN(n2416) );
  CLKBUF_X3 U2251 ( .A(n2355), .Z(n2002) );
  NAND2_X1 U2252 ( .A1(n2367), .A2(n2839), .ZN(n2364) );
  INV_X1 U2253 ( .A(n2784), .ZN(n2355) );
  NAND2_X2 U2254 ( .A1(n3028), .A2(IR_REG_31__SCAN_IN), .ZN(n2346) );
  XNOR2_X2 U2255 ( .A(n2361), .B(IR_REG_22__SCAN_IN), .ZN(n2838) );
  OAI21_X1 U2256 ( .B1(n3717), .B2(n2375), .A(n2374), .ZN(n3267) );
  OAI21_X1 U2257 ( .B1(n3717), .B2(n3079), .A(n2338), .ZN(n3270) );
  NAND2_X4 U2258 ( .A1(n2337), .A2(n2336), .ZN(n3717) );
  AOI21_X1 U2259 ( .B1(n3643), .B2(n3646), .A(n3644), .ZN(n3544) );
  AOI21_X1 U2260 ( .B1(n2985), .B2(n4270), .A(n2984), .ZN(n3551) );
  NAND2_X1 U2261 ( .A1(n2120), .A2(n2125), .ZN(n4158) );
  NAND2_X1 U2262 ( .A1(n3442), .A2(n2291), .ZN(n3443) );
  INV_X2 U2263 ( .A(n4535), .ZN(n2003) );
  NAND2_X1 U2264 ( .A1(n2187), .A2(n2014), .ZN(n3442) );
  AOI21_X1 U2265 ( .B1(n2500), .B2(n2113), .A(n2112), .ZN(n2064) );
  AOI22_X1 U2266 ( .A1(n3151), .A2(REG2_REG_6__SCAN_IN), .B1(n4463), .B2(n3150), .ZN(n3153) );
  AND2_X1 U2267 ( .A1(n3796), .A2(n3799), .ZN(n3775) );
  AND2_X1 U2268 ( .A1(n3809), .A2(n3806), .ZN(n3764) );
  INV_X1 U2269 ( .A(n2949), .ZN(n3882) );
  INV_X1 U2270 ( .A(n2896), .ZN(n3883) );
  INV_X4 U2271 ( .A(n2398), .ZN(n2792) );
  AND2_X2 U2272 ( .A1(n2856), .A2(n2364), .ZN(n2398) );
  XNOR2_X1 U2273 ( .A(n3073), .B(n3072), .ZN(n3111) );
  AND3_X1 U2274 ( .A1(n2353), .A2(n2352), .A3(n2351), .ZN(n2357) );
  AOI21_X1 U2275 ( .B1(REG1_REG_3__SCAN_IN), .B2(n3093), .A(n3071), .ZN(n3073)
         );
  XNOR2_X1 U2276 ( .A(n2348), .B(n2347), .ZN(n2354) );
  XNOR2_X1 U2277 ( .A(n2321), .B(IR_REG_26__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U2278 ( .A1(n2861), .A2(IR_REG_31__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U2279 ( .A1(n2083), .A2(n2195), .ZN(n3079) );
  INV_X1 U2280 ( .A(n2409), .ZN(n2083) );
  AND2_X1 U2281 ( .A1(n2063), .A2(n2062), .ZN(n2409) );
  INV_X1 U2282 ( .A(IR_REG_14__SCAN_IN), .ZN(n2601) );
  NOR2_X1 U2283 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2306)
         );
  INV_X1 U2284 ( .A(IR_REG_15__SCAN_IN), .ZN(n2614) );
  INV_X1 U2285 ( .A(IR_REG_16__SCAN_IN), .ZN(n2632) );
  NOR2_X1 U2286 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2313)
         );
  NOR2_X1 U2287 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2314)
         );
  NOR2_X1 U2288 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2315)
         );
  NOR2_X1 U2289 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2303)
         );
  NOR2_X1 U2290 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2316)
         );
  NOR2_X1 U2291 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2302)
         );
  NOR2_X1 U2292 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2301)
         );
  INV_X1 U2293 ( .A(IR_REG_13__SCAN_IN), .ZN(n2585) );
  INV_X1 U2294 ( .A(IR_REG_25__SCAN_IN), .ZN(n2341) );
  OAI211_X1 U2295 ( .C1(n3443), .C2(n2175), .A(n2174), .B(1'b1), .ZN(n3911) );
  AOI21_X1 U2297 ( .B1(n3539), .B2(n3538), .A(n3537), .ZN(n3644) );
  INV_X4 U2298 ( .A(n2390), .ZN(n2349) );
  INV_X2 U2299 ( .A(n2442), .ZN(n3719) );
  INV_X1 U2300 ( .A(n2364), .ZN(n2110) );
  INV_X1 U2301 ( .A(IR_REG_24__SCAN_IN), .ZN(n2814) );
  INV_X1 U2302 ( .A(n2939), .ZN(n2257) );
  AND2_X1 U2303 ( .A1(n3847), .A2(n2972), .ZN(n3740) );
  NAND2_X1 U2304 ( .A1(n4522), .A2(n3270), .ZN(n3799) );
  OR2_X1 U2305 ( .A1(n3255), .A2(n3254), .ZN(n2284) );
  NOR2_X1 U2306 ( .A1(n3667), .A2(n2287), .ZN(n2286) );
  INV_X1 U2307 ( .A(n3587), .ZN(n2287) );
  NAND2_X1 U2308 ( .A1(n2080), .A2(n2024), .ZN(n3070) );
  INV_X1 U2309 ( .A(n3388), .ZN(n2904) );
  NAND2_X1 U2310 ( .A1(n3369), .A2(n3388), .ZN(n3817) );
  INV_X1 U2311 ( .A(n3659), .ZN(n2994) );
  AND2_X1 U2312 ( .A1(n2308), .A2(n2309), .ZN(n2118) );
  OAI22_X1 U2313 ( .A1(n2807), .A2(n2886), .B1(n2887), .B2(n2433), .ZN(n2432)
         );
  NAND2_X1 U2314 ( .A1(n2288), .A2(n2286), .ZN(n3664) );
  OR2_X1 U2315 ( .A1(n3039), .A2(IR_REG_28__SCAN_IN), .ZN(n2337) );
  AOI21_X1 U2316 ( .B1(n3039), .B2(IR_REG_27__SCAN_IN), .A(n2292), .ZN(n2336)
         );
  AND2_X1 U2317 ( .A1(n4454), .A2(n2324), .ZN(n2325) );
  AND2_X1 U2318 ( .A1(n3000), .A2(n2834), .ZN(n2868) );
  INV_X1 U2319 ( .A(n2050), .ZN(n2609) );
  INV_X1 U2321 ( .A(n2410), .ZN(n2442) );
  NOR2_X1 U2322 ( .A1(n3104), .A2(n2185), .ZN(n2184) );
  NAND2_X1 U2323 ( .A1(n2181), .A2(n2180), .ZN(n2179) );
  INV_X1 U2324 ( .A(n3104), .ZN(n2180) );
  INV_X1 U2325 ( .A(n2186), .ZN(n2181) );
  NAND2_X1 U2326 ( .A1(n3911), .A2(n3910), .ZN(n3922) );
  NAND2_X1 U2327 ( .A1(n3950), .A2(n2221), .ZN(n2069) );
  NOR2_X1 U2328 ( .A1(n3967), .A2(n2222), .ZN(n2221) );
  NAND2_X1 U2329 ( .A1(n2220), .A2(n2219), .ZN(n2068) );
  INV_X1 U2330 ( .A(n3967), .ZN(n2219) );
  INV_X1 U2331 ( .A(n3965), .ZN(n2220) );
  NAND2_X1 U2332 ( .A1(n4487), .A2(n4488), .ZN(n4486) );
  OR2_X1 U2333 ( .A1(n2797), .A2(n2848), .ZN(n4025) );
  OR2_X1 U2334 ( .A1(n2770), .A2(n2769), .ZN(n2782) );
  NAND2_X1 U2335 ( .A1(n2051), .A2(REG3_REG_21__SCAN_IN), .ZN(n2726) );
  INV_X1 U2336 ( .A(n2933), .ZN(n2246) );
  AOI21_X1 U2337 ( .B1(n2255), .B2(n2253), .A(n2026), .ZN(n2252) );
  NAND2_X1 U2338 ( .A1(n2938), .A2(n2254), .ZN(n2251) );
  OR2_X1 U2339 ( .A1(n2866), .A2(n2838), .ZN(n4551) );
  NAND2_X1 U2340 ( .A1(n2366), .A2(n3761), .ZN(n2837) );
  INV_X1 U2341 ( .A(IR_REG_19__SCAN_IN), .ZN(n2363) );
  NOR2_X1 U2342 ( .A1(n3846), .A2(n2158), .ZN(n2157) );
  AND2_X1 U2343 ( .A1(n3873), .A2(n4069), .ZN(n3725) );
  INV_X1 U2344 ( .A(n2157), .ZN(n2155) );
  INV_X1 U2345 ( .A(n3600), .ZN(n2275) );
  INV_X1 U2346 ( .A(n4216), .ZN(n2967) );
  OR2_X1 U2347 ( .A1(n3481), .A2(n3482), .ZN(n2280) );
  NAND2_X1 U2348 ( .A1(n2349), .A2(REG2_REG_2__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U2349 ( .A1(n2214), .A2(n2212), .ZN(n3930) );
  INV_X1 U2350 ( .A(n2213), .ZN(n2212) );
  OAI21_X1 U2351 ( .B1(n3452), .B2(n2040), .A(n3913), .ZN(n2213) );
  AND2_X1 U2352 ( .A1(n2160), .A2(n3850), .ZN(n2159) );
  NOR2_X1 U2353 ( .A1(n2123), .A2(n2122), .ZN(n2121) );
  OR2_X1 U2354 ( .A1(n4236), .A2(n2124), .ZN(n2119) );
  AOI21_X1 U2355 ( .B1(n3837), .B2(n3736), .A(n2126), .ZN(n2125) );
  INV_X1 U2356 ( .A(n3737), .ZN(n2126) );
  INV_X1 U2357 ( .A(n2923), .ZN(n2099) );
  INV_X1 U2358 ( .A(n2229), .ZN(n2228) );
  OAI21_X1 U2359 ( .B1(n4251), .B2(n2230), .A(n2926), .ZN(n2229) );
  INV_X1 U2360 ( .A(n2925), .ZN(n2230) );
  NOR2_X1 U2361 ( .A1(n2577), .A2(n2576), .ZN(n2050) );
  INV_X1 U2362 ( .A(n4293), .ZN(n2917) );
  INV_X1 U2363 ( .A(n4290), .ZN(n2918) );
  INV_X1 U2364 ( .A(n2132), .ZN(n2131) );
  OAI21_X1 U2365 ( .B1(n2134), .B2(n2133), .A(n3826), .ZN(n2132) );
  INV_X1 U2366 ( .A(n3821), .ZN(n2133) );
  INV_X1 U2367 ( .A(n3879), .ZN(n2955) );
  NAND2_X1 U2368 ( .A1(n2145), .A2(n3809), .ZN(n2142) );
  AND2_X1 U2369 ( .A1(n3169), .A2(n3213), .ZN(n2897) );
  AND2_X1 U2370 ( .A1(n2892), .A2(n2891), .ZN(n2226) );
  NAND2_X1 U2371 ( .A1(n3213), .A2(n2890), .ZN(n2891) );
  NAND2_X1 U2372 ( .A1(n3798), .A2(n3775), .ZN(n2946) );
  AND2_X1 U2373 ( .A1(n4207), .A2(n3680), .ZN(n2163) );
  INV_X1 U2374 ( .A(n4244), .ZN(n2995) );
  AND2_X1 U2375 ( .A1(n2165), .A2(n2924), .ZN(n2164) );
  INV_X1 U2376 ( .A(IR_REG_27__SCAN_IN), .ZN(n2342) );
  NAND2_X1 U2377 ( .A1(n2654), .A2(n2345), .ZN(n2861) );
  NAND2_X1 U2378 ( .A1(n2812), .A2(IR_REG_31__SCAN_IN), .ZN(n2836) );
  INV_X1 U2379 ( .A(n2811), .ZN(n2812) );
  INV_X1 U2380 ( .A(IR_REG_23__SCAN_IN), .ZN(n2835) );
  INV_X1 U2381 ( .A(IR_REG_1__SCAN_IN), .ZN(n2062) );
  INV_X1 U2382 ( .A(IR_REG_0__SCAN_IN), .ZN(n2063) );
  NAND2_X1 U2383 ( .A1(n3417), .A2(n3418), .ZN(n2269) );
  OR2_X1 U2384 ( .A1(n2477), .A2(n2476), .ZN(n2490) );
  AND2_X1 U2385 ( .A1(n2377), .A2(n2376), .ZN(n2382) );
  NAND2_X1 U2386 ( .A1(n3267), .A2(n2339), .ZN(n2376) );
  AND2_X1 U2387 ( .A1(n3481), .A2(n3482), .ZN(n2278) );
  INV_X1 U2388 ( .A(n2641), .ZN(n2268) );
  XNOR2_X1 U2389 ( .A(n2261), .B(n2398), .ZN(n2419) );
  OAI21_X1 U2390 ( .B1(n2947), .B2(n2433), .A(n2415), .ZN(n2261) );
  INV_X1 U2391 ( .A(n3398), .ZN(n2113) );
  AND2_X1 U2392 ( .A1(n2284), .A2(n3625), .ZN(n2281) );
  NAND2_X1 U2393 ( .A1(n2032), .A2(n2284), .ZN(n2282) );
  NAND2_X1 U2394 ( .A1(n3255), .A2(n3254), .ZN(n2285) );
  OAI211_X1 U2395 ( .C1(n2416), .C2(n3159), .A(n2381), .B(n2380), .ZN(n3115)
         );
  OAI22_X1 U2396 ( .A1(n2805), .A2(n3522), .B1(n3659), .B2(n2794), .ZN(n3655)
         );
  INV_X1 U2397 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U2398 ( .A1(n3005), .A2(n2060), .ZN(n2288) );
  NAND2_X1 U2399 ( .A1(n2526), .A2(REG3_REG_10__SCAN_IN), .ZN(n2543) );
  INV_X1 U2400 ( .A(n2528), .ZN(n2526) );
  AND2_X1 U2401 ( .A1(n2268), .A2(n2043), .ZN(n2265) );
  INV_X1 U2402 ( .A(n3568), .ZN(n2267) );
  INV_X1 U2403 ( .A(n2286), .ZN(n2059) );
  AND2_X1 U2404 ( .A1(n2736), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U2405 ( .A1(n2286), .A2(n2061), .ZN(n2058) );
  AND2_X1 U2406 ( .A1(n2598), .A2(n2597), .ZN(n3705) );
  NAND2_X1 U2407 ( .A1(n3719), .A2(REG0_REG_7__SCAN_IN), .ZN(n2482) );
  AND2_X1 U2408 ( .A1(n2350), .A2(n2354), .ZN(n2410) );
  NAND2_X1 U2409 ( .A1(n2082), .A2(n2081), .ZN(n2080) );
  OAI21_X1 U2410 ( .B1(n3081), .B2(n3082), .A(n2194), .ZN(n3083) );
  XNOR2_X1 U2411 ( .A(n3070), .B(n2203), .ZN(n3093) );
  AND3_X1 U2412 ( .A1(n2182), .A2(n2179), .A3(n2035), .ZN(n3149) );
  XNOR2_X1 U2413 ( .A(n3930), .B(n3931), .ZN(n3915) );
  OAI22_X1 U2414 ( .A1(n3942), .A2(n3941), .B1(n3946), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3954) );
  NOR2_X1 U2415 ( .A1(n4508), .A2(n3986), .ZN(n2201) );
  INV_X1 U2416 ( .A(n2218), .ZN(n2078) );
  INV_X1 U2417 ( .A(n4488), .ZN(n2075) );
  NAND2_X1 U2418 ( .A1(n4475), .A2(n3977), .ZN(n4487) );
  INV_X1 U2419 ( .A(n3976), .ZN(n3975) );
  AND2_X1 U2420 ( .A1(n4025), .A2(n2798), .ZN(n3552) );
  NAND2_X1 U2421 ( .A1(n2780), .A2(REG3_REG_27__SCAN_IN), .ZN(n2797) );
  INV_X1 U2422 ( .A(n2782), .ZN(n2780) );
  INV_X1 U2423 ( .A(n2256), .ZN(n2255) );
  OAI21_X1 U2424 ( .B1(n2259), .B2(n2005), .A(n2941), .ZN(n2256) );
  NAND2_X1 U2425 ( .A1(n2725), .A2(n2724), .ZN(n2740) );
  INV_X1 U2426 ( .A(n2726), .ZN(n2725) );
  NAND2_X1 U2427 ( .A1(n2739), .A2(REG3_REG_24__SCAN_IN), .ZN(n2770) );
  INV_X1 U2428 ( .A(n2740), .ZN(n2739) );
  INV_X1 U2429 ( .A(n2105), .ZN(n2104) );
  OAI21_X1 U2430 ( .B1(n2107), .B2(n2106), .A(n2936), .ZN(n2105) );
  AOI21_X1 U2431 ( .B1(n2241), .B2(n2240), .A(n2031), .ZN(n2239) );
  INV_X1 U2432 ( .A(n2245), .ZN(n2240) );
  NOR2_X1 U2433 ( .A1(n2242), .A2(n2108), .ZN(n2107) );
  INV_X1 U2434 ( .A(n2931), .ZN(n2108) );
  AOI21_X1 U2435 ( .B1(n2245), .B2(n2934), .A(n2028), .ZN(n2244) );
  INV_X1 U2436 ( .A(n4171), .ZN(n2249) );
  NAND2_X1 U2437 ( .A1(n2676), .A2(REG3_REG_19__SCAN_IN), .ZN(n2690) );
  INV_X1 U2438 ( .A(n2676), .ZN(n2678) );
  AND2_X1 U2439 ( .A1(n2630), .A2(n2629), .ZN(n4237) );
  NAND2_X1 U2440 ( .A1(n2622), .A2(REG3_REG_16__SCAN_IN), .ZN(n2664) );
  INV_X1 U2441 ( .A(n2624), .ZN(n2622) );
  AND2_X1 U2442 ( .A1(n3572), .A2(n4277), .ZN(n2165) );
  NAND2_X1 U2443 ( .A1(n3521), .A2(n3759), .ZN(n2153) );
  INV_X1 U2444 ( .A(n2235), .ZN(n2233) );
  INV_X1 U2445 ( .A(n3878), .ZN(n3469) );
  NAND2_X1 U2446 ( .A1(n2048), .A2(REG3_REG_9__SCAN_IN), .ZN(n2528) );
  INV_X1 U2447 ( .A(n2508), .ZN(n2048) );
  OAI21_X1 U2448 ( .B1(n3363), .B2(n2952), .A(n3817), .ZN(n3298) );
  AOI21_X1 U2449 ( .B1(n3378), .B2(n2906), .A(n2905), .ZN(n2907) );
  NOR2_X1 U2450 ( .A1(n2904), .A2(n3369), .ZN(n2905) );
  MUX2_X1 U2451 ( .A(n2441), .B(n3107), .S(n3061), .Z(n3312) );
  NAND2_X1 U2452 ( .A1(n3061), .A2(n3114), .ZN(n2053) );
  INV_X1 U2453 ( .A(n3194), .ZN(n3289) );
  AND2_X1 U2454 ( .A1(n3063), .A2(n3119), .ZN(n4272) );
  AND2_X1 U2455 ( .A1(n3063), .A2(n3087), .ZN(n4273) );
  AND2_X1 U2456 ( .A1(n3267), .A2(n2893), .ZN(n3269) );
  NAND2_X1 U2457 ( .A1(n2979), .A2(n3750), .ZN(n4270) );
  OAI21_X1 U2458 ( .B1(n4044), .B2(n2944), .A(n2943), .ZN(n4012) );
  NOR2_X2 U2459 ( .A1(n4184), .A2(n4163), .ZN(n4164) );
  INV_X1 U2460 ( .A(n3580), .ZN(n4207) );
  OR2_X1 U2461 ( .A1(n3474), .A2(n3603), .ZN(n3513) );
  NAND3_X1 U2462 ( .A1(n4454), .A2(n2818), .A3(n2817), .ZN(n3053) );
  AND2_X1 U2463 ( .A1(n2341), .A2(n2319), .ZN(n2320) );
  NOR2_X1 U2464 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2310)
         );
  INV_X1 U2465 ( .A(IR_REG_20__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2466 ( .A1(n2329), .A2(IR_REG_31__SCAN_IN), .ZN(n2331) );
  AND2_X1 U2467 ( .A1(n2603), .A2(n2613), .ZN(n3963) );
  NAND2_X1 U2468 ( .A1(n3717), .A2(DATAI_1_), .ZN(n2338) );
  AND2_X1 U2469 ( .A1(n2726), .A2(n2708), .ZN(n4166) );
  AND2_X1 U2470 ( .A1(n2776), .A2(n2775), .ZN(n4087) );
  AND2_X1 U2471 ( .A1(n2867), .A2(n4255), .ZN(n3703) );
  NAND2_X1 U2472 ( .A1(n2868), .A2(n2841), .ZN(n3711) );
  INV_X1 U2473 ( .A(n4041), .ZN(n4014) );
  NAND2_X1 U2474 ( .A1(n2696), .A2(n2695), .ZN(n4204) );
  INV_X1 U2475 ( .A(n4237), .ZN(n4274) );
  INV_X1 U2476 ( .A(n3705), .ZN(n4271) );
  NAND2_X1 U2477 ( .A1(n3886), .A2(n3887), .ZN(n3895) );
  XNOR2_X1 U2478 ( .A(n3443), .B(n3462), .ZN(n3457) );
  NAND2_X1 U2479 ( .A1(n2011), .A2(n2038), .ZN(n2174) );
  NOR2_X1 U2480 ( .A1(n2011), .A2(n3462), .ZN(n2175) );
  XNOR2_X1 U2481 ( .A(n3922), .B(n3912), .ZN(n3925) );
  NAND2_X1 U2482 ( .A1(n3950), .A2(REG1_REG_14__SCAN_IN), .ZN(n3966) );
  AND2_X1 U2483 ( .A1(n4489), .A2(n2201), .ZN(n4506) );
  NAND2_X1 U2484 ( .A1(n4489), .A2(n3987), .ZN(n4507) );
  AOI21_X1 U2485 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n4505) );
  NAND2_X1 U2486 ( .A1(n4486), .A2(n2218), .ZN(n4499) );
  OR2_X1 U2487 ( .A1(n4469), .A2(n3119), .ZN(n4514) );
  OAI21_X1 U2488 ( .B1(n4490), .B2(n2200), .A(n2198), .ZN(n2202) );
  INV_X1 U2489 ( .A(n3939), .ZN(n4510) );
  NAND2_X1 U2490 ( .A1(n4030), .A2(n4029), .ZN(n4317) );
  XNOR2_X1 U2491 ( .A(n3872), .B(n4026), .ZN(n4318) );
  AND2_X1 U2492 ( .A1(n2088), .A2(n2092), .ZN(n2087) );
  INV_X1 U2493 ( .A(n2085), .ZN(n2084) );
  OAI21_X1 U2494 ( .B1(n3551), .B2(n4587), .A(n2095), .ZN(n2085) );
  NAND2_X1 U2495 ( .A1(n4587), .A2(REG1_REG_28__SCAN_IN), .ZN(n2095) );
  NAND2_X1 U2496 ( .A1(n4589), .A2(n4570), .ZN(n2086) );
  NAND2_X1 U2497 ( .A1(n3909), .A2(REG1_REG_11__SCAN_IN), .ZN(n3913) );
  NOR2_X1 U2498 ( .A1(n2216), .A2(n4672), .ZN(n2215) );
  INV_X1 U2499 ( .A(n2125), .ZN(n2124) );
  NOR2_X1 U2500 ( .A1(n2124), .A2(n3837), .ZN(n2123) );
  INV_X1 U2501 ( .A(n3843), .ZN(n2122) );
  NAND2_X1 U2502 ( .A1(n2894), .A2(n2993), .ZN(n3796) );
  INV_X1 U2503 ( .A(n2898), .ZN(n2887) );
  NOR2_X1 U2504 ( .A1(n3599), .A2(n2278), .ZN(n2277) );
  NOR2_X1 U2505 ( .A1(n3566), .A2(n3568), .ZN(n3610) );
  INV_X1 U2506 ( .A(n2805), .ZN(n2796) );
  NAND3_X1 U2507 ( .A1(n2069), .A2(n2044), .A3(n2068), .ZN(n3976) );
  NOR2_X1 U2508 ( .A1(n2690), .A2(n3011), .ZN(n2051) );
  NOR2_X1 U2509 ( .A1(n2664), .A2(n2663), .ZN(n2676) );
  INV_X1 U2510 ( .A(n2921), .ZN(n2232) );
  NAND2_X1 U2511 ( .A1(n2919), .A2(n2006), .ZN(n2235) );
  NAND2_X1 U2512 ( .A1(n2236), .A2(n2006), .ZN(n2234) );
  NOR2_X1 U2513 ( .A1(n2543), .A2(n2542), .ZN(n2559) );
  AND2_X1 U2514 ( .A1(n3816), .A2(n2135), .ZN(n2134) );
  AND2_X1 U2515 ( .A1(n3378), .A2(n2295), .ZN(n2903) );
  AND2_X1 U2516 ( .A1(n3881), .A2(n3258), .ZN(n2906) );
  NOR2_X1 U2517 ( .A1(n3309), .A2(n2144), .ZN(n2143) );
  INV_X1 U2518 ( .A(n3809), .ZN(n2144) );
  AND2_X1 U2519 ( .A1(n2899), .A2(n2895), .ZN(n2109) );
  INV_X1 U2520 ( .A(n3806), .ZN(n2145) );
  INV_X1 U2521 ( .A(n2943), .ZN(n2093) );
  AND2_X1 U2522 ( .A1(n2255), .A2(n2020), .ZN(n2254) );
  AND2_X1 U2523 ( .A1(n2005), .A2(n2020), .ZN(n2253) );
  OAI21_X1 U2524 ( .B1(n2156), .B2(n4098), .A(n2154), .ZN(n4017) );
  INV_X1 U2525 ( .A(n2159), .ZN(n2156) );
  AOI21_X1 U2526 ( .B1(n2159), .B2(n2155), .A(n2030), .ZN(n2154) );
  NOR2_X1 U2527 ( .A1(n4050), .A2(n4013), .ZN(n3998) );
  NOR2_X1 U2528 ( .A1(n4130), .A2(n4144), .ZN(n2171) );
  AND2_X1 U2529 ( .A1(n2320), .A2(n2335), .ZN(n2238) );
  OR2_X1 U2530 ( .A1(n2654), .A2(n2327), .ZN(n2115) );
  INV_X1 U2531 ( .A(n2117), .ZN(n2116) );
  OAI21_X1 U2532 ( .B1(n2327), .B2(n2118), .A(n2363), .ZN(n2117) );
  INV_X1 U2533 ( .A(IR_REG_17__SCAN_IN), .ZN(n2308) );
  INV_X1 U2534 ( .A(IR_REG_7__SCAN_IN), .ZN(n2472) );
  INV_X1 U2535 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2476) );
  INV_X1 U2536 ( .A(n2976), .ZN(n4048) );
  NOR2_X1 U2537 ( .A1(n2272), .A2(n2275), .ZN(n2271) );
  INV_X1 U2538 ( .A(n2280), .ZN(n2272) );
  INV_X1 U2539 ( .A(n2274), .ZN(n2273) );
  OAI21_X1 U2540 ( .B1(n2277), .B2(n2275), .A(n3654), .ZN(n2274) );
  AND2_X1 U2541 ( .A1(n2637), .A2(n2638), .ZN(n3568) );
  NOR2_X1 U2542 ( .A1(n3237), .A2(n2067), .ZN(n2066) );
  INV_X1 U2543 ( .A(n2421), .ZN(n2067) );
  NAND2_X1 U2544 ( .A1(n2279), .A2(n2277), .ZN(n2114) );
  INV_X1 U2545 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2542) );
  AND2_X1 U2546 ( .A1(n2759), .A2(n3540), .ZN(n2760) );
  AND4_X1 U2547 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n2949)
         );
  AND4_X1 U2548 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n2947)
         );
  NAND2_X1 U2549 ( .A1(n2002), .A2(REG3_REG_2__SCAN_IN), .ZN(n2395) );
  OR2_X1 U2550 ( .A1(n2443), .A2(n3069), .ZN(n2352) );
  AND2_X1 U2551 ( .A1(n3070), .A2(n4464), .ZN(n3071) );
  AOI22_X1 U2552 ( .A1(n3094), .A2(REG2_REG_3__SCAN_IN), .B1(n4464), .B2(n3084), .ZN(n3085) );
  NAND2_X1 U2553 ( .A1(n3111), .A2(n2209), .ZN(n2207) );
  NOR2_X1 U2554 ( .A1(n3101), .A2(n2210), .ZN(n2209) );
  NAND2_X1 U2555 ( .A1(n2206), .A2(n2205), .ZN(n2204) );
  INV_X1 U2556 ( .A(n3101), .ZN(n2205) );
  INV_X1 U2557 ( .A(n2211), .ZN(n2206) );
  AOI22_X1 U2558 ( .A1(n3204), .A2(n3203), .B1(n4669), .B2(n3202), .ZN(n3326)
         );
  NAND2_X1 U2559 ( .A1(n3329), .A2(n3328), .ZN(n3331) );
  NAND2_X1 U2560 ( .A1(n3326), .A2(n4461), .ZN(n3328) );
  XNOR2_X1 U2561 ( .A(n3451), .B(n3462), .ZN(n3459) );
  INV_X1 U2562 ( .A(IR_REG_11__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U2563 ( .A1(n3459), .A2(REG1_REG_10__SCAN_IN), .ZN(n3458) );
  NAND2_X1 U2564 ( .A1(n3915), .A2(REG1_REG_12__SCAN_IN), .ZN(n3933) );
  NAND2_X1 U2565 ( .A1(n3957), .A2(n3956), .ZN(n3959) );
  XNOR2_X1 U2566 ( .A(n3976), .B(n4543), .ZN(n4477) );
  NAND2_X1 U2567 ( .A1(n2173), .A2(n2172), .ZN(n3983) );
  NAND2_X1 U2568 ( .A1(n3961), .A2(n2289), .ZN(n2172) );
  NAND2_X1 U2569 ( .A1(n3957), .A2(n2021), .ZN(n2173) );
  NAND2_X1 U2570 ( .A1(n4542), .A2(n4367), .ZN(n2218) );
  AOI21_X1 U2571 ( .B1(n2201), .B2(n2199), .A(n2045), .ZN(n2198) );
  INV_X1 U2572 ( .A(n4491), .ZN(n2199) );
  INV_X1 U2573 ( .A(n2201), .ZN(n2200) );
  NAND2_X1 U2574 ( .A1(n2161), .A2(n2159), .ZN(n4038) );
  NAND2_X1 U2575 ( .A1(n3850), .A2(n2161), .ZN(n4036) );
  AND2_X1 U2576 ( .A1(n2804), .A2(n2803), .ZN(n4041) );
  NAND2_X1 U2577 ( .A1(n4236), .A2(n3837), .ZN(n2120) );
  INV_X1 U2578 ( .A(n2051), .ZN(n2707) );
  OR2_X1 U2579 ( .A1(n4236), .A2(n3736), .ZN(n4174) );
  AND2_X1 U2580 ( .A1(n2098), .A2(n2227), .ZN(n2097) );
  AOI21_X1 U2581 ( .B1(n2228), .B2(n2230), .A(n2039), .ZN(n2227) );
  NAND2_X1 U2582 ( .A1(n2100), .A2(n2099), .ZN(n2098) );
  AND2_X1 U2583 ( .A1(n4197), .A2(n4198), .ZN(n4223) );
  NAND2_X1 U2584 ( .A1(n2050), .A2(n2037), .ZN(n2624) );
  AOI21_X1 U2585 ( .B1(n2151), .B2(n2150), .A(n2149), .ZN(n2148) );
  INV_X1 U2586 ( .A(n3727), .ZN(n2149) );
  AND2_X1 U2587 ( .A1(n2653), .A2(n2652), .ZN(n4265) );
  AND2_X1 U2588 ( .A1(n2102), .A2(n2019), .ZN(n4252) );
  NAND2_X1 U2589 ( .A1(n4268), .A2(n2923), .ZN(n2102) );
  NAND2_X1 U2590 ( .A1(n4252), .A2(n4251), .ZN(n4250) );
  NAND2_X1 U2591 ( .A1(n2559), .A2(REG3_REG_12__SCAN_IN), .ZN(n2577) );
  INV_X1 U2592 ( .A(n2559), .ZN(n2561) );
  AND3_X1 U2593 ( .A1(n2581), .A2(n2580), .A3(n2579), .ZN(n3522) );
  AND2_X1 U2594 ( .A1(n3467), .A2(n3466), .ZN(n4293) );
  NAND2_X1 U2595 ( .A1(n2129), .A2(n2127), .ZN(n4287) );
  AOI21_X1 U2596 ( .B1(n2131), .B2(n2133), .A(n2128), .ZN(n2127) );
  INV_X1 U2597 ( .A(n3823), .ZN(n2128) );
  NAND2_X1 U2598 ( .A1(n2130), .A2(n3821), .ZN(n3407) );
  NAND2_X1 U2599 ( .A1(n2954), .A2(n2134), .ZN(n2130) );
  INV_X1 U2600 ( .A(n4272), .ZN(n4288) );
  NAND2_X1 U2601 ( .A1(n2954), .A2(n3816), .ZN(n3353) );
  NAND2_X1 U2602 ( .A1(n2049), .A2(REG3_REG_8__SCAN_IN), .ZN(n2508) );
  INV_X1 U2603 ( .A(n2490), .ZN(n2049) );
  NAND2_X1 U2604 ( .A1(n3817), .A2(n2951), .ZN(n3378) );
  NAND2_X1 U2605 ( .A1(n2146), .A2(n3814), .ZN(n3363) );
  OAI21_X1 U2606 ( .B1(n3223), .B2(n2141), .A(n2136), .ZN(n2146) );
  AOI21_X1 U2607 ( .B1(n2140), .B2(n2138), .A(n2137), .ZN(n2136) );
  INV_X1 U2608 ( .A(n2143), .ZN(n2138) );
  NAND2_X1 U2609 ( .A1(n2458), .A2(REG3_REG_6__SCAN_IN), .ZN(n2477) );
  INV_X1 U2610 ( .A(n2460), .ZN(n2458) );
  NAND2_X1 U2611 ( .A1(n2139), .A2(n2140), .ZN(n3184) );
  NAND2_X1 U2612 ( .A1(n3223), .A2(n2143), .ZN(n2139) );
  NAND2_X1 U2613 ( .A1(n2445), .A2(REG3_REG_5__SCAN_IN), .ZN(n2460) );
  INV_X1 U2614 ( .A(n2447), .ZN(n2445) );
  NAND2_X1 U2615 ( .A1(n2898), .A2(n2888), .ZN(n2899) );
  OAI21_X1 U2616 ( .B1(n3223), .B2(n2145), .A(n3809), .ZN(n3310) );
  NAND2_X1 U2617 ( .A1(n2897), .A2(n3168), .ZN(n2225) );
  NAND2_X1 U2618 ( .A1(n3229), .A2(n2886), .ZN(n3316) );
  NAND2_X1 U2619 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2447) );
  NAND2_X1 U2620 ( .A1(n4525), .A2(n2888), .ZN(n3224) );
  AND2_X1 U2621 ( .A1(n3805), .A2(n3802), .ZN(n3757) );
  NAND2_X1 U2622 ( .A1(n3803), .A2(n3800), .ZN(n3169) );
  INV_X1 U2623 ( .A(n3775), .ZN(n3274) );
  INV_X1 U2624 ( .A(n4273), .ZN(n4521) );
  INV_X1 U2625 ( .A(n4270), .ZN(n4523) );
  NOR2_X1 U2626 ( .A1(n4011), .A2(n2093), .ZN(n2091) );
  NAND2_X1 U2627 ( .A1(n2091), .A2(n2944), .ZN(n2088) );
  NAND2_X1 U2628 ( .A1(n4011), .A2(n2093), .ZN(n2092) );
  NOR2_X1 U2629 ( .A1(n4030), .A2(n4005), .ZN(n4004) );
  INV_X1 U2630 ( .A(n4278), .ZN(n4525) );
  NAND2_X1 U2631 ( .A1(n4047), .A2(n4048), .ZN(n4050) );
  AND2_X1 U2632 ( .A1(n4056), .A2(n4069), .ZN(n4047) );
  NAND2_X1 U2633 ( .A1(n4164), .A2(n2010), .ZN(n4109) );
  INV_X1 U2634 ( .A(n4123), .ZN(n4130) );
  NAND2_X1 U2635 ( .A1(n4164), .A2(n2171), .ZN(n4132) );
  NAND2_X1 U2636 ( .A1(n4224), .A2(n2013), .ZN(n4184) );
  AND2_X1 U2637 ( .A1(n3514), .A2(n3572), .ZN(n4280) );
  NAND2_X1 U2638 ( .A1(n2166), .A2(n2007), .ZN(n3474) );
  NOR2_X1 U2639 ( .A1(n2168), .A2(n3368), .ZN(n4301) );
  NAND2_X1 U2640 ( .A1(n2166), .A2(n2017), .ZN(n3412) );
  NAND2_X1 U2641 ( .A1(n2166), .A2(n2953), .ZN(n3359) );
  NOR2_X1 U2642 ( .A1(n3288), .A2(n2162), .ZN(n3318) );
  AND2_X1 U2643 ( .A1(n3318), .A2(n3374), .ZN(n3370) );
  INV_X1 U2644 ( .A(n3258), .ZN(n3374) );
  AND3_X1 U2645 ( .A1(n2991), .A2(n2990), .A3(n2989), .ZN(n3001) );
  INV_X1 U2646 ( .A(IR_REG_28__SCAN_IN), .ZN(n2340) );
  XNOR2_X1 U2647 ( .A(n2815), .B(n2814), .ZN(n2819) );
  XNOR2_X1 U2648 ( .A(n2836), .B(n2835), .ZN(n3062) );
  OR3_X1 U2649 ( .A1(n2505), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2522) );
  AND2_X1 U2650 ( .A1(n2722), .A2(n2721), .ZN(n4162) );
  AOI21_X1 U2651 ( .B1(n3664), .B2(n3018), .A(n3017), .ZN(n3019) );
  INV_X1 U2652 ( .A(n2971), .ZN(n4163) );
  NAND2_X1 U2653 ( .A1(n3005), .A2(n3588), .ZN(n3593) );
  INV_X1 U2654 ( .A(n2278), .ZN(n2276) );
  INV_X1 U2655 ( .A(n3312), .ZN(n3628) );
  NAND2_X1 U2656 ( .A1(n3626), .A2(n3625), .ZN(n3624) );
  INV_X1 U2657 ( .A(n3643), .ZN(n3645) );
  NAND2_X1 U2658 ( .A1(n3192), .A2(n3193), .ZN(n2111) );
  AOI22_X1 U2659 ( .A1(n3629), .A2(n2888), .B1(n3238), .B2(n3695), .ZN(n3242)
         );
  INV_X1 U2660 ( .A(n3385), .ZN(n2112) );
  NAND2_X1 U2661 ( .A1(n3717), .A2(DATAI_0_), .ZN(n2374) );
  INV_X1 U2662 ( .A(n3703), .ZN(n3629) );
  AND2_X1 U2663 ( .A1(n2714), .A2(n2713), .ZN(n4179) );
  MUX2_X1 U2664 ( .A(n3934), .B(n2587), .S(n3717), .Z(n3659) );
  AND2_X1 U2665 ( .A1(n2732), .A2(n2731), .ZN(n4147) );
  NAND2_X1 U2666 ( .A1(n2288), .A2(n3587), .ZN(n3666) );
  OAI21_X1 U2667 ( .B1(n2266), .B2(n2263), .A(n2043), .ZN(n2262) );
  INV_X1 U2668 ( .A(n3636), .ZN(n2263) );
  NAND2_X1 U2669 ( .A1(n3624), .A2(n2457), .ZN(n3257) );
  INV_X1 U2670 ( .A(n3711), .ZN(n3623) );
  AND2_X1 U2671 ( .A1(n2868), .A2(n2863), .ZN(n3707) );
  INV_X1 U2672 ( .A(n3689), .ZN(n3708) );
  OR3_X1 U2673 ( .A1(n3752), .A2(n3751), .A3(n3750), .ZN(n3864) );
  NAND2_X1 U2674 ( .A1(n2789), .A2(n2788), .ZN(n4065) );
  INV_X1 U2675 ( .A(n4087), .ZN(n3873) );
  NAND2_X1 U2676 ( .A1(n2755), .A2(n2754), .ZN(n4066) );
  INV_X1 U2677 ( .A(n4124), .ZN(n4084) );
  INV_X1 U2678 ( .A(n4147), .ZN(n4103) );
  INV_X1 U2679 ( .A(n4162), .ZN(n3874) );
  INV_X1 U2680 ( .A(n4179), .ZN(n4143) );
  NAND2_X1 U2681 ( .A1(n2684), .A2(n2683), .ZN(n4216) );
  NAND2_X1 U2682 ( .A1(n2670), .A2(n2669), .ZN(n4239) );
  INV_X1 U2683 ( .A(n4265), .ZN(n3677) );
  INV_X1 U2684 ( .A(n3522), .ZN(n3876) );
  NAND4_X1 U2685 ( .A1(n2533), .A2(n2532), .A3(n2531), .A4(n2530), .ZN(n3485)
         );
  OR2_X1 U2686 ( .A1(n2443), .A2(n4672), .ZN(n2532) );
  NAND4_X1 U2687 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n3879)
         );
  NAND4_X1 U2688 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3388)
         );
  INV_X1 U2689 ( .A(n2947), .ZN(n3238) );
  NAND2_X1 U2690 ( .A1(n3895), .A2(n3894), .ZN(n2193) );
  XNOR2_X1 U2691 ( .A(n3085), .B(n3072), .ZN(n3112) );
  NAND2_X1 U2692 ( .A1(n2207), .A2(n2204), .ZN(n3100) );
  AND2_X1 U2693 ( .A1(n2208), .A2(n2211), .ZN(n3102) );
  NAND2_X1 U2694 ( .A1(n3111), .A2(REG1_REG_4__SCAN_IN), .ZN(n2208) );
  NAND2_X1 U2695 ( .A1(n2179), .A2(n2182), .ZN(n3103) );
  AND2_X1 U2696 ( .A1(n2183), .A2(n2186), .ZN(n3105) );
  NAND2_X1 U2697 ( .A1(n3112), .A2(REG2_REG_4__SCAN_IN), .ZN(n2183) );
  XNOR2_X1 U2698 ( .A(n3144), .B(n2073), .ZN(n3146) );
  AOI21_X1 U2699 ( .B1(n3146), .B2(REG1_REG_6__SCAN_IN), .A(n3145), .ZN(n3204)
         );
  AND2_X1 U2700 ( .A1(n3144), .A2(n4463), .ZN(n3145) );
  XNOR2_X1 U2701 ( .A(n3326), .B(n3327), .ZN(n3205) );
  NAND2_X1 U2702 ( .A1(n3205), .A2(REG1_REG_8__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U2703 ( .A1(n3323), .A2(REG2_REG_8__SCAN_IN), .ZN(n2191) );
  INV_X1 U2704 ( .A(n3322), .ZN(n2189) );
  NAND2_X1 U2705 ( .A1(n3458), .A2(n2217), .ZN(n3454) );
  NAND2_X1 U2706 ( .A1(n3451), .A2(n4459), .ZN(n2217) );
  NAND2_X1 U2707 ( .A1(n3454), .A2(n3453), .ZN(n3914) );
  NAND2_X1 U2708 ( .A1(n3443), .A2(n4459), .ZN(n2178) );
  NAND2_X1 U2709 ( .A1(n3457), .A2(REG2_REG_10__SCAN_IN), .ZN(n2176) );
  AOI21_X1 U2710 ( .B1(n3932), .B2(n4626), .A(n2072), .ZN(n2070) );
  INV_X1 U2711 ( .A(n3935), .ZN(n2072) );
  NAND2_X1 U2712 ( .A1(n3933), .A2(n3932), .ZN(n3936) );
  OAI22_X1 U2713 ( .A1(n3925), .A2(n3924), .B1(n3923), .B2(n3931), .ZN(n3942)
         );
  AND2_X1 U2714 ( .A1(n3966), .A2(n3965), .ZN(n3968) );
  NAND2_X1 U2715 ( .A1(n2069), .A2(n2068), .ZN(n3974) );
  XNOR2_X1 U2716 ( .A(n3983), .B(n2634), .ZN(n4480) );
  INV_X1 U2717 ( .A(n2079), .ZN(n3980) );
  OAI21_X1 U2718 ( .B1(n4487), .B2(n2077), .A(n2074), .ZN(n2079) );
  AOI21_X1 U2719 ( .B1(n2076), .B2(n2075), .A(n2047), .ZN(n2074) );
  AND2_X1 U2720 ( .A1(n2771), .A2(n2782), .ZN(n4073) );
  OAI21_X1 U2721 ( .B1(n2938), .B2(n2005), .A(n2255), .ZN(n4055) );
  NAND2_X1 U2722 ( .A1(n2938), .A2(n2259), .ZN(n2258) );
  NAND2_X1 U2723 ( .A1(n2932), .A2(n2107), .ZN(n2103) );
  NAND2_X1 U2724 ( .A1(n2243), .A2(n2241), .ZN(n4139) );
  NAND2_X1 U2725 ( .A1(n4171), .A2(n2245), .ZN(n2243) );
  NAND2_X1 U2726 ( .A1(n2249), .A2(n2248), .ZN(n2247) );
  NAND2_X1 U2727 ( .A1(n3514), .A2(n2165), .ZN(n4254) );
  NAND2_X1 U2728 ( .A1(n2153), .A2(n2151), .ZN(n4269) );
  NAND2_X1 U2729 ( .A1(n4291), .A2(n2919), .ZN(n3473) );
  OR2_X1 U2730 ( .A1(n4229), .A2(n2997), .ZN(n4305) );
  INV_X1 U2731 ( .A(n4530), .ZN(n4255) );
  OR2_X1 U2732 ( .A1(n2003), .A2(n3306), .ZN(n4193) );
  AND2_X1 U2733 ( .A1(n3058), .A2(n2987), .ZN(n4530) );
  INV_X1 U2734 ( .A(n4193), .ZN(n4532) );
  AOI21_X1 U2735 ( .B1(n4321), .B2(n2998), .A(n4320), .ZN(n4322) );
  OAI21_X1 U2736 ( .B1(n3558), .B2(n4577), .A(n3551), .ZN(n3002) );
  AND2_X1 U2737 ( .A1(n4224), .A2(n3680), .ZN(n4208) );
  AND2_X2 U2738 ( .A1(n3221), .A2(n3001), .ZN(n4739) );
  AND2_X1 U2739 ( .A1(n2819), .A2(n2832), .ZN(n3054) );
  INV_X1 U2740 ( .A(n2354), .ZN(n4453) );
  INV_X1 U2741 ( .A(n3087), .ZN(n3119) );
  NAND2_X1 U2742 ( .A1(n2654), .A2(n2320), .ZN(n2334) );
  AND2_X1 U2743 ( .A1(n3062), .A2(STATE_REG_SCAN_IN), .ZN(n4539) );
  NAND2_X1 U2744 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U2745 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2333) );
  OR2_X1 U2746 ( .A1(n2328), .A2(n2327), .ZN(n2362) );
  INV_X1 U2747 ( .A(IR_REG_5__SCAN_IN), .ZN(n2439) );
  OR3_X1 U2748 ( .A1(n2437), .A2(IR_REG_3__SCAN_IN), .A3(IR_REG_4__SCAN_IN), 
        .ZN(n2438) );
  INV_X1 U2749 ( .A(n2196), .ZN(n2195) );
  OAI21_X1 U2750 ( .B1(IR_REG_31__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(n2197), 
        .ZN(n2196) );
  CLKBUF_X1 U2751 ( .A(n3130), .Z(n3131) );
  AOI21_X1 U2752 ( .B1(n2018), .B2(n4505), .A(n4504), .ZN(n4512) );
  OAI21_X1 U2753 ( .B1(n3558), .B2(n2086), .A(n2084), .ZN(n3003) );
  INV_X2 U2754 ( .A(n2422), .ZN(n2339) );
  INV_X1 U2755 ( .A(n2886), .ZN(n2888) );
  NAND2_X1 U2756 ( .A1(n2053), .A2(n2052), .ZN(n2886) );
  OR2_X1 U2757 ( .A1(n2942), .A2(n2257), .ZN(n2005) );
  OR2_X1 U2758 ( .A1(n3603), .A2(n3877), .ZN(n2006) );
  INV_X1 U2759 ( .A(n3495), .ZN(n2169) );
  OAI21_X1 U2760 ( .B1(n2918), .B2(n2235), .A(n2234), .ZN(n3502) );
  INV_X1 U2761 ( .A(n3419), .ZN(n2170) );
  OAI21_X1 U2762 ( .B1(n2641), .B2(n2267), .A(n2294), .ZN(n2266) );
  INV_X1 U2763 ( .A(n3759), .ZN(n2150) );
  INV_X1 U2764 ( .A(n2934), .ZN(n2248) );
  AND2_X1 U2765 ( .A1(n2167), .A2(n4300), .ZN(n2007) );
  OAI21_X1 U2766 ( .B1(n4268), .B2(n2101), .A(n2097), .ZN(n4220) );
  NAND2_X1 U2767 ( .A1(n2918), .A2(n2917), .ZN(n4291) );
  AND2_X1 U2768 ( .A1(n2233), .A2(n2921), .ZN(n2008) );
  AND2_X1 U2769 ( .A1(n3730), .A2(n3727), .ZN(n2009) );
  INV_X1 U2770 ( .A(n3453), .ZN(n2216) );
  AND2_X1 U2771 ( .A1(n2171), .A2(n4110), .ZN(n2010) );
  OR2_X1 U2772 ( .A1(n3444), .A2(n2177), .ZN(n2011) );
  NAND2_X1 U2773 ( .A1(n2654), .A2(n2308), .ZN(n2012) );
  NAND2_X1 U2774 ( .A1(n2111), .A2(n2421), .ZN(n3234) );
  NAND2_X1 U2775 ( .A1(n2269), .A2(n2521), .ZN(n3491) );
  AND2_X1 U2776 ( .A1(n2163), .A2(n4185), .ZN(n2013) );
  NOR2_X1 U2777 ( .A1(n3325), .A2(n2188), .ZN(n2014) );
  OR2_X1 U2778 ( .A1(n3327), .A2(n2190), .ZN(n2015) );
  AND2_X1 U2779 ( .A1(n2010), .A2(n3546), .ZN(n2016) );
  XNOR2_X1 U2780 ( .A(n2331), .B(n2330), .ZN(n2367) );
  INV_X1 U2781 ( .A(IR_REG_31__SCAN_IN), .ZN(n2327) );
  INV_X1 U2782 ( .A(n2858), .ZN(n2808) );
  NAND3_X1 U2783 ( .A1(n2326), .A2(n4455), .A3(n2325), .ZN(n2378) );
  NAND4_X1 U2784 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n2898)
         );
  AND2_X1 U2785 ( .A1(n2953), .A2(n2170), .ZN(n2017) );
  NAND2_X1 U2786 ( .A1(n2888), .A2(n2887), .ZN(n3806) );
  NAND2_X1 U2787 ( .A1(n4486), .A2(n2076), .ZN(n2018) );
  NAND2_X1 U2788 ( .A1(n2247), .A2(n2933), .ZN(n4156) );
  NAND2_X1 U2789 ( .A1(n2103), .A2(n2239), .ZN(n4116) );
  OR2_X1 U2790 ( .A1(n4262), .A2(n4279), .ZN(n2019) );
  NAND4_X1 U2791 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n2893)
         );
  NAND2_X1 U2792 ( .A1(n2258), .A2(n2939), .ZN(n4078) );
  NAND2_X1 U2793 ( .A1(n4250), .A2(n2925), .ZN(n4234) );
  NAND2_X2 U2794 ( .A1(n4453), .A2(n3037), .ZN(n2784) );
  OR2_X1 U2795 ( .A1(n4087), .A2(n4069), .ZN(n2020) );
  XNOR2_X1 U2796 ( .A(n2440), .B(n2439), .ZN(n3107) );
  NAND2_X1 U2797 ( .A1(n3037), .A2(n2354), .ZN(n2390) );
  INV_X1 U2798 ( .A(n4045), .ZN(n2160) );
  AND2_X1 U2799 ( .A1(n2055), .A2(n2054), .ZN(n3577) );
  AND2_X1 U2800 ( .A1(n3956), .A2(n2289), .ZN(n2021) );
  AND2_X1 U2801 ( .A1(n2243), .A2(n2244), .ZN(n2022) );
  AND2_X1 U2802 ( .A1(n2538), .A2(n2521), .ZN(n2023) );
  INV_X1 U2803 ( .A(n2141), .ZN(n2140) );
  NAND2_X1 U2804 ( .A1(n4465), .A2(REG1_REG_2__SCAN_IN), .ZN(n2024) );
  NOR2_X1 U2805 ( .A1(n2935), .A2(n2246), .ZN(n2245) );
  AND2_X1 U2806 ( .A1(n2153), .A2(n3729), .ZN(n2025) );
  INV_X1 U2807 ( .A(n2061), .ZN(n2060) );
  NAND2_X1 U2808 ( .A1(n2036), .A2(n3588), .ZN(n2061) );
  INV_X1 U2809 ( .A(n2242), .ZN(n2241) );
  NAND2_X1 U2810 ( .A1(n2250), .A2(n2244), .ZN(n2242) );
  NOR2_X1 U2811 ( .A1(n2974), .A2(n3873), .ZN(n2026) );
  AND2_X1 U2812 ( .A1(n3959), .A2(n3958), .ZN(n2027) );
  INV_X1 U2813 ( .A(n2944), .ZN(n2096) );
  INV_X1 U2814 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2507) );
  AND2_X2 U2815 ( .A1(n2110), .A2(n2378), .ZN(n2567) );
  NOR2_X1 U2816 ( .A1(n4143), .A2(n4163), .ZN(n2028) );
  NAND2_X1 U2817 ( .A1(n2994), .A2(n3876), .ZN(n2029) );
  NAND2_X1 U2818 ( .A1(n3716), .A2(n3715), .ZN(n2030) );
  AND2_X1 U2819 ( .A1(n3874), .A2(n4144), .ZN(n2031) );
  AND2_X1 U2820 ( .A1(n4164), .A2(n2016), .ZN(n4056) );
  INV_X1 U2821 ( .A(n3079), .ZN(n3888) );
  INV_X1 U2822 ( .A(n2101), .ZN(n2100) );
  NAND2_X1 U2823 ( .A1(n2228), .A2(n2019), .ZN(n2101) );
  INV_X1 U2824 ( .A(n2919), .ZN(n2237) );
  OAI21_X1 U2825 ( .B1(n2234), .B2(n2232), .A(n2029), .ZN(n2231) );
  OAI21_X1 U2826 ( .B1(n2917), .B2(n2237), .A(n2920), .ZN(n2236) );
  NOR2_X1 U2827 ( .A1(n2360), .A2(IR_REG_22__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U2828 ( .A1(n2457), .A2(n2285), .ZN(n2032) );
  AND2_X1 U2829 ( .A1(n3600), .A2(n2590), .ZN(n2033) );
  INV_X1 U2830 ( .A(n4011), .ZN(n2094) );
  OAI21_X1 U2831 ( .B1(n2416), .B2(n4522), .A(n2368), .ZN(n2386) );
  INV_X1 U2832 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3080) );
  OR2_X1 U2833 ( .A1(n3107), .A2(n2444), .ZN(n2034) );
  INV_X1 U2834 ( .A(IR_REG_26__SCAN_IN), .ZN(n2335) );
  INV_X1 U2835 ( .A(n2152), .ZN(n2151) );
  NAND2_X1 U2836 ( .A1(n2009), .A2(n3729), .ZN(n2152) );
  OR2_X1 U2837 ( .A1(n3107), .A2(n3315), .ZN(n2035) );
  INV_X1 U2838 ( .A(IR_REG_29__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U2839 ( .A1(n4164), .A2(n4151), .ZN(n4129) );
  NOR2_X1 U2840 ( .A1(n4242), .A2(n2995), .ZN(n4224) );
  INV_X1 U2841 ( .A(n4589), .ZN(n4587) );
  AND2_X2 U2842 ( .A1(n3001), .A2(n3000), .ZN(n4589) );
  AND2_X1 U2843 ( .A1(n3268), .A2(n2895), .ZN(n3168) );
  INV_X1 U2844 ( .A(n4142), .ZN(n2250) );
  XNOR2_X1 U2845 ( .A(n2333), .B(IR_REG_21__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U2846 ( .A1(n2283), .A2(n2282), .ZN(n3397) );
  NAND2_X1 U2847 ( .A1(n2114), .A2(n3600), .ZN(n3653) );
  AOI21_X1 U2848 ( .B1(n3566), .B2(n2268), .A(n2266), .ZN(n3635) );
  NAND2_X1 U2849 ( .A1(n2264), .A2(n2262), .ZN(n3674) );
  NAND2_X1 U2850 ( .A1(n2065), .A2(n2064), .ZN(n3417) );
  NAND2_X1 U2851 ( .A1(n2279), .A2(n2276), .ZN(n3598) );
  INV_X1 U2852 ( .A(n3811), .ZN(n2137) );
  OR2_X1 U2853 ( .A1(n2717), .A2(n2716), .ZN(n2036) );
  AOI21_X1 U2854 ( .B1(n4290), .B2(n2008), .A(n2231), .ZN(n3528) );
  NAND2_X1 U2855 ( .A1(n2916), .A2(n2915), .ZN(n4290) );
  NAND2_X1 U2856 ( .A1(n3397), .A2(n3398), .ZN(n3383) );
  AND2_X1 U2857 ( .A1(n3756), .A2(n4097), .ZN(n3845) );
  INV_X1 U2858 ( .A(n3845), .ZN(n2158) );
  AND2_X1 U2859 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2037) );
  NAND2_X1 U2860 ( .A1(n2269), .A2(n2023), .ZN(n3492) );
  INV_X1 U2861 ( .A(n4144), .ZN(n4151) );
  AND2_X1 U2862 ( .A1(n3723), .A2(DATAI_22_), .ZN(n4144) );
  NOR2_X1 U2863 ( .A1(n3513), .A2(n2994), .ZN(n3514) );
  OR2_X1 U2864 ( .A1(n3444), .A2(n3462), .ZN(n2038) );
  AND2_X1 U2865 ( .A1(n3677), .A2(n2995), .ZN(n2039) );
  OR2_X1 U2866 ( .A1(n2216), .A2(n3462), .ZN(n2040) );
  NAND2_X1 U2867 ( .A1(n3450), .A2(n2290), .ZN(n3451) );
  NAND2_X1 U2868 ( .A1(n4224), .A2(n2163), .ZN(n4183) );
  INV_X1 U2869 ( .A(n3824), .ZN(n2135) );
  AND2_X1 U2870 ( .A1(n2191), .A2(n2192), .ZN(n2041) );
  AND2_X1 U2871 ( .A1(n2176), .A2(n2178), .ZN(n2042) );
  NAND2_X1 U2872 ( .A1(n4524), .A2(n2367), .ZN(n2997) );
  INV_X1 U2873 ( .A(n3368), .ZN(n2166) );
  NAND2_X1 U2874 ( .A1(n2859), .A2(IR_REG_31__SCAN_IN), .ZN(n3039) );
  OR2_X1 U2875 ( .A1(n2661), .A2(n2660), .ZN(n2043) );
  NAND2_X1 U2876 ( .A1(n2111), .A2(n2066), .ZN(n3235) );
  AND2_X1 U2877 ( .A1(n3717), .A2(DATAI_20_), .ZN(n4177) );
  AND2_X1 U2878 ( .A1(n3717), .A2(DATAI_25_), .ZN(n4088) );
  NAND2_X1 U2879 ( .A1(n3290), .A2(n3289), .ZN(n3288) );
  INV_X1 U2880 ( .A(n2168), .ZN(n2167) );
  NAND2_X1 U2881 ( .A1(n2017), .A2(n2169), .ZN(n2168) );
  INV_X1 U2882 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2190) );
  NAND2_X1 U2883 ( .A1(n4457), .A2(REG1_REG_15__SCAN_IN), .ZN(n2044) );
  INV_X1 U2884 ( .A(n2077), .ZN(n2076) );
  OR2_X1 U2885 ( .A1(n4498), .A2(n2078), .ZN(n2077) );
  INV_X1 U2886 ( .A(IR_REG_0__SCAN_IN), .ZN(n2375) );
  INV_X1 U2887 ( .A(n4463), .ZN(n2073) );
  INV_X1 U2888 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2185) );
  AND2_X1 U2889 ( .A1(n4540), .A2(REG2_REG_18__SCAN_IN), .ZN(n2045) );
  INV_X1 U2890 ( .A(n3985), .ZN(n4542) );
  NAND2_X1 U2891 ( .A1(n3081), .A2(n2193), .ZN(n2046) );
  AND2_X1 U2892 ( .A1(n4540), .A2(REG1_REG_18__SCAN_IN), .ZN(n2047) );
  INV_X1 U2893 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2177) );
  XNOR2_X1 U2894 ( .A(n2424), .B(IR_REG_3__SCAN_IN), .ZN(n4464) );
  INV_X1 U2895 ( .A(n4464), .ZN(n2203) );
  INV_X1 U2896 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2210) );
  INV_X1 U2897 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2222) );
  NAND2_X1 U2898 ( .A1(n3717), .A2(n3031), .ZN(n2052) );
  NAND2_X1 U2899 ( .A1(n3674), .A2(n2056), .ZN(n2054) );
  OAI21_X1 U2900 ( .B1(n3674), .B2(n2056), .A(n2675), .ZN(n2055) );
  INV_X1 U2901 ( .A(n2674), .ZN(n2056) );
  OAI21_X2 U2902 ( .B1(n3005), .B2(n2059), .A(n2057), .ZN(n3539) );
  AND3_X2 U2903 ( .A1(n2409), .A2(n2305), .A3(n2306), .ZN(n2584) );
  NAND3_X1 U2904 ( .A1(n2282), .A2(n2500), .A3(n2283), .ZN(n2065) );
  INV_X1 U2905 ( .A(n3932), .ZN(n2071) );
  OAI21_X1 U2906 ( .B1(n3915), .B2(n2071), .A(n2070), .ZN(n3948) );
  NAND3_X1 U2907 ( .A1(n2207), .A2(n2034), .A3(n2204), .ZN(n3144) );
  INV_X1 U2908 ( .A(n2080), .ZN(n3902) );
  NAND2_X1 U2909 ( .A1(n3900), .A2(n3899), .ZN(n2081) );
  INV_X1 U2910 ( .A(n3898), .ZN(n2082) );
  NAND2_X1 U2911 ( .A1(n2083), .A2(IR_REG_31__SCAN_IN), .ZN(n2396) );
  OAI211_X1 U2912 ( .C1(n4044), .C2(n2090), .A(n2089), .B(n2087), .ZN(n3558)
         );
  NAND2_X1 U2913 ( .A1(n4044), .A2(n2091), .ZN(n2089) );
  NAND2_X1 U2914 ( .A1(n4011), .A2(n2096), .ZN(n2090) );
  INV_X1 U2915 ( .A(n4220), .ZN(n2928) );
  INV_X1 U2916 ( .A(n2239), .ZN(n2106) );
  NAND2_X1 U2917 ( .A1(n2932), .A2(n2931), .ZN(n4171) );
  OAI21_X2 U2918 ( .B1(n2932), .B2(n2106), .A(n2104), .ZN(n2938) );
  NAND2_X1 U2919 ( .A1(n3274), .A2(n3269), .ZN(n3268) );
  NAND3_X1 U2920 ( .A1(n2897), .A2(n2109), .A3(n3268), .ZN(n2223) );
  AND2_X2 U2921 ( .A1(n2307), .A2(n2584), .ZN(n2654) );
  NAND2_X1 U2922 ( .A1(n2114), .A2(n2033), .ZN(n2591) );
  NAND2_X1 U2923 ( .A1(n2115), .A2(n2116), .ZN(n2329) );
  AND2_X1 U2924 ( .A1(n2654), .A2(n2118), .ZN(n2328) );
  NAND2_X1 U2925 ( .A1(n2119), .A2(n2121), .ZN(n2973) );
  NAND2_X1 U2926 ( .A1(n2954), .A2(n2131), .ZN(n2129) );
  OAI21_X1 U2927 ( .B1(n3309), .B2(n2142), .A(n3812), .ZN(n2141) );
  NAND2_X1 U2928 ( .A1(n2654), .A2(n2147), .ZN(n3028) );
  AND2_X1 U2929 ( .A1(n2345), .A2(n2347), .ZN(n2147) );
  OAI21_X1 U2930 ( .B1(n3521), .B2(n2152), .A(n2148), .ZN(n4260) );
  NAND2_X1 U2931 ( .A1(n4098), .A2(n2157), .ZN(n2161) );
  NAND2_X1 U2932 ( .A1(n4098), .A2(n3845), .ZN(n4080) );
  NAND2_X1 U2933 ( .A1(n2886), .A2(n3312), .ZN(n2162) );
  NAND2_X1 U2934 ( .A1(n3514), .A2(n2164), .ZN(n4242) );
  NAND2_X1 U2935 ( .A1(n3112), .A2(n2184), .ZN(n2182) );
  NAND2_X1 U2936 ( .A1(n3086), .A2(n3072), .ZN(n2186) );
  NAND2_X1 U2937 ( .A1(n3322), .A2(n2015), .ZN(n2187) );
  NAND2_X1 U2938 ( .A1(n2189), .A2(n4461), .ZN(n2192) );
  NOR2_X1 U2939 ( .A1(n4461), .A2(REG2_REG_8__SCAN_IN), .ZN(n2188) );
  XNOR2_X1 U2940 ( .A(n3322), .B(n4461), .ZN(n3323) );
  NAND3_X1 U2941 ( .A1(n3077), .A2(n3895), .A3(n3894), .ZN(n2194) );
  NAND3_X1 U2942 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2197) );
  NAND2_X1 U2943 ( .A1(n4490), .A2(n4491), .ZN(n4489) );
  INV_X1 U2944 ( .A(n2202), .ZN(n3991) );
  NAND2_X1 U2945 ( .A1(n3074), .A2(n3072), .ZN(n2211) );
  NAND2_X1 U2946 ( .A1(n3459), .A2(n2215), .ZN(n2214) );
  XNOR2_X1 U2947 ( .A(n3964), .B(n3949), .ZN(n3950) );
  NAND2_X1 U2948 ( .A1(n3210), .A2(n2899), .ZN(n3308) );
  NAND2_X1 U2949 ( .A1(n2226), .A2(n2225), .ZN(n3210) );
  OAI211_X1 U2950 ( .C1(n2226), .C2(n2224), .A(n2223), .B(n2900), .ZN(n2902)
         );
  INV_X1 U2951 ( .A(n2899), .ZN(n2224) );
  MUX2_X1 U2952 ( .A(n2475), .B(n3202), .S(n3061), .Z(n3369) );
  NAND2_X1 U2953 ( .A1(n2654), .A2(n2238), .ZN(n2859) );
  NAND2_X1 U2954 ( .A1(n2251), .A2(n2252), .ZN(n4044) );
  NAND2_X1 U2955 ( .A1(n2938), .A2(n2937), .ZN(n4096) );
  NOR2_X1 U2956 ( .A1(n2940), .A2(n2260), .ZN(n2259) );
  INV_X1 U2957 ( .A(n2937), .ZN(n2260) );
  NAND2_X1 U2958 ( .A1(n3566), .A2(n2265), .ZN(n2264) );
  NAND2_X1 U2959 ( .A1(n3480), .A2(n2280), .ZN(n2279) );
  NAND2_X1 U2960 ( .A1(n2270), .A2(n2273), .ZN(n2589) );
  NAND2_X1 U2961 ( .A1(n3480), .A2(n2271), .ZN(n2270) );
  NAND2_X1 U2962 ( .A1(n3626), .A2(n2281), .ZN(n2283) );
  INV_X1 U2963 ( .A(n3893), .ZN(n3081) );
  NAND2_X1 U2964 ( .A1(n3078), .A2(n3077), .ZN(n3893) );
  NAND2_X1 U2965 ( .A1(n4465), .A2(REG2_REG_2__SCAN_IN), .ZN(n3077) );
  OR2_X1 U2966 ( .A1(n4465), .A2(REG2_REG_2__SCAN_IN), .ZN(n3078) );
  INV_X1 U2967 ( .A(IR_REG_6__SCAN_IN), .ZN(n2471) );
  OR3_X1 U2968 ( .A1(n4316), .A2(n4577), .A3(n4318), .ZN(n4325) );
  XNOR2_X1 U2969 ( .A(n2365), .B(n2398), .ZN(n2385) );
  XNOR2_X1 U2970 ( .A(n2399), .B(n2792), .ZN(n2404) );
  XNOR2_X1 U2971 ( .A(n2385), .B(n2386), .ZN(n3161) );
  INV_X1 U2972 ( .A(n3270), .ZN(n2993) );
  XNOR2_X1 U2973 ( .A(n2435), .B(n2434), .ZN(n3237) );
  OR2_X1 U2974 ( .A1(n4108), .A2(n2784), .ZN(n2746) );
  OR2_X1 U2975 ( .A1(n4133), .A2(n2784), .ZN(n2732) );
  OR2_X1 U2976 ( .A1(n4210), .A2(n2784), .ZN(n2684) );
  OAI211_X1 U2977 ( .C1(n3606), .C2(n2784), .A(n2566), .B(n2565), .ZN(n3877)
         );
  OR2_X1 U2978 ( .A1(n2784), .A2(n2369), .ZN(n2372) );
  INV_X1 U2979 ( .A(n3037), .ZN(n2350) );
  INV_X1 U2980 ( .A(n3998), .ZN(n4028) );
  INV_X1 U2981 ( .A(n2894), .ZN(n4522) );
  NAND2_X1 U2982 ( .A1(n3539), .A2(n3536), .ZN(n3643) );
  INV_X1 U2983 ( .A(n3114), .ZN(n3072) );
  OR2_X1 U2984 ( .A1(n3982), .A2(n3981), .ZN(n2289) );
  OR2_X1 U2985 ( .A1(n3449), .A2(n3448), .ZN(n2290) );
  OR2_X1 U2986 ( .A1(n3449), .A2(n3441), .ZN(n2291) );
  AND2_X1 U2987 ( .A1(n2342), .A2(IR_REG_28__SCAN_IN), .ZN(n2292) );
  NAND2_X1 U2988 ( .A1(n2955), .A2(n2170), .ZN(n2911) );
  INV_X1 U2989 ( .A(IR_REG_30__SCAN_IN), .ZN(n3029) );
  AND3_X1 U2990 ( .A1(n2847), .A2(n2846), .A3(n3623), .ZN(n2293) );
  NAND2_X1 U2991 ( .A1(n2647), .A2(n3615), .ZN(n2294) );
  INV_X1 U2992 ( .A(n3880), .ZN(n3354) );
  INV_X1 U2993 ( .A(n4458), .ZN(n3909) );
  OR2_X1 U2994 ( .A1(n3258), .A2(n3881), .ZN(n2295) );
  NAND2_X2 U2995 ( .A1(n3222), .A2(n4255), .ZN(n4535) );
  AND2_X1 U2996 ( .A1(n4120), .A2(n2970), .ZN(n4142) );
  AND2_X1 U2997 ( .A1(n3419), .A2(n3879), .ZN(n2296) );
  OR2_X1 U2998 ( .A1(n3389), .A2(n3880), .ZN(n2297) );
  NAND2_X1 U2999 ( .A1(n2502), .A2(n2501), .ZN(n2298) );
  MUX2_X1 U3000 ( .A(n4461), .B(DATAI_8_), .S(n3723), .Z(n3389) );
  OR2_X1 U3001 ( .A1(n3554), .A2(n4391), .ZN(n2299) );
  OR2_X1 U3002 ( .A1(n3554), .A2(n4451), .ZN(n2300) );
  INV_X1 U3003 ( .A(n2654), .ZN(n2655) );
  NAND2_X1 U3004 ( .A1(n2378), .A2(n2364), .ZN(n2422) );
  INV_X1 U3005 ( .A(n3485), .ZN(n2913) );
  NAND2_X1 U3006 ( .A1(n3495), .A2(n3485), .ZN(n2915) );
  INV_X1 U3007 ( .A(n4223), .ZN(n2927) );
  NOR2_X1 U3008 ( .A1(n2344), .A2(n2343), .ZN(n2345) );
  AND2_X1 U3009 ( .A1(n3017), .A2(n3018), .ZN(n2736) );
  OR2_X1 U3010 ( .A1(n2761), .A2(n3542), .ZN(n2765) );
  AND2_X1 U3011 ( .A1(n4465), .A2(REG2_REG_2__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U3012 ( .A1(n3909), .A2(REG2_REG_11__SCAN_IN), .ZN(n3910) );
  INV_X1 U3013 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2489) );
  AND2_X1 U3014 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  INV_X1 U3015 ( .A(n2567), .ZN(n2433) );
  OR2_X1 U3016 ( .A1(n2784), .A2(n3243), .ZN(n2428) );
  AND2_X1 U3017 ( .A1(n3729), .A2(n3726), .ZN(n3759) );
  NAND2_X1 U3018 ( .A1(n3289), .A2(n2947), .ZN(n3214) );
  NOR2_X1 U3019 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2305)
         );
  OR2_X1 U3020 ( .A1(n4046), .A2(n2784), .ZN(n2789) );
  OR2_X1 U3021 ( .A1(n4187), .A2(n2784), .ZN(n2696) );
  OR2_X1 U3022 ( .A1(n2442), .A2(n2391), .ZN(n2392) );
  XNOR2_X1 U3023 ( .A(n3149), .B(n4463), .ZN(n3151) );
  INV_X1 U3024 ( .A(n4501), .ZN(n4502) );
  INV_X1 U3025 ( .A(n4279), .ZN(n4277) );
  OR2_X1 U3026 ( .A1(n2837), .A2(n2367), .ZN(n4278) );
  INV_X1 U3027 ( .A(n3525), .ZN(n3572) );
  INV_X1 U3028 ( .A(n2997), .ZN(n2998) );
  AND2_X1 U3029 ( .A1(n2875), .A2(n3136), .ZN(n3689) );
  AND2_X1 U3030 ( .A1(n2868), .A2(n2864), .ZN(n3695) );
  INV_X1 U3031 ( .A(n4526), .ZN(n3978) );
  AND2_X1 U3032 ( .A1(n2746), .A2(n2745), .ZN(n4124) );
  NAND3_X1 U3033 ( .A1(n3884), .A2(REG1_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3900) );
  INV_X1 U3034 ( .A(n4497), .ZN(n4494) );
  INV_X1 U3035 ( .A(n4286), .ZN(n4231) );
  INV_X1 U3036 ( .A(n4305), .ZN(n4516) );
  AOI21_X1 U3037 ( .B1(n2820), .B2(n3055), .A(n3054), .ZN(n3000) );
  AND2_X1 U3038 ( .A1(n4528), .A2(n4551), .ZN(n4577) );
  INV_X1 U3039 ( .A(n4577), .ZN(n4570) );
  AND2_X1 U3040 ( .A1(n4539), .A2(n2378), .ZN(n3058) );
  NAND2_X1 U3041 ( .A1(n2557), .A2(n2554), .ZN(n4458) );
  AND2_X1 U3042 ( .A1(n3076), .A2(n3064), .ZN(n4500) );
  NAND2_X1 U3043 ( .A1(n2855), .A2(n2854), .ZN(n3872) );
  OR2_X1 U3044 ( .A1(n4469), .A2(n3866), .ZN(n3939) );
  OR2_X1 U3045 ( .A1(n4469), .A2(n4467), .ZN(n4497) );
  NAND2_X1 U3046 ( .A1(n4535), .A2(n3307), .ZN(n4286) );
  NAND2_X1 U3047 ( .A1(n4589), .A2(n2998), .ZN(n4391) );
  NAND2_X1 U3048 ( .A1(n4739), .A2(n2998), .ZN(n4451) );
  INV_X1 U3049 ( .A(n4739), .ZN(n4737) );
  INV_X1 U3050 ( .A(n4537), .ZN(n4538) );
  NAND2_X1 U3051 ( .A1(n3053), .A2(n3058), .ZN(n4537) );
  XNOR2_X1 U3052 ( .A(n2318), .B(IR_REG_25__SCAN_IN), .ZN(n4455) );
  AND2_X1 U3053 ( .A1(n2631), .A2(n2616), .ZN(n4457) );
  NAND4_X1 U3054 ( .A1(n2303), .A2(n2302), .A3(n2301), .A4(n2471), .ZN(n2582)
         );
  NAND4_X1 U3055 ( .A1(n2614), .A2(n2601), .A3(n2585), .A4(n2632), .ZN(n2304)
         );
  NOR2_X1 U3056 ( .A1(n2582), .A2(n2304), .ZN(n2307) );
  INV_X1 U3057 ( .A(IR_REG_18__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U3058 ( .A1(n2328), .A2(n2310), .ZN(n2332) );
  INV_X1 U3059 ( .A(n2332), .ZN(n2312) );
  INV_X1 U3060 ( .A(IR_REG_21__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U3061 ( .A1(n2312), .A2(n2311), .ZN(n2360) );
  NAND2_X1 U3062 ( .A1(n2811), .A2(n2814), .ZN(n2326) );
  NAND4_X1 U3063 ( .A1(n2316), .A2(n2315), .A3(n2314), .A4(n2313), .ZN(n2344)
         );
  INV_X1 U3064 ( .A(n2344), .ZN(n2319) );
  NAND2_X1 U3065 ( .A1(n2654), .A2(n2319), .ZN(n2317) );
  NAND2_X1 U3066 ( .A1(n2317), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U3067 ( .A1(n2334), .A2(IR_REG_31__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U3068 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U3069 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .ZN(n2323) );
  OAI21_X1 U3070 ( .B1(n2814), .B2(IR_REG_31__SCAN_IN), .A(n2323), .ZN(n2324)
         );
  NAND2_X1 U3071 ( .A1(n2339), .A2(n3270), .ZN(n2359) );
  NAND4_X1 U3072 ( .A1(n2335), .A2(n2342), .A3(n2341), .A4(n2340), .ZN(n2343)
         );
  XNOR2_X2 U3073 ( .A(n2346), .B(IR_REG_30__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3074 ( .A1(n2349), .A2(REG2_REG_1__SCAN_IN), .ZN(n2353) );
  OR2_X2 U3075 ( .A1(n3037), .A2(n2354), .ZN(n2443) );
  INV_X1 U3076 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U3077 ( .A1(n2410), .A2(REG0_REG_1__SCAN_IN), .ZN(n2351) );
  INV_X1 U3078 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U3079 ( .A1(n2355), .A2(REG3_REG_1__SCAN_IN), .ZN(n2356) );
  NAND2_X2 U3080 ( .A1(n2357), .A2(n2356), .ZN(n2894) );
  NAND2_X1 U3081 ( .A1(n2894), .A2(n2567), .ZN(n2358) );
  NAND2_X1 U3082 ( .A1(n2359), .A2(n2358), .ZN(n2365) );
  XNOR2_X2 U3083 ( .A(n2362), .B(n2363), .ZN(n4526) );
  NAND2_X1 U3084 ( .A1(n2838), .A2(n4526), .ZN(n2856) );
  INV_X1 U3085 ( .A(n2838), .ZN(n2366) );
  INV_X1 U3086 ( .A(n2839), .ZN(n3761) );
  INV_X1 U3087 ( .A(n2837), .ZN(n4524) );
  NAND2_X1 U3088 ( .A1(n3270), .A2(n2567), .ZN(n2368) );
  INV_X2 U3089 ( .A(n2443), .ZN(n2850) );
  NAND2_X1 U3090 ( .A1(n2850), .A2(REG1_REG_0__SCAN_IN), .ZN(n2373) );
  INV_X1 U3091 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3092 ( .A1(n2349), .A2(REG2_REG_0__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3093 ( .A1(n2410), .A2(REG0_REG_0__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3094 ( .A1(n2567), .A2(n2893), .ZN(n2377) );
  INV_X1 U3095 ( .A(n2378), .ZN(n3016) );
  NAND2_X1 U3096 ( .A1(n3016), .A2(REG1_REG_0__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3097 ( .A1(n2382), .A2(n2379), .ZN(n3116) );
  INV_X1 U3098 ( .A(n2893), .ZN(n3159) );
  NAND2_X1 U3099 ( .A1(n3016), .A2(IR_REG_0__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3100 ( .A1(n3267), .A2(n2567), .ZN(n2380) );
  NAND2_X1 U3101 ( .A1(n3116), .A2(n3115), .ZN(n2384) );
  NAND2_X1 U3102 ( .A1(n2382), .A2(n2398), .ZN(n2383) );
  NAND2_X1 U3103 ( .A1(n2384), .A2(n2383), .ZN(n3164) );
  NAND2_X1 U3104 ( .A1(n3161), .A2(n3164), .ZN(n3162) );
  INV_X1 U3105 ( .A(n2385), .ZN(n2387) );
  NAND2_X1 U3106 ( .A1(n2387), .A2(n2386), .ZN(n2388) );
  NAND2_X1 U3107 ( .A1(n3162), .A2(n2388), .ZN(n3130) );
  INV_X1 U3108 ( .A(n3130), .ZN(n2402) );
  INV_X1 U3109 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2389) );
  OR2_X1 U3110 ( .A1(n2443), .A2(n2389), .ZN(n2394) );
  INV_X1 U3111 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2391) );
  AND4_X2 U3112 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n2896)
         );
  XNOR2_X2 U3113 ( .A(n2396), .B(IR_REG_2__SCAN_IN), .ZN(n4465) );
  MUX2_X1 U3114 ( .A(n4465), .B(DATAI_2_), .S(n3717), .Z(n3179) );
  NAND2_X1 U3115 ( .A1(n3179), .A2(n2339), .ZN(n2397) );
  OAI21_X1 U3116 ( .B1(n2433), .B2(n2896), .A(n2397), .ZN(n2399) );
  NAND2_X1 U3117 ( .A1(n3179), .A2(n2567), .ZN(n2400) );
  OAI21_X1 U3118 ( .B1(n2416), .B2(n2896), .A(n2400), .ZN(n2403) );
  XNOR2_X1 U3119 ( .A(n2404), .B(n2403), .ZN(n3129) );
  INV_X1 U3120 ( .A(n3129), .ZN(n2401) );
  NAND2_X1 U3121 ( .A1(n2402), .A2(n2401), .ZN(n3132) );
  INV_X1 U3122 ( .A(n2403), .ZN(n2406) );
  INV_X1 U3123 ( .A(n2404), .ZN(n2405) );
  NAND2_X1 U3124 ( .A1(n2406), .A2(n2405), .ZN(n2407) );
  NAND2_X1 U3125 ( .A1(n3132), .A2(n2407), .ZN(n3192) );
  INV_X1 U3126 ( .A(IR_REG_2__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3127 ( .A1(n2409), .A2(n2408), .ZN(n2437) );
  NAND2_X1 U3128 ( .A1(n2437), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  MUX2_X1 U3129 ( .A(n4464), .B(DATAI_3_), .S(n3717), .Z(n3194) );
  NAND2_X1 U3130 ( .A1(n3194), .A2(n2339), .ZN(n2415) );
  NAND2_X1 U3131 ( .A1(n2850), .A2(REG1_REG_3__SCAN_IN), .ZN(n2414) );
  OR2_X1 U3132 ( .A1(n2784), .A2(REG3_REG_3__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3133 ( .A1(n2349), .A2(REG2_REG_3__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3134 ( .A1(n2410), .A2(REG0_REG_3__SCAN_IN), .ZN(n2411) );
  INV_X4 U3135 ( .A(n2433), .ZN(n2858) );
  NAND2_X1 U3136 ( .A1(n3194), .A2(n2858), .ZN(n2417) );
  OAI21_X1 U3137 ( .B1(n2805), .B2(n2947), .A(n2417), .ZN(n2418) );
  XNOR2_X1 U3138 ( .A(n2419), .B(n2418), .ZN(n3193) );
  INV_X1 U3139 ( .A(n2418), .ZN(n2420) );
  NAND2_X1 U3140 ( .A1(n2420), .A2(n2419), .ZN(n2421) );
  INV_X1 U3141 ( .A(IR_REG_3__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3142 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  NAND2_X1 U3143 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2427) );
  INV_X1 U3144 ( .A(IR_REG_4__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3145 ( .A(n2427), .B(n2426), .ZN(n3114) );
  INV_X1 U3146 ( .A(DATAI_4_), .ZN(n3031) );
  NAND2_X1 U3147 ( .A1(n2850), .A2(REG1_REG_4__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U31480 ( .A1(n2410), .A2(REG0_REG_4__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U31490 ( .A1(n2349), .A2(REG2_REG_4__SCAN_IN), .ZN(n2429) );
  OAI21_X1 U3150 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2447), .ZN(n3243) );
  XNOR2_X1 U3151 ( .A(n2432), .B(n2792), .ZN(n2435) );
  OAI22_X1 U3152 ( .A1(n2805), .A2(n2887), .B1(n2886), .B2(n2433), .ZN(n2434)
         );
  NAND2_X1 U3153 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3154 ( .A1(n3235), .A2(n2436), .ZN(n3626) );
  NAND2_X1 U3155 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2440) );
  INV_X1 U3156 ( .A(DATAI_5_), .ZN(n2441) );
  NAND2_X1 U3157 ( .A1(n3719), .A2(REG0_REG_5__SCAN_IN), .ZN(n2452) );
  INV_X1 U3158 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2444) );
  OR2_X1 U3159 ( .A1(n2443), .A2(n2444), .ZN(n2451) );
  INV_X1 U3160 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3161 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NAND2_X1 U3162 ( .A1(n2460), .A2(n2448), .ZN(n3630) );
  OR2_X1 U3163 ( .A1(n2784), .A2(n3630), .ZN(n2450) );
  INV_X1 U3164 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3315) );
  OR2_X1 U3165 ( .A1(n3722), .A2(n3315), .ZN(n2449) );
  OAI22_X1 U3166 ( .A1(n3312), .A2(n2807), .B1(n2949), .B2(n2433), .ZN(n2453)
         );
  XNOR2_X1 U3167 ( .A(n2453), .B(n2398), .ZN(n2454) );
  OAI22_X1 U3168 ( .A1(n2805), .A2(n2949), .B1(n3312), .B2(n2794), .ZN(n2455)
         );
  XNOR2_X1 U3169 ( .A(n2454), .B(n2455), .ZN(n3625) );
  INV_X1 U3170 ( .A(n2454), .ZN(n2456) );
  NAND2_X1 U3171 ( .A1(n2456), .A2(n2455), .ZN(n2457) );
  NAND2_X1 U3172 ( .A1(n3719), .A2(REG0_REG_6__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3173 ( .A1(n2850), .A2(REG1_REG_6__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3174 ( .A1(n2349), .A2(REG2_REG_6__SCAN_IN), .ZN(n2463) );
  INV_X1 U3175 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3176 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  NAND2_X1 U3177 ( .A1(n2477), .A2(n2461), .ZN(n3338) );
  OR2_X1 U3178 ( .A1(n2784), .A2(n3338), .ZN(n2462) );
  NAND4_X1 U3179 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3881)
         );
  INV_X1 U3180 ( .A(n3881), .ZN(n2950) );
  OR2_X1 U3181 ( .A1(n2584), .A2(n2327), .ZN(n2466) );
  XNOR2_X1 U3182 ( .A(n2466), .B(IR_REG_6__SCAN_IN), .ZN(n4463) );
  MUX2_X1 U3183 ( .A(n4463), .B(DATAI_6_), .S(n3717), .Z(n3258) );
  NAND2_X1 U3184 ( .A1(n3258), .A2(n2858), .ZN(n2467) );
  OAI21_X1 U3185 ( .B1(n2805), .B2(n2950), .A(n2467), .ZN(n3254) );
  NAND2_X1 U3186 ( .A1(n3258), .A2(n2339), .ZN(n2469) );
  NAND2_X1 U3187 ( .A1(n2858), .A2(n3881), .ZN(n2468) );
  NAND2_X1 U3188 ( .A1(n2469), .A2(n2468), .ZN(n2470) );
  XNOR2_X1 U3189 ( .A(n2470), .B(n2792), .ZN(n3255) );
  NAND2_X1 U3190 ( .A1(n2584), .A2(n2471), .ZN(n2505) );
  NAND2_X1 U3191 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3192 ( .A1(n2473), .A2(n2472), .ZN(n2487) );
  OR2_X1 U3193 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  NAND2_X1 U3194 ( .A1(n2487), .A2(n2474), .ZN(n3202) );
  INV_X1 U3195 ( .A(DATAI_7_), .ZN(n2475) );
  NAND2_X1 U3196 ( .A1(n2850), .A2(REG1_REG_7__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3197 ( .A1(n2349), .A2(REG2_REG_7__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3198 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
  NAND2_X1 U3199 ( .A1(n2490), .A2(n2478), .ZN(n3403) );
  OR2_X1 U3200 ( .A1(n2784), .A2(n3403), .ZN(n2479) );
  OAI22_X1 U3201 ( .A1(n3369), .A2(n2807), .B1(n2904), .B2(n2794), .ZN(n2483)
         );
  XNOR2_X1 U3202 ( .A(n2483), .B(n2398), .ZN(n2484) );
  OAI22_X1 U3203 ( .A1(n2805), .A2(n2904), .B1(n3369), .B2(n2794), .ZN(n2485)
         );
  XNOR2_X1 U3204 ( .A(n2484), .B(n2485), .ZN(n3398) );
  INV_X1 U3205 ( .A(n2484), .ZN(n2486) );
  NAND2_X1 U3206 ( .A1(n2486), .A2(n2485), .ZN(n3384) );
  NAND2_X1 U3207 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  XNOR2_X1 U3208 ( .A(n2488), .B(IR_REG_8__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U3209 ( .A1(n3389), .A2(n2339), .ZN(n2497) );
  NAND2_X1 U32100 ( .A1(n3719), .A2(REG0_REG_8__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U32110 ( .A1(n2850), .A2(REG1_REG_8__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U32120 ( .A1(n2349), .A2(REG2_REG_8__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U32130 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U32140 ( .A1(n2508), .A2(n2491), .ZN(n3393) );
  OR2_X1 U32150 ( .A1(n2784), .A2(n3393), .ZN(n2492) );
  NAND4_X1 U32160 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3880)
         );
  NAND2_X1 U32170 ( .A1(n2567), .A2(n3880), .ZN(n2496) );
  NAND2_X1 U32180 ( .A1(n2497), .A2(n2496), .ZN(n2498) );
  XNOR2_X1 U32190 ( .A(n2498), .B(n2792), .ZN(n2502) );
  NAND2_X1 U32200 ( .A1(n3389), .A2(n2858), .ZN(n2499) );
  OAI21_X1 U32210 ( .B1(n2805), .B2(n3354), .A(n2499), .ZN(n2501) );
  AND2_X1 U32220 ( .A1(n3384), .A2(n2298), .ZN(n2500) );
  INV_X1 U32230 ( .A(n2501), .ZN(n2504) );
  INV_X1 U32240 ( .A(n2502), .ZN(n2503) );
  NAND2_X1 U32250 ( .A1(n2504), .A2(n2503), .ZN(n3385) );
  NAND2_X1 U32260 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U32270 ( .A(n2506), .B(IR_REG_9__SCAN_IN), .ZN(n4460) );
  MUX2_X1 U32280 ( .A(n4460), .B(DATAI_9_), .S(n3723), .Z(n3419) );
  NAND2_X1 U32290 ( .A1(n3419), .A2(n2339), .ZN(n2515) );
  INV_X1 U32300 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4675) );
  OR2_X1 U32310 ( .A1(n2442), .A2(n4675), .ZN(n2513) );
  NAND2_X1 U32320 ( .A1(n2850), .A2(REG1_REG_9__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32330 ( .A1(n2349), .A2(REG2_REG_9__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U32340 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  NAND2_X1 U32350 ( .A1(n2528), .A2(n2509), .ZN(n3434) );
  OR2_X1 U32360 ( .A1(n2784), .A2(n3434), .ZN(n2510) );
  NAND2_X1 U32370 ( .A1(n2858), .A2(n3879), .ZN(n2514) );
  NAND2_X1 U32380 ( .A1(n2515), .A2(n2514), .ZN(n2516) );
  XNOR2_X1 U32390 ( .A(n2516), .B(n2398), .ZN(n2519) );
  NAND2_X1 U32400 ( .A1(n3419), .A2(n2858), .ZN(n2517) );
  OAI21_X1 U32410 ( .B1(n2805), .B2(n2955), .A(n2517), .ZN(n2518) );
  XNOR2_X1 U32420 ( .A(n2519), .B(n2518), .ZN(n3418) );
  INV_X1 U32430 ( .A(n2518), .ZN(n2520) );
  NAND2_X1 U32440 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  INV_X1 U32450 ( .A(n2522), .ZN(n2524) );
  INV_X1 U32460 ( .A(IR_REG_9__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32470 ( .A1(n2524), .A2(n2523), .ZN(n2549) );
  NAND2_X1 U32480 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2525) );
  XNOR2_X1 U32490 ( .A(n2525), .B(IR_REG_10__SCAN_IN), .ZN(n4459) );
  MUX2_X1 U32500 ( .A(n4459), .B(DATAI_10_), .S(n3723), .Z(n3495) );
  NAND2_X1 U32510 ( .A1(n3495), .A2(n2339), .ZN(n2535) );
  INV_X1 U32520 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4674) );
  OR2_X1 U32530 ( .A1(n2442), .A2(n4674), .ZN(n2533) );
  INV_X1 U32540 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U32550 ( .A1(n2349), .A2(REG2_REG_10__SCAN_IN), .ZN(n2531) );
  INV_X1 U32560 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U32570 ( .A1(n2528), .A2(n2527), .ZN(n2529) );
  NAND2_X1 U32580 ( .A1(n2543), .A2(n2529), .ZN(n3499) );
  OR2_X1 U32590 ( .A1(n2784), .A2(n3499), .ZN(n2530) );
  NAND2_X1 U32600 ( .A1(n2858), .A2(n3485), .ZN(n2534) );
  NAND2_X1 U32610 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  XNOR2_X1 U32620 ( .A(n2536), .B(n2792), .ZN(n2540) );
  NAND2_X1 U32630 ( .A1(n3495), .A2(n2858), .ZN(n2537) );
  OAI21_X1 U32640 ( .B1(n2805), .B2(n2913), .A(n2537), .ZN(n2539) );
  XNOR2_X1 U32650 ( .A(n2540), .B(n2539), .ZN(n3494) );
  INV_X1 U32660 ( .A(n3494), .ZN(n2538) );
  NAND2_X1 U32670 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  NAND2_X1 U32680 ( .A1(n3492), .A2(n2541), .ZN(n3480) );
  NAND2_X1 U32690 ( .A1(n2850), .A2(REG1_REG_11__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32700 ( .A1(n2543), .A2(n2542), .ZN(n2544) );
  AND2_X1 U32710 ( .A1(n2561), .A2(n2544), .ZN(n4303) );
  NAND2_X1 U32720 ( .A1(n2002), .A2(n4303), .ZN(n2547) );
  NAND2_X1 U32730 ( .A1(n2349), .A2(REG2_REG_11__SCAN_IN), .ZN(n2546) );
  INV_X1 U32740 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4625) );
  OR2_X1 U32750 ( .A1(n2442), .A2(n4625), .ZN(n2545) );
  NAND4_X1 U32760 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n3878)
         );
  INV_X1 U32770 ( .A(n2549), .ZN(n2551) );
  INV_X1 U32780 ( .A(IR_REG_10__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32790 ( .A1(n2551), .A2(n2550), .ZN(n2552) );
  NAND2_X1 U32800 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32810 ( .A1(n2553), .A2(n4718), .ZN(n2557) );
  OR2_X1 U32820 ( .A1(n2553), .A2(n4718), .ZN(n2554) );
  INV_X1 U32830 ( .A(DATAI_11_), .ZN(n2555) );
  MUX2_X1 U32840 ( .A(n4458), .B(n2555), .S(n3723), .Z(n4300) );
  OAI22_X1 U32850 ( .A1(n2805), .A2(n3469), .B1(n4300), .B2(n2808), .ZN(n3482)
         );
  OAI22_X1 U32860 ( .A1(n4300), .A2(n2807), .B1(n3469), .B2(n2808), .ZN(n2556)
         );
  XNOR2_X1 U32870 ( .A(n2556), .B(n2792), .ZN(n3481) );
  NAND2_X1 U32880 ( .A1(n2557), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  XNOR2_X1 U32890 ( .A(n2558), .B(IR_REG_12__SCAN_IN), .ZN(n3912) );
  MUX2_X1 U32900 ( .A(n3912), .B(DATAI_12_), .S(n3723), .Z(n3603) );
  NAND2_X1 U32910 ( .A1(n3603), .A2(n2339), .ZN(n2569) );
  INV_X1 U32920 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32930 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND2_X1 U32940 ( .A1(n2577), .A2(n2562), .ZN(n3606) );
  NAND2_X1 U32950 ( .A1(n3719), .A2(REG0_REG_12__SCAN_IN), .ZN(n2564) );
  INV_X1 U32960 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4626) );
  OR2_X1 U32970 ( .A1(n2443), .A2(n4626), .ZN(n2563) );
  AND2_X1 U32980 ( .A1(n2564), .A2(n2563), .ZN(n2566) );
  NAND2_X1 U32990 ( .A1(n2349), .A2(REG2_REG_12__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U33000 ( .A1(n2567), .A2(n3877), .ZN(n2568) );
  NAND2_X1 U33010 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  XNOR2_X1 U33020 ( .A(n2570), .B(n2792), .ZN(n2573) );
  INV_X1 U33030 ( .A(n3877), .ZN(n4289) );
  NAND2_X1 U33040 ( .A1(n3603), .A2(n2858), .ZN(n2571) );
  OAI21_X1 U33050 ( .B1(n2805), .B2(n4289), .A(n2571), .ZN(n2572) );
  AND2_X1 U33060 ( .A1(n2573), .A2(n2572), .ZN(n3599) );
  INV_X1 U33070 ( .A(n2572), .ZN(n2575) );
  INV_X1 U33080 ( .A(n2573), .ZN(n2574) );
  NAND2_X1 U33090 ( .A1(n2575), .A2(n2574), .ZN(n3600) );
  NAND2_X1 U33100 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
  AND2_X1 U33110 ( .A1(n2609), .A2(n2578), .ZN(n3661) );
  NAND2_X1 U33120 ( .A1(n3661), .A2(n2002), .ZN(n2581) );
  AOI22_X1 U33130 ( .A1(n3719), .A2(REG0_REG_13__SCAN_IN), .B1(n2850), .B2(
        REG1_REG_13__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U33140 ( .A1(n2349), .A2(REG2_REG_13__SCAN_IN), .ZN(n2579) );
  INV_X1 U33150 ( .A(n2582), .ZN(n2583) );
  NAND2_X1 U33160 ( .A1(n2584), .A2(n2583), .ZN(n2599) );
  NAND2_X1 U33170 ( .A1(n2599), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U33180 ( .A(n2586), .B(n2585), .ZN(n3934) );
  INV_X1 U33190 ( .A(DATAI_13_), .ZN(n2587) );
  OAI22_X1 U33200 ( .A1(n3522), .A2(n2808), .B1(n3659), .B2(n2807), .ZN(n2588)
         );
  XNOR2_X1 U33210 ( .A(n2588), .B(n2398), .ZN(n3654) );
  NAND2_X1 U33220 ( .A1(n2589), .A2(n3655), .ZN(n2592) );
  INV_X1 U33230 ( .A(n3654), .ZN(n2590) );
  NAND2_X1 U33240 ( .A1(n2592), .A2(n2591), .ZN(n3566) );
  XNOR2_X1 U33250 ( .A(n2609), .B(REG3_REG_14__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U33260 ( .A1(n3574), .A2(n2002), .ZN(n2598) );
  INV_X1 U33270 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33280 ( .A1(n3719), .A2(REG0_REG_14__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U33290 ( .A1(n2850), .A2(REG1_REG_14__SCAN_IN), .ZN(n2593) );
  OAI211_X1 U33300 ( .C1(n2595), .C2(n3722), .A(n2594), .B(n2593), .ZN(n2596)
         );
  INV_X1 U33310 ( .A(n2596), .ZN(n2597) );
  NOR2_X1 U33320 ( .A1(n2599), .A2(IR_REG_13__SCAN_IN), .ZN(n2602) );
  OR2_X1 U33330 ( .A1(n2602), .A2(n2327), .ZN(n2600) );
  MUX2_X1 U33340 ( .A(n2600), .B(IR_REG_31__SCAN_IN), .S(n2601), .Z(n2603) );
  NAND2_X1 U33350 ( .A1(n2602), .A2(n2601), .ZN(n2613) );
  MUX2_X1 U33360 ( .A(n3963), .B(DATAI_14_), .S(n3723), .Z(n3525) );
  NAND2_X1 U33370 ( .A1(n3525), .A2(n2339), .ZN(n2604) );
  OAI21_X1 U33380 ( .B1(n3705), .B2(n2794), .A(n2604), .ZN(n2605) );
  XNOR2_X1 U33390 ( .A(n2605), .B(n2792), .ZN(n2637) );
  NAND2_X1 U33400 ( .A1(n3525), .A2(n2858), .ZN(n2606) );
  OAI21_X1 U33410 ( .B1(n2805), .B2(n3705), .A(n2606), .ZN(n2638) );
  INV_X1 U33420 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3981) );
  INV_X1 U33430 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2608) );
  INV_X1 U33440 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2607) );
  OAI21_X1 U33450 ( .B1(n2609), .B2(n2608), .A(n2607), .ZN(n2610) );
  AND2_X1 U33460 ( .A1(n2610), .A2(n2624), .ZN(n4281) );
  NAND2_X1 U33470 ( .A1(n4281), .A2(n2002), .ZN(n2612) );
  AOI22_X1 U33480 ( .A1(n3719), .A2(REG0_REG_15__SCAN_IN), .B1(n2850), .B2(
        REG1_REG_15__SCAN_IN), .ZN(n2611) );
  OAI211_X1 U33490 ( .C1(n3722), .C2(n3981), .A(n2612), .B(n2611), .ZN(n4262)
         );
  NAND2_X1 U33500 ( .A1(n2796), .A2(n4262), .ZN(n2618) );
  NAND2_X1 U33510 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U33520 ( .A1(n2615), .A2(n2614), .ZN(n2631) );
  OR2_X1 U3353 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  MUX2_X1 U33540 ( .A(n4457), .B(DATAI_15_), .S(n3717), .Z(n4279) );
  NAND2_X1 U3355 ( .A1(n4279), .A2(n2858), .ZN(n2617) );
  NAND2_X1 U3356 ( .A1(n2618), .A2(n2617), .ZN(n2642) );
  NAND2_X1 U3357 ( .A1(n4262), .A2(n2858), .ZN(n2620) );
  NAND2_X1 U3358 ( .A1(n4279), .A2(n2339), .ZN(n2619) );
  NAND2_X1 U3359 ( .A1(n2620), .A2(n2619), .ZN(n2621) );
  XNOR2_X1 U3360 ( .A(n2621), .B(n2792), .ZN(n3612) );
  INV_X1 U3361 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3362 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  NAND2_X1 U3363 ( .A1(n2664), .A2(n2625), .ZN(n4256) );
  OR2_X1 U3364 ( .A1(n4256), .A2(n2784), .ZN(n2630) );
  INV_X1 U3365 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U3366 ( .A1(n3719), .A2(REG0_REG_16__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U3367 ( .A1(n2349), .A2(REG2_REG_16__SCAN_IN), .ZN(n2626) );
  OAI211_X1 U3368 ( .C1(n2443), .C2(n4476), .A(n2627), .B(n2626), .ZN(n2628)
         );
  INV_X1 U3369 ( .A(n2628), .ZN(n2629) );
  NAND2_X1 U3370 ( .A1(n2631), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  XNOR2_X1 U3371 ( .A(n2633), .B(n2632), .ZN(n4543) );
  INV_X1 U3372 ( .A(n4543), .ZN(n2634) );
  MUX2_X1 U3373 ( .A(n2634), .B(DATAI_16_), .S(n3723), .Z(n4261) );
  INV_X1 U3374 ( .A(n4261), .ZN(n2924) );
  OAI22_X1 U3375 ( .A1(n4237), .A2(n2808), .B1(n2924), .B2(n2807), .ZN(n2635)
         );
  XNOR2_X1 U3376 ( .A(n2635), .B(n2398), .ZN(n2643) );
  OAI22_X1 U3377 ( .A1(n4237), .A2(n2805), .B1(n2924), .B2(n2794), .ZN(n2644)
         );
  INV_X1 U3378 ( .A(n2644), .ZN(n2636) );
  NAND2_X1 U3379 ( .A1(n2643), .A2(n2636), .ZN(n3615) );
  INV_X1 U3380 ( .A(n2637), .ZN(n2640) );
  INV_X1 U3381 ( .A(n2638), .ZN(n2639) );
  NAND2_X1 U3382 ( .A1(n2640), .A2(n2639), .ZN(n3567) );
  OAI211_X1 U3383 ( .C1(n2642), .C2(n3612), .A(n3615), .B(n3567), .ZN(n2641)
         );
  INV_X1 U3384 ( .A(n2642), .ZN(n3701) );
  INV_X1 U3385 ( .A(n3612), .ZN(n2646) );
  INV_X1 U3386 ( .A(n2643), .ZN(n2645) );
  NAND2_X1 U3387 ( .A1(n2645), .A2(n2644), .ZN(n3614) );
  OAI21_X1 U3388 ( .B1(n3701), .B2(n2646), .A(n3614), .ZN(n2647) );
  XNOR2_X1 U3389 ( .A(n2664), .B(REG3_REG_17__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U3390 ( .A1(n4245), .A2(n2002), .ZN(n2653) );
  INV_X1 U3391 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U3392 ( .A1(n3719), .A2(REG0_REG_17__SCAN_IN), .ZN(n2649) );
  INV_X1 U3393 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4367) );
  OR2_X1 U3394 ( .A1(n2443), .A2(n4367), .ZN(n2648) );
  OAI211_X1 U3395 ( .C1(n2650), .C2(n3722), .A(n2649), .B(n2648), .ZN(n2651)
         );
  INV_X1 U3396 ( .A(n2651), .ZN(n2652) );
  NAND2_X1 U3397 ( .A1(n2655), .A2(IR_REG_31__SCAN_IN), .ZN(n2656) );
  MUX2_X1 U3398 ( .A(IR_REG_31__SCAN_IN), .B(n2656), .S(IR_REG_17__SCAN_IN), 
        .Z(n2657) );
  AND2_X1 U3399 ( .A1(n2657), .A2(n2012), .ZN(n3985) );
  INV_X1 U3400 ( .A(DATAI_17_), .ZN(n2658) );
  MUX2_X1 U3401 ( .A(n4542), .B(n2658), .S(n3723), .Z(n4244) );
  OAI22_X1 U3402 ( .A1(n4265), .A2(n2808), .B1(n4244), .B2(n2807), .ZN(n2659)
         );
  XNOR2_X1 U3403 ( .A(n2659), .B(n2792), .ZN(n2661) );
  OAI22_X1 U3404 ( .A1(n4265), .A2(n2805), .B1(n4244), .B2(n2794), .ZN(n2660)
         );
  NAND2_X1 U3405 ( .A1(n2661), .A2(n2660), .ZN(n3636) );
  INV_X1 U3406 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4623) );
  INV_X1 U3407 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2662) );
  OAI21_X1 U3408 ( .B1(n2664), .B2(n4623), .A(n2662), .ZN(n2665) );
  NAND2_X1 U3409 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2663) );
  AND2_X1 U3410 ( .A1(n2665), .A2(n2678), .ZN(n4227) );
  NAND2_X1 U3411 ( .A1(n4227), .A2(n2002), .ZN(n2670) );
  INV_X1 U3412 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U3413 ( .A1(n2349), .A2(REG2_REG_18__SCAN_IN), .ZN(n2667) );
  INV_X1 U3414 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3973) );
  OR2_X1 U3415 ( .A1(n2443), .A2(n3973), .ZN(n2666) );
  OAI211_X1 U3416 ( .C1(n2442), .C2(n4641), .A(n2667), .B(n2666), .ZN(n2668)
         );
  INV_X1 U3417 ( .A(n2668), .ZN(n2669) );
  NAND2_X1 U3418 ( .A1(n2012), .A2(IR_REG_31__SCAN_IN), .ZN(n2671) );
  XNOR2_X1 U3419 ( .A(n2671), .B(IR_REG_18__SCAN_IN), .ZN(n4540) );
  INV_X1 U3420 ( .A(n4540), .ZN(n4513) );
  INV_X1 U3421 ( .A(DATAI_18_), .ZN(n2672) );
  MUX2_X1 U3422 ( .A(n4513), .B(n2672), .S(n3717), .Z(n3680) );
  INV_X1 U3423 ( .A(n3680), .ZN(n4225) );
  AOI22_X1 U3424 ( .A1(n4239), .A2(n2796), .B1(n2858), .B2(n4225), .ZN(n2674)
         );
  INV_X1 U3425 ( .A(n4239), .ZN(n4202) );
  OAI22_X1 U3426 ( .A1(n4202), .A2(n2808), .B1(n2807), .B2(n3680), .ZN(n2673)
         );
  XOR2_X1 U3427 ( .A(n2792), .B(n2673), .Z(n3675) );
  INV_X1 U3428 ( .A(n3675), .ZN(n2675) );
  INV_X1 U3429 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3430 ( .A1(n2678), .A2(n2677), .ZN(n2679) );
  NAND2_X1 U3431 ( .A1(n2690), .A2(n2679), .ZN(n4210) );
  INV_X1 U3432 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U3433 ( .A1(n2349), .A2(REG2_REG_19__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3434 ( .A1(n2850), .A2(REG1_REG_19__SCAN_IN), .ZN(n2680) );
  OAI211_X1 U3435 ( .C1(n2442), .C2(n4640), .A(n2681), .B(n2680), .ZN(n2682)
         );
  INV_X1 U3436 ( .A(n2682), .ZN(n2683) );
  MUX2_X1 U3437 ( .A(n3978), .B(DATAI_19_), .S(n3717), .Z(n3580) );
  OAI22_X1 U3438 ( .A1(n2967), .A2(n2808), .B1(n4207), .B2(n2807), .ZN(n2685)
         );
  XNOR2_X1 U3439 ( .A(n2685), .B(n2792), .ZN(n2687) );
  OAI22_X1 U3440 ( .A1(n2967), .A2(n2805), .B1(n4207), .B2(n2794), .ZN(n2686)
         );
  NOR2_X1 U3441 ( .A1(n2687), .A2(n2686), .ZN(n2688) );
  AOI21_X1 U3442 ( .B1(n2687), .B2(n2686), .A(n2688), .ZN(n3579) );
  NAND2_X1 U3443 ( .A1(n3577), .A2(n3579), .ZN(n3578) );
  INV_X1 U3444 ( .A(n2688), .ZN(n2689) );
  NAND2_X1 U3445 ( .A1(n3578), .A2(n2689), .ZN(n3006) );
  INV_X1 U3446 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3011) );
  NAND2_X1 U3447 ( .A1(n2690), .A2(n3011), .ZN(n2691) );
  NAND2_X1 U3448 ( .A1(n2707), .A2(n2691), .ZN(n4187) );
  INV_X1 U3449 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U3450 ( .A1(n3719), .A2(REG0_REG_20__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3451 ( .A1(n2850), .A2(REG1_REG_20__SCAN_IN), .ZN(n2692) );
  OAI211_X1 U3452 ( .C1(n4188), .C2(n3722), .A(n2693), .B(n2692), .ZN(n2694)
         );
  INV_X1 U3453 ( .A(n2694), .ZN(n2695) );
  NAND2_X1 U3454 ( .A1(n4204), .A2(n2858), .ZN(n2698) );
  NAND2_X1 U3455 ( .A1(n2339), .A2(n4177), .ZN(n2697) );
  NAND2_X1 U3456 ( .A1(n2698), .A2(n2697), .ZN(n2699) );
  XNOR2_X1 U3457 ( .A(n2699), .B(n2792), .ZN(n2702) );
  NAND2_X1 U34580 ( .A1(n4204), .A2(n2796), .ZN(n2701) );
  NAND2_X1 U34590 ( .A1(n2858), .A2(n4177), .ZN(n2700) );
  NAND2_X1 U3460 ( .A1(n2701), .A2(n2700), .ZN(n2703) );
  NAND2_X1 U3461 ( .A1(n2702), .A2(n2703), .ZN(n3589) );
  NAND2_X1 U3462 ( .A1(n3006), .A2(n3589), .ZN(n3005) );
  INV_X1 U3463 ( .A(n2702), .ZN(n2705) );
  INV_X1 U3464 ( .A(n2703), .ZN(n2704) );
  NAND2_X1 U3465 ( .A1(n2705), .A2(n2704), .ZN(n3588) );
  INV_X1 U3466 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U34670 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  NAND2_X1 U3468 ( .A1(n4166), .A2(n2002), .ZN(n2714) );
  INV_X1 U34690 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3470 ( .A1(n3719), .A2(REG0_REG_21__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U34710 ( .A1(n2850), .A2(REG1_REG_21__SCAN_IN), .ZN(n2709) );
  OAI211_X1 U3472 ( .C1(n2711), .C2(n3722), .A(n2710), .B(n2709), .ZN(n2712)
         );
  INV_X1 U34730 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3474 ( .A1(n3723), .A2(DATAI_21_), .ZN(n2971) );
  OAI22_X1 U34750 ( .A1(n4179), .A2(n2808), .B1(n2971), .B2(n2807), .ZN(n2715)
         );
  XNOR2_X1 U3476 ( .A(n2715), .B(n2792), .ZN(n2717) );
  OAI22_X1 U34770 ( .A1(n4179), .A2(n2805), .B1(n2971), .B2(n2808), .ZN(n2716)
         );
  NAND2_X1 U3478 ( .A1(n2717), .A2(n2716), .ZN(n3587) );
  XNOR2_X1 U34790 ( .A(n2726), .B(REG3_REG_22__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U3480 ( .A1(n4150), .A2(n2002), .ZN(n2722) );
  INV_X1 U34810 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U3482 ( .A1(n3719), .A2(REG0_REG_22__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U34830 ( .A1(n2349), .A2(REG2_REG_22__SCAN_IN), .ZN(n2718) );
  OAI211_X1 U3484 ( .C1(n2443), .C2(n4717), .A(n2719), .B(n2718), .ZN(n2720)
         );
  INV_X1 U34850 ( .A(n2720), .ZN(n2721) );
  OAI22_X1 U3486 ( .A1(n4162), .A2(n2808), .B1(n4151), .B2(n2807), .ZN(n2723)
         );
  XNOR2_X1 U34870 ( .A(n2723), .B(n2792), .ZN(n2735) );
  OAI22_X1 U3488 ( .A1(n4162), .A2(n2805), .B1(n4151), .B2(n2794), .ZN(n2734)
         );
  XNOR2_X1 U34890 ( .A(n2735), .B(n2734), .ZN(n3667) );
  AND2_X1 U3490 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2724) );
  INV_X1 U34910 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3668) );
  INV_X1 U3492 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3021) );
  OAI21_X1 U34930 ( .B1(n2726), .B2(n3668), .A(n3021), .ZN(n2727) );
  NAND2_X1 U3494 ( .A1(n2740), .A2(n2727), .ZN(n4133) );
  INV_X1 U34950 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U3496 ( .A1(n3719), .A2(REG0_REG_23__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U34970 ( .A1(n2349), .A2(REG2_REG_23__SCAN_IN), .ZN(n2728) );
  OAI211_X1 U3498 ( .C1(n2443), .C2(n4715), .A(n2729), .B(n2728), .ZN(n2730)
         );
  INV_X1 U34990 ( .A(n2730), .ZN(n2731) );
  NAND2_X1 U3500 ( .A1(n3723), .A2(DATAI_23_), .ZN(n4123) );
  OAI22_X1 U35010 ( .A1(n4147), .A2(n2805), .B1(n4123), .B2(n2808), .ZN(n2737)
         );
  OAI22_X1 U3502 ( .A1(n4147), .A2(n2808), .B1(n4123), .B2(n2807), .ZN(n2733)
         );
  XNOR2_X1 U35030 ( .A(n2733), .B(n2792), .ZN(n2738) );
  XOR2_X1 U3504 ( .A(n2737), .B(n2738), .Z(n3017) );
  OR2_X1 U35050 ( .A1(n2735), .A2(n2734), .ZN(n3018) );
  NAND2_X1 U35060 ( .A1(n2738), .A2(n2737), .ZN(n3538) );
  INV_X1 U35070 ( .A(n3538), .ZN(n2749) );
  INV_X1 U35080 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U35090 ( .A1(n2740), .A2(n4612), .ZN(n2741) );
  NAND2_X1 U35100 ( .A1(n2770), .A2(n2741), .ZN(n4108) );
  INV_X1 U35110 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4107) );
  NAND2_X1 U35120 ( .A1(n3719), .A2(REG0_REG_24__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U35130 ( .A1(n2850), .A2(REG1_REG_24__SCAN_IN), .ZN(n2742) );
  OAI211_X1 U35140 ( .C1(n4107), .C2(n3722), .A(n2743), .B(n2742), .ZN(n2744)
         );
  INV_X1 U35150 ( .A(n2744), .ZN(n2745) );
  NAND2_X1 U35160 ( .A1(n3717), .A2(DATAI_24_), .ZN(n4110) );
  OAI22_X1 U35170 ( .A1(n4124), .A2(n2808), .B1(n4110), .B2(n2807), .ZN(n2747)
         );
  XNOR2_X1 U35180 ( .A(n2747), .B(n2792), .ZN(n3646) );
  NOR2_X1 U35190 ( .A1(n2794), .A2(n4110), .ZN(n2748) );
  AOI21_X1 U35200 ( .B1(n4084), .B2(n2796), .A(n2748), .ZN(n3537) );
  NAND2_X1 U35210 ( .A1(n3538), .A2(n3537), .ZN(n3535) );
  OAI21_X1 U35220 ( .B1(n2749), .B2(n3646), .A(n3535), .ZN(n2759) );
  XNOR2_X1 U35230 ( .A(n2770), .B(REG3_REG_25__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U35240 ( .A1(n4091), .A2(n2002), .ZN(n2755) );
  INV_X1 U35250 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U35260 ( .A1(n3719), .A2(REG0_REG_25__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U35270 ( .A1(n2850), .A2(REG1_REG_25__SCAN_IN), .ZN(n2750) );
  OAI211_X1 U35280 ( .C1(n2752), .C2(n3722), .A(n2751), .B(n2750), .ZN(n2753)
         );
  INV_X1 U35290 ( .A(n2753), .ZN(n2754) );
  NAND2_X1 U35300 ( .A1(n4066), .A2(n2858), .ZN(n2757) );
  NAND2_X1 U35310 ( .A1(n2339), .A2(n4088), .ZN(n2756) );
  NAND2_X1 U35320 ( .A1(n2757), .A2(n2756), .ZN(n2758) );
  XNOR2_X1 U35330 ( .A(n2758), .B(n2792), .ZN(n3542) );
  INV_X1 U35340 ( .A(n4066), .ZN(n4106) );
  INV_X1 U35350 ( .A(n4088), .ZN(n3546) );
  OAI22_X1 U35360 ( .A1(n4106), .A2(n2805), .B1(n2794), .B2(n3546), .ZN(n3541)
         );
  NAND2_X1 U35370 ( .A1(n3542), .A2(n3541), .ZN(n3540) );
  NAND2_X1 U35380 ( .A1(n3539), .A2(n2760), .ZN(n2767) );
  INV_X1 U35390 ( .A(n3646), .ZN(n2763) );
  INV_X1 U35400 ( .A(n3541), .ZN(n2762) );
  AOI21_X1 U35410 ( .B1(n2763), .B2(n3537), .A(n2762), .ZN(n2761) );
  NAND3_X1 U35420 ( .A1(n2763), .A2(n3537), .A3(n2762), .ZN(n2764) );
  NAND2_X1 U35430 ( .A1(n2767), .A2(n2766), .ZN(n3684) );
  INV_X1 U35440 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3545) );
  INV_X1 U35450 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2768) );
  OAI21_X1 U35460 ( .B1(n2770), .B2(n3545), .A(n2768), .ZN(n2771) );
  NAND2_X1 U35470 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2769) );
  NAND2_X1 U35480 ( .A1(n4073), .A2(n2002), .ZN(n2776) );
  INV_X1 U35490 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4687) );
  NAND2_X1 U35500 ( .A1(n3719), .A2(REG0_REG_26__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U35510 ( .A1(n2850), .A2(REG1_REG_26__SCAN_IN), .ZN(n2772) );
  OAI211_X1 U35520 ( .C1(n4687), .C2(n3722), .A(n2773), .B(n2772), .ZN(n2774)
         );
  INV_X1 U35530 ( .A(n2774), .ZN(n2775) );
  NAND2_X1 U35540 ( .A1(n3723), .A2(DATAI_26_), .ZN(n4069) );
  OAI22_X1 U35550 ( .A1(n4087), .A2(n2808), .B1(n2807), .B2(n4069), .ZN(n2777)
         );
  XNOR2_X1 U35560 ( .A(n2777), .B(n2792), .ZN(n2779) );
  OAI22_X1 U35570 ( .A1(n4087), .A2(n2805), .B1(n2794), .B2(n4069), .ZN(n2778)
         );
  NAND2_X1 U35580 ( .A1(n2779), .A2(n2778), .ZN(n3686) );
  NOR2_X1 U35590 ( .A1(n2779), .A2(n2778), .ZN(n3685) );
  AOI21_X2 U35600 ( .B1(n3684), .B2(n3686), .A(n3685), .ZN(n3560) );
  INV_X1 U35610 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2781) );
  NAND2_X1 U35620 ( .A1(n2782), .A2(n2781), .ZN(n2783) );
  NAND2_X1 U35630 ( .A1(n2797), .A2(n2783), .ZN(n4046) );
  INV_X1 U35640 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U35650 ( .A1(n3719), .A2(REG0_REG_27__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U35660 ( .A1(n2349), .A2(REG2_REG_27__SCAN_IN), .ZN(n2785) );
  OAI211_X1 U35670 ( .C1(n2443), .C2(n4714), .A(n2786), .B(n2785), .ZN(n2787)
         );
  INV_X1 U35680 ( .A(n2787), .ZN(n2788) );
  NAND2_X1 U35690 ( .A1(n4065), .A2(n2858), .ZN(n2791) );
  AND2_X1 U35700 ( .A1(n3717), .A2(DATAI_27_), .ZN(n2976) );
  NAND2_X1 U35710 ( .A1(n2339), .A2(n2976), .ZN(n2790) );
  NAND2_X1 U35720 ( .A1(n2791), .A2(n2790), .ZN(n2793) );
  XNOR2_X1 U35730 ( .A(n2793), .B(n2792), .ZN(n2845) );
  NOR2_X1 U35740 ( .A1(n4048), .A2(n2794), .ZN(n2795) );
  AOI21_X1 U35750 ( .B1(n4065), .B2(n2796), .A(n2795), .ZN(n2843) );
  XNOR2_X1 U35760 ( .A(n2845), .B(n2843), .ZN(n3559) );
  NAND2_X1 U35770 ( .A1(n3560), .A2(n3559), .ZN(n2885) );
  INV_X1 U35780 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U35790 ( .A1(n2797), .A2(n2848), .ZN(n2798) );
  NAND2_X1 U35800 ( .A1(n3552), .A2(n2002), .ZN(n2804) );
  INV_X1 U35810 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U3582 ( .A1(n3719), .A2(REG0_REG_28__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U3583 ( .A1(n2349), .A2(REG2_REG_28__SCAN_IN), .ZN(n2799) );
  OAI211_X1 U3584 ( .C1(n2801), .C2(n2443), .A(n2800), .B(n2799), .ZN(n2802)
         );
  INV_X1 U3585 ( .A(n2802), .ZN(n2803) );
  AND2_X1 U3586 ( .A1(n3717), .A2(DATAI_28_), .ZN(n4013) );
  INV_X1 U3587 ( .A(n4013), .ZN(n2983) );
  OAI22_X1 U3588 ( .A1(n4041), .A2(n2805), .B1(n2808), .B2(n2983), .ZN(n2806)
         );
  XNOR2_X1 U3589 ( .A(n2806), .B(n2398), .ZN(n2810) );
  OAI22_X1 U3590 ( .A1(n4041), .A2(n2808), .B1(n2807), .B2(n2983), .ZN(n2809)
         );
  XNOR2_X1 U3591 ( .A(n2810), .B(n2809), .ZN(n2847) );
  INV_X1 U3592 ( .A(n2847), .ZN(n2842) );
  NAND2_X1 U3593 ( .A1(n2836), .A2(n2835), .ZN(n2813) );
  NAND2_X1 U3594 ( .A1(n2813), .A2(IR_REG_31__SCAN_IN), .ZN(n2815) );
  INV_X1 U3595 ( .A(n4455), .ZN(n2831) );
  NAND3_X1 U3596 ( .A1(n2819), .A2(B_REG_SCAN_IN), .A3(n2831), .ZN(n2818) );
  INV_X1 U3597 ( .A(n2819), .ZN(n4456) );
  INV_X1 U3598 ( .A(B_REG_SCAN_IN), .ZN(n2816) );
  NAND2_X1 U3599 ( .A1(n4456), .A2(n2816), .ZN(n2817) );
  INV_X1 U3600 ( .A(n3053), .ZN(n2820) );
  INV_X1 U3601 ( .A(D_REG_0__SCAN_IN), .ZN(n3055) );
  INV_X1 U3602 ( .A(n4454), .ZN(n2832) );
  INV_X1 U3603 ( .A(D_REG_2__SCAN_IN), .ZN(n4638) );
  INV_X1 U3604 ( .A(D_REG_12__SCAN_IN), .ZN(n4635) );
  INV_X1 U3605 ( .A(D_REG_27__SCAN_IN), .ZN(n4653) );
  INV_X1 U3606 ( .A(D_REG_25__SCAN_IN), .ZN(n4656) );
  NAND4_X1 U3607 ( .A1(n4638), .A2(n4635), .A3(n4653), .A4(n4656), .ZN(n2821)
         );
  NOR3_X1 U3608 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(n2821), 
        .ZN(n4605) );
  NOR4_X1 U3609 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2823) );
  NOR4_X1 U3610 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2822) );
  NAND3_X1 U3611 ( .A1(n4605), .A2(n2823), .A3(n2822), .ZN(n2829) );
  NOR4_X1 U3612 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2827) );
  NOR4_X1 U3613 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2826) );
  NOR4_X1 U3614 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2825) );
  NOR4_X1 U3615 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2824) );
  NAND4_X1 U3616 ( .A1(n2827), .A2(n2826), .A3(n2825), .A4(n2824), .ZN(n2828)
         );
  NOR2_X1 U3617 ( .A1(n2829), .A2(n2828), .ZN(n2988) );
  AND2_X1 U3618 ( .A1(n2988), .A2(D_REG_1__SCAN_IN), .ZN(n2830) );
  OR2_X1 U3619 ( .A1(n3053), .A2(n2830), .ZN(n2833) );
  NAND2_X1 U3620 ( .A1(n2832), .A2(n2831), .ZN(n3056) );
  NAND2_X1 U3621 ( .A1(n2833), .A2(n3056), .ZN(n3219) );
  INV_X1 U3622 ( .A(n3219), .ZN(n2834) );
  NAND2_X1 U3623 ( .A1(n2838), .A2(n2839), .ZN(n2980) );
  OAI211_X1 U3624 ( .C1(n2837), .C2(n4526), .A(n4278), .B(n2980), .ZN(n2869)
         );
  INV_X1 U3625 ( .A(n2869), .ZN(n2840) );
  AND2_X1 U3626 ( .A1(n3058), .A2(n2840), .ZN(n2841) );
  NAND2_X1 U3627 ( .A1(n2842), .A2(n3623), .ZN(n2884) );
  INV_X1 U3628 ( .A(n2843), .ZN(n2844) );
  NAND2_X1 U3629 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  NAND2_X1 U3630 ( .A1(n2885), .A2(n2293), .ZN(n2883) );
  NOR2_X1 U3631 ( .A1(n2847), .A2(n2846), .ZN(n2881) );
  NOR2_X1 U3632 ( .A1(n2848), .A2(STATE_REG_SCAN_IN), .ZN(n2880) );
  INV_X1 U3633 ( .A(n4025), .ZN(n2849) );
  NAND2_X1 U3634 ( .A1(n2849), .A2(n2002), .ZN(n2855) );
  INV_X1 U3635 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U3636 ( .A1(n2850), .A2(REG1_REG_29__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U3637 ( .A1(n2349), .A2(REG2_REG_29__SCAN_IN), .ZN(n2851) );
  OAI211_X1 U3638 ( .C1(n2442), .C2(n4724), .A(n2852), .B(n2851), .ZN(n2853)
         );
  INV_X1 U3639 ( .A(n2853), .ZN(n2854) );
  INV_X1 U3640 ( .A(n3872), .ZN(n2878) );
  INV_X1 U3641 ( .A(n2856), .ZN(n2857) );
  NAND3_X1 U3642 ( .A1(n4539), .A2(n2858), .A3(n2857), .ZN(n3867) );
  OAI21_X1 U3643 ( .B1(n2859), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2860) );
  MUX2_X1 U3644 ( .A(IR_REG_31__SCAN_IN), .B(n2860), .S(IR_REG_28__SCAN_IN), 
        .Z(n2862) );
  NAND2_X1 U3645 ( .A1(n2862), .A2(n2861), .ZN(n3087) );
  NOR2_X1 U3646 ( .A1(n3867), .A2(n3119), .ZN(n2863) );
  INV_X1 U3647 ( .A(n3707), .ZN(n3669) );
  NOR2_X1 U3648 ( .A1(n3867), .A2(n3087), .ZN(n2864) );
  AND2_X1 U3649 ( .A1(n3058), .A2(n4525), .ZN(n2865) );
  NAND2_X1 U3650 ( .A1(n2868), .A2(n2865), .ZN(n2867) );
  NAND2_X1 U3651 ( .A1(n2367), .A2(n3978), .ZN(n2866) );
  NOR2_X1 U3652 ( .A1(n4551), .A2(n2839), .ZN(n2987) );
  AOI22_X1 U3653 ( .A1(n4065), .A2(n3695), .B1(n4013), .B2(n3629), .ZN(n2877)
         );
  INV_X1 U3654 ( .A(n2868), .ZN(n2874) );
  NAND2_X1 U3655 ( .A1(n2869), .A2(n4278), .ZN(n2870) );
  NAND2_X1 U3656 ( .A1(n2874), .A2(n2870), .ZN(n3135) );
  AND2_X1 U3657 ( .A1(n2367), .A2(n4526), .ZN(n2871) );
  OR2_X1 U3658 ( .A1(n2980), .A2(n2871), .ZN(n2986) );
  NAND4_X1 U3659 ( .A1(n3135), .A2(n2986), .A3(n3062), .A4(n2378), .ZN(n2872)
         );
  NAND2_X1 U3660 ( .A1(n2872), .A2(STATE_REG_SCAN_IN), .ZN(n2875) );
  INV_X1 U3661 ( .A(n3867), .ZN(n2873) );
  NAND2_X1 U3662 ( .A1(n2874), .A2(n2873), .ZN(n3136) );
  NAND2_X1 U3663 ( .A1(n3552), .A2(n3708), .ZN(n2876) );
  OAI211_X1 U3664 ( .C1(n2878), .C2(n3669), .A(n2877), .B(n2876), .ZN(n2879)
         );
  AOI211_X1 U3665 ( .C1(n2881), .C2(n3623), .A(n2880), .B(n2879), .ZN(n2882)
         );
  OAI211_X1 U3666 ( .C1(n2885), .C2(n2884), .A(n2883), .B(n2882), .ZN(U3217)
         );
  NAND2_X1 U3667 ( .A1(n2886), .A2(n2898), .ZN(n3809) );
  INV_X1 U3668 ( .A(n3214), .ZN(n2889) );
  NOR2_X1 U3669 ( .A1(n3764), .A2(n2889), .ZN(n2892) );
  NAND2_X1 U3670 ( .A1(n3194), .A2(n3238), .ZN(n3213) );
  INV_X1 U3671 ( .A(n3179), .ZN(n3175) );
  NAND2_X1 U3672 ( .A1(n3175), .A2(n2896), .ZN(n3211) );
  INV_X1 U3673 ( .A(n3211), .ZN(n2890) );
  NAND2_X1 U3674 ( .A1(n3270), .A2(n2894), .ZN(n2895) );
  NAND2_X1 U3675 ( .A1(n3883), .A2(n3175), .ZN(n3803) );
  NAND2_X1 U3676 ( .A1(n3179), .A2(n2896), .ZN(n3800) );
  NAND2_X1 U3677 ( .A1(n3312), .A2(n2949), .ZN(n2900) );
  NAND2_X1 U3678 ( .A1(n3628), .A2(n3882), .ZN(n2901) );
  NAND2_X1 U3679 ( .A1(n2902), .A2(n2901), .ZN(n3183) );
  INV_X1 U3680 ( .A(n3369), .ZN(n3399) );
  NAND2_X1 U3681 ( .A1(n3399), .A2(n2904), .ZN(n2951) );
  NAND2_X1 U3682 ( .A1(n3183), .A2(n2903), .ZN(n2908) );
  NAND2_X1 U3683 ( .A1(n2908), .A2(n2907), .ZN(n3297) );
  NAND2_X1 U3684 ( .A1(n3297), .A2(n2297), .ZN(n2910) );
  INV_X1 U3685 ( .A(n3389), .ZN(n2953) );
  NAND2_X1 U3686 ( .A1(n3389), .A2(n3880), .ZN(n2909) );
  NAND2_X1 U3687 ( .A1(n2910), .A2(n2909), .ZN(n3352) );
  OAI21_X1 U3688 ( .B1(n3352), .B2(n2296), .A(n2911), .ZN(n2912) );
  INV_X1 U3689 ( .A(n2912), .ZN(n3411) );
  NAND2_X1 U3690 ( .A1(n2169), .A2(n2913), .ZN(n2914) );
  NAND2_X1 U3691 ( .A1(n3411), .A2(n2914), .ZN(n2916) );
  NAND2_X1 U3692 ( .A1(n4300), .A2(n3878), .ZN(n3467) );
  INV_X1 U3693 ( .A(n4300), .ZN(n4296) );
  NAND2_X1 U3694 ( .A1(n4296), .A2(n3469), .ZN(n3466) );
  NAND2_X1 U3695 ( .A1(n4300), .A2(n3469), .ZN(n2919) );
  NAND2_X1 U3696 ( .A1(n3603), .A2(n3877), .ZN(n2920) );
  NAND2_X1 U3697 ( .A1(n3522), .A2(n3659), .ZN(n2921) );
  NAND2_X1 U3698 ( .A1(n3705), .A2(n3525), .ZN(n3729) );
  NAND2_X1 U3699 ( .A1(n4271), .A2(n3572), .ZN(n3726) );
  NAND2_X1 U3700 ( .A1(n3528), .A2(n2150), .ZN(n3529) );
  NAND2_X1 U3701 ( .A1(n3705), .A2(n3572), .ZN(n2922) );
  NAND2_X1 U3702 ( .A1(n3529), .A2(n2922), .ZN(n4268) );
  NAND2_X1 U3703 ( .A1(n4262), .A2(n4279), .ZN(n2923) );
  NAND2_X1 U3704 ( .A1(n4237), .A2(n4261), .ZN(n3836) );
  NAND2_X1 U3705 ( .A1(n4274), .A2(n2924), .ZN(n3833) );
  NAND2_X1 U3706 ( .A1(n3836), .A2(n3833), .ZN(n4251) );
  NAND2_X1 U3707 ( .A1(n4274), .A2(n4261), .ZN(n2925) );
  NAND2_X1 U3708 ( .A1(n4265), .A2(n4244), .ZN(n2926) );
  OR2_X1 U3709 ( .A1(n4239), .A2(n3680), .ZN(n4197) );
  NAND2_X1 U3710 ( .A1(n4239), .A2(n3680), .ZN(n4198) );
  NAND2_X1 U3711 ( .A1(n2928), .A2(n2927), .ZN(n4221) );
  NAND2_X1 U3712 ( .A1(n4202), .A2(n3680), .ZN(n2929) );
  NAND2_X1 U3713 ( .A1(n4221), .A2(n2929), .ZN(n4194) );
  NAND2_X1 U3714 ( .A1(n4216), .A2(n3580), .ZN(n2930) );
  NAND2_X1 U3715 ( .A1(n4194), .A2(n2930), .ZN(n2932) );
  NAND2_X1 U3716 ( .A1(n2967), .A2(n4207), .ZN(n2931) );
  NOR2_X1 U3717 ( .A1(n4204), .A2(n4177), .ZN(n2934) );
  NAND2_X1 U3718 ( .A1(n4204), .A2(n4177), .ZN(n2933) );
  NOR2_X1 U3719 ( .A1(n4179), .A2(n2971), .ZN(n2935) );
  NAND2_X1 U3720 ( .A1(n4162), .A2(n4144), .ZN(n4120) );
  NAND2_X1 U3721 ( .A1(n3874), .A2(n4151), .ZN(n2970) );
  NAND2_X1 U3722 ( .A1(n4147), .A2(n4123), .ZN(n2936) );
  NAND2_X1 U3723 ( .A1(n4103), .A2(n4130), .ZN(n2937) );
  NOR2_X1 U3724 ( .A1(n4124), .A2(n4110), .ZN(n2940) );
  NAND2_X1 U3725 ( .A1(n4124), .A2(n4110), .ZN(n2939) );
  NOR2_X1 U3726 ( .A1(n4066), .A2(n4088), .ZN(n2942) );
  NAND2_X1 U3727 ( .A1(n4066), .A2(n4088), .ZN(n2941) );
  INV_X1 U3728 ( .A(n4069), .ZN(n2974) );
  NOR2_X1 U3729 ( .A1(n4065), .A2(n2976), .ZN(n2944) );
  NAND2_X1 U3730 ( .A1(n4065), .A2(n2976), .ZN(n2943) );
  NAND2_X1 U3731 ( .A1(n4041), .A2(n4013), .ZN(n3716) );
  NAND2_X1 U3732 ( .A1(n4014), .A2(n2983), .ZN(n4016) );
  NAND2_X1 U3733 ( .A1(n3716), .A2(n4016), .ZN(n4011) );
  XNOR2_X1 U3734 ( .A(n2364), .B(n2838), .ZN(n2945) );
  NAND2_X1 U3735 ( .A1(n2945), .A2(n4526), .ZN(n4528) );
  AND2_X1 U3736 ( .A1(n3267), .A2(n3159), .ZN(n3798) );
  NAND2_X1 U3737 ( .A1(n2946), .A2(n3799), .ZN(n3171) );
  INV_X1 U3738 ( .A(n3169), .ZN(n3758) );
  NAND2_X1 U3739 ( .A1(n3171), .A2(n3758), .ZN(n3170) );
  NAND2_X1 U3740 ( .A1(n3170), .A2(n3800), .ZN(n3283) );
  NAND2_X1 U3741 ( .A1(n3194), .A2(n2947), .ZN(n3805) );
  NAND2_X1 U3742 ( .A1(n3289), .A2(n3238), .ZN(n3802) );
  NAND2_X1 U3743 ( .A1(n3283), .A2(n3757), .ZN(n2948) );
  NAND2_X1 U3744 ( .A1(n2948), .A2(n3805), .ZN(n3223) );
  AND2_X1 U3745 ( .A1(n3312), .A2(n3882), .ZN(n3309) );
  NAND2_X1 U3746 ( .A1(n3628), .A2(n2949), .ZN(n3812) );
  NAND2_X1 U3747 ( .A1(n3374), .A2(n3881), .ZN(n3811) );
  NAND2_X1 U3748 ( .A1(n3258), .A2(n2950), .ZN(n3814) );
  INV_X1 U3749 ( .A(n2951), .ZN(n2952) );
  NAND2_X1 U3750 ( .A1(n3389), .A2(n3354), .ZN(n3820) );
  NAND2_X1 U3751 ( .A1(n3298), .A2(n3820), .ZN(n2954) );
  NAND2_X1 U3752 ( .A1(n2953), .A2(n3880), .ZN(n3816) );
  AND2_X1 U3753 ( .A1(n2170), .A2(n3879), .ZN(n3824) );
  NAND2_X1 U3754 ( .A1(n3419), .A2(n2955), .ZN(n3821) );
  NAND2_X1 U3755 ( .A1(n2169), .A2(n3485), .ZN(n3826) );
  NAND2_X1 U3756 ( .A1(n3495), .A2(n2913), .ZN(n3823) );
  INV_X1 U3757 ( .A(n3603), .ZN(n2956) );
  NAND2_X1 U3758 ( .A1(n2956), .A2(n3877), .ZN(n3503) );
  NAND2_X1 U3759 ( .A1(n3659), .A2(n3876), .ZN(n2957) );
  NAND2_X1 U3760 ( .A1(n3503), .A2(n2957), .ZN(n2959) );
  INV_X1 U3761 ( .A(n3467), .ZN(n2958) );
  NOR2_X1 U3762 ( .A1(n2959), .A2(n2958), .ZN(n3827) );
  NAND2_X1 U3763 ( .A1(n4287), .A2(n3827), .ZN(n2963) );
  INV_X1 U3764 ( .A(n2959), .ZN(n2962) );
  NAND2_X1 U3765 ( .A1(n3603), .A2(n4289), .ZN(n3505) );
  NAND2_X1 U3766 ( .A1(n3466), .A2(n3505), .ZN(n2961) );
  NOR2_X1 U3767 ( .A1(n3659), .A2(n3876), .ZN(n2960) );
  AOI21_X1 U3768 ( .B1(n2962), .B2(n2961), .A(n2960), .ZN(n3830) );
  NAND2_X1 U3769 ( .A1(n2963), .A2(n3830), .ZN(n3521) );
  INV_X1 U3770 ( .A(n4262), .ZN(n3523) );
  NAND2_X1 U3771 ( .A1(n3523), .A2(n4279), .ZN(n3730) );
  NAND2_X1 U3772 ( .A1(n4262), .A2(n4277), .ZN(n3727) );
  INV_X1 U3773 ( .A(n4251), .ZN(n4259) );
  NAND2_X1 U3774 ( .A1(n4260), .A2(n4259), .ZN(n4258) );
  NAND2_X1 U3775 ( .A1(n4258), .A2(n3833), .ZN(n4236) );
  NAND2_X1 U3776 ( .A1(n4216), .A2(n4207), .ZN(n3769) );
  NAND2_X1 U3777 ( .A1(n3769), .A2(n4198), .ZN(n2964) );
  AND2_X1 U3778 ( .A1(n3677), .A2(n4244), .ZN(n4196) );
  OR2_X1 U3779 ( .A1(n2964), .A2(n4196), .ZN(n3736) );
  INV_X1 U3780 ( .A(n2964), .ZN(n2966) );
  OR2_X1 U3781 ( .A1(n3677), .A2(n4244), .ZN(n4195) );
  NAND2_X1 U3782 ( .A1(n4197), .A2(n4195), .ZN(n2965) );
  NAND2_X1 U3783 ( .A1(n2966), .A2(n2965), .ZN(n2968) );
  NAND2_X1 U3784 ( .A1(n2967), .A2(n3580), .ZN(n3770) );
  NAND2_X1 U3785 ( .A1(n2968), .A2(n3770), .ZN(n4172) );
  INV_X1 U3786 ( .A(n4177), .ZN(n4185) );
  NOR2_X1 U3787 ( .A1(n4204), .A2(n4185), .ZN(n2969) );
  NOR2_X1 U3788 ( .A1(n4172), .A2(n2969), .ZN(n3837) );
  NAND2_X1 U3789 ( .A1(n4204), .A2(n4185), .ZN(n3737) );
  OR2_X1 U3790 ( .A1(n4143), .A2(n2971), .ZN(n4118) );
  AND2_X1 U3791 ( .A1(n4120), .A2(n4118), .ZN(n3843) );
  NAND2_X1 U3792 ( .A1(n4103), .A2(n4123), .ZN(n3768) );
  AND2_X1 U3793 ( .A1(n3768), .A2(n2970), .ZN(n3847) );
  AND2_X1 U3794 ( .A1(n4143), .A2(n2971), .ZN(n4117) );
  NAND2_X1 U3795 ( .A1(n4120), .A2(n4117), .ZN(n2972) );
  NAND2_X1 U3796 ( .A1(n2973), .A2(n3740), .ZN(n4098) );
  INV_X1 U3797 ( .A(n4110), .ZN(n4102) );
  NAND2_X1 U3798 ( .A1(n4124), .A2(n4102), .ZN(n3756) );
  NAND2_X1 U3799 ( .A1(n4147), .A2(n4130), .ZN(n4097) );
  NAND2_X1 U3800 ( .A1(n4087), .A2(n2974), .ZN(n3754) );
  OR2_X1 U3801 ( .A1(n4066), .A2(n3546), .ZN(n4059) );
  NAND2_X1 U3802 ( .A1(n3754), .A2(n4059), .ZN(n3846) );
  INV_X1 U3803 ( .A(n3846), .ZN(n2975) );
  NAND2_X1 U3804 ( .A1(n4066), .A2(n3546), .ZN(n3753) );
  NAND2_X1 U3805 ( .A1(n4084), .A2(n4110), .ZN(n4079) );
  NAND2_X1 U3806 ( .A1(n3753), .A2(n4079), .ZN(n4058) );
  AOI21_X1 U3807 ( .B1(n2975), .B2(n4058), .A(n3725), .ZN(n3850) );
  INV_X1 U3808 ( .A(n4065), .ZN(n2977) );
  NAND2_X1 U3809 ( .A1(n2977), .A2(n2976), .ZN(n3715) );
  NAND2_X1 U3810 ( .A1(n4065), .A2(n4048), .ZN(n3849) );
  NAND2_X1 U3811 ( .A1(n3715), .A2(n3849), .ZN(n4045) );
  NAND2_X1 U3812 ( .A1(n4038), .A2(n3715), .ZN(n2978) );
  XNOR2_X1 U3813 ( .A(n2978), .B(n2094), .ZN(n2985) );
  NAND2_X1 U3814 ( .A1(n2838), .A2(n3978), .ZN(n2979) );
  INV_X1 U3815 ( .A(n2367), .ZN(n3047) );
  NAND2_X1 U3816 ( .A1(n3047), .A2(n2839), .ZN(n3750) );
  INV_X1 U3817 ( .A(n2980), .ZN(n3063) );
  NAND2_X1 U3818 ( .A1(n3872), .A2(n4273), .ZN(n2982) );
  NAND2_X1 U3819 ( .A1(n4065), .A2(n4272), .ZN(n2981) );
  OAI211_X1 U3820 ( .C1(n2983), .C2(n4278), .A(n2982), .B(n2981), .ZN(n2984)
         );
  INV_X1 U3821 ( .A(n3000), .ZN(n3221) );
  NAND2_X1 U3822 ( .A1(n3058), .A2(n2986), .ZN(n3218) );
  NOR2_X1 U3823 ( .A1(n3218), .A2(n2987), .ZN(n2991) );
  OAI21_X1 U3824 ( .B1(n3053), .B2(D_REG_1__SCAN_IN), .A(n3056), .ZN(n2990) );
  OR2_X1 U3825 ( .A1(n3053), .A2(n2988), .ZN(n2989) );
  MUX2_X1 U3826 ( .A(REG0_REG_28__SCAN_IN), .B(n3002), .S(n4739), .Z(n2992) );
  INV_X1 U3827 ( .A(n2992), .ZN(n2999) );
  NAND2_X1 U3828 ( .A1(n2993), .A2(n4576), .ZN(n3265) );
  NOR2_X2 U3829 ( .A1(n3265), .A2(n3179), .ZN(n3290) );
  NAND2_X1 U3830 ( .A1(n3370), .A2(n3369), .ZN(n3368) );
  NAND2_X1 U3831 ( .A1(n4050), .A2(n4013), .ZN(n2996) );
  NAND2_X1 U3832 ( .A1(n4028), .A2(n2996), .ZN(n3554) );
  NAND2_X1 U3833 ( .A1(n2999), .A2(n2300), .ZN(U3514) );
  INV_X1 U3834 ( .A(n3003), .ZN(n3004) );
  NAND2_X1 U3835 ( .A1(n3004), .A2(n2299), .ZN(U3546) );
  INV_X1 U3836 ( .A(n3005), .ZN(n3008) );
  AOI21_X1 U3837 ( .B1(n3589), .B2(n3588), .A(n3006), .ZN(n3007) );
  AOI21_X1 U3838 ( .B1(n3008), .B2(n3588), .A(n3007), .ZN(n3009) );
  NOR2_X1 U3839 ( .A1(n3009), .A2(n3711), .ZN(n3015) );
  NOR2_X1 U3840 ( .A1(n3689), .A2(n4187), .ZN(n3014) );
  NAND2_X1 U3841 ( .A1(n3695), .A2(n4216), .ZN(n3010) );
  OAI21_X1 U3842 ( .B1(STATE_REG_SCAN_IN), .B2(n3011), .A(n3010), .ZN(n3013)
         );
  OAI22_X1 U3843 ( .A1(n4179), .A2(n3669), .B1(n3703), .B2(n4185), .ZN(n3012)
         );
  OR4_X1 U3844 ( .A1(n3015), .A2(n3014), .A3(n3013), .A4(n3012), .ZN(U3230) );
  AND2_X2 U3845 ( .A1(n4539), .A2(n3016), .ZN(U4043) );
  INV_X2 U3846 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3847 ( .A(n3539), .ZN(n3020) );
  NOR3_X1 U3848 ( .A1(n3020), .A2(n3019), .A3(n3711), .ZN(n3025) );
  NOR2_X1 U3849 ( .A1(n3689), .A2(n4133), .ZN(n3024) );
  OAI22_X1 U3850 ( .A1(n4124), .A2(n3669), .B1(STATE_REG_SCAN_IN), .B2(n3021), 
        .ZN(n3023) );
  INV_X1 U3851 ( .A(n3695), .ZN(n3704) );
  OAI22_X1 U3852 ( .A1(n4162), .A2(n3704), .B1(n3703), .B2(n4123), .ZN(n3022)
         );
  OR4_X1 U3853 ( .A1(n3025), .A2(n3024), .A3(n3023), .A4(n3022), .ZN(U3213) );
  INV_X1 U3854 ( .A(DATAI_1_), .ZN(n3026) );
  MUX2_X1 U3855 ( .A(n3079), .B(n3026), .S(U3149), .Z(n3027) );
  INV_X1 U3856 ( .A(n3027), .ZN(U3351) );
  NAND3_X1 U3857 ( .A1(n3029), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3030) );
  INV_X1 U3858 ( .A(DATAI_31_), .ZN(n4685) );
  OAI22_X1 U3859 ( .A1(n3028), .A2(n3030), .B1(STATE_REG_SCAN_IN), .B2(n4685), 
        .ZN(U3321) );
  MUX2_X1 U3860 ( .A(n3031), .B(n3114), .S(STATE_REG_SCAN_IN), .Z(n3032) );
  INV_X1 U3861 ( .A(n3032), .ZN(U3348) );
  INV_X1 U3862 ( .A(n3934), .ZN(n3946) );
  NAND2_X1 U3863 ( .A1(n3946), .A2(STATE_REG_SCAN_IN), .ZN(n3033) );
  OAI21_X1 U3864 ( .B1(STATE_REG_SCAN_IN), .B2(n2587), .A(n3033), .ZN(U3339)
         );
  MUX2_X1 U3865 ( .A(n3107), .B(n2441), .S(U3149), .Z(n3034) );
  INV_X1 U3866 ( .A(n3034), .ZN(U3347) );
  INV_X1 U3867 ( .A(n3963), .ZN(n3949) );
  INV_X1 U3868 ( .A(DATAI_14_), .ZN(n3035) );
  MUX2_X1 U3869 ( .A(n3949), .B(n3035), .S(U3149), .Z(n3036) );
  INV_X1 U3870 ( .A(n3036), .ZN(U3338) );
  INV_X1 U3871 ( .A(DATAI_30_), .ZN(n4634) );
  NAND2_X1 U3872 ( .A1(n3037), .A2(STATE_REG_SCAN_IN), .ZN(n3038) );
  OAI21_X1 U3873 ( .B1(STATE_REG_SCAN_IN), .B2(n4634), .A(n3038), .ZN(U3322)
         );
  INV_X1 U3874 ( .A(DATAI_27_), .ZN(n3041) );
  XNOR2_X1 U3875 ( .A(n3039), .B(IR_REG_27__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U3876 ( .A1(n4467), .A2(STATE_REG_SCAN_IN), .ZN(n3040) );
  OAI21_X1 U3877 ( .B1(STATE_REG_SCAN_IN), .B2(n3041), .A(n3040), .ZN(U3325)
         );
  INV_X1 U3878 ( .A(DATAI_28_), .ZN(n3043) );
  NAND2_X1 U3879 ( .A1(n3119), .A2(STATE_REG_SCAN_IN), .ZN(n3042) );
  OAI21_X1 U3880 ( .B1(STATE_REG_SCAN_IN), .B2(n3043), .A(n3042), .ZN(U3324)
         );
  INV_X1 U3881 ( .A(DATAI_21_), .ZN(n3045) );
  NAND2_X1 U3882 ( .A1(n2839), .A2(STATE_REG_SCAN_IN), .ZN(n3044) );
  OAI21_X1 U3883 ( .B1(STATE_REG_SCAN_IN), .B2(n3045), .A(n3044), .ZN(U3331)
         );
  INV_X1 U3884 ( .A(DATAI_19_), .ZN(n4689) );
  MUX2_X1 U3885 ( .A(n4689), .B(n4526), .S(STATE_REG_SCAN_IN), .Z(n3046) );
  INV_X1 U3886 ( .A(n3046), .ZN(U3333) );
  INV_X1 U3887 ( .A(DATAI_20_), .ZN(n3049) );
  NAND2_X1 U3888 ( .A1(n3047), .A2(STATE_REG_SCAN_IN), .ZN(n3048) );
  OAI21_X1 U3889 ( .B1(STATE_REG_SCAN_IN), .B2(n3049), .A(n3048), .ZN(U3332)
         );
  INV_X1 U3890 ( .A(DATAI_22_), .ZN(n4684) );
  NAND2_X1 U3891 ( .A1(n2838), .A2(STATE_REG_SCAN_IN), .ZN(n3050) );
  OAI21_X1 U3892 ( .B1(STATE_REG_SCAN_IN), .B2(n4684), .A(n3050), .ZN(U3330)
         );
  INV_X1 U3893 ( .A(DATAI_12_), .ZN(n3051) );
  INV_X1 U3894 ( .A(n3912), .ZN(n3931) );
  MUX2_X1 U3895 ( .A(n3051), .B(n3931), .S(STATE_REG_SCAN_IN), .Z(n3052) );
  INV_X1 U3896 ( .A(n3052), .ZN(U3340) );
  AOI22_X1 U3897 ( .A1(n4537), .A2(n3055), .B1(n3054), .B2(n4539), .ZN(U3458)
         );
  INV_X1 U3898 ( .A(D_REG_1__SCAN_IN), .ZN(n4637) );
  INV_X1 U3899 ( .A(n3056), .ZN(n3057) );
  AOI22_X1 U3900 ( .A1(n4537), .A2(n4637), .B1(n3057), .B2(n4539), .ZN(U3459)
         );
  INV_X1 U3901 ( .A(n3058), .ZN(n3060) );
  INV_X1 U3902 ( .A(n3062), .ZN(n3059) );
  NAND2_X1 U3903 ( .A1(n3059), .A2(STATE_REG_SCAN_IN), .ZN(n3870) );
  NAND2_X1 U3904 ( .A1(n3060), .A2(n3870), .ZN(n3076) );
  AOI21_X1 U3905 ( .B1(n3063), .B2(n3062), .A(n3061), .ZN(n3075) );
  INV_X1 U3906 ( .A(n3075), .ZN(n3064) );
  INV_X1 U3907 ( .A(U4043), .ZN(n3875) );
  NOR2_X1 U3908 ( .A1(n4500), .A2(U4043), .ZN(U3148) );
  INV_X1 U3909 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U3910 ( .A1(U4043), .A2(n3238), .ZN(n3065) );
  OAI21_X1 U3911 ( .B1(U4043), .B2(n4723), .A(n3065), .ZN(U3553) );
  INV_X1 U3912 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U3913 ( .A1(U4043), .A2(n3388), .ZN(n3066) );
  OAI21_X1 U3914 ( .B1(U4043), .B2(n4699), .A(n3066), .ZN(U3557) );
  INV_X1 U3915 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U3916 ( .A1(U4043), .A2(n3485), .ZN(n3067) );
  OAI21_X1 U3917 ( .B1(U4043), .B2(n4720), .A(n3067), .ZN(U3560) );
  INV_X1 U3918 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U3919 ( .A1(n3677), .A2(U4043), .ZN(n3068) );
  OAI21_X1 U3920 ( .B1(U4043), .B2(n4655), .A(n3068), .ZN(U3567) );
  MUX2_X1 U3921 ( .A(n3069), .B(REG1_REG_1__SCAN_IN), .S(n3079), .Z(n3884) );
  NAND2_X1 U3922 ( .A1(n3888), .A2(REG1_REG_1__SCAN_IN), .ZN(n3899) );
  MUX2_X1 U3923 ( .A(n2389), .B(REG1_REG_2__SCAN_IN), .S(n4465), .Z(n3898) );
  INV_X1 U3924 ( .A(n3073), .ZN(n3074) );
  MUX2_X1 U3925 ( .A(REG1_REG_5__SCAN_IN), .B(n2444), .S(n3107), .Z(n3101) );
  XNOR2_X1 U3926 ( .A(n3146), .B(REG1_REG_6__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U3927 ( .A1(n3076), .A2(n3075), .ZN(n4469) );
  MUX2_X1 U3928 ( .A(n3080), .B(REG2_REG_1__SCAN_IN), .S(n3079), .Z(n3886) );
  AND2_X1 U3929 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3887)
         );
  NAND2_X1 U3930 ( .A1(n3888), .A2(REG2_REG_1__SCAN_IN), .ZN(n3894) );
  XNOR2_X1 U3931 ( .A(n3083), .B(n4464), .ZN(n3094) );
  INV_X1 U3932 ( .A(n3083), .ZN(n3084) );
  INV_X1 U3933 ( .A(n3085), .ZN(n3086) );
  MUX2_X1 U3934 ( .A(REG2_REG_5__SCAN_IN), .B(n3315), .S(n3107), .Z(n3104) );
  INV_X1 U3935 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3339) );
  XNOR2_X1 U3936 ( .A(n3151), .B(n3339), .ZN(n3090) );
  INV_X1 U3937 ( .A(n4467), .ZN(n3117) );
  OR2_X1 U3938 ( .A1(n3117), .A2(n3087), .ZN(n3866) );
  AND2_X1 U3939 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3259) );
  AOI21_X1 U3940 ( .B1(n4500), .B2(ADDR_REG_6__SCAN_IN), .A(n3259), .ZN(n3088)
         );
  OAI21_X1 U3941 ( .B1(n4514), .B2(n2073), .A(n3088), .ZN(n3089) );
  AOI21_X1 U3942 ( .B1(n3090), .B2(n4510), .A(n3089), .ZN(n3091) );
  OAI21_X1 U3943 ( .B1(n3092), .B2(n4497), .A(n3091), .ZN(U3246) );
  XOR2_X1 U3944 ( .A(REG1_REG_3__SCAN_IN), .B(n3093), .Z(n3096) );
  XOR2_X1 U3945 ( .A(n3094), .B(REG2_REG_3__SCAN_IN), .Z(n3095) );
  AOI22_X1 U3946 ( .A1(n4494), .A2(n3096), .B1(n4510), .B2(n3095), .ZN(n3098)
         );
  INV_X1 U3947 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3291) );
  NOR2_X1 U3948 ( .A1(STATE_REG_SCAN_IN), .A2(n3291), .ZN(n3195) );
  AOI21_X1 U3949 ( .B1(n4500), .B2(ADDR_REG_3__SCAN_IN), .A(n3195), .ZN(n3097)
         );
  OAI211_X1 U3950 ( .C1(n2203), .C2(n4514), .A(n3098), .B(n3097), .ZN(U3243)
         );
  INV_X1 U3951 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U3952 ( .A1(n4204), .A2(U4043), .ZN(n3099) );
  OAI21_X1 U3953 ( .B1(U4043), .B2(n4701), .A(n3099), .ZN(U3570) );
  AOI211_X1 U3954 ( .C1(n3102), .C2(n3101), .A(n4497), .B(n3100), .ZN(n3110)
         );
  AOI211_X1 U3955 ( .C1(n3105), .C2(n3104), .A(n3939), .B(n3103), .ZN(n3109)
         );
  AND2_X1 U3956 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3627) );
  AOI21_X1 U3957 ( .B1(n4500), .B2(ADDR_REG_5__SCAN_IN), .A(n3627), .ZN(n3106)
         );
  OAI21_X1 U3958 ( .B1(n4514), .B2(n3107), .A(n3106), .ZN(n3108) );
  OR3_X1 U3959 ( .A1(n3110), .A2(n3109), .A3(n3108), .ZN(U3245) );
  XNOR2_X1 U3960 ( .A(n3111), .B(REG1_REG_4__SCAN_IN), .ZN(n3128) );
  XOR2_X1 U3961 ( .A(REG2_REG_4__SCAN_IN), .B(n3112), .Z(n3126) );
  NAND2_X1 U3962 ( .A1(n4500), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3963 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3239) );
  OAI211_X1 U3964 ( .C1(n4514), .C2(n3114), .A(n3113), .B(n3239), .ZN(n3125)
         );
  XNOR2_X1 U3965 ( .A(n3116), .B(n3115), .ZN(n3143) );
  NAND3_X1 U3966 ( .A1(n3143), .A2(n3119), .A3(n3117), .ZN(n3123) );
  INV_X1 U3967 ( .A(n3866), .ZN(n3121) );
  INV_X1 U3968 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4534) );
  NAND2_X1 U3969 ( .A1(n4467), .A2(n4534), .ZN(n3118) );
  AND2_X1 U3970 ( .A1(n3119), .A2(n3118), .ZN(n4468) );
  NOR2_X1 U3971 ( .A1(n4468), .A2(IR_REG_0__SCAN_IN), .ZN(n3120) );
  AOI211_X1 U3972 ( .C1(n3121), .C2(n3887), .A(n3120), .B(n3875), .ZN(n3122)
         );
  NAND2_X1 U3973 ( .A1(n3123), .A2(n3122), .ZN(n3906) );
  INV_X1 U3974 ( .A(n3906), .ZN(n3124) );
  AOI211_X1 U3975 ( .C1(n4510), .C2(n3126), .A(n3125), .B(n3124), .ZN(n3127)
         );
  OAI21_X1 U3976 ( .B1(n3128), .B2(n4497), .A(n3127), .ZN(U3244) );
  INV_X1 U3977 ( .A(n3132), .ZN(n3133) );
  AOI21_X1 U3978 ( .B1(n3129), .B2(n3131), .A(n3133), .ZN(n3140) );
  INV_X1 U3979 ( .A(n3218), .ZN(n3134) );
  NAND3_X1 U3980 ( .A1(n3136), .A2(n3135), .A3(n3134), .ZN(n3158) );
  AOI22_X1 U3981 ( .A1(n3707), .A2(n3238), .B1(n3695), .B2(n2894), .ZN(n3137)
         );
  OAI21_X1 U3982 ( .B1(n3703), .B2(n3175), .A(n3137), .ZN(n3138) );
  AOI21_X1 U3983 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3158), .A(n3138), .ZN(n3139)
         );
  OAI21_X1 U3984 ( .B1(n3140), .B2(n3711), .A(n3139), .ZN(U3234) );
  AOI22_X1 U3985 ( .A1(n3629), .A2(n3267), .B1(n3707), .B2(n2894), .ZN(n3142)
         );
  NAND2_X1 U3986 ( .A1(n3158), .A2(REG3_REG_0__SCAN_IN), .ZN(n3141) );
  OAI211_X1 U3987 ( .C1(n3143), .C2(n3711), .A(n3142), .B(n3141), .ZN(U3229)
         );
  INV_X1 U3988 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4669) );
  MUX2_X1 U3989 ( .A(REG1_REG_7__SCAN_IN), .B(n4669), .S(n3202), .Z(n3147) );
  XOR2_X1 U3990 ( .A(n3147), .B(n3204), .Z(n3156) );
  AND2_X1 U3991 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3400) );
  AOI21_X1 U3992 ( .B1(n4500), .B2(ADDR_REG_7__SCAN_IN), .A(n3400), .ZN(n3148)
         );
  OAI21_X1 U3993 ( .B1(n4514), .B2(n3202), .A(n3148), .ZN(n3155) );
  INV_X1 U3994 ( .A(n3149), .ZN(n3150) );
  INV_X1 U3995 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4668) );
  MUX2_X1 U3996 ( .A(REG2_REG_7__SCAN_IN), .B(n4668), .S(n3202), .Z(n3152) );
  NOR2_X1 U3997 ( .A1(n3153), .A2(n3152), .ZN(n3201) );
  AOI211_X1 U3998 ( .C1(n3153), .C2(n3152), .A(n3939), .B(n3201), .ZN(n3154)
         );
  AOI211_X1 U3999 ( .C1(n3156), .C2(n4494), .A(n3155), .B(n3154), .ZN(n3157)
         );
  INV_X1 U4000 ( .A(n3157), .ZN(U3247) );
  INV_X1 U4001 ( .A(n3158), .ZN(n3167) );
  OAI22_X1 U4002 ( .A1(n3159), .A2(n3704), .B1(n3669), .B2(n2896), .ZN(n3160)
         );
  AOI21_X1 U4003 ( .B1(n3270), .B2(n3629), .A(n3160), .ZN(n3166) );
  CLKBUF_X1 U4004 ( .A(n3162), .Z(n3163) );
  OAI211_X1 U4005 ( .C1(n3161), .C2(n3164), .A(n3623), .B(n3163), .ZN(n3165)
         );
  OAI211_X1 U4006 ( .C1(n3167), .C2(n3278), .A(n3166), .B(n3165), .ZN(U3219)
         );
  NAND2_X1 U4007 ( .A1(n3168), .A2(n3169), .ZN(n3212) );
  OAI21_X1 U4008 ( .B1(n3168), .B2(n3169), .A(n3212), .ZN(n4517) );
  INV_X1 U4009 ( .A(n4517), .ZN(n3178) );
  INV_X1 U4010 ( .A(n4528), .ZN(n3177) );
  OAI21_X1 U4011 ( .B1(n3758), .B2(n3171), .A(n3170), .ZN(n3172) );
  NAND2_X1 U4012 ( .A1(n3172), .A2(n4270), .ZN(n3174) );
  AOI22_X1 U4013 ( .A1(n4272), .A2(n2894), .B1(n4273), .B2(n3238), .ZN(n3173)
         );
  OAI211_X1 U4014 ( .C1(n4278), .C2(n3175), .A(n3174), .B(n3173), .ZN(n3176)
         );
  AOI21_X1 U4015 ( .B1(n3177), .B2(n4517), .A(n3176), .ZN(n4520) );
  OAI21_X1 U4016 ( .B1(n3178), .B2(n4551), .A(n4520), .ZN(n3250) );
  NAND2_X1 U4017 ( .A1(n3250), .A2(n4739), .ZN(n3182) );
  INV_X1 U4018 ( .A(n4451), .ZN(n3429) );
  AND2_X1 U4019 ( .A1(n3265), .A2(n3179), .ZN(n3180) );
  NOR2_X1 U4020 ( .A1(n3290), .A2(n3180), .ZN(n4515) );
  NAND2_X1 U4021 ( .A1(n3429), .A2(n4515), .ZN(n3181) );
  OAI211_X1 U4022 ( .C1(n4739), .C2(n2391), .A(n3182), .B(n3181), .ZN(U3471)
         );
  AND2_X1 U4023 ( .A1(n3814), .A2(n3811), .ZN(n3774) );
  XOR2_X1 U4024 ( .A(n3183), .B(n3774), .Z(n3336) );
  XNOR2_X1 U4025 ( .A(n3184), .B(n3774), .ZN(n3187) );
  AOI22_X1 U4026 ( .A1(n4272), .A2(n3882), .B1(n4273), .B2(n3388), .ZN(n3185)
         );
  OAI21_X1 U4027 ( .B1(n3374), .B2(n4278), .A(n3185), .ZN(n3186) );
  AOI21_X1 U4028 ( .B1(n3187), .B2(n4270), .A(n3186), .ZN(n3344) );
  OAI21_X1 U4029 ( .B1(n3336), .B2(n4577), .A(n3344), .ZN(n3248) );
  NOR2_X1 U4030 ( .A1(n3318), .A2(n3374), .ZN(n3188) );
  OR2_X1 U4031 ( .A1(n3370), .A2(n3188), .ZN(n3337) );
  INV_X1 U4032 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3189) );
  OAI22_X1 U4033 ( .A1(n3337), .A2(n4451), .B1(n4739), .B2(n3189), .ZN(n3190)
         );
  AOI21_X1 U4034 ( .B1(n3248), .B2(n4739), .A(n3190), .ZN(n3191) );
  INV_X1 U4035 ( .A(n3191), .ZN(U3479) );
  XNOR2_X1 U4036 ( .A(n3193), .B(n3192), .ZN(n3199) );
  AOI22_X1 U4037 ( .A1(n3629), .A2(n3194), .B1(n3695), .B2(n3883), .ZN(n3197)
         );
  AOI21_X1 U4038 ( .B1(n3707), .B2(n2898), .A(n3195), .ZN(n3196) );
  OAI211_X1 U4039 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3689), .A(n3197), .B(n3196), 
        .ZN(n3198) );
  AOI21_X1 U4040 ( .B1(n3623), .B2(n3199), .A(n3198), .ZN(n3200) );
  INV_X1 U4041 ( .A(n3200), .ZN(U3215) );
  INV_X1 U4042 ( .A(n3202), .ZN(n4462) );
  AOI21_X1 U40430 ( .B1(n4462), .B2(REG2_REG_7__SCAN_IN), .A(n3201), .ZN(n3322) );
  XNOR2_X1 U4044 ( .A(n3323), .B(REG2_REG_8__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4045 ( .A1(n4462), .A2(REG1_REG_7__SCAN_IN), .ZN(n3203) );
  OAI211_X1 U4046 ( .C1(n3205), .C2(REG1_REG_8__SCAN_IN), .A(n3329), .B(n4494), 
        .ZN(n3208) );
  AND2_X1 U4047 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3390) );
  INV_X1 U4048 ( .A(n4461), .ZN(n3327) );
  NOR2_X1 U4049 ( .A1(n4514), .A2(n3327), .ZN(n3206) );
  AOI211_X1 U4050 ( .C1(n4500), .C2(ADDR_REG_8__SCAN_IN), .A(n3390), .B(n3206), 
        .ZN(n3207) );
  OAI211_X1 U4051 ( .C1(n3209), .C2(n3939), .A(n3208), .B(n3207), .ZN(U3248)
         );
  NAND2_X1 U4052 ( .A1(n3212), .A2(n3211), .ZN(n3282) );
  NAND2_X1 U4053 ( .A1(n3282), .A2(n3213), .ZN(n3215) );
  NAND2_X1 U4054 ( .A1(n3215), .A2(n3214), .ZN(n3216) );
  NAND2_X1 U4055 ( .A1(n3216), .A2(n3764), .ZN(n3217) );
  NAND2_X1 U4056 ( .A1(n3210), .A2(n3217), .ZN(n4556) );
  NOR2_X1 U4057 ( .A1(n3219), .A2(n3218), .ZN(n3220) );
  NAND2_X1 U4058 ( .A1(n3221), .A2(n3220), .ZN(n3222) );
  OR2_X1 U4059 ( .A1(n2364), .A2(n4526), .ZN(n3306) );
  XNOR2_X1 U4060 ( .A(n3764), .B(n3223), .ZN(n3227) );
  AOI22_X1 U4061 ( .A1(n4273), .A2(n3882), .B1(n4272), .B2(n3238), .ZN(n3225)
         );
  OAI211_X1 U4062 ( .C1(n4556), .C2(n4528), .A(n3225), .B(n3224), .ZN(n3226)
         );
  AOI21_X1 U4063 ( .B1(n3227), .B2(n4270), .A(n3226), .ZN(n3228) );
  INV_X1 U4064 ( .A(n3228), .ZN(n4558) );
  INV_X1 U4065 ( .A(n3288), .ZN(n3229) );
  OAI211_X1 U4066 ( .C1(n3229), .C2(n2886), .A(n2998), .B(n3316), .ZN(n4557)
         );
  OAI22_X1 U4067 ( .A1(n4557), .A2(n3978), .B1(n4255), .B2(n3243), .ZN(n3230)
         );
  OAI21_X1 U4068 ( .B1(n4558), .B2(n3230), .A(n4535), .ZN(n3232) );
  NAND2_X1 U4069 ( .A1(n2003), .A2(REG2_REG_4__SCAN_IN), .ZN(n3231) );
  OAI211_X1 U4070 ( .C1(n4556), .C2(n4193), .A(n3232), .B(n3231), .ZN(U3286)
         );
  INV_X1 U4071 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U4072 ( .A1(n4066), .A2(U4043), .ZN(n3233) );
  OAI21_X1 U4073 ( .B1(U4043), .B2(n4649), .A(n3233), .ZN(U3575) );
  INV_X1 U4074 ( .A(n3235), .ZN(n3236) );
  AOI211_X1 U4075 ( .C1(n3237), .C2(n3234), .A(n3711), .B(n3236), .ZN(n3245)
         );
  INV_X1 U4076 ( .A(n3239), .ZN(n3240) );
  AOI21_X1 U4077 ( .B1(n3707), .B2(n3882), .A(n3240), .ZN(n3241) );
  OAI211_X1 U4078 ( .C1(n3689), .C2(n3243), .A(n3242), .B(n3241), .ZN(n3244)
         );
  OR2_X1 U4079 ( .A1(n3245), .A2(n3244), .ZN(U3227) );
  INV_X1 U4080 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3246) );
  OAI22_X1 U4081 ( .A1(n3337), .A2(n4391), .B1(n4589), .B2(n3246), .ZN(n3247)
         );
  AOI21_X1 U4082 ( .B1(n3248), .B2(n4589), .A(n3247), .ZN(n3249) );
  INV_X1 U4083 ( .A(n3249), .ZN(U3524) );
  NAND2_X1 U4084 ( .A1(n3250), .A2(n4589), .ZN(n3252) );
  INV_X1 U4085 ( .A(n4391), .ZN(n4312) );
  NAND2_X1 U4086 ( .A1(n4312), .A2(n4515), .ZN(n3251) );
  OAI211_X1 U4087 ( .C1(n4589), .C2(n2389), .A(n3252), .B(n3251), .ZN(U3520)
         );
  INV_X1 U4088 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U4089 ( .A1(n4065), .A2(U4043), .ZN(n3253) );
  OAI21_X1 U4090 ( .B1(U4043), .B2(n4705), .A(n3253), .ZN(U3577) );
  XNOR2_X1 U4091 ( .A(n3255), .B(n3254), .ZN(n3256) );
  XNOR2_X1 U4092 ( .A(n3257), .B(n3256), .ZN(n3263) );
  AOI22_X1 U4093 ( .A1(n3629), .A2(n3258), .B1(n3695), .B2(n3882), .ZN(n3261)
         );
  AOI21_X1 U4094 ( .B1(n3707), .B2(n3388), .A(n3259), .ZN(n3260) );
  OAI211_X1 U4095 ( .C1(n3689), .C2(n3338), .A(n3261), .B(n3260), .ZN(n3262)
         );
  AOI21_X1 U4096 ( .B1(n3263), .B2(n3623), .A(n3262), .ZN(n3264) );
  INV_X1 U4097 ( .A(n3264), .ZN(U3236) );
  NAND2_X1 U4098 ( .A1(n4535), .A2(n4526), .ZN(n4229) );
  INV_X1 U4099 ( .A(n3265), .ZN(n3266) );
  AOI21_X1 U4100 ( .B1(n3267), .B2(n3270), .A(n3266), .ZN(n4548) );
  OAI21_X1 U4101 ( .B1(n3274), .B2(n3269), .A(n3268), .ZN(n4545) );
  NAND2_X1 U4102 ( .A1(n3270), .A2(n4525), .ZN(n3273) );
  NAND2_X1 U4103 ( .A1(n4273), .A2(n3883), .ZN(n3272) );
  NAND2_X1 U4104 ( .A1(n4272), .A2(n2893), .ZN(n3271) );
  AND3_X1 U4105 ( .A1(n3273), .A2(n3272), .A3(n3271), .ZN(n3277) );
  INV_X1 U4106 ( .A(n3798), .ZN(n3782) );
  XNOR2_X1 U4107 ( .A(n3274), .B(n3782), .ZN(n3275) );
  NAND2_X1 U4108 ( .A1(n3275), .A2(n4270), .ZN(n3276) );
  OAI211_X1 U4109 ( .C1(n4545), .C2(n4528), .A(n3277), .B(n3276), .ZN(n4546)
         );
  MUX2_X1 U4110 ( .A(REG2_REG_1__SCAN_IN), .B(n4546), .S(n4535), .Z(n3280) );
  OAI22_X1 U4111 ( .A1(n4193), .A2(n4545), .B1(n3278), .B2(n4255), .ZN(n3279)
         );
  AOI211_X1 U4112 ( .C1(n4516), .C2(n4548), .A(n3280), .B(n3279), .ZN(n3281)
         );
  INV_X1 U4113 ( .A(n3281), .ZN(U3289) );
  XNOR2_X1 U4114 ( .A(n3282), .B(n3757), .ZN(n4552) );
  XNOR2_X1 U4115 ( .A(n3283), .B(n3757), .ZN(n3286) );
  AOI22_X1 U4116 ( .A1(n4272), .A2(n3883), .B1(n4273), .B2(n2898), .ZN(n3284)
         );
  OAI21_X1 U4117 ( .B1(n3289), .B2(n4278), .A(n3284), .ZN(n3285) );
  AOI21_X1 U4118 ( .B1(n3286), .B2(n4270), .A(n3285), .ZN(n3287) );
  OAI21_X1 U4119 ( .B1(n4552), .B2(n4528), .A(n3287), .ZN(n4554) );
  INV_X1 U4120 ( .A(n4554), .ZN(n3296) );
  INV_X1 U4121 ( .A(n4552), .ZN(n3294) );
  OAI21_X1 U4122 ( .B1(n3290), .B2(n3289), .A(n3288), .ZN(n4550) );
  AOI22_X1 U4123 ( .A1(n2003), .A2(REG2_REG_3__SCAN_IN), .B1(n4530), .B2(n3291), .ZN(n3292) );
  OAI21_X1 U4124 ( .B1(n4305), .B2(n4550), .A(n3292), .ZN(n3293) );
  AOI21_X1 U4125 ( .B1(n4532), .B2(n3294), .A(n3293), .ZN(n3295) );
  OAI21_X1 U4126 ( .B1(n2003), .B2(n3296), .A(n3295), .ZN(U3287) );
  AND2_X1 U4127 ( .A1(n3816), .A2(n3820), .ZN(n3773) );
  XNOR2_X1 U4128 ( .A(n3297), .B(n3773), .ZN(n3348) );
  XNOR2_X1 U4129 ( .A(n3298), .B(n3773), .ZN(n3301) );
  AOI22_X1 U4130 ( .A1(n4272), .A2(n3388), .B1(n4273), .B2(n3879), .ZN(n3300)
         );
  NAND2_X1 U4131 ( .A1(n3389), .A2(n4525), .ZN(n3299) );
  OAI211_X1 U4132 ( .C1(n3301), .C2(n4523), .A(n3300), .B(n3299), .ZN(n3345)
         );
  AOI21_X1 U4133 ( .B1(n3348), .B2(n4570), .A(n3345), .ZN(n3305) );
  INV_X1 U4134 ( .A(n3359), .ZN(n3302) );
  AOI21_X1 U4135 ( .B1(n3389), .B2(n3368), .A(n3302), .ZN(n3347) );
  AOI22_X1 U4136 ( .A1(n3347), .A2(n4312), .B1(REG1_REG_8__SCAN_IN), .B2(n4587), .ZN(n3303) );
  OAI21_X1 U4137 ( .B1(n3305), .B2(n4587), .A(n3303), .ZN(U3526) );
  AOI22_X1 U4138 ( .A1(n3347), .A2(n3429), .B1(REG0_REG_8__SCAN_IN), .B2(n4737), .ZN(n3304) );
  OAI21_X1 U4139 ( .B1(n3305), .B2(n4737), .A(n3304), .ZN(U3483) );
  NAND2_X1 U4140 ( .A1(n4528), .A2(n3306), .ZN(n3307) );
  INV_X1 U4141 ( .A(n3309), .ZN(n3808) );
  NAND2_X1 U4142 ( .A1(n3808), .A2(n3812), .ZN(n3772) );
  XNOR2_X1 U4143 ( .A(n3308), .B(n3772), .ZN(n4563) );
  XNOR2_X1 U4144 ( .A(n3310), .B(n3772), .ZN(n3314) );
  AOI22_X1 U4145 ( .A1(n4273), .A2(n3881), .B1(n4272), .B2(n2898), .ZN(n3311)
         );
  OAI21_X1 U4146 ( .B1(n3312), .B2(n4278), .A(n3311), .ZN(n3313) );
  AOI21_X1 U4147 ( .B1(n3314), .B2(n4270), .A(n3313), .ZN(n4564) );
  MUX2_X1 U4148 ( .A(n4564), .B(n3315), .S(n2003), .Z(n3321) );
  AND2_X1 U4149 ( .A1(n3316), .A2(n3628), .ZN(n3317) );
  NOR2_X1 U4150 ( .A1(n3318), .A2(n3317), .ZN(n4567) );
  INV_X1 U4151 ( .A(n3630), .ZN(n3319) );
  AOI22_X1 U4152 ( .A1(n4516), .A2(n4567), .B1(n3319), .B2(n4530), .ZN(n3320)
         );
  OAI211_X1 U4153 ( .C1(n4286), .C2(n4563), .A(n3321), .B(n3320), .ZN(U3285)
         );
  INV_X1 U4154 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3441) );
  MUX2_X1 U4155 ( .A(n3441), .B(REG2_REG_9__SCAN_IN), .S(n4460), .Z(n3325) );
  INV_X1 U4156 ( .A(n3442), .ZN(n3324) );
  AOI211_X1 U4157 ( .C1(n2041), .C2(n3325), .A(n3939), .B(n3324), .ZN(n3335)
         );
  INV_X1 U4158 ( .A(n4460), .ZN(n3449) );
  XOR2_X1 U4159 ( .A(REG1_REG_9__SCAN_IN), .B(n4460), .Z(n3330) );
  NAND2_X1 U4160 ( .A1(n3331), .A2(n3330), .ZN(n3450) );
  OAI211_X1 U4161 ( .C1(n3331), .C2(n3330), .A(n3450), .B(n4494), .ZN(n3333)
         );
  AND2_X1 U4162 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3420) );
  AOI21_X1 U4163 ( .B1(n4500), .B2(ADDR_REG_9__SCAN_IN), .A(n3420), .ZN(n3332)
         );
  OAI211_X1 U4164 ( .C1(n4514), .C2(n3449), .A(n3333), .B(n3332), .ZN(n3334)
         );
  OR2_X1 U4165 ( .A1(n3335), .A2(n3334), .ZN(U3249) );
  INV_X1 U4166 ( .A(n3336), .ZN(n3342) );
  NOR2_X1 U4167 ( .A1(n3337), .A2(n4305), .ZN(n3341) );
  OAI22_X1 U4168 ( .A1(n4535), .A2(n3339), .B1(n3338), .B2(n4255), .ZN(n3340)
         );
  AOI211_X1 U4169 ( .C1(n3342), .C2(n4231), .A(n3341), .B(n3340), .ZN(n3343)
         );
  OAI21_X1 U4170 ( .B1(n2003), .B2(n3344), .A(n3343), .ZN(U3284) );
  INV_X1 U4171 ( .A(n3345), .ZN(n3351) );
  OAI22_X1 U4172 ( .A1(n4535), .A2(n2190), .B1(n3393), .B2(n4255), .ZN(n3346)
         );
  AOI21_X1 U4173 ( .B1(n3347), .B2(n4516), .A(n3346), .ZN(n3350) );
  NAND2_X1 U4174 ( .A1(n3348), .A2(n4231), .ZN(n3349) );
  OAI211_X1 U4175 ( .C1(n3351), .C2(n2003), .A(n3350), .B(n3349), .ZN(U3282)
         );
  AND2_X1 U4176 ( .A1(n2135), .A2(n3821), .ZN(n3776) );
  XNOR2_X1 U4177 ( .A(n3352), .B(n3776), .ZN(n3439) );
  XNOR2_X1 U4178 ( .A(n3353), .B(n3776), .ZN(n3357) );
  OAI22_X1 U4179 ( .A1(n3354), .A2(n4288), .B1(n4521), .B2(n2913), .ZN(n3355)
         );
  AOI21_X1 U4180 ( .B1(n3419), .B2(n4525), .A(n3355), .ZN(n3356) );
  OAI21_X1 U4181 ( .B1(n3357), .B2(n4523), .A(n3356), .ZN(n3436) );
  AOI21_X1 U4182 ( .B1(n3439), .B2(n4570), .A(n3436), .ZN(n3362) );
  INV_X1 U4183 ( .A(n3412), .ZN(n3358) );
  AOI21_X1 U4184 ( .B1(n3419), .B2(n3359), .A(n3358), .ZN(n3433) );
  AOI22_X1 U4185 ( .A1(n3433), .A2(n4312), .B1(REG1_REG_9__SCAN_IN), .B2(n4587), .ZN(n3360) );
  OAI21_X1 U4186 ( .B1(n3362), .B2(n4587), .A(n3360), .ZN(U3527) );
  AOI22_X1 U4187 ( .A1(n3433), .A2(n3429), .B1(REG0_REG_9__SCAN_IN), .B2(n4737), .ZN(n3361) );
  OAI21_X1 U4188 ( .B1(n3362), .B2(n4737), .A(n3361), .ZN(U3485) );
  INV_X1 U4189 ( .A(n3378), .ZN(n3815) );
  XNOR2_X1 U4190 ( .A(n3363), .B(n3815), .ZN(n3367) );
  NAND2_X1 U4191 ( .A1(n4272), .A2(n3881), .ZN(n3365) );
  NAND2_X1 U4192 ( .A1(n4273), .A2(n3880), .ZN(n3364) );
  OAI211_X1 U4193 ( .C1(n3369), .C2(n4278), .A(n3365), .B(n3364), .ZN(n3366)
         );
  AOI21_X1 U4194 ( .B1(n3367), .B2(n4270), .A(n3366), .ZN(n4574) );
  OAI211_X1 U4195 ( .C1(n3370), .C2(n3369), .A(n2998), .B(n3368), .ZN(n4573)
         );
  INV_X1 U4196 ( .A(n4573), .ZN(n3373) );
  INV_X1 U4197 ( .A(n4229), .ZN(n3372) );
  OAI22_X1 U4198 ( .A1(n4535), .A2(n4668), .B1(n3403), .B2(n4255), .ZN(n3371)
         );
  AOI21_X1 U4199 ( .B1(n3373), .B2(n3372), .A(n3371), .ZN(n3382) );
  NAND2_X1 U4200 ( .A1(n3183), .A2(n3881), .ZN(n3375) );
  NAND2_X1 U4201 ( .A1(n3375), .A2(n3374), .ZN(n3377) );
  OR2_X1 U4202 ( .A1(n3183), .A2(n3881), .ZN(n3376) );
  AND2_X1 U4203 ( .A1(n3377), .A2(n3376), .ZN(n3379) );
  NAND2_X1 U4204 ( .A1(n3379), .A2(n3378), .ZN(n4571) );
  INV_X1 U4205 ( .A(n3379), .ZN(n3380) );
  NAND2_X1 U4206 ( .A1(n3380), .A2(n3815), .ZN(n4569) );
  NAND3_X1 U4207 ( .A1(n4571), .A2(n4231), .A3(n4569), .ZN(n3381) );
  OAI211_X1 U4208 ( .C1(n4574), .C2(n2003), .A(n3382), .B(n3381), .ZN(U3283)
         );
  NAND2_X1 U4209 ( .A1(n3383), .A2(n3384), .ZN(n3387) );
  NAND2_X1 U4210 ( .A1(n2298), .A2(n3385), .ZN(n3386) );
  XNOR2_X1 U4211 ( .A(n3387), .B(n3386), .ZN(n3395) );
  AOI22_X1 U4212 ( .A1(n3629), .A2(n3389), .B1(n3695), .B2(n3388), .ZN(n3392)
         );
  AOI21_X1 U4213 ( .B1(n3707), .B2(n3879), .A(n3390), .ZN(n3391) );
  OAI211_X1 U4214 ( .C1(n3689), .C2(n3393), .A(n3392), .B(n3391), .ZN(n3394)
         );
  AOI21_X1 U4215 ( .B1(n3395), .B2(n3623), .A(n3394), .ZN(n3396) );
  INV_X1 U4216 ( .A(n3396), .ZN(U3218) );
  XOR2_X1 U4217 ( .A(n3398), .B(n3397), .Z(n3405) );
  AOI22_X1 U4218 ( .A1(n3629), .A2(n3399), .B1(n3695), .B2(n3881), .ZN(n3402)
         );
  AOI21_X1 U4219 ( .B1(n3707), .B2(n3880), .A(n3400), .ZN(n3401) );
  OAI211_X1 U4220 ( .C1(n3689), .C2(n3403), .A(n3402), .B(n3401), .ZN(n3404)
         );
  AOI21_X1 U4221 ( .B1(n3405), .B2(n3623), .A(n3404), .ZN(n3406) );
  INV_X1 U4222 ( .A(n3406), .ZN(U3210) );
  NAND2_X1 U4223 ( .A1(n3823), .A2(n3826), .ZN(n3771) );
  XNOR2_X1 U4224 ( .A(n3407), .B(n3771), .ZN(n3410) );
  AOI22_X1 U4225 ( .A1(n4272), .A2(n3879), .B1(n4273), .B2(n3878), .ZN(n3409)
         );
  NAND2_X1 U4226 ( .A1(n3495), .A2(n4525), .ZN(n3408) );
  OAI211_X1 U4227 ( .C1(n3410), .C2(n4523), .A(n3409), .B(n3408), .ZN(n3426)
         );
  INV_X1 U4228 ( .A(n3426), .ZN(n3416) );
  XOR2_X1 U4229 ( .A(n3411), .B(n3771), .Z(n3427) );
  NAND2_X1 U4230 ( .A1(n3427), .A2(n4231), .ZN(n3415) );
  AOI21_X1 U4231 ( .B1(n3495), .B2(n3412), .A(n4301), .ZN(n3430) );
  OAI22_X1 U4232 ( .A1(n4535), .A2(n2177), .B1(n3499), .B2(n4255), .ZN(n3413)
         );
  AOI21_X1 U4233 ( .B1(n3430), .B2(n4516), .A(n3413), .ZN(n3414) );
  OAI211_X1 U4234 ( .C1(n2003), .C2(n3416), .A(n3415), .B(n3414), .ZN(U3280)
         );
  XNOR2_X1 U4235 ( .A(n3417), .B(n3418), .ZN(n3424) );
  AOI22_X1 U4236 ( .A1(n3629), .A2(n3419), .B1(n3695), .B2(n3880), .ZN(n3422)
         );
  AOI21_X1 U4237 ( .B1(n3707), .B2(n3485), .A(n3420), .ZN(n3421) );
  OAI211_X1 U4238 ( .C1(n3689), .C2(n3434), .A(n3422), .B(n3421), .ZN(n3423)
         );
  AOI21_X1 U4239 ( .B1(n3424), .B2(n3623), .A(n3423), .ZN(n3425) );
  INV_X1 U4240 ( .A(n3425), .ZN(U3228) );
  AOI21_X1 U4241 ( .B1(n3427), .B2(n4570), .A(n3426), .ZN(n3432) );
  AOI22_X1 U4242 ( .A1(n3430), .A2(n4312), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4587), .ZN(n3428) );
  OAI21_X1 U4243 ( .B1(n3432), .B2(n4587), .A(n3428), .ZN(U3528) );
  AOI22_X1 U4244 ( .A1(n3430), .A2(n3429), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4737), .ZN(n3431) );
  OAI21_X1 U4245 ( .B1(n3432), .B2(n4737), .A(n3431), .ZN(U3487) );
  INV_X1 U4246 ( .A(n3433), .ZN(n3435) );
  OAI22_X1 U4247 ( .A1(n3435), .A2(n4305), .B1(n3434), .B2(n4255), .ZN(n3438)
         );
  MUX2_X1 U4248 ( .A(REG2_REG_9__SCAN_IN), .B(n3436), .S(n4535), .Z(n3437) );
  AOI211_X1 U4249 ( .C1(n4231), .C2(n3439), .A(n3438), .B(n3437), .ZN(n3440)
         );
  INV_X1 U4250 ( .A(n3440), .ZN(U3281) );
  INV_X1 U4251 ( .A(n4459), .ZN(n3462) );
  INV_X1 U4252 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4676) );
  MUX2_X1 U4253 ( .A(REG2_REG_11__SCAN_IN), .B(n4676), .S(n4458), .Z(n3444) );
  AOI21_X1 U4254 ( .B1(n2042), .B2(n3444), .A(n3939), .ZN(n3447) );
  AND2_X1 U4255 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3484) );
  AOI21_X1 U4256 ( .B1(n4500), .B2(ADDR_REG_11__SCAN_IN), .A(n3484), .ZN(n3445) );
  OAI21_X1 U4257 ( .B1(n4514), .B2(n4458), .A(n3445), .ZN(n3446) );
  AOI21_X1 U4258 ( .B1(n3447), .B2(n3911), .A(n3446), .ZN(n3456) );
  INV_X1 U4259 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3448) );
  INV_X1 U4260 ( .A(n3451), .ZN(n3452) );
  XNOR2_X1 U4261 ( .A(n4458), .B(REG1_REG_11__SCAN_IN), .ZN(n3453) );
  OAI211_X1 U4262 ( .C1(n3454), .C2(n3453), .A(n3914), .B(n4494), .ZN(n3455)
         );
  NAND2_X1 U4263 ( .A1(n3456), .A2(n3455), .ZN(U3251) );
  XNOR2_X1 U4264 ( .A(n3457), .B(n2177), .ZN(n3464) );
  OAI211_X1 U4265 ( .C1(n3459), .C2(REG1_REG_10__SCAN_IN), .A(n3458), .B(n4494), .ZN(n3461) );
  AND2_X1 U4266 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3496) );
  AOI21_X1 U4267 ( .B1(n4500), .B2(ADDR_REG_10__SCAN_IN), .A(n3496), .ZN(n3460) );
  OAI211_X1 U4268 ( .C1(n4514), .C2(n3462), .A(n3461), .B(n3460), .ZN(n3463)
         );
  AOI21_X1 U4269 ( .B1(n4510), .B2(n3464), .A(n3463), .ZN(n3465) );
  INV_X1 U4270 ( .A(n3465), .ZN(U3250) );
  NAND2_X1 U4271 ( .A1(n3503), .A2(n3505), .ZN(n3783) );
  INV_X1 U4272 ( .A(n3466), .ZN(n3468) );
  OAI21_X1 U4273 ( .B1(n4287), .B2(n3468), .A(n3467), .ZN(n3506) );
  XOR2_X1 U4274 ( .A(n3783), .B(n3506), .Z(n3472) );
  OAI22_X1 U4275 ( .A1(n3522), .A2(n4521), .B1(n4288), .B2(n3469), .ZN(n3470)
         );
  AOI21_X1 U4276 ( .B1(n3603), .B2(n4525), .A(n3470), .ZN(n3471) );
  OAI21_X1 U4277 ( .B1(n3472), .B2(n4523), .A(n3471), .ZN(n4384) );
  INV_X1 U4278 ( .A(n4384), .ZN(n3479) );
  XNOR2_X1 U4279 ( .A(n3473), .B(n3783), .ZN(n4385) );
  NAND2_X1 U4280 ( .A1(n3474), .A2(n3603), .ZN(n3475) );
  NAND2_X1 U4281 ( .A1(n3513), .A2(n3475), .ZN(n4448) );
  NOR2_X1 U4282 ( .A1(n4448), .A2(n4305), .ZN(n3477) );
  INV_X1 U4283 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3924) );
  OAI22_X1 U4284 ( .A1(n4535), .A2(n3924), .B1(n3606), .B2(n4255), .ZN(n3476)
         );
  AOI211_X1 U4285 ( .C1(n4385), .C2(n4231), .A(n3477), .B(n3476), .ZN(n3478)
         );
  OAI21_X1 U4286 ( .B1(n2003), .B2(n3479), .A(n3478), .ZN(U3278) );
  XOR2_X1 U4287 ( .A(n3482), .B(n3481), .Z(n3483) );
  XNOR2_X1 U4288 ( .A(n3480), .B(n3483), .ZN(n3490) );
  AOI21_X1 U4289 ( .B1(n3695), .B2(n3485), .A(n3484), .ZN(n3487) );
  NAND2_X1 U4290 ( .A1(n3707), .A2(n3877), .ZN(n3486) );
  OAI211_X1 U4291 ( .C1(n3703), .C2(n4300), .A(n3487), .B(n3486), .ZN(n3488)
         );
  AOI21_X1 U4292 ( .B1(n3708), .B2(n4303), .A(n3488), .ZN(n3489) );
  OAI21_X1 U4293 ( .B1(n3490), .B2(n3711), .A(n3489), .ZN(U3233) );
  INV_X1 U4294 ( .A(n3492), .ZN(n3493) );
  AOI211_X1 U4295 ( .C1(n3494), .C2(n3491), .A(n3711), .B(n3493), .ZN(n3501)
         );
  AOI22_X1 U4296 ( .A1(n3629), .A2(n3495), .B1(n3707), .B2(n3878), .ZN(n3498)
         );
  AOI21_X1 U4297 ( .B1(n3695), .B2(n3879), .A(n3496), .ZN(n3497) );
  OAI211_X1 U4298 ( .C1(n3689), .C2(n3499), .A(n3498), .B(n3497), .ZN(n3500)
         );
  OR2_X1 U4299 ( .A1(n3501), .A2(n3500), .ZN(U3214) );
  XNOR2_X1 U4300 ( .A(n3522), .B(n3659), .ZN(n3779) );
  XOR2_X1 U4301 ( .A(n3779), .B(n3502), .Z(n3512) );
  INV_X1 U4302 ( .A(n3503), .ZN(n3504) );
  AOI21_X1 U4303 ( .B1(n3506), .B2(n3505), .A(n3504), .ZN(n3507) );
  XNOR2_X1 U4304 ( .A(n3507), .B(n3779), .ZN(n3510) );
  AOI22_X1 U4305 ( .A1(n4271), .A2(n4273), .B1(n4272), .B2(n3877), .ZN(n3508)
         );
  OAI21_X1 U4306 ( .B1(n3659), .B2(n4278), .A(n3508), .ZN(n3509) );
  AOI21_X1 U4307 ( .B1(n3510), .B2(n4270), .A(n3509), .ZN(n3511) );
  OAI21_X1 U4308 ( .B1(n3512), .B2(n4528), .A(n3511), .ZN(n4380) );
  INV_X1 U4309 ( .A(n4380), .ZN(n3520) );
  INV_X1 U4310 ( .A(n3512), .ZN(n4381) );
  INV_X1 U4311 ( .A(n3513), .ZN(n3516) );
  INV_X1 U4312 ( .A(n3514), .ZN(n3515) );
  OAI21_X1 U4313 ( .B1(n3516), .B2(n3659), .A(n3515), .ZN(n4444) );
  AOI22_X1 U4314 ( .A1(n2003), .A2(REG2_REG_13__SCAN_IN), .B1(n3661), .B2(
        n4530), .ZN(n3517) );
  OAI21_X1 U4315 ( .B1(n4444), .B2(n4305), .A(n3517), .ZN(n3518) );
  AOI21_X1 U4316 ( .B1(n4381), .B2(n4532), .A(n3518), .ZN(n3519) );
  OAI21_X1 U4317 ( .B1(n3520), .B2(n2003), .A(n3519), .ZN(U3277) );
  INV_X1 U4318 ( .A(n3521), .ZN(n3733) );
  XNOR2_X1 U4319 ( .A(n3733), .B(n3759), .ZN(n3527) );
  OAI22_X1 U4320 ( .A1(n3523), .A2(n4521), .B1(n3522), .B2(n4288), .ZN(n3524)
         );
  AOI21_X1 U4321 ( .B1(n3525), .B2(n4525), .A(n3524), .ZN(n3526) );
  OAI21_X1 U4322 ( .B1(n3527), .B2(n4523), .A(n3526), .ZN(n4377) );
  INV_X1 U4323 ( .A(n4377), .ZN(n3534) );
  OAI21_X1 U4324 ( .B1(n3528), .B2(n2150), .A(n3529), .ZN(n4378) );
  NOR2_X1 U4325 ( .A1(n3514), .A2(n3572), .ZN(n3530) );
  OR2_X1 U4326 ( .A1(n4280), .A2(n3530), .ZN(n4441) );
  AOI22_X1 U4327 ( .A1(n2003), .A2(REG2_REG_14__SCAN_IN), .B1(n3574), .B2(
        n4530), .ZN(n3531) );
  OAI21_X1 U4328 ( .B1(n4441), .B2(n4305), .A(n3531), .ZN(n3532) );
  AOI21_X1 U4329 ( .B1(n4378), .B2(n4231), .A(n3532), .ZN(n3533) );
  OAI21_X1 U4330 ( .B1(n2003), .B2(n3534), .A(n3533), .ZN(U3276) );
  INV_X1 U4331 ( .A(n3535), .ZN(n3536) );
  OAI21_X1 U4332 ( .B1(n3542), .B2(n3541), .A(n3540), .ZN(n3543) );
  XNOR2_X1 U4333 ( .A(n3544), .B(n3543), .ZN(n3550) );
  OAI22_X1 U4334 ( .A1(n4124), .A2(n3704), .B1(STATE_REG_SCAN_IN), .B2(n3545), 
        .ZN(n3548) );
  OAI22_X1 U4335 ( .A1(n4087), .A2(n3669), .B1(n3703), .B2(n3546), .ZN(n3547)
         );
  AOI211_X1 U4336 ( .C1(n4091), .C2(n3708), .A(n3548), .B(n3547), .ZN(n3549)
         );
  OAI21_X1 U4337 ( .B1(n3550), .B2(n3711), .A(n3549), .ZN(U3222) );
  INV_X1 U4338 ( .A(n3551), .ZN(n3556) );
  AOI22_X1 U4339 ( .A1(n3552), .A2(n4530), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2003), .ZN(n3553) );
  OAI21_X1 U4340 ( .B1(n3554), .B2(n4305), .A(n3553), .ZN(n3555) );
  AOI21_X1 U4341 ( .B1(n3556), .B2(n4535), .A(n3555), .ZN(n3557) );
  OAI21_X1 U4342 ( .B1(n3558), .B2(n4286), .A(n3557), .ZN(U3262) );
  XNOR2_X1 U4343 ( .A(n3560), .B(n3559), .ZN(n3565) );
  NOR2_X1 U4344 ( .A1(n4046), .A2(n3689), .ZN(n3563) );
  AOI22_X1 U4345 ( .A1(n3873), .A2(n3695), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3561) );
  OAI21_X1 U4346 ( .B1(n3703), .B2(n4048), .A(n3561), .ZN(n3562) );
  AOI211_X1 U4347 ( .C1(n3707), .C2(n4014), .A(n3563), .B(n3562), .ZN(n3564)
         );
  OAI21_X1 U4348 ( .B1(n3565), .B2(n3711), .A(n3564), .ZN(U3211) );
  INV_X1 U4349 ( .A(n3567), .ZN(n3611) );
  NOR2_X1 U4350 ( .A1(n3611), .A2(n3568), .ZN(n3569) );
  XNOR2_X1 U4351 ( .A(n3566), .B(n3569), .ZN(n3576) );
  AND2_X1 U4352 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n3945) );
  AOI21_X1 U4353 ( .B1(n3695), .B2(n3876), .A(n3945), .ZN(n3571) );
  NAND2_X1 U4354 ( .A1(n3707), .A2(n4262), .ZN(n3570) );
  OAI211_X1 U4355 ( .C1(n3703), .C2(n3572), .A(n3571), .B(n3570), .ZN(n3573)
         );
  AOI21_X1 U4356 ( .B1(n3708), .B2(n3574), .A(n3573), .ZN(n3575) );
  OAI21_X1 U4357 ( .B1(n3576), .B2(n3711), .A(n3575), .ZN(U3212) );
  OAI21_X1 U4358 ( .B1(n3579), .B2(n3577), .A(n3578), .ZN(n3585) );
  AOI22_X1 U4359 ( .A1(n3629), .A2(n3580), .B1(n3695), .B2(n4239), .ZN(n3583)
         );
  NAND2_X1 U4360 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3993) );
  INV_X1 U4361 ( .A(n3993), .ZN(n3581) );
  AOI21_X1 U4362 ( .B1(n3707), .B2(n4204), .A(n3581), .ZN(n3582) );
  OAI211_X1 U4363 ( .C1(n3689), .C2(n4210), .A(n3583), .B(n3582), .ZN(n3584)
         );
  AOI21_X1 U4364 ( .B1(n3585), .B2(n3623), .A(n3584), .ZN(n3586) );
  INV_X1 U4365 ( .A(n3586), .ZN(U3216) );
  NAND2_X1 U4366 ( .A1(n2036), .A2(n3587), .ZN(n3592) );
  INV_X1 U4367 ( .A(n3588), .ZN(n3590) );
  OAI211_X1 U4368 ( .C1(n3006), .C2(n3590), .A(n3589), .B(n3592), .ZN(n3591)
         );
  OAI211_X1 U4369 ( .C1(n3593), .C2(n3592), .A(n3623), .B(n3591), .ZN(n3597)
         );
  AOI22_X1 U4370 ( .A1(n3695), .A2(n4204), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3596) );
  AOI22_X1 U4371 ( .A1(n3874), .A2(n3707), .B1(n3629), .B2(n4163), .ZN(n3595)
         );
  NAND2_X1 U4372 ( .A1(n3708), .A2(n4166), .ZN(n3594) );
  NAND4_X1 U4373 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(U3220)
         );
  INV_X1 U4374 ( .A(n3599), .ZN(n3601) );
  NAND2_X1 U4375 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  XNOR2_X1 U4376 ( .A(n3598), .B(n3602), .ZN(n3608) );
  AOI22_X1 U4377 ( .A1(n3629), .A2(n3603), .B1(n3707), .B2(n3876), .ZN(n3605)
         );
  AND2_X1 U4378 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3916) );
  AOI21_X1 U4379 ( .B1(n3695), .B2(n3878), .A(n3916), .ZN(n3604) );
  OAI211_X1 U4380 ( .C1(n3689), .C2(n3606), .A(n3605), .B(n3604), .ZN(n3607)
         );
  AOI21_X1 U4381 ( .B1(n3608), .B2(n3623), .A(n3607), .ZN(n3609) );
  INV_X1 U4382 ( .A(n3609), .ZN(U3221) );
  NOR2_X1 U4383 ( .A1(n3610), .A2(n3611), .ZN(n3613) );
  NAND2_X1 U4384 ( .A1(n3613), .A2(n3612), .ZN(n3699) );
  NOR2_X1 U4385 ( .A1(n3613), .A2(n3612), .ZN(n3698) );
  AOI21_X1 U4386 ( .B1(n3701), .B2(n3699), .A(n3698), .ZN(n3617) );
  NAND2_X1 U4387 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  XNOR2_X1 U4388 ( .A(n3617), .B(n3616), .ZN(n3621) );
  AOI22_X1 U4389 ( .A1(n3629), .A2(n4261), .B1(n3695), .B2(n4262), .ZN(n3619)
         );
  AND2_X1 U4390 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4474) );
  AOI21_X1 U4391 ( .B1(n3707), .B2(n3677), .A(n4474), .ZN(n3618) );
  OAI211_X1 U4392 ( .C1(n3689), .C2(n4256), .A(n3619), .B(n3618), .ZN(n3620)
         );
  AOI21_X1 U4393 ( .B1(n3621), .B2(n3623), .A(n3620), .ZN(n3622) );
  INV_X1 U4394 ( .A(n3622), .ZN(U3223) );
  OAI211_X1 U4395 ( .C1(n3626), .C2(n3625), .A(n3624), .B(n3623), .ZN(n3634)
         );
  AOI21_X1 U4396 ( .B1(n3707), .B2(n3881), .A(n3627), .ZN(n3633) );
  AOI22_X1 U4397 ( .A1(n3629), .A2(n3628), .B1(n3695), .B2(n2898), .ZN(n3632)
         );
  OR2_X1 U4398 ( .A1(n3689), .A2(n3630), .ZN(n3631) );
  NAND4_X1 U4399 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(U3224)
         );
  NAND2_X1 U4400 ( .A1(n2043), .A2(n3636), .ZN(n3637) );
  XNOR2_X1 U4401 ( .A(n3635), .B(n3637), .ZN(n3642) );
  AND2_X1 U4402 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4485) );
  AOI21_X1 U4403 ( .B1(n3695), .B2(n4274), .A(n4485), .ZN(n3639) );
  NAND2_X1 U4404 ( .A1(n3707), .A2(n4239), .ZN(n3638) );
  OAI211_X1 U4405 ( .C1(n3703), .C2(n4244), .A(n3639), .B(n3638), .ZN(n3640)
         );
  AOI21_X1 U4406 ( .B1(n3708), .B2(n4245), .A(n3640), .ZN(n3641) );
  OAI21_X1 U4407 ( .B1(n3642), .B2(n3711), .A(n3641), .ZN(U3225) );
  NOR2_X1 U4408 ( .A1(n3645), .A2(n3644), .ZN(n3647) );
  XNOR2_X1 U4409 ( .A(n3647), .B(n3646), .ZN(n3652) );
  NOR2_X1 U4410 ( .A1(n3689), .A2(n4108), .ZN(n3650) );
  AOI22_X1 U4411 ( .A1(n4103), .A2(n3695), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3648) );
  OAI21_X1 U4412 ( .B1(n3703), .B2(n4110), .A(n3648), .ZN(n3649) );
  AOI211_X1 U4413 ( .C1(n3707), .C2(n4066), .A(n3650), .B(n3649), .ZN(n3651)
         );
  OAI21_X1 U4414 ( .B1(n3652), .B2(n3711), .A(n3651), .ZN(U3226) );
  XOR2_X1 U4415 ( .A(n3655), .B(n3654), .Z(n3656) );
  XNOR2_X1 U4416 ( .A(n3653), .B(n3656), .ZN(n3663) );
  AND2_X1 U4417 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3929) );
  AOI21_X1 U4418 ( .B1(n3695), .B2(n3877), .A(n3929), .ZN(n3658) );
  NAND2_X1 U4419 ( .A1(n3707), .A2(n4271), .ZN(n3657) );
  OAI211_X1 U4420 ( .C1(n3703), .C2(n3659), .A(n3658), .B(n3657), .ZN(n3660)
         );
  AOI21_X1 U4421 ( .B1(n3708), .B2(n3661), .A(n3660), .ZN(n3662) );
  OAI21_X1 U4422 ( .B1(n3663), .B2(n3711), .A(n3662), .ZN(U3231) );
  INV_X1 U4423 ( .A(n3664), .ZN(n3665) );
  AOI21_X1 U4424 ( .B1(n3667), .B2(n3666), .A(n3665), .ZN(n3673) );
  OAI22_X1 U4425 ( .A1(n4179), .A2(n3704), .B1(n3703), .B2(n4151), .ZN(n3671)
         );
  OAI22_X1 U4426 ( .A1(n4147), .A2(n3669), .B1(STATE_REG_SCAN_IN), .B2(n3668), 
        .ZN(n3670) );
  AOI211_X1 U4427 ( .C1(n4150), .C2(n3708), .A(n3671), .B(n3670), .ZN(n3672)
         );
  OAI21_X1 U4428 ( .B1(n3673), .B2(n3711), .A(n3672), .ZN(U3232) );
  XNOR2_X1 U4429 ( .A(n3675), .B(n2056), .ZN(n3676) );
  XNOR2_X1 U4430 ( .A(n3674), .B(n3676), .ZN(n3683) );
  AND2_X1 U4431 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4501) );
  AOI21_X1 U4432 ( .B1(n3695), .B2(n3677), .A(n4501), .ZN(n3679) );
  NAND2_X1 U4433 ( .A1(n3707), .A2(n4216), .ZN(n3678) );
  OAI211_X1 U4434 ( .C1(n3703), .C2(n3680), .A(n3679), .B(n3678), .ZN(n3681)
         );
  AOI21_X1 U4435 ( .B1(n3708), .B2(n4227), .A(n3681), .ZN(n3682) );
  OAI21_X1 U4436 ( .B1(n3683), .B2(n3711), .A(n3682), .ZN(U3235) );
  INV_X1 U4437 ( .A(n3685), .ZN(n3687) );
  NAND2_X1 U4438 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  XNOR2_X1 U4439 ( .A(n3684), .B(n3688), .ZN(n3697) );
  INV_X1 U4440 ( .A(n4073), .ZN(n3690) );
  NOR2_X1 U4441 ( .A1(n3690), .A2(n3689), .ZN(n3694) );
  NAND2_X1 U4442 ( .A1(n4065), .A2(n3707), .ZN(n3692) );
  NAND2_X1 U4443 ( .A1(U3149), .A2(REG3_REG_26__SCAN_IN), .ZN(n3691) );
  OAI211_X1 U4444 ( .C1(n3703), .C2(n4069), .A(n3692), .B(n3691), .ZN(n3693)
         );
  AOI211_X1 U4445 ( .C1(n3695), .C2(n4066), .A(n3694), .B(n3693), .ZN(n3696)
         );
  OAI21_X1 U4446 ( .B1(n3697), .B2(n3711), .A(n3696), .ZN(U3237) );
  INV_X1 U4447 ( .A(n3698), .ZN(n3700) );
  NAND2_X1 U4448 ( .A1(n3700), .A2(n3699), .ZN(n3702) );
  XNOR2_X1 U4449 ( .A(n3702), .B(n3701), .ZN(n3712) );
  AND2_X1 U4450 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n3970) );
  OAI22_X1 U4451 ( .A1(n3705), .A2(n3704), .B1(n3703), .B2(n4277), .ZN(n3706)
         );
  AOI211_X1 U4452 ( .C1(n3707), .C2(n4274), .A(n3970), .B(n3706), .ZN(n3710)
         );
  NAND2_X1 U4453 ( .A1(n3708), .A2(n4281), .ZN(n3709) );
  OAI211_X1 U4454 ( .C1(n3712), .C2(n3711), .A(n3710), .B(n3709), .ZN(U3238)
         );
  AND2_X1 U4455 ( .A1(n3717), .A2(DATAI_30_), .ZN(n4005) );
  INV_X1 U4456 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4688) );
  INV_X1 U4457 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4309) );
  OR2_X1 U4458 ( .A1(n2443), .A2(n4309), .ZN(n3714) );
  NAND2_X1 U4459 ( .A1(n3719), .A2(REG0_REG_31__SCAN_IN), .ZN(n3713) );
  OAI211_X1 U4460 ( .C1(n3722), .C2(n4688), .A(n3714), .B(n3713), .ZN(n4000)
         );
  INV_X1 U4461 ( .A(n4000), .ZN(n3748) );
  NAND2_X1 U4462 ( .A1(n3717), .A2(DATAI_29_), .ZN(n4026) );
  NAND2_X1 U4463 ( .A1(n3872), .A2(n4026), .ZN(n3718) );
  AND2_X1 U4464 ( .A1(n4016), .A2(n3718), .ZN(n3851) );
  INV_X1 U4465 ( .A(n4005), .ZN(n3749) );
  INV_X1 U4466 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4010) );
  INV_X1 U4467 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4315) );
  OR2_X1 U4468 ( .A1(n2443), .A2(n4315), .ZN(n3721) );
  NAND2_X1 U4469 ( .A1(n3719), .A2(REG0_REG_30__SCAN_IN), .ZN(n3720) );
  OAI211_X1 U4470 ( .C1(n3722), .C2(n4010), .A(n3721), .B(n3720), .ZN(n4020)
         );
  OR2_X1 U4471 ( .A1(n3872), .A2(n4026), .ZN(n3724) );
  NAND2_X1 U4472 ( .A1(n3723), .A2(DATAI_31_), .ZN(n4001) );
  NAND2_X1 U4473 ( .A1(n4001), .A2(n4000), .ZN(n3856) );
  OAI211_X1 U4474 ( .C1(n3749), .C2(n4020), .A(n3724), .B(n3856), .ZN(n3743)
         );
  AOI21_X1 U4475 ( .B1(n2030), .B2(n3851), .A(n3743), .ZN(n3852) );
  INV_X1 U4476 ( .A(n3725), .ZN(n3755) );
  NAND3_X1 U4477 ( .A1(n3851), .A2(n2160), .A3(n3755), .ZN(n3746) );
  NAND2_X1 U4478 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  NAND2_X1 U4479 ( .A1(n3728), .A2(n3730), .ZN(n3732) );
  INV_X1 U4480 ( .A(n3732), .ZN(n3829) );
  NAND2_X1 U4481 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  NAND2_X1 U4482 ( .A1(n3732), .A2(n3731), .ZN(n3832) );
  OAI211_X1 U4483 ( .C1(n3733), .C2(n3829), .A(n3836), .B(n3832), .ZN(n3735)
         );
  INV_X1 U4484 ( .A(n3837), .ZN(n3734) );
  AOI21_X1 U4485 ( .B1(n3735), .B2(n3833), .A(n3734), .ZN(n3739) );
  NAND2_X1 U4486 ( .A1(n3837), .A2(n3736), .ZN(n3738) );
  NAND2_X1 U4487 ( .A1(n3738), .A2(n3737), .ZN(n3839) );
  OAI21_X1 U4488 ( .B1(n3739), .B2(n3839), .A(n3843), .ZN(n3741) );
  NAND2_X1 U4489 ( .A1(n3741), .A2(n3740), .ZN(n3742) );
  AOI21_X1 U4490 ( .B1(n3742), .B2(n3845), .A(n4058), .ZN(n3744) );
  NOR4_X1 U4491 ( .A1(n3744), .A2(n2030), .A3(n3846), .A4(n3743), .ZN(n3745)
         );
  AOI21_X1 U4492 ( .B1(n3852), .B2(n3746), .A(n3745), .ZN(n3747) );
  AOI21_X1 U4493 ( .B1(n4005), .B2(n3748), .A(n3747), .ZN(n3752) );
  NAND2_X1 U4494 ( .A1(n3749), .A2(n4020), .ZN(n3855) );
  AOI21_X1 U4495 ( .B1(n3855), .B2(n4000), .A(n4001), .ZN(n3751) );
  NAND2_X1 U4496 ( .A1(n4059), .A2(n3753), .ZN(n4081) );
  NOR2_X1 U4497 ( .A1(n4011), .A2(n4081), .ZN(n3795) );
  INV_X1 U4498 ( .A(n4318), .ZN(n3794) );
  NAND2_X1 U4499 ( .A1(n3755), .A2(n3754), .ZN(n4062) );
  NOR2_X1 U4500 ( .A1(n4062), .A2(n2250), .ZN(n3793) );
  NAND2_X1 U4501 ( .A1(n3756), .A2(n4079), .ZN(n4100) );
  INV_X1 U4502 ( .A(n4100), .ZN(n3790) );
  INV_X1 U4503 ( .A(n4117), .ZN(n3840) );
  NAND2_X1 U4504 ( .A1(n3840), .A2(n4118), .ZN(n4157) );
  XNOR2_X1 U4505 ( .A(n4204), .B(n4177), .ZN(n4175) );
  INV_X1 U4506 ( .A(n4175), .ZN(n3767) );
  NAND4_X1 U4507 ( .A1(n2009), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  XNOR2_X1 U4508 ( .A(n4005), .B(n4020), .ZN(n3762) );
  NOR2_X1 U4509 ( .A1(n4001), .A2(n4000), .ZN(n3857) );
  INV_X1 U4510 ( .A(n3857), .ZN(n3760) );
  AND4_X1 U4511 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3856), .ZN(n3763)
         );
  NAND4_X1 U4512 ( .A1(n3764), .A2(n4293), .A3(n3815), .A4(n3763), .ZN(n3765)
         );
  NOR4_X1 U4513 ( .A1(n4157), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3789)
         );
  NAND2_X1 U4514 ( .A1(n4097), .A2(n3768), .ZN(n4122) );
  INV_X1 U4515 ( .A(n4122), .ZN(n3788) );
  NAND2_X1 U4516 ( .A1(n3770), .A2(n3769), .ZN(n4201) );
  INV_X1 U4517 ( .A(n4201), .ZN(n3780) );
  NOR2_X1 U4518 ( .A1(n3772), .A2(n3771), .ZN(n3778) );
  AND4_X1 U4519 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3777)
         );
  NAND4_X1 U4520 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3786)
         );
  INV_X1 U4521 ( .A(n4196), .ZN(n3781) );
  AND2_X1 U4522 ( .A1(n3781), .A2(n4195), .ZN(n4235) );
  NAND2_X1 U4523 ( .A1(n4576), .A2(n2893), .ZN(n3797) );
  AND2_X1 U4524 ( .A1(n3782), .A2(n3797), .ZN(n4578) );
  NOR2_X1 U4525 ( .A1(n4251), .A2(n3783), .ZN(n3784) );
  NAND4_X1 U4526 ( .A1(n4235), .A2(n4223), .A3(n4578), .A4(n3784), .ZN(n3785)
         );
  NOR2_X1 U4527 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  NAND4_X1 U4528 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3791)
         );
  NOR2_X1 U4529 ( .A1(n4045), .A2(n3791), .ZN(n3792) );
  NAND4_X1 U4530 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3862)
         );
  OAI211_X1 U4531 ( .C1(n3798), .C2(n2839), .A(n3797), .B(n3796), .ZN(n3801)
         );
  NAND3_X1 U4532 ( .A1(n3801), .A2(n3800), .A3(n3799), .ZN(n3804) );
  NAND3_X1 U4533 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3807) );
  NAND3_X1 U4534 ( .A1(n3807), .A2(n3806), .A3(n3805), .ZN(n3810) );
  NAND3_X1 U4535 ( .A1(n3810), .A2(n3809), .A3(n3808), .ZN(n3813) );
  AOI21_X1 U4536 ( .B1(n3813), .B2(n3812), .A(n2137), .ZN(n3819) );
  NAND2_X1 U4537 ( .A1(n3815), .A2(n3814), .ZN(n3818) );
  OAI211_X1 U4538 ( .C1(n3819), .C2(n3818), .A(n3817), .B(n3816), .ZN(n3822)
         );
  AND3_X1 U4539 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3825) );
  OAI21_X1 U4540 ( .B1(n3825), .B2(n3824), .A(n3823), .ZN(n3828) );
  NAND3_X1 U4541 ( .A1(n3828), .A2(n3827), .A3(n3826), .ZN(n3831) );
  AOI21_X1 U4542 ( .B1(n3831), .B2(n3830), .A(n3829), .ZN(n3835) );
  INV_X1 U4543 ( .A(n3832), .ZN(n3834) );
  OAI21_X1 U4544 ( .B1(n3835), .B2(n3834), .A(n3833), .ZN(n3838) );
  NAND3_X1 U4545 ( .A1(n3838), .A2(n3837), .A3(n3836), .ZN(n3842) );
  INV_X1 U4546 ( .A(n3839), .ZN(n3841) );
  NAND3_X1 U4547 ( .A1(n3842), .A2(n3841), .A3(n3840), .ZN(n3844) );
  NAND2_X1 U4548 ( .A1(n3844), .A2(n3843), .ZN(n3848) );
  AOI211_X1 U4549 ( .C1(n3848), .C2(n3847), .A(n3846), .B(n2158), .ZN(n3854)
         );
  NAND3_X1 U4550 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(n3853) );
  OAI21_X1 U4551 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n3860) );
  INV_X1 U4552 ( .A(n3855), .ZN(n3858) );
  OAI21_X1 U4553 ( .B1(n3858), .B2(n3857), .A(n3856), .ZN(n3859) );
  NAND2_X1 U4554 ( .A1(n3860), .A2(n3859), .ZN(n3861) );
  MUX2_X1 U4555 ( .A(n3862), .B(n3861), .S(n2367), .Z(n3863) );
  NAND2_X1 U4556 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  XNOR2_X1 U4557 ( .A(n3865), .B(n3978), .ZN(n3871) );
  NOR2_X1 U4558 ( .A1(n3867), .A2(n3866), .ZN(n3869) );
  OAI21_X1 U4559 ( .B1(n3870), .B2(n2838), .A(B_REG_SCAN_IN), .ZN(n3868) );
  OAI22_X1 U4560 ( .A1(n3871), .A2(n3870), .B1(n3869), .B2(n3868), .ZN(U3239)
         );
  MUX2_X1 U4561 ( .A(DATAO_REG_31__SCAN_IN), .B(n4000), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4562 ( .A(DATAO_REG_30__SCAN_IN), .B(n4020), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4563 ( .A(DATAO_REG_29__SCAN_IN), .B(n3872), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4564 ( .A(DATAO_REG_28__SCAN_IN), .B(n4014), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4565 ( .A(DATAO_REG_26__SCAN_IN), .B(n3873), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4566 ( .A(DATAO_REG_24__SCAN_IN), .B(n4084), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4567 ( .A(DATAO_REG_23__SCAN_IN), .B(n4103), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4568 ( .A(DATAO_REG_22__SCAN_IN), .B(n3874), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4569 ( .A(n4143), .B(DATAO_REG_21__SCAN_IN), .S(n3875), .Z(U3571)
         );
  MUX2_X1 U4570 ( .A(n4216), .B(DATAO_REG_19__SCAN_IN), .S(n3875), .Z(U3569)
         );
  MUX2_X1 U4571 ( .A(n4239), .B(DATAO_REG_18__SCAN_IN), .S(n3875), .Z(U3568)
         );
  MUX2_X1 U4572 ( .A(DATAO_REG_16__SCAN_IN), .B(n4274), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4573 ( .A(DATAO_REG_15__SCAN_IN), .B(n4262), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4574 ( .A(DATAO_REG_14__SCAN_IN), .B(n4271), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4575 ( .A(DATAO_REG_13__SCAN_IN), .B(n3876), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4576 ( .A(DATAO_REG_12__SCAN_IN), .B(n3877), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4577 ( .A(DATAO_REG_11__SCAN_IN), .B(n3878), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4578 ( .A(DATAO_REG_9__SCAN_IN), .B(n3879), .S(U4043), .Z(U3559) );
  MUX2_X1 U4579 ( .A(DATAO_REG_8__SCAN_IN), .B(n3880), .S(U4043), .Z(U3558) );
  MUX2_X1 U4580 ( .A(DATAO_REG_6__SCAN_IN), .B(n3881), .S(U4043), .Z(U3556) );
  MUX2_X1 U4581 ( .A(DATAO_REG_5__SCAN_IN), .B(n3882), .S(U4043), .Z(U3555) );
  MUX2_X1 U4582 ( .A(DATAO_REG_4__SCAN_IN), .B(n2898), .S(U4043), .Z(U3554) );
  MUX2_X1 U4583 ( .A(DATAO_REG_2__SCAN_IN), .B(n3883), .S(U4043), .Z(U3552) );
  MUX2_X1 U4584 ( .A(DATAO_REG_1__SCAN_IN), .B(n2894), .S(U4043), .Z(U3551) );
  MUX2_X1 U4585 ( .A(DATAO_REG_0__SCAN_IN), .B(n2893), .S(U4043), .Z(U3550) );
  AND2_X1 U4586 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3885)
         );
  OAI211_X1 U4587 ( .C1(n3885), .C2(n3884), .A(n4494), .B(n3900), .ZN(n3892)
         );
  OAI211_X1 U4588 ( .C1(n3887), .C2(n3886), .A(n4510), .B(n3895), .ZN(n3891)
         );
  AOI22_X1 U4589 ( .A1(n4500), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3890) );
  INV_X1 U4590 ( .A(n4514), .ZN(n3905) );
  NAND2_X1 U4591 ( .A1(n3905), .A2(n3888), .ZN(n3889) );
  NAND4_X1 U4592 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(U3241)
         );
  NAND3_X1 U4593 ( .A1(n3895), .A2(n3894), .A3(n3893), .ZN(n3896) );
  NAND2_X1 U4594 ( .A1(n2046), .A2(n3896), .ZN(n3897) );
  NOR2_X1 U4595 ( .A1(n3939), .A2(n3897), .ZN(n3904) );
  AND3_X1 U4596 ( .A1(n3900), .A2(n3899), .A3(n3898), .ZN(n3901) );
  NOR3_X1 U4597 ( .A1(n4497), .A2(n3902), .A3(n3901), .ZN(n3903) );
  AOI211_X1 U4598 ( .C1(n3905), .C2(n4465), .A(n3904), .B(n3903), .ZN(n3908)
         );
  AOI22_X1 U4599 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4500), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3907) );
  NAND3_X1 U4600 ( .A1(n3908), .A2(n3907), .A3(n3906), .ZN(U3242) );
  XNOR2_X1 U4601 ( .A(n3925), .B(REG2_REG_12__SCAN_IN), .ZN(n3920) );
  INV_X1 U4602 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4389) );
  OAI211_X1 U4603 ( .C1(n3915), .C2(REG1_REG_12__SCAN_IN), .A(n3933), .B(n4494), .ZN(n3918) );
  AOI21_X1 U4604 ( .B1(n4500), .B2(ADDR_REG_12__SCAN_IN), .A(n3916), .ZN(n3917) );
  OAI211_X1 U4605 ( .C1(n4514), .C2(n3931), .A(n3918), .B(n3917), .ZN(n3919)
         );
  AOI21_X1 U4606 ( .B1(n4510), .B2(n3920), .A(n3919), .ZN(n3921) );
  INV_X1 U4607 ( .A(n3921), .ZN(U3252) );
  INV_X1 U4608 ( .A(n3922), .ZN(n3923) );
  INV_X1 U4609 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3926) );
  NOR2_X1 U4610 ( .A1(n3934), .A2(n3926), .ZN(n3941) );
  AOI21_X1 U4611 ( .B1(n3926), .B2(n3934), .A(n3941), .ZN(n3927) );
  XNOR2_X1 U4612 ( .A(n3942), .B(n3927), .ZN(n3940) );
  NOR2_X1 U4613 ( .A1(n4514), .A2(n3934), .ZN(n3928) );
  AOI211_X1 U4614 ( .C1(n4500), .C2(ADDR_REG_13__SCAN_IN), .A(n3929), .B(n3928), .ZN(n3938) );
  NAND2_X1 U4615 ( .A1(n3930), .A2(n3912), .ZN(n3932) );
  XNOR2_X1 U4616 ( .A(n3934), .B(REG1_REG_13__SCAN_IN), .ZN(n3935) );
  OAI211_X1 U4617 ( .C1(n3936), .C2(n3935), .A(n3948), .B(n4494), .ZN(n3937)
         );
  OAI211_X1 U4618 ( .C1(n3940), .C2(n3939), .A(n3938), .B(n3937), .ZN(U3253)
         );
  XNOR2_X1 U4619 ( .A(n3954), .B(n3963), .ZN(n3943) );
  NAND2_X1 U4620 ( .A1(n3943), .A2(REG2_REG_14__SCAN_IN), .ZN(n3957) );
  OAI211_X1 U4621 ( .C1(n3943), .C2(REG2_REG_14__SCAN_IN), .A(n3957), .B(n4510), .ZN(n3953) );
  NOR2_X1 U4622 ( .A1(n4514), .A2(n3949), .ZN(n3944) );
  AOI211_X1 U4623 ( .C1(n4500), .C2(ADDR_REG_14__SCAN_IN), .A(n3945), .B(n3944), .ZN(n3952) );
  NAND2_X1 U4624 ( .A1(n3946), .A2(REG1_REG_13__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U4625 ( .A1(n3948), .A2(n3947), .ZN(n3964) );
  OAI211_X1 U4626 ( .C1(n3950), .C2(REG1_REG_14__SCAN_IN), .A(n3966), .B(n4494), .ZN(n3951) );
  NAND3_X1 U4627 ( .A1(n3953), .A2(n3952), .A3(n3951), .ZN(U3254) );
  INV_X1 U4628 ( .A(n4457), .ZN(n3982) );
  XNOR2_X1 U4629 ( .A(n4457), .B(REG2_REG_15__SCAN_IN), .ZN(n3961) );
  INV_X1 U4630 ( .A(n3954), .ZN(n3955) );
  NAND2_X1 U4631 ( .A1(n3955), .A2(n3963), .ZN(n3956) );
  INV_X1 U4632 ( .A(n3959), .ZN(n3960) );
  INV_X1 U4633 ( .A(n3961), .ZN(n3958) );
  AOI21_X1 U4634 ( .B1(n3961), .B2(n3960), .A(n2027), .ZN(n3962) );
  NAND2_X1 U4635 ( .A1(n4510), .A2(n3962), .ZN(n3972) );
  NAND2_X1 U4636 ( .A1(n3964), .A2(n3963), .ZN(n3965) );
  XNOR2_X1 U4637 ( .A(n4457), .B(REG1_REG_15__SCAN_IN), .ZN(n3967) );
  AOI211_X1 U4638 ( .C1(n3968), .C2(n3967), .A(n3974), .B(n4497), .ZN(n3969)
         );
  AOI211_X1 U4639 ( .C1(n4500), .C2(ADDR_REG_15__SCAN_IN), .A(n3970), .B(n3969), .ZN(n3971) );
  OAI211_X1 U4640 ( .C1(n3982), .C2(n4514), .A(n3972), .B(n3971), .ZN(U3255)
         );
  AOI22_X1 U4641 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4513), .B1(n4540), .B2(
        n3973), .ZN(n4498) );
  AOI22_X1 U4642 ( .A1(n3985), .A2(REG1_REG_17__SCAN_IN), .B1(n4367), .B2(
        n4542), .ZN(n4488) );
  NAND2_X1 U4643 ( .A1(n3975), .A2(n4543), .ZN(n3977) );
  NAND2_X1 U4644 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  XNOR2_X1 U4645 ( .A(n3978), .B(REG1_REG_19__SCAN_IN), .ZN(n3979) );
  XNOR2_X1 U4646 ( .A(n3980), .B(n3979), .ZN(n3997) );
  NAND2_X1 U4647 ( .A1(n3983), .A2(n4543), .ZN(n3984) );
  INV_X1 U4648 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U4649 ( .A1(n4480), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U4650 ( .A1(n3984), .A2(n4478), .ZN(n4490) );
  NOR2_X1 U4651 ( .A1(n3985), .A2(REG2_REG_17__SCAN_IN), .ZN(n3986) );
  AOI21_X1 U4652 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3985), .A(n3986), .ZN(n4491) );
  INV_X1 U4653 ( .A(n3986), .ZN(n3987) );
  NAND2_X1 U4654 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4540), .ZN(n3988) );
  OAI21_X1 U4655 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4540), .A(n3988), .ZN(n4508) );
  INV_X1 U4656 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3989) );
  MUX2_X1 U4657 ( .A(n3989), .B(REG2_REG_19__SCAN_IN), .S(n4526), .Z(n3990) );
  XNOR2_X1 U4658 ( .A(n3991), .B(n3990), .ZN(n3995) );
  NAND2_X1 U4659 ( .A1(n4500), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3992) );
  OAI211_X1 U4660 ( .C1(n4514), .C2(n4526), .A(n3993), .B(n3992), .ZN(n3994)
         );
  AOI21_X1 U4661 ( .B1(n3995), .B2(n4510), .A(n3994), .ZN(n3996) );
  OAI21_X1 U4662 ( .B1(n3997), .B2(n4497), .A(n3996), .ZN(U3259) );
  NAND2_X1 U4663 ( .A1(n3998), .A2(n4026), .ZN(n4030) );
  XNOR2_X1 U4664 ( .A(n4004), .B(n4001), .ZN(n4395) );
  NAND2_X1 U4665 ( .A1(n4467), .A2(B_REG_SCAN_IN), .ZN(n3999) );
  AND2_X1 U4666 ( .A1(n4273), .A2(n3999), .ZN(n4021) );
  NAND2_X1 U4667 ( .A1(n4021), .A2(n4000), .ZN(n4007) );
  OAI21_X1 U4668 ( .B1(n4001), .B2(n4278), .A(n4007), .ZN(n4392) );
  NAND2_X1 U4669 ( .A1(n4535), .A2(n4392), .ZN(n4003) );
  NAND2_X1 U4670 ( .A1(n2003), .A2(REG2_REG_31__SCAN_IN), .ZN(n4002) );
  OAI211_X1 U4671 ( .C1(n4395), .C2(n4305), .A(n4003), .B(n4002), .ZN(U3260)
         );
  AOI21_X1 U4672 ( .B1(n4005), .B2(n4030), .A(n4004), .ZN(n4396) );
  NAND2_X1 U4673 ( .A1(n4396), .A2(n4516), .ZN(n4009) );
  NAND2_X1 U4674 ( .A1(n4525), .A2(n4005), .ZN(n4006) );
  NAND2_X1 U4675 ( .A1(n4007), .A2(n4006), .ZN(n4397) );
  NAND2_X1 U4676 ( .A1(n4535), .A2(n4397), .ZN(n4008) );
  OAI211_X1 U4677 ( .C1(n4535), .C2(n4010), .A(n4009), .B(n4008), .ZN(U3261)
         );
  NAND2_X1 U4678 ( .A1(n4012), .A2(n4011), .ZN(n4316) );
  NAND2_X1 U4679 ( .A1(n4014), .A2(n4013), .ZN(n4319) );
  NAND2_X1 U4680 ( .A1(n4316), .A2(n4319), .ZN(n4015) );
  XNOR2_X1 U4681 ( .A(n4015), .B(n4318), .ZN(n4035) );
  NAND2_X1 U4682 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  XNOR2_X1 U4683 ( .A(n4018), .B(n4318), .ZN(n4024) );
  NOR2_X1 U4684 ( .A1(n4278), .A2(n4026), .ZN(n4019) );
  AOI21_X1 U4685 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4022) );
  OAI21_X1 U4686 ( .B1(n4041), .B2(n4288), .A(n4022), .ZN(n4023) );
  AOI21_X1 U4687 ( .B1(n4024), .B2(n4270), .A(n4023), .ZN(n4323) );
  OAI21_X1 U4688 ( .B1(n4025), .B2(n4255), .A(n4323), .ZN(n4033) );
  INV_X1 U4689 ( .A(n4026), .ZN(n4027) );
  NAND2_X1 U4690 ( .A1(n4028), .A2(n4027), .ZN(n4029) );
  INV_X1 U4691 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4031) );
  OAI22_X1 U4692 ( .A1(n4317), .A2(n4305), .B1(n4031), .B2(n4535), .ZN(n4032)
         );
  AOI21_X1 U4693 ( .B1(n4535), .B2(n4033), .A(n4032), .ZN(n4034) );
  OAI21_X1 U4694 ( .B1(n4035), .B2(n4286), .A(n4034), .ZN(U3354) );
  NAND2_X1 U4695 ( .A1(n4036), .A2(n4045), .ZN(n4037) );
  NAND2_X1 U4696 ( .A1(n4038), .A2(n4037), .ZN(n4043) );
  OAI22_X1 U4697 ( .A1(n4087), .A2(n4288), .B1(n4048), .B2(n4278), .ZN(n4039)
         );
  INV_X1 U4698 ( .A(n4039), .ZN(n4040) );
  OAI21_X1 U4699 ( .B1(n4041), .B2(n4521), .A(n4040), .ZN(n4042) );
  AOI21_X1 U4700 ( .B1(n4043), .B2(n4270), .A(n4042), .ZN(n4327) );
  XNOR2_X1 U4701 ( .A(n4044), .B(n4045), .ZN(n4326) );
  NAND2_X1 U4702 ( .A1(n4326), .A2(n4231), .ZN(n4054) );
  NOR2_X1 U4703 ( .A1(n4046), .A2(n4255), .ZN(n4052) );
  OR2_X1 U4704 ( .A1(n4047), .A2(n4048), .ZN(n4049) );
  NAND2_X1 U4705 ( .A1(n4050), .A2(n4049), .ZN(n4329) );
  NOR2_X1 U4706 ( .A1(n4329), .A2(n4305), .ZN(n4051) );
  AOI211_X1 U4707 ( .C1(n2003), .C2(REG2_REG_27__SCAN_IN), .A(n4052), .B(n4051), .ZN(n4053) );
  OAI211_X1 U4708 ( .C1(n4327), .C2(n2003), .A(n4054), .B(n4053), .ZN(U3263)
         );
  XOR2_X1 U4709 ( .A(n4062), .B(n4055), .Z(n4331) );
  NOR2_X1 U4710 ( .A1(n4056), .A2(n4069), .ZN(n4057) );
  OR2_X1 U4711 ( .A1(n4047), .A2(n4057), .ZN(n4406) );
  INV_X1 U4712 ( .A(n4058), .ZN(n4061) );
  INV_X1 U4713 ( .A(n4059), .ZN(n4060) );
  AOI21_X1 U4714 ( .B1(n4080), .B2(n4061), .A(n4060), .ZN(n4063) );
  XNOR2_X1 U4715 ( .A(n4063), .B(n4062), .ZN(n4064) );
  NAND2_X1 U4716 ( .A1(n4064), .A2(n4270), .ZN(n4072) );
  NAND2_X1 U4717 ( .A1(n4065), .A2(n4273), .ZN(n4068) );
  NAND2_X1 U4718 ( .A1(n4066), .A2(n4272), .ZN(n4067) );
  OAI211_X1 U4719 ( .C1(n4278), .C2(n4069), .A(n4068), .B(n4067), .ZN(n4070)
         );
  INV_X1 U4720 ( .A(n4070), .ZN(n4071) );
  NAND2_X1 U4721 ( .A1(n4072), .A2(n4071), .ZN(n4330) );
  NAND2_X1 U4722 ( .A1(n4330), .A2(n4535), .ZN(n4075) );
  AOI22_X1 U4723 ( .A1(n4073), .A2(n4530), .B1(REG2_REG_26__SCAN_IN), .B2(
        n2003), .ZN(n4074) );
  OAI211_X1 U4724 ( .C1(n4305), .C2(n4406), .A(n4075), .B(n4074), .ZN(n4076)
         );
  AOI21_X1 U4725 ( .B1(n4331), .B2(n4231), .A(n4076), .ZN(n4077) );
  INV_X1 U4726 ( .A(n4077), .ZN(U3264) );
  XNOR2_X1 U4727 ( .A(n4078), .B(n4081), .ZN(n4335) );
  INV_X1 U4728 ( .A(n4335), .ZN(n4095) );
  NAND2_X1 U4729 ( .A1(n4080), .A2(n4079), .ZN(n4082) );
  XNOR2_X1 U4730 ( .A(n4082), .B(n4081), .ZN(n4083) );
  NAND2_X1 U4731 ( .A1(n4083), .A2(n4270), .ZN(n4086) );
  AOI22_X1 U4732 ( .A1(n4084), .A2(n4272), .B1(n4088), .B2(n4525), .ZN(n4085)
         );
  OAI211_X1 U4733 ( .C1(n4087), .C2(n4521), .A(n4086), .B(n4085), .ZN(n4334)
         );
  INV_X1 U4734 ( .A(n4056), .ZN(n4090) );
  NAND2_X1 U4735 ( .A1(n4109), .A2(n4088), .ZN(n4089) );
  NAND2_X1 U4736 ( .A1(n4090), .A2(n4089), .ZN(n4410) );
  AOI22_X1 U4737 ( .A1(n4091), .A2(n4530), .B1(REG2_REG_25__SCAN_IN), .B2(
        n2003), .ZN(n4092) );
  OAI21_X1 U4738 ( .B1(n4410), .B2(n4305), .A(n4092), .ZN(n4093) );
  AOI21_X1 U4739 ( .B1(n4535), .B2(n4334), .A(n4093), .ZN(n4094) );
  OAI21_X1 U4740 ( .B1(n4095), .B2(n4286), .A(n4094), .ZN(U3265) );
  XOR2_X1 U4741 ( .A(n4100), .B(n4096), .Z(n4339) );
  INV_X1 U4742 ( .A(n4339), .ZN(n4115) );
  NAND2_X1 U4743 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  XOR2_X1 U4744 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND2_X1 U4745 ( .A1(n4101), .A2(n4270), .ZN(n4105) );
  AOI22_X1 U4746 ( .A1(n4103), .A2(n4272), .B1(n4102), .B2(n4525), .ZN(n4104)
         );
  OAI211_X1 U4747 ( .C1(n4106), .C2(n4521), .A(n4105), .B(n4104), .ZN(n4338)
         );
  OAI22_X1 U4748 ( .A1(n4108), .A2(n4255), .B1(n4107), .B2(n4535), .ZN(n4113)
         );
  INV_X1 U4749 ( .A(n4132), .ZN(n4111) );
  OAI21_X1 U4750 ( .B1(n4111), .B2(n4110), .A(n4109), .ZN(n4414) );
  NOR2_X1 U4751 ( .A1(n4414), .A2(n4305), .ZN(n4112) );
  AOI211_X1 U4752 ( .C1(n4338), .C2(n4535), .A(n4113), .B(n4112), .ZN(n4114)
         );
  OAI21_X1 U4753 ( .B1(n4115), .B2(n4286), .A(n4114), .ZN(U3266) );
  XOR2_X1 U4754 ( .A(n4122), .B(n4116), .Z(n4343) );
  INV_X1 U4755 ( .A(n4343), .ZN(n4138) );
  OR2_X1 U4756 ( .A1(n4158), .A2(n4117), .ZN(n4119) );
  NAND2_X1 U4757 ( .A1(n4119), .A2(n4118), .ZN(n4141) );
  NAND2_X1 U4758 ( .A1(n4141), .A2(n4142), .ZN(n4140) );
  NAND2_X1 U4759 ( .A1(n4140), .A2(n4120), .ZN(n4121) );
  XOR2_X1 U4760 ( .A(n4122), .B(n4121), .Z(n4127) );
  NOR2_X1 U4761 ( .A1(n4162), .A2(n4288), .ZN(n4126) );
  OAI22_X1 U4762 ( .A1(n4124), .A2(n4521), .B1(n4278), .B2(n4123), .ZN(n4125)
         );
  AOI211_X1 U4763 ( .C1(n4127), .C2(n4270), .A(n4126), .B(n4125), .ZN(n4128)
         );
  INV_X1 U4764 ( .A(n4128), .ZN(n4342) );
  NAND2_X1 U4765 ( .A1(n4129), .A2(n4130), .ZN(n4131) );
  NAND2_X1 U4766 ( .A1(n4132), .A2(n4131), .ZN(n4418) );
  INV_X1 U4767 ( .A(n4133), .ZN(n4134) );
  AOI22_X1 U4768 ( .A1(REG2_REG_23__SCAN_IN), .A2(n2003), .B1(n4134), .B2(
        n4530), .ZN(n4135) );
  OAI21_X1 U4769 ( .B1(n4418), .B2(n4305), .A(n4135), .ZN(n4136) );
  AOI21_X1 U4770 ( .B1(n4342), .B2(n4535), .A(n4136), .ZN(n4137) );
  OAI21_X1 U4771 ( .B1(n4138), .B2(n4286), .A(n4137), .ZN(U3267) );
  OAI21_X1 U4772 ( .B1(n2022), .B2(n2250), .A(n4139), .ZN(n4348) );
  OAI21_X1 U4773 ( .B1(n4142), .B2(n4141), .A(n4140), .ZN(n4149) );
  NAND2_X1 U4774 ( .A1(n4143), .A2(n4272), .ZN(n4146) );
  NAND2_X1 U4775 ( .A1(n4525), .A2(n4144), .ZN(n4145) );
  OAI211_X1 U4776 ( .C1(n4147), .C2(n4521), .A(n4146), .B(n4145), .ZN(n4148)
         );
  AOI21_X1 U4777 ( .B1(n4149), .B2(n4270), .A(n4148), .ZN(n4347) );
  AOI22_X1 U4778 ( .A1(n2003), .A2(REG2_REG_22__SCAN_IN), .B1(n4150), .B2(
        n4530), .ZN(n4153) );
  OR2_X1 U4779 ( .A1(n4164), .A2(n4151), .ZN(n4345) );
  NAND3_X1 U4780 ( .A1(n4129), .A2(n4345), .A3(n4516), .ZN(n4152) );
  OAI211_X1 U4781 ( .C1(n4347), .C2(n2003), .A(n4153), .B(n4152), .ZN(n4154)
         );
  INV_X1 U4782 ( .A(n4154), .ZN(n4155) );
  OAI21_X1 U4783 ( .B1(n4348), .B2(n4286), .A(n4155), .ZN(U3268) );
  XOR2_X1 U4784 ( .A(n4157), .B(n4156), .Z(n4350) );
  INV_X1 U4785 ( .A(n4350), .ZN(n4170) );
  XNOR2_X1 U4786 ( .A(n4158), .B(n4157), .ZN(n4159) );
  NAND2_X1 U4787 ( .A1(n4159), .A2(n4270), .ZN(n4161) );
  AOI22_X1 U4788 ( .A1(n4204), .A2(n4272), .B1(n4163), .B2(n4525), .ZN(n4160)
         );
  OAI211_X1 U4789 ( .C1(n4162), .C2(n4521), .A(n4161), .B(n4160), .ZN(n4349)
         );
  AND2_X1 U4790 ( .A1(n4184), .A2(n4163), .ZN(n4165) );
  OR2_X1 U4791 ( .A1(n4165), .A2(n4164), .ZN(n4423) );
  AOI22_X1 U4792 ( .A1(n2003), .A2(REG2_REG_21__SCAN_IN), .B1(n4166), .B2(
        n4530), .ZN(n4167) );
  OAI21_X1 U4793 ( .B1(n4423), .B2(n4305), .A(n4167), .ZN(n4168) );
  AOI21_X1 U4794 ( .B1(n4349), .B2(n4535), .A(n4168), .ZN(n4169) );
  OAI21_X1 U4795 ( .B1(n4170), .B2(n4286), .A(n4169), .ZN(U3269) );
  XNOR2_X1 U4796 ( .A(n4171), .B(n4175), .ZN(n4353) );
  INV_X1 U4797 ( .A(n4172), .ZN(n4173) );
  NAND2_X1 U4798 ( .A1(n4174), .A2(n4173), .ZN(n4176) );
  XNOR2_X1 U4799 ( .A(n4176), .B(n4175), .ZN(n4181) );
  AOI22_X1 U4800 ( .A1(n4216), .A2(n4272), .B1(n4177), .B2(n4525), .ZN(n4178)
         );
  OAI21_X1 U4801 ( .B1(n4179), .B2(n4521), .A(n4178), .ZN(n4180) );
  AOI21_X1 U4802 ( .B1(n4181), .B2(n4270), .A(n4180), .ZN(n4182) );
  OAI21_X1 U4803 ( .B1(n4353), .B2(n4528), .A(n4182), .ZN(n4354) );
  NAND2_X1 U4804 ( .A1(n4354), .A2(n4535), .ZN(n4192) );
  INV_X1 U4805 ( .A(n4183), .ZN(n4186) );
  OAI21_X1 U4806 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4427) );
  INV_X1 U4807 ( .A(n4427), .ZN(n4190) );
  OAI22_X1 U4808 ( .A1(n4535), .A2(n4188), .B1(n4187), .B2(n4255), .ZN(n4189)
         );
  AOI21_X1 U4809 ( .B1(n4190), .B2(n4516), .A(n4189), .ZN(n4191) );
  OAI211_X1 U4810 ( .C1(n4353), .C2(n4193), .A(n4192), .B(n4191), .ZN(U3270)
         );
  XNOR2_X1 U4811 ( .A(n4194), .B(n4201), .ZN(n4359) );
  INV_X1 U4812 ( .A(n4359), .ZN(n4214) );
  OAI21_X1 U4813 ( .B1(n4236), .B2(n4196), .A(n4195), .ZN(n4215) );
  INV_X1 U4814 ( .A(n4197), .ZN(n4199) );
  OAI21_X1 U4815 ( .B1(n4215), .B2(n4199), .A(n4198), .ZN(n4200) );
  XOR2_X1 U4816 ( .A(n4201), .B(n4200), .Z(n4206) );
  OAI22_X1 U4817 ( .A1(n4202), .A2(n4288), .B1(n4278), .B2(n4207), .ZN(n4203)
         );
  AOI21_X1 U4818 ( .B1(n4273), .B2(n4204), .A(n4203), .ZN(n4205) );
  OAI21_X1 U4819 ( .B1(n4206), .B2(n4523), .A(n4205), .ZN(n4358) );
  OR2_X1 U4820 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  NAND2_X1 U4821 ( .A1(n4183), .A2(n4209), .ZN(n4430) );
  NOR2_X1 U4822 ( .A1(n4430), .A2(n4305), .ZN(n4212) );
  OAI22_X1 U4823 ( .A1(n4535), .A2(n3989), .B1(n4210), .B2(n4255), .ZN(n4211)
         );
  AOI211_X1 U4824 ( .C1(n4358), .C2(n4535), .A(n4212), .B(n4211), .ZN(n4213)
         );
  OAI21_X1 U4825 ( .B1(n4214), .B2(n4286), .A(n4213), .ZN(U3271) );
  XNOR2_X1 U4826 ( .A(n4215), .B(n4223), .ZN(n4219) );
  AOI22_X1 U4827 ( .A1(n4216), .A2(n4273), .B1(n4225), .B2(n4525), .ZN(n4217)
         );
  OAI21_X1 U4828 ( .B1(n4265), .B2(n4288), .A(n4217), .ZN(n4218) );
  AOI21_X1 U4829 ( .B1(n4219), .B2(n4270), .A(n4218), .ZN(n4363) );
  INV_X1 U4830 ( .A(n4221), .ZN(n4222) );
  AOI21_X1 U4831 ( .B1(n4223), .B2(n4220), .A(n4222), .ZN(n4364) );
  INV_X1 U4832 ( .A(n4364), .ZN(n4232) );
  XNOR2_X1 U4833 ( .A(n4224), .B(n4225), .ZN(n4226) );
  NAND2_X1 U4834 ( .A1(n4226), .A2(n2998), .ZN(n4362) );
  AOI22_X1 U4835 ( .A1(n2003), .A2(REG2_REG_18__SCAN_IN), .B1(n4227), .B2(
        n4530), .ZN(n4228) );
  OAI21_X1 U4836 ( .B1(n4362), .B2(n4229), .A(n4228), .ZN(n4230) );
  AOI21_X1 U4837 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(n4233) );
  OAI21_X1 U4838 ( .B1(n2003), .B2(n4363), .A(n4233), .ZN(U3272) );
  XNOR2_X1 U4839 ( .A(n4234), .B(n4235), .ZN(n4366) );
  INV_X1 U4840 ( .A(n4366), .ZN(n4249) );
  XNOR2_X1 U4841 ( .A(n4236), .B(n4235), .ZN(n4241) );
  OAI22_X1 U4842 ( .A1(n4237), .A2(n4288), .B1(n4278), .B2(n4244), .ZN(n4238)
         );
  AOI21_X1 U4843 ( .B1(n4273), .B2(n4239), .A(n4238), .ZN(n4240) );
  OAI21_X1 U4844 ( .B1(n4241), .B2(n4523), .A(n4240), .ZN(n4365) );
  INV_X1 U4845 ( .A(n4242), .ZN(n4253) );
  INV_X1 U4846 ( .A(n4224), .ZN(n4243) );
  OAI21_X1 U4847 ( .B1(n4253), .B2(n4244), .A(n4243), .ZN(n4435) );
  AOI22_X1 U4848 ( .A1(n2003), .A2(REG2_REG_17__SCAN_IN), .B1(n4245), .B2(
        n4530), .ZN(n4246) );
  OAI21_X1 U4849 ( .B1(n4435), .B2(n4305), .A(n4246), .ZN(n4247) );
  AOI21_X1 U4850 ( .B1(n4365), .B2(n4535), .A(n4247), .ZN(n4248) );
  OAI21_X1 U4851 ( .B1(n4249), .B2(n4286), .A(n4248), .ZN(U3273) );
  OAI21_X1 U4852 ( .B1(n4252), .B2(n4251), .A(n4250), .ZN(n4372) );
  AOI21_X1 U4853 ( .B1(n4261), .B2(n4254), .A(n4253), .ZN(n4370) );
  OAI22_X1 U4854 ( .A1(n4535), .A2(n4479), .B1(n4256), .B2(n4255), .ZN(n4257)
         );
  AOI21_X1 U4855 ( .B1(n4370), .B2(n4516), .A(n4257), .ZN(n4267) );
  OAI211_X1 U4856 ( .C1(n4260), .C2(n4259), .A(n4258), .B(n4270), .ZN(n4264)
         );
  AOI22_X1 U4857 ( .A1(n4262), .A2(n4272), .B1(n4261), .B2(n4525), .ZN(n4263)
         );
  OAI211_X1 U4858 ( .C1(n4265), .C2(n4521), .A(n4264), .B(n4263), .ZN(n4369)
         );
  NAND2_X1 U4859 ( .A1(n4369), .A2(n4535), .ZN(n4266) );
  OAI211_X1 U4860 ( .C1(n4372), .C2(n4286), .A(n4267), .B(n4266), .ZN(U3274)
         );
  XNOR2_X1 U4861 ( .A(n4268), .B(n2009), .ZN(n4376) );
  OAI211_X1 U4862 ( .C1(n2025), .C2(n2009), .A(n4270), .B(n4269), .ZN(n4276)
         );
  AOI22_X1 U4863 ( .A1(n4274), .A2(n4273), .B1(n4272), .B2(n4271), .ZN(n4275)
         );
  OAI211_X1 U4864 ( .C1(n4278), .C2(n4277), .A(n4276), .B(n4275), .ZN(n4373)
         );
  XNOR2_X1 U4865 ( .A(n4280), .B(n4279), .ZN(n4374) );
  INV_X1 U4866 ( .A(n4374), .ZN(n4283) );
  AOI22_X1 U4867 ( .A1(n2003), .A2(REG2_REG_15__SCAN_IN), .B1(n4281), .B2(
        n4530), .ZN(n4282) );
  OAI21_X1 U4868 ( .B1(n4283), .B2(n4305), .A(n4282), .ZN(n4284) );
  AOI21_X1 U4869 ( .B1(n4373), .B2(n4535), .A(n4284), .ZN(n4285) );
  OAI21_X1 U4870 ( .B1(n4376), .B2(n4286), .A(n4285), .ZN(U3275) );
  XOR2_X1 U4871 ( .A(n4287), .B(n4293), .Z(n4298) );
  OAI22_X1 U4872 ( .A1(n4289), .A2(n4521), .B1(n4288), .B2(n2913), .ZN(n4295)
         );
  INV_X1 U4873 ( .A(n4291), .ZN(n4292) );
  AOI21_X1 U4874 ( .B1(n4293), .B2(n4290), .A(n4292), .ZN(n4299) );
  NOR2_X1 U4875 ( .A1(n4299), .A2(n4528), .ZN(n4294) );
  AOI211_X1 U4876 ( .C1(n4525), .C2(n4296), .A(n4295), .B(n4294), .ZN(n4297)
         );
  OAI21_X1 U4877 ( .B1(n4523), .B2(n4298), .A(n4297), .ZN(n4387) );
  INV_X1 U4878 ( .A(n4387), .ZN(n4308) );
  INV_X1 U4879 ( .A(n4299), .ZN(n4388) );
  OR2_X1 U4880 ( .A1(n4301), .A2(n4300), .ZN(n4302) );
  NAND2_X1 U4881 ( .A1(n3474), .A2(n4302), .ZN(n4452) );
  AOI22_X1 U4882 ( .A1(n2003), .A2(REG2_REG_11__SCAN_IN), .B1(n4303), .B2(
        n4530), .ZN(n4304) );
  OAI21_X1 U4883 ( .B1(n4452), .B2(n4305), .A(n4304), .ZN(n4306) );
  AOI21_X1 U4884 ( .B1(n4388), .B2(n4532), .A(n4306), .ZN(n4307) );
  OAI21_X1 U4885 ( .B1(n4308), .B2(n2003), .A(n4307), .ZN(U3279) );
  NOR2_X1 U4886 ( .A1(n4589), .A2(n4309), .ZN(n4310) );
  AOI21_X1 U4887 ( .B1(n4589), .B2(n4392), .A(n4310), .ZN(n4311) );
  OAI21_X1 U4888 ( .B1(n4395), .B2(n4391), .A(n4311), .ZN(U3549) );
  NAND2_X1 U4889 ( .A1(n4396), .A2(n4312), .ZN(n4314) );
  NAND2_X1 U4890 ( .A1(n4589), .A2(n4397), .ZN(n4313) );
  OAI211_X1 U4891 ( .C1(n4589), .C2(n4315), .A(n4314), .B(n4313), .ZN(U3548)
         );
  NAND4_X1 U4892 ( .A1(n4316), .A2(n4570), .A3(n4318), .A4(n4319), .ZN(n4324)
         );
  INV_X1 U4893 ( .A(n4317), .ZN(n4321) );
  NOR3_X1 U4894 ( .A1(n4319), .A2(n4318), .A3(n4577), .ZN(n4320) );
  NAND4_X1 U4895 ( .A1(n4325), .A2(n4324), .A3(n4323), .A4(n4322), .ZN(n4401)
         );
  MUX2_X1 U4896 ( .A(REG1_REG_29__SCAN_IN), .B(n4401), .S(n4589), .Z(U3547) );
  NAND2_X1 U4897 ( .A1(n4326), .A2(n4570), .ZN(n4328) );
  OAI211_X1 U4898 ( .C1(n2997), .C2(n4329), .A(n4328), .B(n4327), .ZN(n4402)
         );
  MUX2_X1 U4899 ( .A(REG1_REG_27__SCAN_IN), .B(n4402), .S(n4589), .Z(U3545) );
  INV_X1 U4900 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4332) );
  AOI21_X1 U4901 ( .B1(n4331), .B2(n4570), .A(n4330), .ZN(n4403) );
  MUX2_X1 U4902 ( .A(n4332), .B(n4403), .S(n4589), .Z(n4333) );
  OAI21_X1 U4903 ( .B1(n4391), .B2(n4406), .A(n4333), .ZN(U3544) );
  INV_X1 U4904 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4336) );
  AOI21_X1 U4905 ( .B1(n4335), .B2(n4570), .A(n4334), .ZN(n4407) );
  MUX2_X1 U4906 ( .A(n4336), .B(n4407), .S(n4589), .Z(n4337) );
  OAI21_X1 U4907 ( .B1(n4391), .B2(n4410), .A(n4337), .ZN(U3543) );
  INV_X1 U4908 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U4909 ( .B1(n4339), .B2(n4570), .A(n4338), .ZN(n4411) );
  MUX2_X1 U4910 ( .A(n4340), .B(n4411), .S(n4589), .Z(n4341) );
  OAI21_X1 U4911 ( .B1(n4391), .B2(n4414), .A(n4341), .ZN(U3542) );
  AOI21_X1 U4912 ( .B1(n4343), .B2(n4570), .A(n4342), .ZN(n4415) );
  MUX2_X1 U4913 ( .A(n4715), .B(n4415), .S(n4589), .Z(n4344) );
  OAI21_X1 U4914 ( .B1(n4391), .B2(n4418), .A(n4344), .ZN(U3541) );
  NAND3_X1 U4915 ( .A1(n4345), .A2(n2998), .A3(n4129), .ZN(n4346) );
  OAI211_X1 U4916 ( .C1(n4348), .C2(n4577), .A(n4347), .B(n4346), .ZN(n4419)
         );
  MUX2_X1 U4917 ( .A(REG1_REG_22__SCAN_IN), .B(n4419), .S(n4589), .Z(U3540) );
  INV_X1 U4918 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4351) );
  AOI21_X1 U4919 ( .B1(n4350), .B2(n4570), .A(n4349), .ZN(n4420) );
  MUX2_X1 U4920 ( .A(n4351), .B(n4420), .S(n4589), .Z(n4352) );
  OAI21_X1 U4921 ( .B1(n4391), .B2(n4423), .A(n4352), .ZN(U3539) );
  INV_X1 U4922 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4356) );
  INV_X1 U4923 ( .A(n4551), .ZN(n4560) );
  INV_X1 U4924 ( .A(n4353), .ZN(n4355) );
  AOI21_X1 U4925 ( .B1(n4560), .B2(n4355), .A(n4354), .ZN(n4424) );
  MUX2_X1 U4926 ( .A(n4356), .B(n4424), .S(n4589), .Z(n4357) );
  OAI21_X1 U4927 ( .B1(n4391), .B2(n4427), .A(n4357), .ZN(U3538) );
  INV_X1 U4928 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4360) );
  AOI21_X1 U4929 ( .B1(n4359), .B2(n4570), .A(n4358), .ZN(n4428) );
  MUX2_X1 U4930 ( .A(n4360), .B(n4428), .S(n4589), .Z(n4361) );
  OAI21_X1 U4931 ( .B1(n4391), .B2(n4430), .A(n4361), .ZN(U3537) );
  OAI211_X1 U4932 ( .C1(n4364), .C2(n4577), .A(n4363), .B(n4362), .ZN(n4431)
         );
  MUX2_X1 U4933 ( .A(REG1_REG_18__SCAN_IN), .B(n4431), .S(n4589), .Z(U3536) );
  AOI21_X1 U4934 ( .B1(n4366), .B2(n4570), .A(n4365), .ZN(n4432) );
  MUX2_X1 U4935 ( .A(n4367), .B(n4432), .S(n4589), .Z(n4368) );
  OAI21_X1 U4936 ( .B1(n4391), .B2(n4435), .A(n4368), .ZN(U3535) );
  AOI21_X1 U4937 ( .B1(n2998), .B2(n4370), .A(n4369), .ZN(n4371) );
  OAI21_X1 U4938 ( .B1(n4372), .B2(n4577), .A(n4371), .ZN(n4436) );
  MUX2_X1 U4939 ( .A(REG1_REG_16__SCAN_IN), .B(n4436), .S(n4589), .Z(U3534) );
  AOI21_X1 U4940 ( .B1(n2998), .B2(n4374), .A(n4373), .ZN(n4375) );
  OAI21_X1 U4941 ( .B1(n4376), .B2(n4577), .A(n4375), .ZN(n4437) );
  MUX2_X1 U4942 ( .A(REG1_REG_15__SCAN_IN), .B(n4437), .S(n4589), .Z(U3533) );
  AOI21_X1 U4943 ( .B1(n4378), .B2(n4570), .A(n4377), .ZN(n4438) );
  MUX2_X1 U4944 ( .A(n2222), .B(n4438), .S(n4589), .Z(n4379) );
  OAI21_X1 U4945 ( .B1(n4391), .B2(n4441), .A(n4379), .ZN(U3532) );
  INV_X1 U4946 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4382) );
  AOI21_X1 U4947 ( .B1(n4560), .B2(n4381), .A(n4380), .ZN(n4442) );
  MUX2_X1 U4948 ( .A(n4382), .B(n4442), .S(n4589), .Z(n4383) );
  OAI21_X1 U4949 ( .B1(n4391), .B2(n4444), .A(n4383), .ZN(U3531) );
  AOI21_X1 U4950 ( .B1(n4385), .B2(n4570), .A(n4384), .ZN(n4445) );
  MUX2_X1 U4951 ( .A(n4626), .B(n4445), .S(n4589), .Z(n4386) );
  OAI21_X1 U4952 ( .B1(n4391), .B2(n4448), .A(n4386), .ZN(U3530) );
  AOI21_X1 U4953 ( .B1(n4560), .B2(n4388), .A(n4387), .ZN(n4449) );
  MUX2_X1 U4954 ( .A(n4389), .B(n4449), .S(n4589), .Z(n4390) );
  OAI21_X1 U4955 ( .B1(n4391), .B2(n4452), .A(n4390), .ZN(U3529) );
  NAND2_X1 U4956 ( .A1(n4739), .A2(n4392), .ZN(n4394) );
  NAND2_X1 U4957 ( .A1(n4737), .A2(REG0_REG_31__SCAN_IN), .ZN(n4393) );
  OAI211_X1 U4958 ( .C1(n4395), .C2(n4451), .A(n4394), .B(n4393), .ZN(U3517)
         );
  INV_X1 U4959 ( .A(n4396), .ZN(n4400) );
  NAND2_X1 U4960 ( .A1(n4739), .A2(n4397), .ZN(n4399) );
  NAND2_X1 U4961 ( .A1(n4737), .A2(REG0_REG_30__SCAN_IN), .ZN(n4398) );
  OAI211_X1 U4962 ( .C1(n4400), .C2(n4451), .A(n4399), .B(n4398), .ZN(U3516)
         );
  MUX2_X1 U4963 ( .A(REG0_REG_29__SCAN_IN), .B(n4401), .S(n4739), .Z(U3515) );
  MUX2_X1 U4964 ( .A(REG0_REG_27__SCAN_IN), .B(n4402), .S(n4739), .Z(U3513) );
  INV_X1 U4965 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U4966 ( .A(n4404), .B(n4403), .S(n4739), .Z(n4405) );
  OAI21_X1 U4967 ( .B1(n4406), .B2(n4451), .A(n4405), .ZN(U3512) );
  INV_X1 U4968 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4408) );
  MUX2_X1 U4969 ( .A(n4408), .B(n4407), .S(n4739), .Z(n4409) );
  OAI21_X1 U4970 ( .B1(n4410), .B2(n4451), .A(n4409), .ZN(U3511) );
  INV_X1 U4971 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4412) );
  MUX2_X1 U4972 ( .A(n4412), .B(n4411), .S(n4739), .Z(n4413) );
  OAI21_X1 U4973 ( .B1(n4414), .B2(n4451), .A(n4413), .ZN(U3510) );
  INV_X1 U4974 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4416) );
  MUX2_X1 U4975 ( .A(n4416), .B(n4415), .S(n4739), .Z(n4417) );
  OAI21_X1 U4976 ( .B1(n4418), .B2(n4451), .A(n4417), .ZN(U3509) );
  MUX2_X1 U4977 ( .A(REG0_REG_22__SCAN_IN), .B(n4419), .S(n4739), .Z(U3508) );
  INV_X1 U4978 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4421) );
  MUX2_X1 U4979 ( .A(n4421), .B(n4420), .S(n4739), .Z(n4422) );
  OAI21_X1 U4980 ( .B1(n4423), .B2(n4451), .A(n4422), .ZN(U3507) );
  INV_X1 U4981 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4425) );
  MUX2_X1 U4982 ( .A(n4425), .B(n4424), .S(n4739), .Z(n4426) );
  OAI21_X1 U4983 ( .B1(n4427), .B2(n4451), .A(n4426), .ZN(U3506) );
  MUX2_X1 U4984 ( .A(n4640), .B(n4428), .S(n4739), .Z(n4429) );
  OAI21_X1 U4985 ( .B1(n4430), .B2(n4451), .A(n4429), .ZN(U3505) );
  MUX2_X1 U4986 ( .A(REG0_REG_18__SCAN_IN), .B(n4431), .S(n4739), .Z(U3503) );
  INV_X1 U4987 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4433) );
  MUX2_X1 U4988 ( .A(n4433), .B(n4432), .S(n4739), .Z(n4434) );
  OAI21_X1 U4989 ( .B1(n4435), .B2(n4451), .A(n4434), .ZN(U3501) );
  MUX2_X1 U4990 ( .A(REG0_REG_16__SCAN_IN), .B(n4436), .S(n4739), .Z(U3499) );
  MUX2_X1 U4991 ( .A(REG0_REG_15__SCAN_IN), .B(n4437), .S(n4739), .Z(U3497) );
  INV_X1 U4992 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4439) );
  MUX2_X1 U4993 ( .A(n4439), .B(n4438), .S(n4739), .Z(n4440) );
  OAI21_X1 U4994 ( .B1(n4441), .B2(n4451), .A(n4440), .ZN(U3495) );
  INV_X1 U4995 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4671) );
  MUX2_X1 U4996 ( .A(n4671), .B(n4442), .S(n4739), .Z(n4443) );
  OAI21_X1 U4997 ( .B1(n4444), .B2(n4451), .A(n4443), .ZN(U3493) );
  INV_X1 U4998 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4446) );
  MUX2_X1 U4999 ( .A(n4446), .B(n4445), .S(n4739), .Z(n4447) );
  OAI21_X1 U5000 ( .B1(n4448), .B2(n4451), .A(n4447), .ZN(U3491) );
  MUX2_X1 U5001 ( .A(n4625), .B(n4449), .S(n4739), .Z(n4450) );
  OAI21_X1 U5002 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(U3489) );
  MUX2_X1 U5003 ( .A(DATAI_29_), .B(n4453), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5004 ( .A(n4454), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5005 ( .A(n4455), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5006 ( .A(DATAI_24_), .B(n4456), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5007 ( .A(n4457), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5008 ( .A(n3909), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5009 ( .A(n4459), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5010 ( .A(n4460), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5011 ( .A(DATAI_8_), .B(n4461), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5012 ( .A(DATAI_7_), .B(n4462), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5013 ( .A(n4463), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5014 ( .A(DATAI_3_), .B(n4464), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5015 ( .A(n4465), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5016 ( .A(n4469), .ZN(n4466) );
  OAI211_X1 U5017 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4467), .A(n4466), .B(n4468), 
        .ZN(n4473) );
  OAI22_X1 U5018 ( .A1(n4469), .A2(n4468), .B1(n4497), .B2(REG1_REG_0__SCAN_IN), .ZN(n4470) );
  INV_X1 U5019 ( .A(n4470), .ZN(n4472) );
  AOI22_X1 U5020 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4500), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4471) );
  OAI221_X1 U5021 ( .B1(IR_REG_0__SCAN_IN), .B2(n4473), .C1(n2375), .C2(n4472), 
        .A(n4471), .ZN(U3240) );
  AOI21_X1 U5022 ( .B1(n4500), .B2(ADDR_REG_16__SCAN_IN), .A(n4474), .ZN(n4484) );
  OAI21_X1 U5023 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4482) );
  OAI21_X1 U5024 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4481) );
  AOI22_X1 U5025 ( .A1(n4494), .A2(n4482), .B1(n4510), .B2(n4481), .ZN(n4483)
         );
  OAI211_X1 U5026 ( .C1(n4543), .C2(n4514), .A(n4484), .B(n4483), .ZN(U3256)
         );
  AOI21_X1 U5027 ( .B1(n4500), .B2(ADDR_REG_17__SCAN_IN), .A(n4485), .ZN(n4496) );
  OAI21_X1 U5028 ( .B1(n4488), .B2(n4487), .A(n4486), .ZN(n4493) );
  OAI21_X1 U5029 ( .B1(n4491), .B2(n4490), .A(n4489), .ZN(n4492) );
  AOI22_X1 U5030 ( .A1(n4494), .A2(n4493), .B1(n4510), .B2(n4492), .ZN(n4495)
         );
  OAI211_X1 U5031 ( .C1(n4542), .C2(n4514), .A(n4496), .B(n4495), .ZN(U3257)
         );
  NAND2_X1 U5032 ( .A1(n4500), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5033 ( .A1(n4503), .A2(n4502), .ZN(n4504) );
  AOI21_X1 U5034 ( .B1(n4508), .B2(n4507), .A(n4506), .ZN(n4509) );
  NAND2_X1 U5035 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  OAI211_X1 U5036 ( .C1(n4514), .C2(n4513), .A(n4512), .B(n4511), .ZN(U3258)
         );
  AOI22_X1 U5037 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4530), .B1(
        REG2_REG_2__SCAN_IN), .B2(n2003), .ZN(n4519) );
  AOI22_X1 U5038 ( .A1(n4532), .A2(n4517), .B1(n4516), .B2(n4515), .ZN(n4518)
         );
  OAI211_X1 U5039 ( .C1(n2003), .C2(n4520), .A(n4519), .B(n4518), .ZN(U3288)
         );
  OAI22_X1 U5040 ( .A1(n4578), .A2(n4523), .B1(n4522), .B2(n4521), .ZN(n4580)
         );
  AOI21_X1 U5041 ( .B1(n4524), .B2(n4526), .A(n4525), .ZN(n4527) );
  OAI22_X1 U5042 ( .A1(n4578), .A2(n4528), .B1(n4527), .B2(n4576), .ZN(n4529)
         );
  NOR2_X1 U5043 ( .A1(n4580), .A2(n4529), .ZN(n4536) );
  INV_X1 U5044 ( .A(n4578), .ZN(n4531) );
  AOI22_X1 U5045 ( .A1(n4532), .A2(n4531), .B1(REG3_REG_0__SCAN_IN), .B2(n4530), .ZN(n4533) );
  OAI221_X1 U5046 ( .B1(n2003), .B2(n4536), .C1(n4535), .C2(n4534), .A(n4533), 
        .ZN(U3290) );
  INV_X1 U5047 ( .A(D_REG_31__SCAN_IN), .ZN(n4721) );
  NOR2_X1 U5048 ( .A1(n4538), .A2(n4721), .ZN(U3291) );
  AND2_X1 U5049 ( .A1(D_REG_30__SCAN_IN), .A2(n4537), .ZN(U3292) );
  AND2_X1 U5050 ( .A1(D_REG_29__SCAN_IN), .A2(n4537), .ZN(U3293) );
  AND2_X1 U5051 ( .A1(D_REG_28__SCAN_IN), .A2(n4537), .ZN(U3294) );
  NOR2_X1 U5052 ( .A1(n4538), .A2(n4653), .ZN(U3295) );
  AND2_X1 U5053 ( .A1(D_REG_26__SCAN_IN), .A2(n4537), .ZN(U3296) );
  NOR2_X1 U5054 ( .A1(n4538), .A2(n4656), .ZN(U3297) );
  INV_X1 U5055 ( .A(D_REG_24__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U5056 ( .A1(n4538), .A2(n4698), .ZN(U3298) );
  AND2_X1 U5057 ( .A1(D_REG_23__SCAN_IN), .A2(n4537), .ZN(U3299) );
  AND2_X1 U5058 ( .A1(D_REG_22__SCAN_IN), .A2(n4537), .ZN(U3300) );
  INV_X1 U5059 ( .A(D_REG_21__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U5060 ( .A1(n4538), .A2(n4704), .ZN(U3301) );
  AND2_X1 U5061 ( .A1(D_REG_20__SCAN_IN), .A2(n4537), .ZN(U3302) );
  AND2_X1 U5062 ( .A1(D_REG_19__SCAN_IN), .A2(n4537), .ZN(U3303) );
  INV_X1 U5063 ( .A(D_REG_18__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5064 ( .A1(n4538), .A2(n4650), .ZN(U3304) );
  AND2_X1 U5065 ( .A1(D_REG_17__SCAN_IN), .A2(n4537), .ZN(U3305) );
  AND2_X1 U5066 ( .A1(D_REG_16__SCAN_IN), .A2(n4537), .ZN(U3306) );
  AND2_X1 U5067 ( .A1(D_REG_15__SCAN_IN), .A2(n4537), .ZN(U3307) );
  AND2_X1 U5068 ( .A1(D_REG_14__SCAN_IN), .A2(n4537), .ZN(U3308) );
  AND2_X1 U5069 ( .A1(D_REG_13__SCAN_IN), .A2(n4537), .ZN(U3309) );
  NOR2_X1 U5070 ( .A1(n4538), .A2(n4635), .ZN(U3310) );
  INV_X1 U5071 ( .A(D_REG_11__SCAN_IN), .ZN(n4702) );
  NOR2_X1 U5072 ( .A1(n4538), .A2(n4702), .ZN(U3311) );
  INV_X1 U5073 ( .A(D_REG_10__SCAN_IN), .ZN(n4652) );
  NOR2_X1 U5074 ( .A1(n4538), .A2(n4652), .ZN(U3312) );
  AND2_X1 U5075 ( .A1(D_REG_9__SCAN_IN), .A2(n4537), .ZN(U3313) );
  AND2_X1 U5076 ( .A1(D_REG_8__SCAN_IN), .A2(n4537), .ZN(U3314) );
  AND2_X1 U5077 ( .A1(D_REG_7__SCAN_IN), .A2(n4537), .ZN(U3315) );
  AND2_X1 U5078 ( .A1(D_REG_6__SCAN_IN), .A2(n4537), .ZN(U3316) );
  AND2_X1 U5079 ( .A1(D_REG_5__SCAN_IN), .A2(n4537), .ZN(U3317) );
  AND2_X1 U5080 ( .A1(D_REG_4__SCAN_IN), .A2(n4537), .ZN(U3318) );
  INV_X1 U5081 ( .A(D_REG_3__SCAN_IN), .ZN(n4707) );
  NOR2_X1 U5082 ( .A1(n4538), .A2(n4707), .ZN(U3319) );
  NOR2_X1 U5083 ( .A1(n4538), .A2(n4638), .ZN(U3320) );
  INV_X1 U5084 ( .A(DATAI_23_), .ZN(n4614) );
  AOI21_X1 U5085 ( .B1(U3149), .B2(n4614), .A(n4539), .ZN(U3329) );
  OAI22_X1 U5086 ( .A1(U3149), .A2(n4540), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4541) );
  INV_X1 U5087 ( .A(n4541), .ZN(U3334) );
  AOI22_X1 U5088 ( .A1(STATE_REG_SCAN_IN), .A2(n4542), .B1(n2658), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5089 ( .A(DATAI_16_), .ZN(n4708) );
  AOI22_X1 U5090 ( .A1(STATE_REG_SCAN_IN), .A2(n4543), .B1(n4708), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5091 ( .A(DATAI_0_), .ZN(n4544) );
  AOI22_X1 U5092 ( .A1(STATE_REG_SCAN_IN), .A2(n2375), .B1(n4544), .B2(U3149), 
        .ZN(U3352) );
  NOR2_X1 U5093 ( .A1(n4545), .A2(n4551), .ZN(n4547) );
  AOI211_X1 U5094 ( .C1(n2998), .C2(n4548), .A(n4547), .B(n4546), .ZN(n4582)
         );
  INV_X1 U5095 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5096 ( .A1(n4739), .A2(n4582), .B1(n4549), .B2(n4737), .ZN(U3469)
         );
  OAI22_X1 U5097 ( .A1(n4552), .A2(n4551), .B1(n2997), .B2(n4550), .ZN(n4553)
         );
  NOR2_X1 U5098 ( .A1(n4554), .A2(n4553), .ZN(n4584) );
  INV_X1 U5099 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5100 ( .A1(n4739), .A2(n4584), .B1(n4555), .B2(n4737), .ZN(U3473)
         );
  INV_X1 U5101 ( .A(n4556), .ZN(n4561) );
  INV_X1 U5102 ( .A(n4557), .ZN(n4559) );
  AOI211_X1 U5103 ( .C1(n4561), .C2(n4560), .A(n4559), .B(n4558), .ZN(n4585)
         );
  INV_X1 U5104 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5105 ( .A1(n4739), .A2(n4585), .B1(n4562), .B2(n4737), .ZN(U3475)
         );
  NOR2_X1 U5106 ( .A1(n4563), .A2(n4577), .ZN(n4566) );
  INV_X1 U5107 ( .A(n4564), .ZN(n4565) );
  AOI211_X1 U5108 ( .C1(n2998), .C2(n4567), .A(n4566), .B(n4565), .ZN(n4586)
         );
  INV_X1 U5109 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5110 ( .A1(n4739), .A2(n4586), .B1(n4568), .B2(n4737), .ZN(U3477)
         );
  NAND3_X1 U5111 ( .A1(n4571), .A2(n4570), .A3(n4569), .ZN(n4572) );
  AND3_X1 U5112 ( .A1(n4574), .A2(n4573), .A3(n4572), .ZN(n4588) );
  INV_X1 U5113 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5114 ( .A1(n4739), .A2(n4588), .B1(n4575), .B2(n4737), .ZN(U3481)
         );
  OAI22_X1 U5115 ( .A1(n4578), .A2(n4577), .B1(n2837), .B2(n4576), .ZN(n4579)
         );
  OR2_X1 U5116 ( .A1(n4580), .A2(n4579), .ZN(n4738) );
  OAI22_X1 U5117 ( .A1(n4587), .A2(n4738), .B1(REG1_REG_0__SCAN_IN), .B2(n4589), .ZN(n4581) );
  INV_X1 U5118 ( .A(n4581), .ZN(U3518) );
  AOI22_X1 U5119 ( .A1(n4589), .A2(n4582), .B1(n3069), .B2(n4587), .ZN(U3519)
         );
  INV_X1 U5120 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5121 ( .A1(n4589), .A2(n4584), .B1(n4583), .B2(n4587), .ZN(U3521)
         );
  AOI22_X1 U5122 ( .A1(n4589), .A2(n4585), .B1(n2210), .B2(n4587), .ZN(U3522)
         );
  AOI22_X1 U5123 ( .A1(n4589), .A2(n4586), .B1(n2444), .B2(n4587), .ZN(U3523)
         );
  AOI22_X1 U5124 ( .A1(n4589), .A2(n4588), .B1(n4669), .B2(n4587), .ZN(U3525)
         );
  NAND4_X1 U5125 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4684), .A3(n4689), .A4(n4685), .ZN(n4593) );
  NAND4_X1 U5126 ( .A1(REG2_REG_26__SCAN_IN), .A2(REG2_REG_29__SCAN_IN), .A3(
        REG3_REG_0__SCAN_IN), .A4(n4688), .ZN(n4592) );
  AND4_X1 U5127 ( .A1(REG0_REG_13__SCAN_IN), .A2(REG0_REG_10__SCAN_IN), .A3(
        REG0_REG_9__SCAN_IN), .A4(n4672), .ZN(n4590) );
  NAND4_X1 U5128 ( .A1(n4590), .A2(n4669), .A3(n4676), .A4(n4668), .ZN(n4591)
         );
  NOR4_X1 U5129 ( .A1(IR_REG_15__SCAN_IN), .A2(n4593), .A3(n4592), .A4(n4591), 
        .ZN(n4736) );
  NAND4_X1 U5130 ( .A1(IR_REG_7__SCAN_IN), .A2(DATAI_11_), .A3(DATAI_10_), 
        .A4(n4623), .ZN(n4608) );
  NOR4_X1 U5131 ( .A1(REG3_REG_16__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .A3(
        DATAO_REG_25__SCAN_IN), .A4(n4650), .ZN(n4596) );
  NOR4_X1 U5132 ( .A1(D_REG_1__SCAN_IN), .A2(DATAI_13_), .A3(
        REG0_REG_18__SCAN_IN), .A4(n4640), .ZN(n4594) );
  AND3_X1 U5133 ( .A1(IR_REG_26__SCAN_IN), .A2(n4594), .A3(DATAI_30_), .ZN(
        n4595) );
  NAND4_X1 U5134 ( .A1(n4596), .A2(n4595), .A3(D_REG_10__SCAN_IN), .A4(n4655), 
        .ZN(n4607) );
  NOR4_X1 U5135 ( .A1(REG2_REG_12__SCAN_IN), .A2(DATAI_23_), .A3(
        ADDR_REG_8__SCAN_IN), .A4(n2375), .ZN(n4604) );
  INV_X1 U5136 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4610) );
  NAND4_X1 U5137 ( .A1(REG3_REG_24__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        n4610), .A4(n2185), .ZN(n4598) );
  NAND4_X1 U5138 ( .A1(REG2_REG_14__SCAN_IN), .A2(REG0_REG_11__SCAN_IN), .A3(
        REG1_REG_2__SCAN_IN), .A4(n4626), .ZN(n4597) );
  NOR4_X1 U5139 ( .A1(DATAO_REG_27__SCAN_IN), .A2(n4704), .A3(n4598), .A4(
        n4597), .ZN(n4603) );
  NAND4_X1 U5140 ( .A1(REG1_REG_27__SCAN_IN), .A2(REG1_REG_23__SCAN_IN), .A3(
        n4718), .A4(n4717), .ZN(n4601) );
  NAND3_X1 U5141 ( .A1(REG0_REG_29__SCAN_IN), .A2(DATAO_REG_3__SCAN_IN), .A3(
        DATAO_REG_20__SCAN_IN), .ZN(n4600) );
  NAND4_X1 U5142 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        DATAO_REG_7__SCAN_IN), .A4(n4708), .ZN(n4599) );
  NOR4_X1 U5143 ( .A1(DATAO_REG_10__SCAN_IN), .A2(n4601), .A3(n4600), .A4(
        n4599), .ZN(n4602) );
  NAND4_X1 U5144 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4606)
         );
  NOR3_X1 U5145 ( .A1(n4608), .A2(n4607), .A3(n4606), .ZN(n4735) );
  AOI22_X1 U5146 ( .A1(n4610), .A2(keyinput17), .B1(keyinput10), .B2(n4188), 
        .ZN(n4609) );
  OAI221_X1 U5147 ( .B1(n4610), .B2(keyinput17), .C1(n4188), .C2(keyinput10), 
        .A(n4609), .ZN(n4620) );
  AOI22_X1 U5148 ( .A1(n4612), .A2(keyinput11), .B1(keyinput4), .B2(n2185), 
        .ZN(n4611) );
  OAI221_X1 U5149 ( .B1(n4612), .B2(keyinput11), .C1(n2185), .C2(keyinput4), 
        .A(n4611), .ZN(n4619) );
  AOI22_X1 U5150 ( .A1(n4614), .A2(keyinput2), .B1(n2375), .B2(keyinput9), 
        .ZN(n4613) );
  OAI221_X1 U5151 ( .B1(n4614), .B2(keyinput2), .C1(n2375), .C2(keyinput9), 
        .A(n4613), .ZN(n4618) );
  INV_X1 U5152 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5153 ( .A1(n4616), .A2(keyinput35), .B1(n3924), .B2(keyinput14), 
        .ZN(n4615) );
  OAI221_X1 U5154 ( .B1(n4616), .B2(keyinput35), .C1(n3924), .C2(keyinput14), 
        .A(n4615), .ZN(n4617) );
  NOR4_X1 U5155 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4666)
         );
  AOI22_X1 U5156 ( .A1(n2389), .A2(keyinput6), .B1(n2595), .B2(keyinput27), 
        .ZN(n4621) );
  OAI221_X1 U5157 ( .B1(n2389), .B2(keyinput6), .C1(n2595), .C2(keyinput27), 
        .A(n4621), .ZN(n4632) );
  AOI22_X1 U5158 ( .A1(n2555), .A2(keyinput19), .B1(n4623), .B2(keyinput59), 
        .ZN(n4622) );
  OAI221_X1 U5159 ( .B1(n2555), .B2(keyinput19), .C1(n4623), .C2(keyinput59), 
        .A(n4622), .ZN(n4631) );
  AOI22_X1 U5160 ( .A1(n4626), .A2(keyinput8), .B1(keyinput55), .B2(n4625), 
        .ZN(n4624) );
  OAI221_X1 U5161 ( .B1(n4626), .B2(keyinput8), .C1(n4625), .C2(keyinput55), 
        .A(n4624), .ZN(n4630) );
  XNOR2_X1 U5162 ( .A(IR_REG_7__SCAN_IN), .B(keyinput39), .ZN(n4628) );
  XNOR2_X1 U5163 ( .A(DATAI_10_), .B(keyinput15), .ZN(n4627) );
  NAND2_X1 U5164 ( .A1(n4628), .A2(n4627), .ZN(n4629) );
  NOR4_X1 U5165 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(n4665)
         );
  AOI22_X1 U5166 ( .A1(n4635), .A2(keyinput5), .B1(keyinput1), .B2(n4634), 
        .ZN(n4633) );
  OAI221_X1 U5167 ( .B1(n4635), .B2(keyinput5), .C1(n4634), .C2(keyinput1), 
        .A(n4633), .ZN(n4647) );
  AOI22_X1 U5168 ( .A1(n4638), .A2(keyinput18), .B1(n4637), .B2(keyinput21), 
        .ZN(n4636) );
  OAI221_X1 U5169 ( .B1(n4638), .B2(keyinput18), .C1(n4637), .C2(keyinput21), 
        .A(n4636), .ZN(n4646) );
  AOI22_X1 U5170 ( .A1(n4641), .A2(keyinput23), .B1(n4640), .B2(keyinput13), 
        .ZN(n4639) );
  OAI221_X1 U5171 ( .B1(n4641), .B2(keyinput23), .C1(n4640), .C2(keyinput13), 
        .A(n4639), .ZN(n4645) );
  XOR2_X1 U5172 ( .A(n2587), .B(keyinput16), .Z(n4643) );
  XNOR2_X1 U5173 ( .A(IR_REG_26__SCAN_IN), .B(keyinput12), .ZN(n4642) );
  NAND2_X1 U5174 ( .A1(n4643), .A2(n4642), .ZN(n4644) );
  NOR4_X1 U5175 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4664)
         );
  AOI22_X1 U5176 ( .A1(n4650), .A2(keyinput47), .B1(keyinput31), .B2(n4649), 
        .ZN(n4648) );
  OAI221_X1 U5177 ( .B1(n4650), .B2(keyinput47), .C1(n4649), .C2(keyinput31), 
        .A(n4648), .ZN(n4662) );
  AOI22_X1 U5178 ( .A1(n4653), .A2(keyinput0), .B1(keyinput7), .B2(n4652), 
        .ZN(n4651) );
  OAI221_X1 U5179 ( .B1(n4653), .B2(keyinput0), .C1(n4652), .C2(keyinput7), 
        .A(n4651), .ZN(n4661) );
  AOI22_X1 U5180 ( .A1(n4656), .A2(keyinput43), .B1(keyinput63), .B2(n4655), 
        .ZN(n4654) );
  OAI221_X1 U5181 ( .B1(n4656), .B2(keyinput43), .C1(n4655), .C2(keyinput63), 
        .A(n4654), .ZN(n4660) );
  XNOR2_X1 U5182 ( .A(IR_REG_27__SCAN_IN), .B(keyinput51), .ZN(n4658) );
  XNOR2_X1 U5183 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput3), .ZN(n4657) );
  NAND2_X1 U5184 ( .A1(n4658), .A2(n4657), .ZN(n4659) );
  NOR4_X1 U5185 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4663)
         );
  NAND4_X1 U5186 ( .A1(n4666), .A2(n4665), .A3(n4664), .A4(n4663), .ZN(n4734)
         );
  AOI22_X1 U5187 ( .A1(n4669), .A2(keyinput30), .B1(keyinput26), .B2(n4668), 
        .ZN(n4667) );
  OAI221_X1 U5188 ( .B1(n4669), .B2(keyinput30), .C1(n4668), .C2(keyinput26), 
        .A(n4667), .ZN(n4682) );
  AOI22_X1 U5189 ( .A1(n4672), .A2(keyinput29), .B1(n4671), .B2(keyinput61), 
        .ZN(n4670) );
  OAI221_X1 U5190 ( .B1(n4672), .B2(keyinput29), .C1(n4671), .C2(keyinput61), 
        .A(n4670), .ZN(n4681) );
  AOI22_X1 U5191 ( .A1(n4675), .A2(keyinput25), .B1(n4674), .B2(keyinput52), 
        .ZN(n4673) );
  OAI221_X1 U5192 ( .B1(n4675), .B2(keyinput25), .C1(n4674), .C2(keyinput52), 
        .A(n4673), .ZN(n4680) );
  XOR2_X1 U5193 ( .A(n4676), .B(keyinput28), .Z(n4678) );
  XNOR2_X1 U5194 ( .A(IR_REG_15__SCAN_IN), .B(keyinput40), .ZN(n4677) );
  NAND2_X1 U5195 ( .A1(n4678), .A2(n4677), .ZN(n4679) );
  NOR4_X1 U5196 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4732)
         );
  AOI22_X1 U5197 ( .A1(n4685), .A2(keyinput60), .B1(n4684), .B2(keyinput38), 
        .ZN(n4683) );
  OAI221_X1 U5198 ( .B1(n4685), .B2(keyinput60), .C1(n4684), .C2(keyinput38), 
        .A(n4683), .ZN(n4696) );
  AOI22_X1 U5199 ( .A1(n4688), .A2(keyinput32), .B1(n4687), .B2(keyinput36), 
        .ZN(n4686) );
  OAI221_X1 U5200 ( .B1(n4688), .B2(keyinput32), .C1(n4687), .C2(keyinput36), 
        .A(n4686), .ZN(n4695) );
  XOR2_X1 U5201 ( .A(n4031), .B(keyinput41), .Z(n4693) );
  XOR2_X1 U5202 ( .A(n4689), .B(keyinput34), .Z(n4692) );
  XNOR2_X1 U5203 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput45), .ZN(n4691) );
  XNOR2_X1 U5204 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput42), .ZN(n4690) );
  NAND4_X1 U5205 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4694)
         );
  NOR3_X1 U5206 ( .A1(n4696), .A2(n4695), .A3(n4694), .ZN(n4731) );
  AOI22_X1 U5207 ( .A1(n4699), .A2(keyinput58), .B1(n4698), .B2(keyinput56), 
        .ZN(n4697) );
  OAI221_X1 U5208 ( .B1(n4699), .B2(keyinput58), .C1(n4698), .C2(keyinput56), 
        .A(n4697), .ZN(n4712) );
  AOI22_X1 U5209 ( .A1(n4702), .A2(keyinput44), .B1(keyinput46), .B2(n4701), 
        .ZN(n4700) );
  OAI221_X1 U5210 ( .B1(n4702), .B2(keyinput44), .C1(n4701), .C2(keyinput46), 
        .A(n4700), .ZN(n4711) );
  AOI22_X1 U5211 ( .A1(n4705), .A2(keyinput24), .B1(n4704), .B2(keyinput37), 
        .ZN(n4703) );
  OAI221_X1 U5212 ( .B1(n4705), .B2(keyinput24), .C1(n4704), .C2(keyinput37), 
        .A(n4703), .ZN(n4710) );
  AOI22_X1 U5213 ( .A1(n4708), .A2(keyinput20), .B1(n4707), .B2(keyinput22), 
        .ZN(n4706) );
  OAI221_X1 U5214 ( .B1(n4708), .B2(keyinput20), .C1(n4707), .C2(keyinput22), 
        .A(n4706), .ZN(n4709) );
  NOR4_X1 U5215 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4730)
         );
  AOI22_X1 U5216 ( .A1(n4715), .A2(keyinput62), .B1(n4714), .B2(keyinput54), 
        .ZN(n4713) );
  OAI221_X1 U5217 ( .B1(n4715), .B2(keyinput62), .C1(n4714), .C2(keyinput54), 
        .A(n4713), .ZN(n4728) );
  AOI22_X1 U5218 ( .A1(n4718), .A2(keyinput33), .B1(keyinput49), .B2(n4717), 
        .ZN(n4716) );
  OAI221_X1 U5219 ( .B1(n4718), .B2(keyinput33), .C1(n4717), .C2(keyinput49), 
        .A(n4716), .ZN(n4727) );
  AOI22_X1 U5220 ( .A1(n4721), .A2(keyinput50), .B1(keyinput53), .B2(n4720), 
        .ZN(n4719) );
  OAI221_X1 U5221 ( .B1(n4721), .B2(keyinput50), .C1(n4720), .C2(keyinput53), 
        .A(n4719), .ZN(n4726) );
  AOI22_X1 U5222 ( .A1(n4724), .A2(keyinput57), .B1(keyinput48), .B2(n4723), 
        .ZN(n4722) );
  OAI221_X1 U5223 ( .B1(n4724), .B2(keyinput57), .C1(n4723), .C2(keyinput48), 
        .A(n4722), .ZN(n4725) );
  NOR4_X1 U5224 ( .A1(n4728), .A2(n4727), .A3(n4726), .A4(n4725), .ZN(n4729)
         );
  NAND4_X1 U5225 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4733)
         );
  AOI211_X1 U5226 ( .C1(n4736), .C2(n4735), .A(n4734), .B(n4733), .ZN(n4741)
         );
  AOI22_X1 U5227 ( .A1(n4739), .A2(n4738), .B1(REG0_REG_0__SCAN_IN), .B2(n4737), .ZN(n4740) );
  XNOR2_X1 U5228 ( .A(n4741), .B(n4740), .ZN(U3467) );
  CLKBUF_X1 U2247 ( .A(n2422), .Z(n2807) );
  CLKBUF_X1 U2320 ( .A(n2390), .Z(n3722) );
endmodule

