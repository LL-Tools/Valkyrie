

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11158, n11159,
         n11160, n11163, n11164, n11166, n11167, n11168, n11169, n11171,
         n11172, n11173, n11174, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22730,
         n22731;

  AND4_X1 U11250 ( .A1(n11238), .A2(n11279), .A3(n16265), .A4(n11273), .ZN(
        n11278) );
  CLKBUF_X2 U11251 ( .A(n19024), .Z(n11223) );
  INV_X1 U11253 ( .A(n11152), .ZN(n21573) );
  AND2_X1 U11255 ( .A1(n16881), .A2(n16237), .ZN(n16240) );
  NAND2_X1 U11256 ( .A1(n16496), .A2(n16498), .ZN(n13592) );
  AOI22_X1 U11257 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16423), .B1(n16409), 
        .B2(n19237), .ZN(n19024) );
  NAND2_X1 U11258 ( .A1(n16188), .A2(n17265), .ZN(n17815) );
  AND2_X1 U11259 ( .A1(n18500), .A2(n18499), .ZN(n18522) );
  INV_X1 U11260 ( .A(n21834), .ZN(n21695) );
  OR2_X1 U11261 ( .A1(n21577), .A2(n21575), .ZN(n11152) );
  NAND2_X1 U11262 ( .A1(n21764), .A2(n21756), .ZN(n21727) );
  NAND2_X1 U11263 ( .A1(n18348), .A2(n18466), .ZN(n18404) );
  NAND2_X1 U11264 ( .A1(n14866), .A2(n14931), .ZN(n14930) );
  CLKBUF_X2 U11265 ( .A(n11597), .Z(n16794) );
  CLKBUF_X1 U11266 ( .A(n12955), .Z(n19190) );
  NOR2_X1 U11267 ( .A1(n17550), .A2(n13406), .ZN(n17528) );
  NOR4_X1 U11268 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n18623), .ZN(n18333) );
  AOI21_X1 U11269 ( .B1(n15669), .B2(n13342), .A(n11274), .ZN(n17579) );
  OR2_X1 U11270 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  OR2_X1 U11271 ( .A1(n13738), .A2(n13737), .ZN(n13759) );
  INV_X1 U11272 ( .A(n16415), .ZN(n13980) );
  NAND2_X1 U11273 ( .A1(n18441), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14163) );
  INV_X1 U11274 ( .A(n18263), .ZN(n16062) );
  AND2_X1 U11275 ( .A1(n13302), .A2(n13301), .ZN(n11147) );
  NAND2_X1 U11276 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14327) );
  NOR2_X1 U11277 ( .A1(n17027), .A2(n14183), .ZN(n14186) );
  BUF_X1 U11278 ( .A(n15574), .Z(n11172) );
  NOR2_X1 U11279 ( .A1(n17059), .A2(n14373), .ZN(n14184) );
  NOR2_X2 U11280 ( .A1(n21237), .A2(n15618), .ZN(n18313) );
  CLKBUF_X2 U11281 ( .A(n15556), .Z(n20821) );
  BUF_X2 U11282 ( .A(n18199), .Z(n18265) );
  BUF_X1 U11283 ( .A(n18279), .Z(n18248) );
  BUF_X2 U11284 ( .A(n14043), .Z(n18262) );
  NAND2_X1 U11285 ( .A1(n11493), .A2(n11492), .ZN(n11609) );
  BUF_X2 U11286 ( .A(n14108), .Z(n18272) );
  BUF_X1 U11287 ( .A(n12604), .Z(n16360) );
  NAND2_X1 U11288 ( .A1(n18703), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18690) );
  OR2_X1 U11289 ( .A1(n13295), .A2(n18853), .ZN(n12541) );
  INV_X1 U11290 ( .A(n18697), .ZN(n18703) );
  BUF_X1 U11291 ( .A(n14066), .Z(n18032) );
  CLKBUF_X2 U11292 ( .A(n14087), .Z(n18270) );
  INV_X2 U11293 ( .A(n18063), .ZN(n18051) );
  INV_X1 U11294 ( .A(n13874), .ZN(n13470) );
  BUF_X4 U11295 ( .A(n15563), .Z(n11171) );
  BUF_X2 U11296 ( .A(n14087), .Z(n18157) );
  CLKBUF_X1 U11297 ( .A(n16824), .Z(n13529) );
  CLKBUF_X1 U11298 ( .A(n11443), .Z(n12332) );
  CLKBUF_X1 U11299 ( .A(n11516), .Z(n11442) );
  CLKBUF_X2 U11300 ( .A(n11395), .Z(n12333) );
  CLKBUF_X2 U11301 ( .A(n11360), .Z(n11984) );
  CLKBUF_X2 U11302 ( .A(n11394), .Z(n11179) );
  CLKBUF_X2 U11303 ( .A(n12569), .Z(n16391) );
  CLKBUF_X2 U11304 ( .A(n11955), .Z(n13536) );
  NAND2_X1 U11305 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21851), .ZN(
        n14030) );
  INV_X2 U11306 ( .A(n13232), .ZN(n20179) );
  CLKBUF_X2 U11307 ( .A(n12711), .Z(n13891) );
  NAND2_X2 U11308 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21392), .ZN(
        n14031) );
  AND2_X2 U11310 ( .A1(n19079), .A2(n12519), .ZN(n12712) );
  AND2_X2 U11311 ( .A1(n19079), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12736) );
  NAND2_X2 U11312 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20789) );
  NAND2_X1 U11313 ( .A1(n13953), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13882) );
  OAI21_X1 U11314 ( .B1(n12465), .B2(n12464), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12472) );
  INV_X2 U11316 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12519) );
  INV_X1 U11317 ( .A(n14907), .ZN(n11705) );
  OR2_X1 U11318 ( .A1(n11328), .A2(n11327), .ZN(n14621) );
  OR2_X1 U11319 ( .A1(n11339), .A2(n11338), .ZN(n11410) );
  AND2_X2 U11320 ( .A1(n11300), .A2(n11318), .ZN(n12076) );
  AND4_X1 U11321 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11300) );
  AND2_X1 U11322 ( .A1(n11312), .A2(n14473), .ZN(n11483) );
  AND2_X1 U11323 ( .A1(n14473), .A2(n14474), .ZN(n11360) );
  AND2_X1 U11324 ( .A1(n16829), .A2(n14304), .ZN(n11444) );
  BUF_X1 U11325 ( .A(n11333), .Z(n11169) );
  AND2_X2 U11326 ( .A1(n11309), .A2(n16829), .ZN(n11517) );
  AND2_X2 U11327 ( .A1(n11312), .A2(n14304), .ZN(n13528) );
  AND2_X1 U11328 ( .A1(n16828), .A2(n14473), .ZN(n11394) );
  AND2_X1 U11329 ( .A1(n11313), .A2(n14474), .ZN(n11395) );
  AND2_X1 U11330 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14474) );
  INV_X1 U11331 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11301) );
  CLKBUF_X1 U11332 ( .A(n22092), .Z(n11143) );
  NOR2_X1 U11333 ( .A1(n14916), .A2(n14910), .ZN(n22092) );
  CLKBUF_X1 U11334 ( .A(n19065), .Z(n11144) );
  NOR2_X1 U11335 ( .A1(n14502), .A2(n14267), .ZN(n19065) );
  CLKBUF_X1 U11336 ( .A(n18374), .Z(n11145) );
  NAND2_X1 U11337 ( .A1(n15063), .A2(n15670), .ZN(n11146) );
  AND2_X1 U11338 ( .A1(n13302), .A2(n13301), .ZN(n13502) );
  AOI21_X2 U11339 ( .B1(n16870), .B2(n19154), .A(n16366), .ZN(n16367) );
  NAND2_X1 U11340 ( .A1(n13092), .A2(n11151), .ZN(n11148) );
  AND2_X1 U11341 ( .A1(n11148), .A2(n11149), .ZN(n16169) );
  OR2_X1 U11342 ( .A1(n11150), .A2(n17345), .ZN(n11149) );
  INV_X1 U11343 ( .A(n16154), .ZN(n11150) );
  AND2_X1 U11344 ( .A1(n13091), .A2(n16154), .ZN(n11151) );
  AOI21_X2 U11345 ( .B1(n17230), .B2(n17353), .A(n17216), .ZN(n16206) );
  AND2_X2 U11346 ( .A1(n14854), .A2(n14925), .ZN(n15653) );
  NOR2_X2 U11347 ( .A1(n14213), .A2(n19044), .ZN(n14212) );
  NOR2_X2 U11348 ( .A1(n17297), .A2(n14205), .ZN(n14204) );
  NOR2_X2 U11349 ( .A1(n15765), .A2(n14185), .ZN(n14188) );
  AND2_X1 U11350 ( .A1(n14859), .A2(n14927), .ZN(n11153) );
  BUF_X1 U11351 ( .A(n12580), .Z(n11154) );
  AND2_X1 U11352 ( .A1(n14859), .A2(n14927), .ZN(n14920) );
  NOR2_X4 U11353 ( .A1(n18690), .A2(n20843), .ZN(n18677) );
  NOR2_X2 U11354 ( .A1(n14159), .A2(n21125), .ZN(n14157) );
  NOR2_X2 U11355 ( .A1(n21028), .A2(n11293), .ZN(n21027) );
  NAND2_X2 U11357 ( .A1(n11548), .A2(n14554), .ZN(n11641) );
  AOI21_X2 U11359 ( .B1(n16269), .B2(n20628), .A(n14018), .ZN(n14019) );
  AND2_X2 U11360 ( .A1(n11184), .A2(n15797), .ZN(n15798) );
  AND2_X2 U11361 ( .A1(n21414), .A2(n15609), .ZN(n21764) );
  NAND3_X2 U11362 ( .A1(n14075), .A2(n14074), .A3(n14073), .ZN(n21290) );
  NOR2_X2 U11363 ( .A1(n14030), .A2(n14028), .ZN(n14108) );
  NAND2_X2 U11364 ( .A1(n21403), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14028) );
  NOR2_X2 U11365 ( .A1(n18543), .A2(n18545), .ZN(n18510) );
  NOR2_X2 U11366 ( .A1(n18502), .A2(n21631), .ZN(n18545) );
  AND2_X1 U11367 ( .A1(n14327), .A2(n11625), .ZN(n11156) );
  OAI21_X1 U11370 ( .B1(n12074), .B2(n11704), .A(n11612), .ZN(n11159) );
  NOR2_X1 U11371 ( .A1(n16652), .A2(n16734), .ZN(n11160) );
  OAI21_X1 U11373 ( .B1(n12074), .B2(n11704), .A(n11612), .ZN(n14290) );
  NOR2_X1 U11374 ( .A1(n16652), .A2(n16734), .ZN(n16650) );
  NAND2_X2 U11375 ( .A1(n11697), .A2(n16624), .ZN(n16652) );
  INV_X1 U11377 ( .A(n17125), .ZN(n11163) );
  INV_X1 U11378 ( .A(n17125), .ZN(n11164) );
  INV_X1 U11380 ( .A(n22730), .ZN(n11166) );
  INV_X1 U11381 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11302) );
  AND2_X2 U11382 ( .A1(n11301), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11309) );
  INV_X1 U11383 ( .A(n11986), .ZN(n11458) );
  INV_X1 U11384 ( .A(n13876), .ZN(n13467) );
  INV_X1 U11385 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U11387 ( .A1(n13182), .A2(n16177), .ZN(n17277) );
  NAND2_X1 U11388 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21848), .ZN(
        n14032) );
  INV_X1 U11389 ( .A(n11826), .ZN(n11174) );
  INV_X2 U11392 ( .A(n13093), .ZN(n16393) );
  XNOR2_X1 U11393 ( .A(n13917), .B(n11267), .ZN(n17082) );
  BUF_X1 U11394 ( .A(n12615), .Z(n12634) );
  XNOR2_X1 U11395 ( .A(n12791), .B(n12792), .ZN(n15056) );
  INV_X1 U11396 ( .A(n19142), .ZN(n17323) );
  INV_X1 U11397 ( .A(n21103), .ZN(n21081) );
  INV_X1 U11398 ( .A(n11838), .ZN(n11854) );
  INV_X1 U11400 ( .A(n22016), .ZN(n22040) );
  AOI21_X1 U11402 ( .B1(n16378), .B2(n17321), .A(n16377), .ZN(n16379) );
  INV_X2 U11403 ( .A(n13705), .ZN(n11217) );
  AND2_X1 U11404 ( .A1(n12796), .A2(n13330), .ZN(n11167) );
  OAI21_X2 U11405 ( .B1(n14871), .B2(n14870), .A(n13062), .ZN(n15054) );
  AND2_X2 U11406 ( .A1(n11260), .A2(n12681), .ZN(n12772) );
  NAND2_X1 U11407 ( .A1(n17085), .A2(n11268), .ZN(n13917) );
  INV_X2 U11409 ( .A(n14603), .ZN(n13765) );
  NAND4_X1 U11411 ( .A1(n20081), .A2(n11176), .A3(n12567), .A4(n13313), .ZN(
        n13271) );
  NOR2_X2 U11412 ( .A1(n20922), .A2(n18608), .ZN(n18376) );
  NAND2_X2 U11413 ( .A1(n18677), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18608) );
  NAND2_X2 U11415 ( .A1(n15056), .A2(n15672), .ZN(n15057) );
  INV_X2 U11417 ( .A(n13300), .ZN(n13301) );
  NAND2_X2 U11418 ( .A1(n12510), .A2(n12509), .ZN(n13300) );
  NAND2_X2 U11420 ( .A1(n15657), .A2(n13901), .ZN(n15811) );
  AND2_X2 U11421 ( .A1(n11211), .A2(n11243), .ZN(n15657) );
  AOI211_X2 U11422 ( .C1(n21700), .C2(n21699), .A(n21698), .B(n21697), .ZN(
        n21712) );
  NAND2_X2 U11424 ( .A1(n12770), .A2(n12769), .ZN(n12791) );
  AOI21_X2 U11425 ( .B1(n17293), .B2(n17290), .A(n16163), .ZN(n13182) );
  NOR2_X4 U11426 ( .A1(n18357), .A2(n21817), .ZN(n21521) );
  OAI211_X2 U11427 ( .C1(n17069), .C2(n17077), .A(n17071), .B(n17075), .ZN(
        n13939) );
  NAND3_X2 U11428 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n21391), .ZN(n18268) );
  INV_X2 U11429 ( .A(n21391), .ZN(n21412) );
  NOR2_X2 U11430 ( .A1(n21851), .A2(n21392), .ZN(n21391) );
  BUF_X2 U11431 ( .A(n15574), .Z(n18255) );
  XNOR2_X2 U11432 ( .A(n13080), .B(n15664), .ZN(n15666) );
  NAND2_X2 U11433 ( .A1(n13079), .A2(n17016), .ZN(n13080) );
  NOR2_X4 U11434 ( .A1(n14031), .A2(n21405), .ZN(n14064) );
  NOR2_X1 U11435 ( .A1(n14031), .A2(n14032), .ZN(n16023) );
  NOR2_X2 U11436 ( .A1(n14030), .A2(n14031), .ZN(n14043) );
  NAND2_X2 U11437 ( .A1(n12458), .A2(n12457), .ZN(n13238) );
  NOR2_X2 U11438 ( .A1(n20789), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20790) );
  CLKBUF_X1 U11439 ( .A(n16638), .Z(n16639) );
  BUF_X1 U11440 ( .A(n16221), .Z(n17232) );
  BUF_X1 U11441 ( .A(n16623), .Z(n16678) );
  NOR2_X1 U11442 ( .A1(n11204), .A2(n15922), .ZN(n16543) );
  AND2_X1 U11443 ( .A1(n17327), .A2(n13189), .ZN(n17316) );
  NAND2_X1 U11444 ( .A1(n15689), .A2(n15688), .ZN(n15866) );
  INV_X1 U11445 ( .A(n16935), .ZN(n11194) );
  NAND2_X1 U11446 ( .A1(n15915), .A2(n15813), .ZN(n16935) );
  NOR2_X2 U11447 ( .A1(n16510), .A2(n16511), .ZN(n16496) );
  INV_X2 U11448 ( .A(n11597), .ZN(n11595) );
  INV_X2 U11449 ( .A(n19024), .ZN(n19054) );
  NOR2_X1 U11451 ( .A1(n18664), .A2(n21431), .ZN(n18299) );
  CLKBUF_X2 U11452 ( .A(n12816), .Z(n19746) );
  AND2_X1 U11453 ( .A1(n12651), .A2(n12650), .ZN(n12813) );
  AND2_X2 U11454 ( .A1(n12647), .A2(n12650), .ZN(n19927) );
  OR2_X1 U11455 ( .A1(n14822), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U11456 ( .A1(n12651), .A2(n12645), .ZN(n19892) );
  OR2_X1 U11457 ( .A1(n11613), .A2(n11473), .ZN(n11499) );
  CLKBUF_X1 U11458 ( .A(n12078), .Z(n16804) );
  XNOR2_X1 U11459 ( .A(n11477), .B(n11476), .ZN(n12078) );
  NAND2_X1 U11460 ( .A1(n11427), .A2(n11426), .ZN(n11477) );
  OAI22_X1 U11461 ( .A1(n12608), .A2(n12550), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16360), .ZN(n12559) );
  NOR2_X1 U11462 ( .A1(n14440), .A2(n14799), .ZN(n14819) );
  NOR2_X1 U11464 ( .A1(n11799), .A2(n11418), .ZN(n11432) );
  INV_X1 U11465 ( .A(n13250), .ZN(n13234) );
  AND2_X1 U11466 ( .A1(n12557), .A2(n12556), .ZN(n17602) );
  NOR2_X2 U11467 ( .A1(n13277), .A2(n19237), .ZN(n12604) );
  NAND2_X1 U11468 ( .A1(n11265), .A2(n12512), .ZN(n13250) );
  AND2_X1 U11469 ( .A1(n11265), .A2(n12534), .ZN(n12955) );
  INV_X4 U11470 ( .A(n20227), .ZN(n19096) );
  AND2_X1 U11471 ( .A1(n11713), .A2(n16332), .ZN(n14279) );
  INV_X2 U11473 ( .A(n19189), .ZN(n14261) );
  INV_X1 U11474 ( .A(n12568), .ZN(n13313) );
  BUF_X1 U11475 ( .A(n12563), .Z(n13232) );
  BUF_X2 U11476 ( .A(n12568), .Z(n14347) );
  OR2_X2 U11477 ( .A1(n11830), .A2(n11826), .ZN(n11913) );
  INV_X2 U11478 ( .A(n12076), .ZN(n11703) );
  INV_X1 U11479 ( .A(n21233), .ZN(n18314) );
  NAND2_X1 U11480 ( .A1(n12528), .A2(n12527), .ZN(n12565) );
  INV_X4 U11481 ( .A(n11838), .ZN(n11173) );
  NAND2_X1 U11482 ( .A1(n12472), .A2(n12471), .ZN(n12563) );
  OR2_X1 U11483 ( .A1(n11349), .A2(n11348), .ZN(n11588) );
  NAND4_X1 U11484 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n14907) );
  NAND2_X1 U11485 ( .A1(n11788), .A2(n11603), .ZN(n11830) );
  INV_X1 U11486 ( .A(n13882), .ZN(n13462) );
  INV_X1 U11487 ( .A(n18006), .ZN(n18253) );
  AND4_X1 U11488 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11370) );
  CLKBUF_X2 U11489 ( .A(n14066), .Z(n21408) );
  BUF_X2 U11490 ( .A(n11483), .Z(n12279) );
  CLKBUF_X2 U11491 ( .A(n12231), .Z(n13535) );
  INV_X1 U11492 ( .A(n13707), .ZN(n13953) );
  BUF_X2 U11493 ( .A(n11950), .Z(n11180) );
  NOR2_X2 U11495 ( .A1(n14028), .A2(n21405), .ZN(n15561) );
  INV_X4 U11497 ( .A(n12459), .ZN(n19079) );
  NAND2_X1 U11498 ( .A1(n21403), .A2(n21392), .ZN(n20778) );
  NAND2_X2 U11499 ( .A1(n21851), .A2(n21848), .ZN(n21405) );
  NOR2_X1 U11500 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13616) );
  XNOR2_X1 U11501 ( .A(n16131), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16146) );
  AND2_X1 U11502 ( .A1(n16130), .A2(n16129), .ZN(n16131) );
  OAI21_X1 U11503 ( .B1(n16389), .B2(n16388), .A(n16387), .ZN(n16396) );
  NAND2_X1 U11504 ( .A1(n16350), .A2(n16349), .ZN(n16389) );
  AOI21_X1 U11505 ( .B1(n16429), .B2(n19157), .A(n16428), .ZN(n16430) );
  AOI211_X1 U11506 ( .C1(n17777), .C2(n17253), .A(n17252), .B(n17251), .ZN(
        n17254) );
  NAND2_X1 U11507 ( .A1(n16214), .A2(n11285), .ZN(n16350) );
  XNOR2_X1 U11508 ( .A(n16398), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16429) );
  OAI21_X1 U11509 ( .B1(n16489), .B2(n16491), .A(n16490), .ZN(n16631) );
  OAI21_X1 U11510 ( .B1(n17257), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17250), .ZN(n17382) );
  AOI21_X1 U11511 ( .B1(n16435), .B2(n16432), .A(n16434), .ZN(n13964) );
  CLKBUF_X1 U11512 ( .A(n17249), .Z(n17257) );
  CLKBUF_X2 U11513 ( .A(n16218), .Z(n17285) );
  AOI211_X1 U11514 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n17814), .A(
        n16419), .B(n16407), .ZN(n16408) );
  OAI22_X1 U11515 ( .A1(n17815), .A2(n11251), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n11250), .ZN(n17239) );
  BUF_X1 U11516 ( .A(n16422), .Z(n16858) );
  OR2_X1 U11517 ( .A1(n13923), .A2(n13922), .ZN(n11213) );
  XNOR2_X1 U11518 ( .A(n16364), .B(n16363), .ZN(n16373) );
  OR2_X2 U11519 ( .A1(n16240), .A2(n14260), .ZN(n17358) );
  OAI21_X1 U11520 ( .B1(n16240), .B2(n16239), .A(n16364), .ZN(n17207) );
  AND2_X1 U11521 ( .A1(n16543), .A2(n16604), .ZN(n16568) );
  NAND2_X1 U11522 ( .A1(n15866), .A2(n11687), .ZN(n15827) );
  AND2_X1 U11523 ( .A1(n11295), .A2(n16899), .ZN(n16400) );
  AND2_X1 U11524 ( .A1(n16899), .A2(n16879), .ZN(n16881) );
  XNOR2_X1 U11525 ( .A(n16256), .B(n16255), .ZN(n16267) );
  AND2_X1 U11526 ( .A1(n15822), .A2(n15963), .ZN(n15920) );
  AOI211_X1 U11527 ( .C1(n21158), .C2(n21157), .A(n21177), .B(n21156), .ZN(
        n21162) );
  AND2_X2 U11528 ( .A1(n11206), .A2(n15721), .ZN(n15822) );
  CLKBUF_X1 U11529 ( .A(n15721), .Z(n15790) );
  OR2_X1 U11530 ( .A1(n16251), .A2(n11838), .ZN(n16252) );
  OR2_X1 U11531 ( .A1(n16353), .A2(n16352), .ZN(n16390) );
  NAND2_X1 U11532 ( .A1(n15100), .A2(n15695), .ZN(n15694) );
  OR2_X1 U11533 ( .A1(n16203), .A2(n14226), .ZN(n16353) );
  NAND2_X1 U11534 ( .A1(n12886), .A2(n12885), .ZN(n15761) );
  AND2_X1 U11537 ( .A1(n15099), .A2(n15103), .ZN(n15100) );
  CLKBUF_X1 U11538 ( .A(n16510), .Z(n16521) );
  AND2_X1 U11539 ( .A1(n15832), .A2(n11594), .ZN(n15930) );
  OR3_X1 U11540 ( .A1(n16910), .A2(n13093), .A3(n17213), .ZN(n16213) );
  AND2_X1 U11541 ( .A1(n11253), .A2(n17416), .ZN(n11252) );
  NOR2_X1 U11542 ( .A1(n12126), .A2(n14930), .ZN(n15099) );
  AOI21_X1 U11543 ( .B1(n12888), .B2(n15664), .A(n12880), .ZN(n12875) );
  NAND2_X1 U11544 ( .A1(n16530), .A2(n16522), .ZN(n16510) );
  NOR2_X1 U11545 ( .A1(n15976), .A2(n11593), .ZN(n15832) );
  NAND2_X1 U11546 ( .A1(n13088), .A2(n18875), .ZN(n13090) );
  OR2_X1 U11547 ( .A1(n11597), .A2(n21921), .ZN(n15830) );
  AND2_X1 U11548 ( .A1(n14222), .A2(n16189), .ZN(n16194) );
  AND2_X1 U11549 ( .A1(n14754), .A2(n14867), .ZN(n14866) );
  NOR2_X1 U11550 ( .A1(n16545), .A2(n16758), .ZN(n11898) );
  NOR2_X1 U11551 ( .A1(n14757), .A2(n14756), .ZN(n14754) );
  CLKBUF_X1 U11552 ( .A(n16545), .Z(n11183) );
  NAND2_X1 U11553 ( .A1(n11587), .A2(n11586), .ZN(n11672) );
  AND2_X1 U11554 ( .A1(n16947), .A2(n16393), .ZN(n16177) );
  CLKBUF_X1 U11555 ( .A(n17171), .Z(n17179) );
  NOR3_X1 U11556 ( .A1(n18473), .A2(n18479), .A3(n18467), .ZN(n18501) );
  AOI211_X1 U11557 ( .C1(n16951), .C2(n16949), .A(n19015), .B(n16948), .ZN(
        n16950) );
  AND2_X1 U11558 ( .A1(n16158), .A2(n11233), .ZN(n19014) );
  NAND2_X1 U11559 ( .A1(n21572), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21732) );
  AND2_X1 U11560 ( .A1(n12105), .A2(n12104), .ZN(n14756) );
  NOR2_X1 U11561 ( .A1(n21755), .A2(n18646), .ZN(n18586) );
  NAND2_X1 U11562 ( .A1(n12094), .A2(n12093), .ZN(n14798) );
  INV_X1 U11563 ( .A(n13177), .ZN(n13180) );
  NAND2_X1 U11564 ( .A1(n14625), .A2(n12085), .ZN(n14797) );
  NAND2_X1 U11565 ( .A1(n18584), .A2(n21770), .ZN(n18583) );
  NOR2_X1 U11566 ( .A1(n19872), .A2(n19925), .ZN(n20355) );
  NAND2_X1 U11567 ( .A1(n13761), .A2(n13760), .ZN(n14427) );
  CLKBUF_X1 U11568 ( .A(n12057), .Z(n14760) );
  NOR2_X1 U11569 ( .A1(n12818), .A2(n12817), .ZN(n12822) );
  CLKBUF_X1 U11570 ( .A(n14479), .Z(n16807) );
  XNOR2_X1 U11571 ( .A(n11599), .B(n11598), .ZN(n12057) );
  NAND2_X1 U11572 ( .A1(n14382), .A2(n13757), .ZN(n14462) );
  NOR2_X2 U11573 ( .A1(n16852), .A2(n19062), .ZN(n16851) );
  XNOR2_X1 U11574 ( .A(n12067), .B(n12068), .ZN(n14479) );
  AND2_X1 U11575 ( .A1(n15842), .A2(n11874), .ZN(n11184) );
  NAND2_X1 U11576 ( .A1(n11500), .A2(n11499), .ZN(n11599) );
  OR2_X1 U11577 ( .A1(n14217), .A2(n14176), .ZN(n16852) );
  AOI22_X1 U11579 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19962), .B1(
        n19927), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12698) );
  OR2_X1 U11580 ( .A1(n14215), .A2(n16886), .ZN(n14217) );
  XNOR2_X1 U11581 ( .A(n11623), .B(n11624), .ZN(n14326) );
  AND2_X1 U11582 ( .A1(n14376), .A2(n13748), .ZN(n14383) );
  NAND2_X1 U11583 ( .A1(n11529), .A2(n11528), .ZN(n11598) );
  NAND2_X1 U11584 ( .A1(n11547), .A2(n11546), .ZN(n14554) );
  NAND2_X1 U11585 ( .A1(n11919), .A2(n11793), .ZN(n22033) );
  NAND2_X1 U11586 ( .A1(n11239), .A2(n11264), .ZN(n19762) );
  NAND2_X1 U11587 ( .A1(n14377), .A2(n14378), .ZN(n14376) );
  NAND2_X2 U11588 ( .A1(n20556), .A2(n14621), .ZN(n16572) );
  XNOR2_X1 U11589 ( .A(n17645), .B(n14631), .ZN(n16842) );
  NAND2_X1 U11590 ( .A1(n14290), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11623) );
  NAND2_X2 U11591 ( .A1(n17690), .A2(n14286), .ZN(n22203) );
  NAND2_X1 U11592 ( .A1(n21871), .A2(n21872), .ZN(n21900) );
  NAND2_X1 U11593 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  AOI21_X1 U11594 ( .B1(n11609), .B2(n11608), .A(n11589), .ZN(n12068) );
  CLKBUF_X1 U11595 ( .A(n12074), .Z(n12075) );
  OR2_X1 U11596 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NAND2_X1 U11597 ( .A1(n11514), .A2(n11513), .ZN(n17645) );
  NOR2_X2 U11598 ( .A1(n19970), .A2(n20286), .ZN(n19971) );
  NOR2_X2 U11599 ( .A1(n20026), .A2(n20288), .ZN(n20027) );
  NOR2_X2 U11600 ( .A1(n19741), .A2(n20286), .ZN(n19742) );
  INV_X2 U11601 ( .A(n18532), .ZN(n21151) );
  XNOR2_X1 U11602 ( .A(n12965), .B(n12966), .ZN(n12962) );
  INV_X1 U11603 ( .A(n21822), .ZN(n21805) );
  NAND2_X1 U11604 ( .A1(n18692), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18691) );
  AND2_X1 U11605 ( .A1(n18289), .A2(n18288), .ZN(n18686) );
  NAND2_X1 U11606 ( .A1(n12616), .A2(n12617), .ZN(n12615) );
  OR2_X1 U11607 ( .A1(n12600), .A2(n12599), .ZN(n12601) );
  XNOR2_X1 U11608 ( .A(n18318), .B(n18317), .ZN(n18692) );
  INV_X1 U11609 ( .A(n18312), .ZN(n18318) );
  AND2_X1 U11610 ( .A1(n15541), .A2(n21388), .ZN(n16121) );
  OAI211_X1 U11612 ( .C1(n12985), .C2(n15058), .A(n12607), .B(n12606), .ZN(
        n12965) );
  NAND2_X1 U11613 ( .A1(n14157), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18568) );
  NAND2_X1 U11614 ( .A1(n12591), .A2(n12590), .ZN(n12592) );
  CLKBUF_X1 U11615 ( .A(n21773), .Z(n21668) );
  OR2_X1 U11616 ( .A1(n13326), .A2(n13323), .ZN(n14407) );
  OAI21_X2 U11617 ( .B1(n20227), .B2(n22264), .A(n14501), .ZN(n14545) );
  AND2_X1 U11618 ( .A1(n11437), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11503) );
  AOI21_X1 U11619 ( .B1(n14488), .B2(n13322), .A(n13321), .ZN(n13326) );
  INV_X2 U11620 ( .A(n20727), .ZN(n20777) );
  NAND2_X1 U11621 ( .A1(n14228), .A2(n18855), .ZN(n12605) );
  AND2_X1 U11622 ( .A1(n14230), .A2(n12571), .ZN(n12585) );
  AND2_X2 U11623 ( .A1(n13234), .A2(n13230), .ZN(n14228) );
  NAND2_X1 U11624 ( .A1(n17602), .A2(n13267), .ZN(n12572) );
  MUX2_X1 U11625 ( .A(n13271), .B(n13262), .S(n12564), .Z(n12580) );
  AND2_X1 U11626 ( .A1(n14396), .A2(n14395), .ZN(n14398) );
  NOR2_X2 U11627 ( .A1(n21439), .A2(n21705), .ZN(n18511) );
  NAND2_X1 U11628 ( .A1(n14025), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14168) );
  AND2_X1 U11629 ( .A1(n11414), .A2(n11412), .ZN(n11711) );
  INV_X1 U11630 ( .A(n13065), .ZN(n13066) );
  XOR2_X1 U11631 ( .A(n18314), .B(n18313), .Z(n18309) );
  AND2_X1 U11632 ( .A1(n12537), .A2(n13301), .ZN(n13266) );
  INV_X1 U11633 ( .A(n12532), .ZN(n12562) );
  MUX2_X1 U11634 ( .A(n13236), .B(n13243), .S(n13238), .Z(n12544) );
  NAND2_X1 U11635 ( .A1(n11235), .A2(n11829), .ZN(n11832) );
  AND2_X1 U11636 ( .A1(n13265), .A2(n12555), .ZN(n12556) );
  AND2_X1 U11637 ( .A1(n14261), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12546) );
  NAND2_X1 U11638 ( .A1(n18326), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18327) );
  OAI21_X1 U11639 ( .B1(n13243), .B2(n12531), .A(n12530), .ZN(n12532) );
  CLKBUF_X2 U11640 ( .A(n13310), .Z(n16414) );
  CLKBUF_X1 U11641 ( .A(n11713), .Z(n14317) );
  NOR2_X1 U11642 ( .A1(n11703), .A2(n22476), .ZN(n12239) );
  AND2_X1 U11643 ( .A1(n11703), .A2(n14621), .ZN(n12058) );
  INV_X2 U11644 ( .A(n21290), .ZN(n21366) );
  AND2_X1 U11645 ( .A1(n12473), .A2(n13239), .ZN(n11265) );
  AND2_X2 U11646 ( .A1(n12529), .A2(n12569), .ZN(n13243) );
  OAI21_X1 U11647 ( .B1(n13238), .B2(n12529), .A(n12554), .ZN(n12530) );
  AND2_X1 U11648 ( .A1(n14559), .A2(n16825), .ZN(n13588) );
  AND2_X1 U11649 ( .A1(n16391), .A2(n19834), .ZN(n13302) );
  AND2_X1 U11650 ( .A1(n11299), .A2(n11805), .ZN(n11713) );
  AND2_X1 U11651 ( .A1(n11717), .A2(n11603), .ZN(n11805) );
  NAND2_X1 U11652 ( .A1(n14587), .A2(n11705), .ZN(n14898) );
  NAND2_X1 U11653 ( .A1(n21000), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18578) );
  INV_X1 U11654 ( .A(n12511), .ZN(n12529) );
  NAND2_X1 U11655 ( .A1(n12076), .A2(n11588), .ZN(n11420) );
  AND2_X1 U11656 ( .A1(n12568), .A2(n12564), .ZN(n13239) );
  NAND3_X1 U11657 ( .A1(n14097), .A2(n14096), .A3(n14095), .ZN(n19358) );
  INV_X2 U11658 ( .A(n11705), .ZN(n16332) );
  BUF_X2 U11659 ( .A(n12511), .Z(n12567) );
  NAND2_X1 U11660 ( .A1(n11408), .A2(n11588), .ZN(n11794) );
  INV_X1 U11662 ( .A(n11410), .ZN(n11717) );
  AND2_X2 U11663 ( .A1(n14587), .A2(n14907), .ZN(n14909) );
  INV_X2 U11664 ( .A(n12569), .ZN(n11176) );
  INV_X1 U11665 ( .A(n11830), .ZN(n11838) );
  OAI21_X2 U11666 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n14669) );
  OAI21_X2 U11667 ( .B1(n14668), .B2(n16004), .A(n14556), .ZN(n14557) );
  INV_X1 U11668 ( .A(n11603), .ZN(n14580) );
  NAND2_X1 U11669 ( .A1(n12456), .A2(n12519), .ZN(n12457) );
  INV_X2 U11670 ( .A(U212), .ZN(n11177) );
  NAND2_X2 U11671 ( .A1(U214), .A2(n20640), .ZN(n20706) );
  INV_X2 U11672 ( .A(n12753), .ZN(n11219) );
  AND4_X1 U11673 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11390) );
  AND4_X1 U11674 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11392) );
  INV_X2 U11675 ( .A(n18006), .ZN(n18271) );
  CLKBUF_X3 U11676 ( .A(n13953), .Z(n13940) );
  AOI22_X1 U11677 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11320) );
  NAND2_X2 U11678 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17942), .ZN(n17936) );
  AND4_X1 U11679 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11391) );
  AND4_X1 U11680 ( .A1(n11377), .A2(n11376), .A3(n11375), .A4(n11374), .ZN(
        n11393) );
  AND2_X2 U11681 ( .A1(n12663), .A2(n13616), .ZN(n12701) );
  INV_X2 U11682 ( .A(n20500), .ZN(n11178) );
  NAND2_X1 U11683 ( .A1(n13615), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12753) );
  BUF_X2 U11684 ( .A(n16023), .Z(n18254) );
  INV_X2 U11685 ( .A(n18834), .ZN(n18841) );
  CLKBUF_X3 U11686 ( .A(n14064), .Z(n18244) );
  INV_X2 U11687 ( .A(n20402), .ZN(n20449) );
  NAND2_X2 U11688 ( .A1(n22270), .A2(n17855), .ZN(n17939) );
  OR2_X1 U11690 ( .A1(n14028), .A2(n21404), .ZN(n18063) );
  NOR2_X1 U11691 ( .A1(n18746), .A2(n18744), .ZN(n21886) );
  AND2_X2 U11692 ( .A1(n12420), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12664) );
  AND2_X1 U11693 ( .A1(n11304), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11313) );
  AND2_X2 U11694 ( .A1(n11303), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16828) );
  INV_X1 U11695 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17059) );
  INV_X2 U11696 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12420) );
  INV_X1 U11697 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11303) );
  OAI21_X1 U11698 ( .B1(n18511), .B2(n21817), .A(n18374), .ZN(n18623) );
  AOI21_X1 U11700 ( .B1(n12608), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12595), .ZN(n12600) );
  NOR2_X1 U11701 ( .A1(n17279), .A2(n17278), .ZN(n17283) );
  NOR2_X1 U11702 ( .A1(n13184), .A2(n17279), .ZN(n13261) );
  OAI21_X1 U11703 ( .B1(n17212), .B2(n16208), .A(n16207), .ZN(n16210) );
  NAND2_X1 U11704 ( .A1(n13163), .A2(n13164), .ZN(n13171) );
  CLKBUF_X1 U11705 ( .A(n17747), .Z(n11181) );
  NAND2_X1 U11706 ( .A1(n15057), .A2(n12794), .ZN(n11182) );
  NAND2_X1 U11707 ( .A1(n15057), .A2(n12794), .ZN(n12879) );
  AOI21_X2 U11708 ( .B1(n18521), .B2(n18619), .A(n11269), .ZN(n18502) );
  NOR2_X1 U11709 ( .A1(n15908), .A2(n15895), .ZN(n11185) );
  NOR2_X1 U11710 ( .A1(n15120), .A2(n15119), .ZN(n11186) );
  NAND2_X1 U11711 ( .A1(n16546), .A2(n16547), .ZN(n16545) );
  NOR2_X1 U11712 ( .A1(n15908), .A2(n15895), .ZN(n15842) );
  NAND2_X1 U11713 ( .A1(n15697), .A2(n15906), .ZN(n15908) );
  NOR2_X1 U11714 ( .A1(n15120), .A2(n15119), .ZN(n15122) );
  BUF_X1 U11715 ( .A(n19794), .Z(n19798) );
  NAND2_X1 U11716 ( .A1(n11788), .A2(n11224), .ZN(n11826) );
  OR2_X2 U11717 ( .A1(n13122), .A2(n13123), .ZN(n13125) );
  NAND2_X1 U11718 ( .A1(n12796), .A2(n13330), .ZN(n11187) );
  NAND2_X1 U11720 ( .A1(n17785), .A2(n17786), .ZN(n11189) );
  INV_X1 U11721 ( .A(n19877), .ZN(n11190) );
  INV_X1 U11722 ( .A(n11190), .ZN(n11191) );
  AND2_X1 U11724 ( .A1(n12651), .A2(n12649), .ZN(n19877) );
  NAND2_X1 U11725 ( .A1(n11712), .A2(n14587), .ZN(n11192) );
  AND2_X1 U11727 ( .A1(n16916), .A2(n11195), .ZN(n11196) );
  INV_X1 U11728 ( .A(n16936), .ZN(n11195) );
  AND2_X1 U11729 ( .A1(n11194), .A2(n11195), .ZN(n16934) );
  NOR2_X2 U11730 ( .A1(n17090), .A2(n16900), .ZN(n16899) );
  NOR2_X1 U11731 ( .A1(n11701), .A2(n16127), .ZN(n16129) );
  NOR2_X1 U11732 ( .A1(n11263), .A2(n11262), .ZN(n11261) );
  INV_X1 U11733 ( .A(n14874), .ZN(n11197) );
  AND2_X1 U11734 ( .A1(n11198), .A2(n14875), .ZN(n15063) );
  NOR2_X1 U11735 ( .A1(n13334), .A2(n11197), .ZN(n11198) );
  AND2_X1 U11736 ( .A1(n18927), .A2(n11199), .ZN(n17476) );
  AND2_X1 U11737 ( .A1(n18928), .A2(n17504), .ZN(n11199) );
  NOR2_X1 U11738 ( .A1(n16999), .A2(n13364), .ZN(n11200) );
  NOR2_X1 U11739 ( .A1(n15732), .A2(n15733), .ZN(n17196) );
  NOR2_X1 U11740 ( .A1(n16999), .A2(n13364), .ZN(n17002) );
  NOR2_X1 U11741 ( .A1(n13326), .A2(n13325), .ZN(n14875) );
  NOR2_X1 U11742 ( .A1(n12126), .A2(n14930), .ZN(n11202) );
  AND2_X1 U11743 ( .A1(n11561), .A2(n11640), .ZN(n11203) );
  OR2_X1 U11744 ( .A1(n16544), .A2(n16002), .ZN(n11204) );
  OR2_X1 U11745 ( .A1(n15922), .A2(n16002), .ZN(n16001) );
  INV_X1 U11746 ( .A(n12262), .ZN(n11205) );
  NOR2_X1 U11747 ( .A1(n15821), .A2(n11205), .ZN(n11206) );
  OAI21_X1 U11748 ( .B1(n14932), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11455), 
        .ZN(n11207) );
  XNOR2_X1 U11749 ( .A(n13556), .B(n13555), .ZN(n11208) );
  OAI21_X1 U11750 ( .B1(n14932), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11455), 
        .ZN(n11613) );
  XNOR2_X1 U11751 ( .A(n13556), .B(n13555), .ZN(n16269) );
  XNOR2_X1 U11752 ( .A(n11672), .B(n11671), .ZN(n12054) );
  XNOR2_X1 U11753 ( .A(n11832), .B(n11831), .ZN(n14325) );
  NAND2_X1 U11754 ( .A1(n14999), .A2(n14998), .ZN(n11209) );
  NAND2_X1 U11755 ( .A1(n14999), .A2(n14998), .ZN(n14997) );
  INV_X1 U11757 ( .A(n15130), .ZN(n11210) );
  NOR2_X1 U11758 ( .A1(n13767), .A2(n11210), .ZN(n11211) );
  AND2_X1 U11760 ( .A1(n11416), .A2(n14621), .ZN(n11371) );
  CLKBUF_X1 U11761 ( .A(n17095), .Z(n11214) );
  NOR2_X1 U11762 ( .A1(n13923), .A2(n13922), .ZN(n17069) );
  AND2_X2 U11763 ( .A1(n17122), .A2(n17111), .ZN(n13034) );
  OR2_X2 U11764 ( .A1(n16882), .A2(n16883), .ZN(n16885) );
  AND2_X1 U11765 ( .A1(n13759), .A2(n13758), .ZN(n13760) );
  OAI21_X2 U11766 ( .B1(n14411), .B2(n19215), .A(n13753), .ZN(n13756) );
  AND2_X2 U11767 ( .A1(n11312), .A2(n14304), .ZN(n11215) );
  AND2_X2 U11768 ( .A1(n12614), .A2(n12613), .ZN(n14411) );
  NAND2_X1 U11769 ( .A1(n13021), .A2(n13020), .ZN(n15716) );
  NOR2_X2 U11770 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NOR2_X2 U11771 ( .A1(n11233), .A2(n14221), .ZN(n16182) );
  OR2_X2 U11772 ( .A1(n16157), .A2(n16156), .ZN(n11233) );
  AND2_X2 U11773 ( .A1(n13739), .A2(n13759), .ZN(n14461) );
  AND2_X1 U11774 ( .A1(n11313), .A2(n11312), .ZN(n11950) );
  AND2_X2 U11775 ( .A1(n14920), .A2(n14921), .ZN(n11243) );
  XNOR2_X1 U11776 ( .A(n14398), .B(n13312), .ZN(n14483) );
  AND2_X2 U11777 ( .A1(n15991), .A2(n15990), .ZN(n15989) );
  AND2_X1 U11778 ( .A1(n16829), .A2(n14304), .ZN(n11216) );
  AND2_X2 U11779 ( .A1(n15989), .A2(n16773), .ZN(n16546) );
  INV_X1 U11780 ( .A(n13647), .ZN(n11218) );
  INV_X2 U11781 ( .A(n13707), .ZN(n11220) );
  NAND2_X1 U11782 ( .A1(n13299), .A2(n11283), .ZN(n13983) );
  INV_X4 U11783 ( .A(n13715), .ZN(n13941) );
  AOI211_X2 U11784 ( .C1(n16378), .C2(n19157), .A(n16369), .B(n16368), .ZN(
        n16370) );
  NOR2_X4 U11785 ( .A1(n17475), .A2(n12922), .ZN(n17797) );
  OR2_X2 U11786 ( .A1(n17472), .A2(n17473), .ZN(n17475) );
  NOR2_X4 U11787 ( .A1(n15108), .A2(n15107), .ZN(n15699) );
  OR2_X2 U11788 ( .A1(n15093), .A2(n15713), .ZN(n15108) );
  AND2_X2 U11789 ( .A1(n15699), .A2(n15698), .ZN(n15697) );
  OAI21_X2 U11790 ( .B1(n15811), .B2(n17100), .A(n13905), .ZN(n17097) );
  AOI21_X2 U11791 ( .B1(n15827), .B2(n11690), .A(n11240), .ZN(n11692) );
  INV_X2 U11792 ( .A(n11416), .ZN(n11408) );
  NAND4_X1 U11793 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11224) );
  AND2_X1 U11794 ( .A1(n16828), .A2(n11309), .ZN(n11225) );
  AND2_X1 U11795 ( .A1(n16828), .A2(n11309), .ZN(n11226) );
  AND2_X1 U11796 ( .A1(n16828), .A2(n11309), .ZN(n11361) );
  INV_X1 U11797 ( .A(n11174), .ZN(n11228) );
  INV_X1 U11798 ( .A(n11174), .ZN(n11229) );
  AND2_X4 U11799 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14304) );
  INV_X1 U11800 ( .A(n11984), .ZN(n11230) );
  NOR2_X2 U11801 ( .A1(n15750), .A2(n15751), .ZN(n15749) );
  OR2_X1 U11802 ( .A1(n16267), .A2(n22017), .ZN(n11238) );
  NAND2_X1 U11803 ( .A1(n14580), .A2(n14907), .ZN(n11231) );
  NAND2_X1 U11804 ( .A1(n14580), .A2(n14907), .ZN(n11907) );
  AOI22_X1 U11805 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16423), .B1(n16409), 
        .B2(n19237), .ZN(n11232) );
  OR2_X2 U11806 ( .A1(n12411), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22016) );
  AND3_X1 U11807 ( .A1(n13247), .A2(n13246), .A3(n13263), .ZN(n13281) );
  OR2_X1 U11808 ( .A1(n11489), .A2(n11488), .ZN(n11610) );
  NAND2_X1 U11809 ( .A1(n11456), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11736) );
  INV_X1 U11810 ( .A(n11803), .ZN(n11456) );
  NOR2_X1 U11811 ( .A1(n13238), .A2(n12563), .ZN(n12473) );
  NAND2_X1 U11812 ( .A1(n18686), .A2(n21426), .ZN(n18293) );
  NAND2_X1 U11813 ( .A1(n11416), .A2(n16332), .ZN(n11803) );
  AND2_X1 U11814 ( .A1(n11803), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11744) );
  INV_X1 U11815 ( .A(n13338), .ZN(n13084) );
  INV_X1 U11816 ( .A(n12893), .ZN(n12895) );
  NAND2_X1 U11817 ( .A1(n18865), .A2(n13743), .ZN(n13745) );
  OAI21_X1 U11818 ( .B1(n12552), .B2(n13298), .A(n12551), .ZN(n12557) );
  NAND2_X1 U11819 ( .A1(n12564), .A2(n13243), .ZN(n12551) );
  NAND2_X1 U11820 ( .A1(n12562), .A2(n12561), .ZN(n14230) );
  AOI21_X1 U11821 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19905), .A(
        n12932), .ZN(n12934) );
  INV_X1 U11822 ( .A(n12936), .ZN(n12931) );
  AND2_X1 U11823 ( .A1(n14127), .A2(n21389), .ZN(n16013) );
  AOI21_X1 U11824 ( .B1(n14138), .B2(n14137), .A(n14136), .ZN(n15535) );
  INV_X1 U11825 ( .A(n21836), .ZN(n18307) );
  NAND2_X1 U11826 ( .A1(n22095), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14916) );
  AND2_X1 U11827 ( .A1(n16461), .A2(n14278), .ZN(n14286) );
  AND2_X1 U11828 ( .A1(n11783), .A2(n14278), .ZN(n11919) );
  NOR2_X1 U11829 ( .A1(n19129), .A2(n13186), .ZN(n17757) );
  INV_X1 U11830 ( .A(n20015), .ZN(n19883) );
  NAND2_X1 U11831 ( .A1(n19749), .A2(n19775), .ZN(n19904) );
  NAND2_X1 U11832 ( .A1(n19749), .A2(n20282), .ZN(n19884) );
  NOR2_X1 U11833 ( .A1(n16413), .A2(n16412), .ZN(n16417) );
  INV_X1 U11834 ( .A(n21773), .ZN(n21685) );
  INV_X1 U11835 ( .A(n11168), .ZN(n11982) );
  NAND2_X1 U11836 ( .A1(n13238), .A2(n12568), .ZN(n12554) );
  AND2_X1 U11837 ( .A1(n11585), .A2(n11584), .ZN(n11659) );
  AND2_X2 U11838 ( .A1(n11302), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11312) );
  OR2_X1 U11839 ( .A1(n11545), .A2(n11544), .ZN(n11642) );
  INV_X1 U11840 ( .A(n11736), .ZN(n11760) );
  OR3_X1 U11841 ( .A1(n17469), .A2(n17493), .A3(n13127), .ZN(n16160) );
  AND3_X1 U11842 ( .A1(n12698), .A2(n12699), .A3(n12700), .ZN(n11258) );
  NAND2_X1 U11843 ( .A1(n11176), .A2(n13301), .ZN(n13298) );
  AND3_X1 U11844 ( .A1(n12568), .A2(n12563), .A3(n12569), .ZN(n12533) );
  AOI22_X1 U11845 ( .A1(n13615), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12429) );
  AND2_X1 U11846 ( .A1(n19856), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12940) );
  INV_X1 U11847 ( .A(n21242), .ZN(n15615) );
  NOR2_X1 U11848 ( .A1(n15519), .A2(n15518), .ZN(n14132) );
  AND2_X1 U11849 ( .A1(n12261), .A2(n15722), .ZN(n12262) );
  NOR2_X1 U11850 ( .A1(n11422), .A2(n22210), .ZN(n13545) );
  AND2_X1 U11851 ( .A1(n15724), .A2(n15723), .ZN(n15722) );
  NOR2_X1 U11852 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12312) );
  OR2_X1 U11853 ( .A1(n14621), .A2(n22476), .ZN(n12405) );
  INV_X1 U11854 ( .A(n12312), .ZN(n12400) );
  OR2_X1 U11855 ( .A1(n20593), .A2(n21977), .ZN(n11687) );
  NAND2_X1 U11856 ( .A1(n14287), .A2(n15726), .ZN(n11704) );
  NAND2_X1 U11857 ( .A1(n12078), .A2(n22210), .ZN(n11493) );
  OAI21_X1 U11858 ( .B1(n11736), .B2(n11497), .A(n11496), .ZN(n11608) );
  NAND2_X1 U11859 ( .A1(n11439), .A2(n14561), .ZN(n11505) );
  INV_X1 U11860 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14307) );
  NOR2_X2 U11861 ( .A1(n13162), .A2(n13161), .ZN(n13163) );
  NOR2_X2 U11862 ( .A1(n13125), .A2(n13118), .ZN(n13119) );
  CLKBUF_X3 U11863 ( .A(n12711), .Z(n13865) );
  AND2_X1 U11864 ( .A1(n12874), .A2(n12873), .ZN(n12894) );
  OR2_X1 U11865 ( .A1(n12855), .A2(n12854), .ZN(n12874) );
  NAND2_X1 U11866 ( .A1(n13730), .A2(n19834), .ZN(n13752) );
  INV_X1 U11867 ( .A(n14228), .ZN(n13294) );
  NOR3_X1 U11868 ( .A1(n13270), .A2(n13996), .A3(n16391), .ZN(n12570) );
  NAND2_X1 U11869 ( .A1(n12439), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12446) );
  NAND2_X1 U11870 ( .A1(n12444), .A2(n12519), .ZN(n12445) );
  AOI221_X1 U11871 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12934), 
        .C1(n19101), .C2(n12934), .A(n12933), .ZN(n13228) );
  NOR2_X1 U11872 ( .A1(n14030), .A2(n20778), .ZN(n15574) );
  NOR2_X1 U11873 ( .A1(n14032), .A2(n20778), .ZN(n14087) );
  NOR2_X1 U11874 ( .A1(n14028), .A2(n14032), .ZN(n15563) );
  OR2_X1 U11875 ( .A1(n18224), .A2(n15542), .ZN(n16117) );
  OR2_X1 U11876 ( .A1(n21492), .A2(n18321), .ZN(n18322) );
  NAND2_X1 U11877 ( .A1(n18293), .A2(n18292), .ZN(n18295) );
  OR2_X1 U11878 ( .A1(n18686), .A2(n21426), .ZN(n18294) );
  INV_X1 U11879 ( .A(n18687), .ZN(n18292) );
  INV_X1 U11880 ( .A(n21228), .ZN(n18316) );
  NOR2_X1 U11881 ( .A1(n21366), .A2(n19476), .ZN(n15545) );
  OAI22_X1 U11882 ( .A1(n21392), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n21855), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15519) );
  INV_X1 U11883 ( .A(n19476), .ZN(n14126) );
  INV_X1 U11884 ( .A(n12058), .ZN(n13577) );
  INV_X1 U11885 ( .A(n22220), .ZN(n14278) );
  INV_X1 U11886 ( .A(n12405), .ZN(n13553) );
  NAND2_X1 U11887 ( .A1(n12389), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12401) );
  NAND2_X1 U11888 ( .A1(n12065), .A2(n12064), .ZN(n14624) );
  NAND2_X1 U11889 ( .A1(n11535), .A2(n11534), .ZN(n14631) );
  AND2_X1 U11890 ( .A1(n11770), .A2(n11769), .ZN(n16461) );
  NAND2_X1 U11891 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  XNOR2_X1 U11892 ( .A(n17095), .B(n13910), .ZN(n17087) );
  NAND2_X1 U11893 ( .A1(n17002), .A2(n16991), .ZN(n17550) );
  NAND2_X1 U11894 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n14206), .ZN(
        n14210) );
  NOR2_X2 U11895 ( .A1(n19005), .A2(n14207), .ZN(n14206) );
  NAND2_X1 U11896 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n14192), .ZN(
        n14197) );
  NOR2_X2 U11897 ( .A1(n18930), .A2(n14197), .ZN(n14196) );
  AND2_X1 U11898 ( .A1(n13507), .A2(n13506), .ZN(n15733) );
  AND2_X1 U11899 ( .A1(n13259), .A2(n18852), .ZN(n13523) );
  INV_X1 U11900 ( .A(n13746), .ZN(n14350) );
  AND2_X1 U11901 ( .A1(n17614), .A2(n17613), .ZN(n19184) );
  INV_X1 U11902 ( .A(n19892), .ZN(n19897) );
  INV_X1 U11903 ( .A(n19953), .ZN(n19939) );
  NAND2_X1 U11904 ( .A1(n11237), .A2(n11264), .ZN(n19787) );
  NAND2_X1 U11905 ( .A1(n19814), .A2(n19775), .ZN(n19946) );
  AND2_X1 U11906 ( .A1(n19959), .A2(n19939), .ZN(n19955) );
  NAND2_X1 U11907 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19959), .ZN(n20288) );
  INV_X1 U11908 ( .A(n19959), .ZN(n20286) );
  NAND4_X1 U11909 ( .A1(n21252), .A2(n15545), .A3(n14129), .A4(n18802), .ZN(
        n18223) );
  CLKBUF_X2 U11910 ( .A(n15561), .Z(n18269) );
  NAND2_X1 U11911 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21848), .ZN(
        n14033) );
  BUF_X1 U11912 ( .A(n15561), .Z(n18245) );
  BUF_X1 U11913 ( .A(n14087), .Z(n18246) );
  AOI21_X1 U11914 ( .B1(n16013), .B2(n16012), .A(n16119), .ZN(n21194) );
  OR2_X1 U11915 ( .A1(n18308), .A2(n21225), .ZN(n21705) );
  OR2_X1 U11916 ( .A1(n21903), .A2(n14896), .ZN(n22095) );
  XNOR2_X1 U11917 ( .A(n11702), .B(n16127), .ZN(n12418) );
  INV_X1 U11918 ( .A(n19775), .ZN(n20282) );
  INV_X1 U11919 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18930) );
  NOR2_X1 U11920 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  OR2_X1 U11921 ( .A1(n17757), .A2(n13187), .ZN(n17515) );
  AND2_X1 U11922 ( .A1(n17789), .A2(n14341), .ZN(n17777) );
  INV_X1 U11923 ( .A(n17789), .ZN(n17814) );
  OAI21_X1 U11924 ( .B1(n16858), .B2(n19130), .A(n11272), .ZN(n16425) );
  AOI21_X1 U11925 ( .B1(n19707), .B2(n19154), .A(n16421), .ZN(n16427) );
  OR2_X1 U11926 ( .A1(n16420), .A2(n16419), .ZN(n16421) );
  INV_X1 U11927 ( .A(n19134), .ZN(n19154) );
  INV_X1 U11928 ( .A(n19159), .ZN(n19130) );
  NAND2_X1 U11929 ( .A1(n19835), .A2(n19834), .ZN(n19953) );
  INV_X1 U11930 ( .A(n14461), .ZN(n14463) );
  INV_X1 U11931 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19905) );
  INV_X1 U11932 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19181) );
  NAND2_X1 U11933 ( .A1(n14376), .A2(n14379), .ZN(n19749) );
  OR2_X1 U11934 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  INV_X1 U11935 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18267) );
  INV_X1 U11936 ( .A(n21735), .ZN(n21700) );
  INV_X1 U11937 ( .A(n21813), .ZN(n21828) );
  AOI21_X1 U11938 ( .B1(n15539), .B2(n15538), .A(n21897), .ZN(n21773) );
  AND2_X1 U11939 ( .A1(n16829), .A2(n14473), .ZN(n11333) );
  OR2_X1 U11940 ( .A1(n11454), .A2(n11453), .ZN(n11614) );
  OR2_X1 U11941 ( .A1(n11588), .A2(n12076), .ZN(n11415) );
  OAI21_X1 U11942 ( .B1(n19794), .B2(n12693), .A(n19096), .ZN(n12694) );
  NAND2_X1 U11943 ( .A1(n12569), .A2(n12567), .ZN(n12542) );
  OAI21_X1 U11944 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21851), .A(
        n14133), .ZN(n14134) );
  OR2_X1 U11945 ( .A1(n14137), .A2(n14138), .ZN(n14133) );
  NAND2_X1 U11946 ( .A1(n11373), .A2(n11422), .ZN(n11414) );
  NOR2_X1 U11947 ( .A1(n11794), .A2(n14907), .ZN(n11412) );
  NAND2_X1 U11948 ( .A1(n15694), .A2(n12161), .ZN(n15721) );
  NAND2_X1 U11949 ( .A1(n11203), .A2(n11649), .ZN(n11660) );
  OR2_X1 U11950 ( .A1(n11468), .A2(n11467), .ZN(n11681) );
  OR2_X1 U11951 ( .A1(n11583), .A2(n11582), .ZN(n11674) );
  NOR2_X1 U11952 ( .A1(n11416), .A2(n22210), .ZN(n11490) );
  INV_X1 U11953 ( .A(n11681), .ZN(n11669) );
  NAND2_X1 U11954 ( .A1(n11760), .A2(n11746), .ZN(n11761) );
  AOI22_X1 U11955 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11216), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11315) );
  NOR2_X2 U11956 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12659) );
  AND2_X2 U11957 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U11958 ( .A1(n11167), .A2(n12838), .ZN(n12893) );
  XNOR2_X1 U11959 ( .A(n12893), .B(n12894), .ZN(n13083) );
  XNOR2_X1 U11960 ( .A(n11187), .B(n12838), .ZN(n13072) );
  NAND2_X1 U11961 ( .A1(n12657), .A2(n12639), .ZN(n11262) );
  NOR2_X1 U11962 ( .A1(n12633), .A2(n12632), .ZN(n12642) );
  OAI22_X1 U11963 ( .A1(n12636), .A2(n19762), .B1(n19787), .B2(n13678), .ZN(
        n12637) );
  NAND2_X1 U11964 ( .A1(n12531), .A2(n13736), .ZN(n12552) );
  INV_X2 U11965 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17630) );
  AND2_X1 U11966 ( .A1(n14399), .A2(n14411), .ZN(n12644) );
  AOI22_X1 U11967 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U11968 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U11969 ( .A1(n12930), .A2(n12929), .ZN(n12936) );
  INV_X1 U11970 ( .A(n12400), .ZN(n13548) );
  AND2_X1 U11971 ( .A1(n12260), .A2(n15789), .ZN(n15723) );
  AND2_X1 U11972 ( .A1(n12096), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12107) );
  NOR2_X1 U11973 ( .A1(n12086), .A2(n11922), .ZN(n12087) );
  INV_X1 U11974 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11922) );
  NOR2_X1 U11975 ( .A1(n11669), .A2(n11498), .ZN(n11589) );
  OAI211_X1 U11976 ( .C1(n15930), .C2(n20617), .A(n15933), .B(n15932), .ZN(
        n20615) );
  INV_X1 U11977 ( .A(n11704), .ZN(n11746) );
  AND2_X1 U11978 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  OR2_X1 U11979 ( .A1(n11761), .A2(n11777), .ZN(n11768) );
  INV_X1 U11980 ( .A(n11588), .ZN(n11407) );
  NAND3_X1 U11981 ( .A1(n22207), .A2(n17722), .A3(n16845), .ZN(n14558) );
  INV_X1 U11982 ( .A(n12075), .ZN(n14630) );
  INV_X1 U11983 ( .A(n22469), .ZN(n14934) );
  NAND2_X1 U11984 ( .A1(n16842), .A2(n22210), .ZN(n11547) );
  NOR2_X2 U11985 ( .A1(n13171), .A2(n13170), .ZN(n13177) );
  NAND2_X1 U11986 ( .A1(n13104), .A2(n11244), .ZN(n13109) );
  INV_X1 U11987 ( .A(n13103), .ZN(n13104) );
  NAND2_X1 U11988 ( .A1(n12610), .A2(n12609), .ZN(n12966) );
  INV_X1 U11989 ( .A(n13057), .ZN(n13051) );
  AND2_X1 U11990 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  INV_X1 U11991 ( .A(n12592), .ZN(n12622) );
  AOI21_X1 U11992 ( .B1(n12603), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12598), .ZN(n12599) );
  NAND2_X2 U11993 ( .A1(n12660), .A2(n17630), .ZN(n13713) );
  OR2_X1 U11994 ( .A1(n19193), .A2(n13965), .ZN(n19202) );
  AND2_X1 U11995 ( .A1(n18855), .A2(n13736), .ZN(n13918) );
  AND2_X1 U11996 ( .A1(n16152), .A2(n16151), .ZN(n17463) );
  NAND2_X1 U11997 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n14190), .ZN(
        n14189) );
  NOR2_X1 U11998 ( .A1(n17816), .A2(n19112), .ZN(n11251) );
  INV_X1 U11999 ( .A(n17816), .ZN(n11250) );
  AND2_X1 U12000 ( .A1(n13510), .A2(n13509), .ZN(n18985) );
  NOR2_X1 U12001 ( .A1(n16160), .A2(n13133), .ZN(n13134) );
  NAND2_X1 U12002 ( .A1(n17745), .A2(n12921), .ZN(n13185) );
  NAND2_X1 U12003 ( .A1(n12837), .A2(n12836), .ZN(n12888) );
  INV_X1 U12004 ( .A(n11182), .ZN(n12837) );
  OR2_X1 U12005 ( .A1(n12872), .A2(n12871), .ZN(n13338) );
  NAND2_X1 U12006 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  NAND2_X1 U12007 ( .A1(n12691), .A2(n11234), .ZN(n11259) );
  NAND2_X1 U12008 ( .A1(n12508), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12509) );
  NAND2_X1 U12009 ( .A1(n12724), .A2(n12723), .ZN(n13303) );
  NAND2_X1 U12010 ( .A1(n11154), .A2(n11266), .ZN(n12582) );
  AND2_X2 U12011 ( .A1(n12419), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12663) );
  INV_X2 U12012 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12419) );
  AND2_X1 U12013 ( .A1(n17595), .A2(n14399), .ZN(n12650) );
  NAND2_X1 U12014 ( .A1(n12520), .A2(n12519), .ZN(n12528) );
  NAND2_X1 U12015 ( .A1(n12426), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12434) );
  NOR2_X2 U12016 ( .A1(n18327), .A2(n18400), .ZN(n14025) );
  NOR2_X2 U12017 ( .A1(n18578), .A2(n18577), .ZN(n18326) );
  NAND2_X1 U12018 ( .A1(n18657), .A2(n18658), .ZN(n18374) );
  XNOR2_X1 U12019 ( .A(n15615), .B(n15581), .ZN(n15583) );
  AOI21_X1 U12020 ( .B1(n14130), .B2(n16013), .A(n14131), .ZN(n15608) );
  NOR2_X1 U12021 ( .A1(n14128), .A2(n14126), .ZN(n21389) );
  NOR3_X1 U12022 ( .A1(n18802), .A2(n14126), .A3(n21366), .ZN(n14119) );
  NOR2_X1 U12023 ( .A1(n19358), .A2(n15530), .ZN(n14129) );
  INV_X1 U12024 ( .A(n15525), .ZN(n14127) );
  NOR2_X1 U12025 ( .A1(n15543), .A2(n21195), .ZN(n15524) );
  AND3_X1 U12026 ( .A1(n14120), .A2(n14119), .A3(n15536), .ZN(n15541) );
  CLKBUF_X1 U12027 ( .A(n14279), .Z(n16463) );
  NAND2_X1 U12028 ( .A1(n16834), .A2(n14286), .ZN(n16331) );
  CLKBUF_X1 U12029 ( .A(n11711), .Z(n11712) );
  AND2_X1 U12030 ( .A1(n11873), .A2(n11872), .ZN(n15843) );
  INV_X1 U12031 ( .A(n16461), .ZN(n16459) );
  AND2_X1 U12032 ( .A1(n12314), .A2(n12313), .ZN(n15924) );
  AOI21_X1 U12033 ( .B1(n16331), .B2(n22387), .A(n22254), .ZN(n20453) );
  OR2_X1 U12034 ( .A1(n12401), .A2(n11926), .ZN(n11928) );
  OR2_X1 U12035 ( .A1(n11928), .A2(n11927), .ZN(n14015) );
  AND2_X1 U12037 ( .A1(n11925), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12389) );
  AND2_X1 U12038 ( .A1(n11924), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12372) );
  CLKBUF_X1 U12039 ( .A(n16514), .Z(n16515) );
  AND2_X1 U12041 ( .A1(n12361), .A2(n12360), .ZN(n16604) );
  OR2_X1 U12042 ( .A1(n22187), .A2(n12400), .ZN(n12360) );
  AOI21_X1 U12043 ( .B1(n11691), .B2(n11277), .A(n11595), .ZN(n16685) );
  CLKBUF_X1 U12044 ( .A(n16543), .Z(n16605) );
  AND2_X1 U12045 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11923), .ZN(
        n12329) );
  CLKBUF_X1 U12046 ( .A(n15922), .Z(n15923) );
  AND2_X1 U12047 ( .A1(n12263), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12294) );
  NAND2_X1 U12048 ( .A1(n12294), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12311) );
  CLKBUF_X1 U12049 ( .A(n15920), .Z(n15921) );
  BUF_X1 U12050 ( .A(n11692), .Z(n16693) );
  NAND2_X1 U12051 ( .A1(n12179), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12162) );
  AND2_X1 U12052 ( .A1(n12210), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12195) );
  NOR2_X1 U12053 ( .A1(n12225), .A2(n12226), .ZN(n12210) );
  NOR2_X1 U12054 ( .A1(n12127), .A2(n12128), .ZN(n12147) );
  NAND2_X1 U12055 ( .A1(n12147), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U12056 ( .A1(n12021), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12127) );
  CLKBUF_X1 U12057 ( .A(n15100), .Z(n15101) );
  AND2_X1 U12058 ( .A1(n12049), .A2(n12048), .ZN(n15633) );
  OR2_X1 U12059 ( .A1(n15632), .A2(n15633), .ZN(n15685) );
  NAND2_X1 U12060 ( .A1(n12116), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12050) );
  AND2_X1 U12061 ( .A1(n12107), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12116) );
  NAND2_X1 U12062 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12086) );
  NAND2_X1 U12063 ( .A1(n14624), .A2(n12084), .ZN(n14625) );
  NAND2_X1 U12064 ( .A1(n15749), .A2(n11885), .ZN(n15984) );
  INV_X1 U12065 ( .A(n15863), .ZN(n11885) );
  NOR2_X2 U12066 ( .A1(n15984), .A2(n15983), .ZN(n15991) );
  AND2_X1 U12067 ( .A1(n11877), .A2(n11876), .ZN(n15797) );
  AND2_X1 U12069 ( .A1(n11861), .A2(n11860), .ZN(n15107) );
  AND2_X1 U12070 ( .A1(n11850), .A2(n11849), .ZN(n14961) );
  AND3_X1 U12071 ( .A1(n11806), .A2(n11805), .A3(n11804), .ZN(n16454) );
  NAND2_X1 U12072 ( .A1(n11505), .A2(n11504), .ZN(n11514) );
  INV_X1 U12073 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17685) );
  AND2_X1 U12074 ( .A1(n11712), .A2(n14287), .ZN(n16834) );
  INV_X1 U12075 ( .A(n14789), .ZN(n14790) );
  OR2_X1 U12076 ( .A1(n14759), .A2(n14760), .ZN(n14789) );
  AND2_X1 U12077 ( .A1(n14615), .A2(n11532), .ZN(n22478) );
  NAND2_X1 U12078 ( .A1(n22210), .A2(n14558), .ZN(n14966) );
  OR2_X1 U12079 ( .A1(n15902), .A2(n20599), .ZN(n14668) );
  NAND2_X1 U12080 ( .A1(n16807), .A2(n14630), .ZN(n15006) );
  AOI21_X1 U12081 ( .B1(n22454), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n14966), 
        .ZN(n14824) );
  INV_X1 U12082 ( .A(n14344), .ZN(n19194) );
  AND2_X1 U12083 ( .A1(n13281), .A2(n13280), .ZN(n19185) );
  AND2_X1 U12084 ( .A1(n14224), .A2(n14223), .ZN(n16198) );
  NAND2_X1 U12085 ( .A1(n16194), .A2(n16195), .ZN(n16192) );
  NAND2_X1 U12086 ( .A1(n14212), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14215) );
  NAND2_X1 U12087 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14198), .ZN(
        n14202) );
  INV_X1 U12088 ( .A(n13149), .ZN(n13151) );
  NAND2_X1 U12089 ( .A1(n13119), .A2(n13116), .ZN(n13149) );
  NAND2_X1 U12090 ( .A1(n12977), .A2(n12976), .ZN(n14432) );
  INV_X1 U12091 ( .A(n14429), .ZN(n12976) );
  INV_X1 U12092 ( .A(n14430), .ZN(n12977) );
  INV_X1 U12093 ( .A(n13983), .ZN(n16415) );
  NAND2_X1 U12094 ( .A1(n17097), .A2(n17096), .ZN(n17095) );
  OR2_X1 U12095 ( .A1(n17134), .A2(n17135), .ZN(n17132) );
  AND2_X1 U12096 ( .A1(n15658), .A2(n15703), .ZN(n15808) );
  NAND2_X1 U12097 ( .A1(n15808), .A2(n15807), .ZN(n17134) );
  AND2_X1 U12098 ( .A1(n17667), .A2(n22272), .ZN(n17883) );
  INV_X1 U12099 ( .A(n14531), .ZN(n19737) );
  NOR2_X2 U12100 ( .A1(n17271), .A2(n14210), .ZN(n14209) );
  NAND2_X1 U12101 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n14204), .ZN(
        n14207) );
  NAND2_X1 U12102 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n14201), .ZN(
        n14205) );
  NOR2_X1 U12103 ( .A1(n17784), .A2(n14199), .ZN(n14198) );
  NAND2_X1 U12104 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n14196), .ZN(
        n14199) );
  NOR2_X1 U12105 ( .A1(n18913), .A2(n14193), .ZN(n14192) );
  INV_X1 U12106 ( .A(n14189), .ZN(n14180) );
  NAND2_X1 U12107 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n14180), .ZN(
        n14193) );
  NOR2_X1 U12108 ( .A1(n17751), .A2(n14187), .ZN(n14190) );
  XNOR2_X1 U12109 ( .A(n12919), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17746) );
  NAND2_X1 U12111 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n14188), .ZN(
        n14187) );
  INV_X1 U12112 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15765) );
  NAND2_X1 U12113 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14184), .ZN(
        n14183) );
  NOR2_X1 U12114 ( .A1(n11288), .A2(n16386), .ZN(n16387) );
  NOR2_X2 U12115 ( .A1(n16885), .A2(n14263), .ZN(n16233) );
  CLKBUF_X1 U12116 ( .A(n17212), .Z(n17244) );
  CLKBUF_X1 U12117 ( .A(n17239), .Z(n17240) );
  OR2_X1 U12118 ( .A1(n16212), .A2(n16211), .ZN(n17259) );
  OR3_X1 U12119 ( .A1(n16946), .A2(n13093), .A3(n17398), .ZN(n17265) );
  NOR2_X1 U12120 ( .A1(n13183), .A2(n13515), .ZN(n17279) );
  INV_X1 U12121 ( .A(n15717), .ZN(n13020) );
  INV_X1 U12122 ( .A(n15704), .ZN(n13021) );
  NAND2_X1 U12123 ( .A1(n13185), .A2(n13514), .ZN(n17472) );
  NAND2_X1 U12124 ( .A1(n12998), .A2(n12997), .ZN(n14856) );
  CLKBUF_X1 U12125 ( .A(n17327), .Z(n17329) );
  NAND2_X1 U12126 ( .A1(n12919), .A2(n12915), .ZN(n17341) );
  XNOR2_X1 U12127 ( .A(n13756), .B(n13754), .ZN(n14384) );
  AND2_X1 U12128 ( .A1(n13276), .A2(n13275), .ZN(n19074) );
  OR2_X1 U12129 ( .A1(n13231), .A2(n13229), .ZN(n19197) );
  BUF_X1 U12130 ( .A(n12827), .Z(n19840) );
  NAND2_X1 U12132 ( .A1(n19814), .A2(n20282), .ZN(n19925) );
  INV_X2 U12133 ( .A(n13238), .ZN(n20081) );
  NAND3_X1 U12134 ( .A1(n19738), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19955), 
        .ZN(n19750) );
  NAND3_X1 U12135 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19737), .A3(n19955), 
        .ZN(n19752) );
  NAND2_X1 U12136 ( .A1(n19909), .A2(n19883), .ZN(n19776) );
  INV_X1 U12137 ( .A(n19750), .ZN(n20292) );
  INV_X1 U12138 ( .A(n19752), .ZN(n20293) );
  AND2_X1 U12139 ( .A1(n12947), .A2(n12946), .ZN(n13212) );
  NOR2_X1 U12140 ( .A1(n16121), .A2(n14131), .ZN(n21838) );
  AOI21_X1 U12141 ( .B1(n15535), .B2(n14142), .A(n15520), .ZN(n21839) );
  NOR2_X1 U12142 ( .A1(n21145), .A2(n21144), .ZN(n21152) );
  NOR2_X1 U12143 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20963), .ZN(n20969) );
  NOR2_X1 U12144 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20878), .ZN(n20893) );
  NOR2_X1 U12145 ( .A1(n21405), .A2(n20778), .ZN(n15562) );
  OAI211_X1 U12146 ( .C1(n16121), .C2(n20725), .A(n21839), .B(n21875), .ZN(
        n21193) );
  INV_X1 U12147 ( .A(n18801), .ZN(n18803) );
  AOI21_X1 U12148 ( .B1(n16117), .B2(n21874), .A(n16116), .ZN(n17655) );
  NOR2_X1 U12149 ( .A1(n19560), .A2(n18223), .ZN(n20725) );
  INV_X1 U12150 ( .A(n20724), .ZN(n20726) );
  NOR2_X1 U12151 ( .A1(n20724), .A2(n21874), .ZN(n20727) );
  NOR2_X2 U12152 ( .A1(n18568), .A2(n21150), .ZN(n18567) );
  INV_X1 U12153 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18577) );
  INV_X1 U12154 ( .A(n21629), .ZN(n21641) );
  NAND2_X1 U12155 ( .A1(n18510), .A2(n18511), .ZN(n18509) );
  NOR2_X1 U12156 ( .A1(n21542), .A2(n18393), .ZN(n18604) );
  XNOR2_X1 U12157 ( .A(n18356), .B(n18323), .ZN(n18668) );
  INV_X1 U12158 ( .A(n18324), .ZN(n18323) );
  NAND2_X1 U12159 ( .A1(n18287), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18288) );
  NAND2_X1 U12160 ( .A1(n18286), .A2(n18285), .ZN(n18289) );
  INV_X1 U12161 ( .A(n21764), .ZN(n21816) );
  AOI211_X1 U12162 ( .C1(n15522), .C2(n15521), .A(n15535), .B(n15520), .ZN(
        n21836) );
  NOR2_X1 U12163 ( .A1(n14053), .A2(n14052), .ZN(n19610) );
  NOR2_X1 U12164 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19279), .ZN(n19607) );
  INV_X1 U12165 ( .A(n14128), .ZN(n19519) );
  NOR2_X1 U12166 ( .A1(n14063), .A2(n14062), .ZN(n19476) );
  NOR2_X1 U12167 ( .A1(n14085), .A2(n14084), .ZN(n21252) );
  INV_X1 U12168 ( .A(n19607), .ZN(n19518) );
  INV_X1 U12169 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21846) );
  INV_X1 U12170 ( .A(n21897), .ZN(n21872) );
  CLKBUF_X1 U12171 ( .A(n14531), .Z(n19738) );
  NOR2_X1 U12172 ( .A1(n16450), .A2(n16297), .ZN(n22139) );
  INV_X1 U12173 ( .A(n22181), .ZN(n22197) );
  NAND2_X1 U12174 ( .A1(n22095), .A2(n14901), .ZN(n22186) );
  INV_X1 U12175 ( .A(n22188), .ZN(n22151) );
  NOR2_X1 U12176 ( .A1(n14916), .A2(n14899), .ZN(n16557) );
  INV_X1 U12177 ( .A(n20551), .ZN(n20544) );
  NAND2_X1 U12178 ( .A1(n16612), .A2(n13576), .ZN(n16614) );
  NOR2_X1 U12179 ( .A1(n15728), .A2(n14623), .ZN(n15903) );
  NAND2_X1 U12180 ( .A1(n14314), .A2(n14278), .ZN(n13564) );
  NOR2_X1 U12181 ( .A1(n20453), .A2(n21905), .ZN(n20469) );
  CLKBUF_X1 U12183 ( .A(n20469), .Z(n20471) );
  CLKBUF_X1 U12184 ( .A(n22385), .Z(n22363) );
  NAND2_X1 U12185 ( .A1(n22299), .A2(n14287), .ZN(n22381) );
  NAND2_X2 U12186 ( .A1(n14286), .A2(n14285), .ZN(n22387) );
  INV_X1 U12187 ( .A(n13583), .ZN(n13584) );
  INV_X1 U12188 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15647) );
  INV_X2 U12189 ( .A(n20599), .ZN(n20628) );
  OR2_X1 U12190 ( .A1(n20627), .A2(n14456), .ZN(n20633) );
  OR2_X1 U12191 ( .A1(n17723), .A2(n22465), .ZN(n20599) );
  NAND2_X1 U12192 ( .A1(n16126), .A2(n16125), .ZN(n16130) );
  NAND2_X1 U12193 ( .A1(n11919), .A2(n16454), .ZN(n15936) );
  INV_X1 U12194 ( .A(n15873), .ZN(n21979) );
  INV_X1 U12195 ( .A(n22033), .ZN(n22038) );
  NAND2_X1 U12196 ( .A1(n22476), .A2(n22211), .ZN(n22465) );
  CLKBUF_X1 U12197 ( .A(n14932), .Z(n14933) );
  OAI21_X1 U12198 ( .B1(n22462), .B2(n22461), .A(n22460), .ZN(n22690) );
  NOR2_X2 U12199 ( .A1(n14789), .A2(n15006), .ZN(n22703) );
  INV_X1 U12200 ( .A(n14954), .ZN(n22711) );
  OR2_X1 U12201 ( .A1(n14706), .A2(n14763), .ZN(n14954) );
  NOR2_X1 U12202 ( .A1(n14966), .A2(n22319), .ZN(n22602) );
  INV_X1 U12203 ( .A(n22644), .ZN(n22647) );
  INV_X1 U12204 ( .A(n22707), .ZN(n22717) );
  OR2_X1 U12205 ( .A1(n22207), .A2(n22210), .ZN(n22220) );
  NAND2_X1 U12206 ( .A1(n17727), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22207) );
  INV_X2 U12207 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22476) );
  INV_X1 U12208 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22210) );
  CLKBUF_X1 U12209 ( .A(n13265), .Z(n14274) );
  INV_X1 U12210 ( .A(n19059), .ZN(n19009) );
  INV_X1 U12211 ( .A(n19072), .ZN(n18916) );
  AND2_X1 U12212 ( .A1(n17731), .A2(n14262), .ZN(n19067) );
  INV_X2 U12213 ( .A(n14411), .ZN(n17054) );
  OR2_X1 U12214 ( .A1(n19193), .A2(n17665), .ZN(n17067) );
  INV_X1 U12215 ( .A(n19067), .ZN(n19011) );
  INV_X1 U12216 ( .A(n18996), .ZN(n19068) );
  INV_X1 U12217 ( .A(n19061), .ZN(n19028) );
  CLKBUF_X1 U12218 ( .A(n15657), .Z(n15658) );
  OR2_X1 U12219 ( .A1(n15128), .A2(n15655), .ZN(n19122) );
  OR2_X1 U12220 ( .A1(n13421), .A2(n13420), .ZN(n14927) );
  OR2_X1 U12221 ( .A1(n13360), .A2(n13359), .ZN(n14604) );
  INV_X1 U12222 ( .A(n14421), .ZN(n13763) );
  INV_X1 U12223 ( .A(n17128), .ZN(n17136) );
  INV_X1 U12224 ( .A(n17595), .ZN(n17621) );
  NOR2_X1 U12225 ( .A1(n16434), .A2(n16433), .ZN(n16436) );
  OR2_X1 U12226 ( .A1(n17153), .A2(n16920), .ZN(n19103) );
  INV_X1 U12227 ( .A(n20277), .ZN(n20172) );
  INV_X1 U12228 ( .A(n20067), .ZN(n20168) );
  NOR2_X1 U12229 ( .A1(n20279), .A2(n20277), .ZN(n20023) );
  AND2_X1 U12230 ( .A1(n20066), .A2(n13313), .ZN(n20277) );
  INV_X1 U12231 ( .A(n20066), .ZN(n20276) );
  INV_X1 U12232 ( .A(n20011), .ZN(n20285) );
  XOR2_X1 U12234 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n14178), .Z(
        n16409) );
  NAND2_X1 U12235 ( .A1(n16851), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14178) );
  NAND2_X1 U12236 ( .A1(n17793), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17792) );
  INV_X1 U12237 ( .A(n17475), .ZN(n17793) );
  INV_X1 U12238 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18913) );
  INV_X1 U12239 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17751) );
  NOR2_X1 U12240 ( .A1(n19250), .A2(n19096), .ZN(n17321) );
  INV_X1 U12241 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14373) );
  AOI21_X1 U12242 ( .B1(n16220), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16222) );
  CLKBUF_X1 U12243 ( .A(n17196), .Z(n17197) );
  CLKBUF_X1 U12244 ( .A(n17472), .Z(n17769) );
  INV_X1 U12245 ( .A(n17515), .ZN(n17516) );
  CLKBUF_X1 U12246 ( .A(n17343), .Z(n17344) );
  CLKBUF_X1 U12247 ( .A(n15763), .Z(n15764) );
  CLKBUF_X1 U12248 ( .A(n15667), .Z(n15668) );
  INV_X1 U12249 ( .A(n13741), .ZN(n17595) );
  AND2_X1 U12250 ( .A1(n13523), .A2(n13520), .ZN(n19159) );
  INV_X1 U12251 ( .A(n18865), .ZN(n14399) );
  NAND2_X1 U12252 ( .A1(n13523), .A2(n13297), .ZN(n19134) );
  INV_X1 U12253 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19856) );
  INV_X1 U12254 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19906) );
  NAND2_X1 U12255 ( .A1(n19909), .A2(n20015), .ZN(n19821) );
  INV_X1 U12256 ( .A(n19749), .ZN(n19814) );
  NAND2_X1 U12257 ( .A1(n14350), .A2(n14349), .ZN(n19775) );
  NOR2_X1 U12258 ( .A1(n19947), .A2(n19925), .ZN(n20262) );
  NAND2_X1 U12259 ( .A1(n19886), .A2(n19885), .ZN(n20368) );
  OAI21_X1 U12260 ( .B1(n19900), .B2(n19899), .A(n19898), .ZN(n20364) );
  INV_X1 U12261 ( .A(n20360), .ZN(n20362) );
  AND2_X1 U12262 ( .A1(n19849), .A2(n19848), .ZN(n19989) );
  NOR2_X1 U12263 ( .A1(n19872), .A2(n19904), .ZN(n20350) );
  INV_X1 U12264 ( .A(n20249), .ZN(n20336) );
  INV_X1 U12265 ( .A(n20334), .ZN(n20243) );
  INV_X1 U12266 ( .A(n20240), .ZN(n20324) );
  OAI21_X1 U12267 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(n20314) );
  INV_X1 U12268 ( .A(n20064), .ZN(n20056) );
  INV_X1 U12269 ( .A(n20261), .ZN(n20269) );
  INV_X1 U12270 ( .A(n20218), .ZN(n20209) );
  INV_X1 U12271 ( .A(n20109), .ZN(n20115) );
  INV_X1 U12272 ( .A(n20232), .ZN(n20298) );
  AND2_X1 U12273 ( .A1(n19213), .A2(n19212), .ZN(n19246) );
  INV_X1 U12274 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17661) );
  INV_X1 U12275 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19834) );
  NOR2_X1 U12276 ( .A1(n21838), .A2(n20724), .ZN(n17656) );
  INV_X1 U12277 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20715) );
  NOR2_X1 U12278 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n21029), .ZN(n21044) );
  NOR2_X1 U12279 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20984), .ZN(n21004) );
  NOR2_X1 U12280 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20934), .ZN(n20946) );
  NOR2_X2 U12281 ( .A1(n21885), .A2(n20879), .ZN(n21092) );
  INV_X1 U12282 ( .A(n21184), .ZN(n20879) );
  INV_X1 U12283 ( .A(n21168), .ZN(n21186) );
  AOI211_X1 U12284 ( .C1(n18051), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14072), .B(n14071), .ZN(n14073) );
  NOR2_X1 U12285 ( .A1(n21099), .A2(n18128), .ZN(n18132) );
  NOR4_X1 U12286 ( .A1(n19610), .A2(n19560), .A3(n21194), .A4(n21897), .ZN(
        n18217) );
  INV_X1 U12287 ( .A(n18217), .ZN(n18218) );
  NOR2_X1 U12288 ( .A1(n21315), .A2(n21309), .ZN(n21308) );
  INV_X1 U12289 ( .A(n21321), .ZN(n21316) );
  NOR2_X1 U12290 ( .A1(n21296), .A2(n21297), .ZN(n21322) );
  INV_X1 U12291 ( .A(n21327), .ZN(n21291) );
  NAND2_X1 U12292 ( .A1(n21291), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21296) );
  NOR3_X1 U12293 ( .A1(n21340), .A2(n21289), .A3(n21288), .ZN(n21334) );
  INV_X1 U12294 ( .A(n21332), .ZN(n21339) );
  NOR2_X1 U12295 ( .A1(n21352), .A2(n21351), .ZN(n21350) );
  AND2_X1 U12296 ( .A1(n21375), .A2(n21290), .ZN(n21359) );
  AND3_X1 U12297 ( .A1(n18282), .A2(n18281), .A3(n18280), .ZN(n21225) );
  NOR2_X1 U12298 ( .A1(n18261), .A2(n18260), .ZN(n21228) );
  NOR2_X1 U12299 ( .A1(n15596), .A2(n15595), .ZN(n21237) );
  NOR2_X1 U12300 ( .A1(n15555), .A2(n15554), .ZN(n21242) );
  NAND2_X1 U12301 ( .A1(n21378), .A2(n21375), .ZN(n21363) );
  INV_X1 U12302 ( .A(n21359), .ZN(n21353) );
  INV_X1 U12303 ( .A(n21375), .ZN(n21365) );
  INV_X1 U12304 ( .A(n21245), .ZN(n21373) );
  NOR2_X1 U12306 ( .A1(n21886), .A2(n18803), .ZN(n18812) );
  NOR2_X1 U12308 ( .A1(n20775), .A2(n20727), .ZN(n20765) );
  INV_X1 U12310 ( .A(n18660), .ZN(n18612) );
  CLKBUF_X1 U12311 ( .A(n18532), .Z(n21018) );
  NAND2_X1 U12312 ( .A1(n18509), .A2(n21708), .ZN(n18503) );
  OAI21_X1 U12313 ( .B1(n20782), .B2(n18579), .A(n19516), .ZN(n18534) );
  INV_X1 U12314 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18400) );
  NAND3_X1 U12315 ( .A1(n22233), .A2(n18745), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18580) );
  INV_X1 U12316 ( .A(n21524), .ZN(n21525) );
  INV_X1 U12317 ( .A(n18634), .ZN(n18661) );
  INV_X1 U12318 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20843) );
  INV_X1 U12319 ( .A(n18750), .ZN(n19516) );
  INV_X2 U12320 ( .A(n19516), .ZN(n19606) );
  INV_X1 U12321 ( .A(n18700), .ZN(n18734) );
  INV_X1 U12322 ( .A(n21793), .ZN(n21803) );
  INV_X1 U12323 ( .A(n21483), .ZN(n21841) );
  INV_X1 U12324 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21861) );
  INV_X1 U12325 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21865) );
  INV_X2 U12326 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21851) );
  INV_X1 U12327 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22288) );
  NAND2_X1 U12328 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22240), .ZN(n18839) );
  AND2_X1 U12329 ( .A1(n13575), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15902)
         );
  CLKBUF_X1 U12330 ( .A(n19275), .Z(n19603) );
  NOR2_X1 U12331 ( .A1(n11920), .A2(n11275), .ZN(n11921) );
  NAND2_X1 U12332 ( .A1(n17809), .A2(n17808), .ZN(n17810) );
  AOI21_X1 U12333 ( .B1(n17765), .B2(n17820), .A(n17764), .ZN(n17766) );
  OAI21_X1 U12334 ( .B1(n19124), .B2(n13196), .A(n17763), .ZN(n17764) );
  AND2_X1 U12335 ( .A1(n13205), .A2(n13204), .ZN(n13206) );
  AOI21_X1 U12336 ( .B1(n17522), .B2(n17818), .A(n13201), .ZN(n13205) );
  NAND2_X1 U12337 ( .A1(n16427), .A2(n16426), .ZN(n16428) );
  INV_X1 U12338 ( .A(n16425), .ZN(n16426) );
  AOI21_X1 U12339 ( .B1(n21659), .B2(n21658), .A(n21657), .ZN(n21660) );
  OR2_X1 U12340 ( .A1(n20640), .A2(n20693), .ZN(U212) );
  NAND2_X2 U12341 ( .A1(n11372), .A2(n11371), .ZN(n11422) );
  AND4_X2 U12342 ( .A1(n11289), .A2(n12913), .A3(n12912), .A4(n12911), .ZN(
        n13093) );
  CLKBUF_X2 U12343 ( .A(n11361), .Z(n12334) );
  NAND2_X2 U12344 ( .A1(n11672), .A2(n11590), .ZN(n11597) );
  AND3_X1 U12345 ( .A1(n12697), .A2(n12696), .A3(n12695), .ZN(n11234) );
  INV_X1 U12346 ( .A(n19941), .ZN(n12825) );
  OR2_X1 U12347 ( .A1(n11913), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11235) );
  AND2_X1 U12348 ( .A1(n13041), .A2(n11292), .ZN(n11236) );
  AND2_X1 U12349 ( .A1(n17054), .A2(n13741), .ZN(n11237) );
  AND2_X1 U12350 ( .A1(n17054), .A2(n17595), .ZN(n11239) );
  OR2_X1 U12351 ( .A1(n15929), .A2(n11689), .ZN(n11240) );
  OR2_X1 U12352 ( .A1(n18306), .A2(n21841), .ZN(n11241) );
  AND2_X1 U12353 ( .A1(n12656), .A2(n12642), .ZN(n11242) );
  NAND2_X1 U12354 ( .A1(n12553), .A2(n19189), .ZN(n13265) );
  NOR2_X2 U12355 ( .A1(n14856), .A2(n14855), .ZN(n14854) );
  NAND2_X1 U12356 ( .A1(n13051), .A2(n13050), .ZN(n13067) );
  XNOR2_X1 U12357 ( .A(n13090), .B(n13089), .ZN(n15762) );
  NAND2_X1 U12358 ( .A1(n15122), .A2(n15094), .ZN(n15093) );
  OR2_X1 U12359 ( .A1(n16391), .A2(n17006), .ZN(n11244) );
  OAI21_X1 U12360 ( .B1(n20227), .B2(n22264), .A(n14501), .ZN(n11245) );
  BUF_X1 U12361 ( .A(n13301), .Z(n20227) );
  INV_X1 U12362 ( .A(n11144), .ZN(n19007) );
  OAI22_X2 U12363 ( .A1(n14579), .A2(n14668), .B1(n20680), .B2(n14665), .ZN(
        n22568) );
  NAND2_X1 U12364 ( .A1(n15902), .A2(n20628), .ZN(n14665) );
  INV_X1 U12365 ( .A(n22510), .ZN(n11246) );
  INV_X1 U12366 ( .A(n11246), .ZN(n11247) );
  INV_X1 U12367 ( .A(n22535), .ZN(n11248) );
  INV_X1 U12368 ( .A(n11248), .ZN(n11249) );
  OAI21_X2 U12369 ( .B1(n14668), .B2(n16599), .A(n14609), .ZN(n22490) );
  NOR3_X2 U12370 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22437), .ZN(n22672) );
  INV_X1 U12371 ( .A(n17239), .ZN(n16197) );
  NAND2_X1 U12372 ( .A1(n16180), .A2(n16179), .ZN(n17415) );
  OAI21_X1 U12373 ( .B1(n16180), .B2(n17411), .A(n11252), .ZN(n11254) );
  OR2_X1 U12374 ( .A1(n16179), .A2(n17411), .ZN(n11253) );
  NAND2_X1 U12375 ( .A1(n11256), .A2(n17411), .ZN(n11255) );
  INV_X1 U12376 ( .A(n17415), .ZN(n11256) );
  OAI21_X2 U12377 ( .B1(n11257), .B2(n11259), .A(n12761), .ZN(n12771) );
  XNOR2_X2 U12378 ( .A(n12772), .B(n12771), .ZN(n14872) );
  NAND3_X1 U12379 ( .A1(n12690), .A2(n12689), .A3(n11258), .ZN(n11257) );
  NAND3_X1 U12380 ( .A1(n11242), .A2(n11261), .A3(n12640), .ZN(n11260) );
  NAND3_X1 U12381 ( .A1(n12641), .A2(n12655), .A3(n12658), .ZN(n11263) );
  NOR2_X1 U12382 ( .A1(n13729), .A2(n18865), .ZN(n11264) );
  NAND2_X1 U12383 ( .A1(n12529), .A2(n11176), .ZN(n12543) );
  INV_X1 U12384 ( .A(n12542), .ZN(n12534) );
  INV_X2 U12385 ( .A(n13713), .ZN(n13621) );
  INV_X1 U12386 ( .A(n14750), .ZN(n12998) );
  NOR2_X2 U12387 ( .A1(n16760), .A2(n16566), .ZN(n16527) );
  NAND2_X1 U12388 ( .A1(n18522), .A2(n18529), .ZN(n18521) );
  AOI21_X1 U12389 ( .B1(n12054), .B2(n12239), .A(n12053), .ZN(n15117) );
  INV_X2 U12390 ( .A(n11595), .ZN(n20593) );
  NOR2_X4 U12391 ( .A1(n17285), .A2(n17269), .ZN(n17422) );
  AND2_X1 U12392 ( .A1(n11835), .A2(n11834), .ZN(n14441) );
  CLKBUF_X1 U12393 ( .A(n14325), .Z(n16299) );
  AND2_X1 U12394 ( .A1(n12683), .A2(n12682), .ZN(n12691) );
  INV_X1 U12395 ( .A(n16468), .ZN(n16384) );
  NAND2_X1 U12396 ( .A1(n16468), .A2(n13591), .ZN(n13598) );
  NAND2_X1 U12397 ( .A1(n15086), .A2(n11686), .ZN(n15689) );
  AOI211_X2 U12398 ( .C1(n17814), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17352), .B(n17220), .ZN(n17221) );
  NAND2_X1 U12399 ( .A1(n12643), .A2(n12644), .ZN(n12654) );
  BUF_X1 U12400 ( .A(n14002), .Z(n11702) );
  AOI22_X1 U12401 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12428) );
  INV_X1 U12402 ( .A(n14442), .ZN(n11837) );
  AOI21_X1 U12403 ( .B1(n16693), .B2(n11693), .A(n20593), .ZN(n16684) );
  XNOR2_X1 U12404 ( .A(n13061), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14871) );
  AOI22_X1 U12405 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11402) );
  XNOR2_X1 U12406 ( .A(n13585), .B(n13584), .ZN(n16468) );
  NAND2_X2 U12407 ( .A1(n12434), .A2(n12433), .ZN(n12568) );
  AND2_X1 U12408 ( .A1(n12581), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11266) );
  INV_X1 U12409 ( .A(n12603), .ZN(n12985) );
  AND2_X1 U12410 ( .A1(n13915), .A2(n13918), .ZN(n11267) );
  OR2_X1 U12411 ( .A1(n17095), .A2(n13913), .ZN(n11268) );
  INV_X1 U12412 ( .A(n12605), .ZN(n12971) );
  INV_X2 U12413 ( .A(n13028), .ZN(n16236) );
  AND2_X1 U12414 ( .A1(n18501), .A2(n21627), .ZN(n11269) );
  OR2_X1 U12415 ( .A1(n21744), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11270) );
  AND2_X1 U12416 ( .A1(n13521), .A2(n11291), .ZN(n11271) );
  OR2_X1 U12417 ( .A1(n16424), .A2(n16423), .ZN(n11272) );
  INV_X1 U12418 ( .A(n17447), .ZN(n17448) );
  AND2_X2 U12419 ( .A1(n22203), .A2(n12412), .ZN(n20627) );
  NAND2_X1 U12420 ( .A1(n13564), .A2(n13563), .ZN(n15817) );
  NAND4_X1 U12421 ( .A1(n16264), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n16263), .ZN(n11273) );
  NOR2_X1 U12422 ( .A1(n13341), .A2(n15778), .ZN(n11274) );
  OAI21_X1 U12423 ( .B1(n13983), .B2(n18862), .A(n13309), .ZN(n14395) );
  AND2_X1 U12424 ( .A1(n16559), .A2(n22037), .ZN(n11275) );
  AND2_X1 U12425 ( .A1(n13917), .A2(n11267), .ZN(n11276) );
  NOR2_X2 U12426 ( .A1(n12409), .A2(n12410), .ZN(n13585) );
  CLKBUF_X3 U12427 ( .A(n16023), .Z(n14088) );
  INV_X1 U12428 ( .A(n15562), .ZN(n16022) );
  AND2_X1 U12429 ( .A1(n22045), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11277) );
  OR3_X1 U12430 ( .A1(n16261), .A2(n16260), .A3(n16263), .ZN(n11279) );
  NOR2_X1 U12431 ( .A1(n14338), .A2(n14339), .ZN(n11280) );
  INV_X1 U12432 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17411) );
  INV_X1 U12433 ( .A(n16010), .ZN(n14120) );
  AND2_X1 U12434 ( .A1(n16226), .A2(n13513), .ZN(n11281) );
  OR2_X1 U12435 ( .A1(n18399), .A2(n20803), .ZN(n11282) );
  INV_X1 U12436 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11626) );
  AND2_X1 U12438 ( .A1(n14347), .A2(n19834), .ZN(n11283) );
  OR2_X1 U12439 ( .A1(n16373), .A2(n13199), .ZN(n11284) );
  AND2_X1 U12440 ( .A1(n16213), .A2(n17259), .ZN(n11285) );
  AND2_X1 U12441 ( .A1(n17242), .A2(n17258), .ZN(n11286) );
  INV_X1 U12443 ( .A(n19230), .ZN(n19055) );
  INV_X2 U12444 ( .A(n18219), .ZN(n18214) );
  NAND2_X1 U12445 ( .A1(n18536), .A2(n18745), .ZN(n18579) );
  AND2_X1 U12446 ( .A1(n21803), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11287) );
  AND2_X1 U12447 ( .A1(n16862), .A2(n16355), .ZN(n11288) );
  OR2_X1 U12448 ( .A1(n16893), .A2(n13093), .ZN(n17215) );
  INV_X1 U12449 ( .A(n17215), .ZN(n16204) );
  NAND2_X2 U12450 ( .A1(n12663), .A2(n17630), .ZN(n13705) );
  INV_X1 U12451 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12226) );
  AND4_X1 U12452 ( .A1(n12899), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n11289) );
  INV_X1 U12453 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16358) );
  INV_X1 U12454 ( .A(n13271), .ZN(n12549) );
  AND2_X1 U12455 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11290) );
  OR2_X1 U12456 ( .A1(n22288), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18842) );
  INV_X1 U12457 ( .A(n19121), .ZN(n17765) );
  INV_X1 U12458 ( .A(n19560), .ZN(n20710) );
  OR2_X1 U12459 ( .A1(n13458), .A2(n13457), .ZN(n15130) );
  NAND2_X1 U12460 ( .A1(n19159), .A2(n17103), .ZN(n11291) );
  AND2_X1 U12461 ( .A1(n13523), .A2(n13522), .ZN(n19157) );
  NOR2_X1 U12462 ( .A1(n13040), .A2(n13039), .ZN(n11292) );
  AND2_X1 U12463 ( .A1(n17789), .A2(n12959), .ZN(n17807) );
  AND2_X1 U12464 ( .A1(n18532), .A2(n11282), .ZN(n11293) );
  NAND2_X1 U12465 ( .A1(n14383), .A2(n14384), .ZN(n14382) );
  NAND2_X1 U12466 ( .A1(n13261), .A2(n17818), .ZN(n11294) );
  INV_X1 U12467 ( .A(n17321), .ZN(n17779) );
  INV_X1 U12468 ( .A(n17779), .ZN(n17820) );
  INV_X2 U12469 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21848) );
  AND2_X1 U12470 ( .A1(n16238), .A2(n16879), .ZN(n11295) );
  NAND2_X1 U12471 ( .A1(n19160), .A2(n13261), .ZN(n11296) );
  AND4_X1 U12472 ( .A1(n11369), .A2(n11368), .A3(n11367), .A4(n11366), .ZN(
        n11297) );
  NAND2_X2 U12473 ( .A1(n13590), .A2(n13589), .ZN(n20556) );
  INV_X1 U12474 ( .A(n16572), .ZN(n13591) );
  AND2_X1 U12475 ( .A1(n11415), .A2(n14621), .ZN(n11298) );
  AND4_X1 U12476 ( .A1(n11408), .A2(n11407), .A3(n12076), .A4(n14621), .ZN(
        n11299) );
  NOR2_X1 U12477 ( .A1(n19892), .A2(n12687), .ZN(n12688) );
  OR2_X1 U12478 ( .A1(n11735), .A2(n11737), .ZN(n11720) );
  NAND2_X1 U12479 ( .A1(n13266), .A2(n13271), .ZN(n12581) );
  AOI21_X1 U12480 ( .B1(n19783), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n12688), .ZN(n12689) );
  OR2_X1 U12481 ( .A1(n11558), .A2(n11557), .ZN(n11651) );
  OR2_X1 U12482 ( .A1(n11571), .A2(n11570), .ZN(n11662) );
  AOI22_X1 U12483 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12462) );
  AND2_X1 U12484 ( .A1(n11755), .A2(n11723), .ZN(n11758) );
  OR2_X1 U12485 ( .A1(n11527), .A2(n11526), .ZN(n11631) );
  OAI211_X1 U12486 ( .C1(n12605), .C2(n14369), .A(n12597), .B(n12596), .ZN(
        n12598) );
  INV_X1 U12487 ( .A(n17318), .ZN(n13133) );
  INV_X1 U12488 ( .A(n12889), .ZN(n12880) );
  AOI22_X1 U12489 ( .A1(n13953), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U12490 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U12491 ( .A1(n11561), .A2(n11640), .ZN(n11650) );
  INV_X1 U12492 ( .A(n15856), .ZN(n12160) );
  INV_X1 U12493 ( .A(n11659), .ZN(n11586) );
  AOI22_X1 U12494 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11363) );
  OR2_X1 U12495 ( .A1(n11412), .A2(n11411), .ZN(n11413) );
  OR2_X1 U12496 ( .A1(n12679), .A2(n12678), .ZN(n13327) );
  XNOR2_X1 U12497 ( .A(n12519), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12935) );
  AOI22_X1 U12498 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12673), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12430) );
  CLKBUF_X1 U12499 ( .A(n13945), .Z(n13647) );
  AND2_X1 U12500 ( .A1(n13955), .A2(n12519), .ZN(n12711) );
  NAND2_X1 U12501 ( .A1(n13616), .A2(n12660), .ZN(n13874) );
  OR2_X1 U12502 ( .A1(n12789), .A2(n12788), .ZN(n13330) );
  AND4_X1 U12503 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n12913) );
  INV_X1 U12504 ( .A(n12572), .ZN(n17629) );
  NAND2_X1 U12505 ( .A1(n12502), .A2(n12519), .ZN(n12510) );
  INV_X1 U12506 ( .A(n11913), .ZN(n11899) );
  AND2_X1 U12507 ( .A1(n16141), .A2(n13548), .ZN(n13549) );
  AND2_X1 U12508 ( .A1(n22196), .A2(n13548), .ZN(n12369) );
  INV_X1 U12509 ( .A(n14627), .ZN(n12084) );
  AND2_X1 U12510 ( .A1(n11698), .A2(n11595), .ZN(n11699) );
  NAND2_X1 U12511 ( .A1(n11174), .A2(n11854), .ZN(n11910) );
  INV_X1 U12512 ( .A(n14441), .ZN(n11836) );
  NOR2_X1 U12513 ( .A1(n12931), .A2(n12935), .ZN(n12932) );
  AND2_X1 U12514 ( .A1(n13621), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13445) );
  INV_X1 U12515 ( .A(n12605), .ZN(n13028) );
  NAND2_X1 U12518 ( .A1(n12497), .A2(n12496), .ZN(n12511) );
  AND2_X1 U12519 ( .A1(n15706), .A2(n15652), .ZN(n13015) );
  INV_X1 U12520 ( .A(n16399), .ZN(n16363) );
  INV_X1 U12521 ( .A(n14751), .ZN(n12997) );
  NAND2_X1 U12522 ( .A1(n12895), .A2(n12894), .ZN(n12914) );
  AND2_X1 U12523 ( .A1(n18865), .A2(n12624), .ZN(n12638) );
  NAND2_X1 U12524 ( .A1(n12526), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12527) );
  AOI22_X1 U12525 ( .A1(n18335), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21780), .B2(n18511), .ZN(n18336) );
  INV_X1 U12526 ( .A(n18319), .ZN(n18317) );
  NAND2_X1 U12527 ( .A1(n15615), .A2(n15581), .ZN(n15618) );
  NAND2_X1 U12528 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  INV_X1 U12529 ( .A(n15843), .ZN(n11874) );
  INV_X1 U12530 ( .A(n14990), .ZN(n11846) );
  INV_X1 U12531 ( .A(n13545), .ZN(n12397) );
  NOR2_X1 U12532 ( .A1(n14015), .A2(n16469), .ZN(n14016) );
  NAND2_X1 U12533 ( .A1(n16568), .A2(n16569), .ZN(n16531) );
  AND2_X1 U12534 ( .A1(n12296), .A2(n12295), .ZN(n15963) );
  AND2_X1 U12535 ( .A1(n22476), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13552) );
  INV_X1 U12536 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U12537 ( .A1(n11597), .A2(n21993), .ZN(n15974) );
  CLKBUF_X1 U12538 ( .A(n20565), .Z(n20566) );
  NAND2_X1 U12539 ( .A1(n11837), .A2(n11836), .ZN(n14440) );
  INV_X1 U12540 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22408) );
  AND2_X1 U12541 ( .A1(n13300), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18855) );
  INV_X1 U12542 ( .A(n16190), .ZN(n14222) );
  OR2_X1 U12543 ( .A1(n12742), .A2(n12741), .ZN(n13315) );
  INV_X1 U12544 ( .A(n12985), .ZN(n16404) );
  INV_X1 U12545 ( .A(n13906), .ZN(n13904) );
  OAI211_X1 U12546 ( .C1(n17789), .C2(n16371), .A(n16374), .B(n11284), .ZN(
        n16375) );
  OR2_X1 U12547 ( .A1(n18911), .A2(n13093), .ZN(n13140) );
  OR2_X1 U12548 ( .A1(n16365), .A2(n16372), .ZN(n16366) );
  NAND2_X1 U12549 ( .A1(n12923), .A2(n11281), .ZN(n16218) );
  AND2_X1 U12550 ( .A1(n13183), .A2(n13515), .ZN(n13184) );
  INV_X1 U12551 ( .A(n12918), .ZN(n17747) );
  OR2_X1 U12552 ( .A1(n12914), .A2(n13093), .ZN(n12919) );
  AND2_X1 U12553 ( .A1(n13523), .A2(n19185), .ZN(n17447) );
  XNOR2_X1 U12554 ( .A(n13746), .B(n13747), .ZN(n14378) );
  NAND2_X1 U12555 ( .A1(n12643), .A2(n12623), .ZN(n12814) );
  AND2_X1 U12556 ( .A1(n14139), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14141) );
  AOI21_X1 U12557 ( .B1(n21855), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14132), .ZN(n14138) );
  NOR2_X1 U12558 ( .A1(n18498), .A2(n18497), .ZN(n18499) );
  NOR2_X1 U12559 ( .A1(n21389), .A2(n21387), .ZN(n15609) );
  INV_X1 U12560 ( .A(n18336), .ZN(n18337) );
  NAND2_X1 U12561 ( .A1(n21521), .A2(n18380), .ZN(n21542) );
  NAND2_X1 U12562 ( .A1(n18691), .A2(n18320), .ZN(n18679) );
  NOR2_X1 U12563 ( .A1(n21252), .A2(n21253), .ZN(n15536) );
  NOR2_X1 U12564 ( .A1(n12348), .A2(n16551), .ZN(n12357) );
  INV_X1 U12565 ( .A(n12311), .ZN(n11923) );
  AND2_X1 U12566 ( .A1(n12195), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12179) );
  INV_X1 U12567 ( .A(n11143), .ZN(n22191) );
  NAND2_X1 U12568 ( .A1(n14905), .A2(n14904), .ZN(n22138) );
  INV_X1 U12569 ( .A(n15101), .ZN(n15102) );
  CLKBUF_X1 U12570 ( .A(n13562), .Z(n14299) );
  NAND2_X1 U12571 ( .A1(n12372), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12382) );
  NOR2_X1 U12572 ( .A1(n12162), .A2(n15753), .ZN(n12263) );
  NAND2_X1 U12573 ( .A1(n12242), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12225) );
  INV_X1 U12574 ( .A(n12146), .ZN(n12242) );
  NOR2_X1 U12575 ( .A1(n12050), .A2(n15647), .ZN(n12021) );
  AND2_X1 U12576 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12087), .ZN(
        n12096) );
  AND2_X1 U12577 ( .A1(n14006), .A2(n14008), .ZN(n14007) );
  AND2_X1 U12578 ( .A1(n16749), .A2(n11821), .ZN(n16764) );
  INV_X1 U12579 ( .A(n21999), .ZN(n21987) );
  AND2_X1 U12580 ( .A1(n11808), .A2(n14329), .ZN(n15873) );
  NOR2_X1 U12581 ( .A1(n16807), .A2(n12075), .ZN(n14827) );
  AND2_X1 U12582 ( .A1(n14759), .A2(n14821), .ZN(n22404) );
  INV_X1 U12583 ( .A(n22404), .ZN(n22419) );
  INV_X1 U12584 ( .A(n22560), .ZN(n14984) );
  INV_X1 U12585 ( .A(n14827), .ZN(n14763) );
  INV_X1 U12586 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22454) );
  INV_X1 U12587 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17709) );
  NAND3_X1 U12588 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22210), .A3(n14558), 
        .ZN(n14670) );
  AND2_X1 U12589 ( .A1(n13228), .A2(n17882), .ZN(n13229) );
  AND2_X1 U12590 ( .A1(n16919), .A2(n16918), .ZN(n17153) );
  OR2_X1 U12591 ( .A1(n17731), .A2(n14234), .ZN(n19059) );
  XNOR2_X1 U12593 ( .A(n16406), .B(n16405), .ZN(n16422) );
  AND3_X1 U12594 ( .A1(n13402), .A2(n13401), .A3(n13400), .ZN(n13766) );
  NAND2_X1 U12595 ( .A1(n13904), .A2(n20227), .ZN(n13905) );
  NAND2_X1 U12596 ( .A1(n17186), .A2(n17187), .ZN(n17188) );
  NAND2_X1 U12597 ( .A1(n20066), .A2(n13985), .ZN(n20067) );
  NAND2_X1 U12598 ( .A1(n17806), .A2(n17818), .ZN(n17809) );
  INV_X1 U12599 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17027) );
  NOR2_X1 U12600 ( .A1(n17798), .A2(n16172), .ZN(n17293) );
  AND2_X1 U12601 ( .A1(n17305), .A2(n13158), .ZN(n17786) );
  AND2_X1 U12602 ( .A1(n13138), .A2(n17511), .ZN(n17493) );
  AND2_X1 U12603 ( .A1(n16225), .A2(n16224), .ZN(n17571) );
  XNOR2_X1 U12604 ( .A(n12879), .B(n12877), .ZN(n12887) );
  OR2_X1 U12605 ( .A1(n14378), .A2(n14377), .ZN(n14379) );
  OR2_X1 U12606 ( .A1(n19909), .A2(n19883), .ZN(n19947) );
  OR2_X1 U12607 ( .A1(n19909), .A2(n20015), .ZN(n19872) );
  BUF_X1 U12608 ( .A(n12814), .Z(n19824) );
  OAI21_X2 U12609 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19236), .A(n19744), 
        .ZN(n19959) );
  NOR2_X2 U12610 ( .A1(n20713), .A2(n16011), .ZN(n21835) );
  NAND2_X1 U12611 ( .A1(n16117), .A2(n18223), .ZN(n14131) );
  NAND2_X1 U12612 ( .A1(n18567), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18552) );
  NOR2_X1 U12613 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n21019), .ZN(n21030) );
  INV_X1 U12614 ( .A(n21049), .ZN(n21052) );
  NOR2_X1 U12615 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20905), .ZN(n20926) );
  NOR2_X1 U12616 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20848), .ZN(n20868) );
  INV_X1 U12617 ( .A(n14144), .ZN(n14146) );
  INV_X1 U12618 ( .A(n19358), .ZN(n21253) );
  NOR2_X1 U12619 ( .A1(n18307), .A2(n16011), .ZN(n16119) );
  NOR2_X1 U12620 ( .A1(n21714), .A2(n18525), .ZN(n18494) );
  INV_X1 U12621 ( .A(n14163), .ZN(n18458) );
  INV_X1 U12622 ( .A(n18534), .ZN(n18486) );
  CLKBUF_X1 U12623 ( .A(n18326), .Z(n18576) );
  INV_X1 U12624 ( .A(n18596), .ZN(n20975) );
  INV_X1 U12625 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18654) );
  OAI21_X2 U12626 ( .B1(n20717), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21900), 
        .ZN(n18745) );
  NAND2_X1 U12627 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18604), .ZN(
        n21575) );
  INV_X1 U12628 ( .A(n21835), .ZN(n21756) );
  NAND2_X1 U12629 ( .A1(n18295), .A2(n18294), .ZN(n18297) );
  NOR2_X1 U12630 ( .A1(n15612), .A2(n16121), .ZN(n21822) );
  INV_X1 U12631 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21855) );
  AOI211_X1 U12632 ( .C1(n18262), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n14094), .B(n14093), .ZN(n14095) );
  OAI211_X1 U12633 ( .C1(n11192), .C2(n14280), .A(n16331), .B(n16451), .ZN(
        n21903) );
  NAND2_X1 U12634 ( .A1(n12357), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U12635 ( .A1(n12329), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12348) );
  INV_X1 U12636 ( .A(n22186), .ZN(n22195) );
  NOR2_X1 U12637 ( .A1(n16614), .A2(n15149), .ZN(n13580) );
  INV_X1 U12638 ( .A(n15817), .ZN(n15728) );
  INV_X1 U12639 ( .A(n22299), .ZN(n22385) );
  AND2_X1 U12640 ( .A1(n16001), .A2(n16003), .ZN(n22171) );
  AND2_X1 U12641 ( .A1(n15859), .A2(n15858), .ZN(n15893) );
  INV_X1 U12642 ( .A(n20633), .ZN(n20623) );
  INV_X1 U12643 ( .A(n22203), .ZN(n20629) );
  INV_X1 U12644 ( .A(n11825), .ZN(n11920) );
  OR2_X1 U12645 ( .A1(n21986), .A2(n15841), .ZN(n21999) );
  OR2_X1 U12646 ( .A1(n15867), .A2(n15877), .ZN(n20591) );
  INV_X1 U12647 ( .A(n15936), .ZN(n21985) );
  CLKBUF_X1 U12648 ( .A(n14435), .Z(n14439) );
  INV_X1 U12649 ( .A(n22017), .ZN(n22037) );
  NAND2_X1 U12650 ( .A1(n16461), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16845) );
  NOR2_X2 U12651 ( .A1(n22419), .A2(n14828), .ZN(n22654) );
  AND2_X1 U12652 ( .A1(n22404), .A2(n14827), .ZN(n22660) );
  AND2_X1 U12653 ( .A1(n22404), .A2(n22403), .ZN(n22666) );
  NOR2_X2 U12654 ( .A1(n22419), .A2(n15006), .ZN(n22667) );
  AND2_X1 U12655 ( .A1(n14760), .A2(n14629), .ZN(n14683) );
  INV_X1 U12656 ( .A(n22431), .ZN(n22673) );
  AND2_X1 U12657 ( .A1(n14683), .A2(n22403), .ZN(n22674) );
  AND2_X1 U12658 ( .A1(n14683), .A2(n14682), .ZN(n22560) );
  INV_X1 U12659 ( .A(n22684), .ZN(n14986) );
  INV_X1 U12660 ( .A(n14828), .ZN(n14764) );
  NOR2_X2 U12661 ( .A1(n14789), .A2(n14763), .ZN(n22689) );
  INV_X1 U12662 ( .A(n22699), .ZN(n22616) );
  AND2_X1 U12663 ( .A1(n16807), .A2(n12075), .ZN(n22403) );
  INV_X1 U12664 ( .A(n22715), .ZN(n22701) );
  OR2_X1 U12665 ( .A1(n16807), .A2(n14630), .ZN(n14828) );
  INV_X1 U12666 ( .A(n22725), .ZN(n14956) );
  INV_X1 U12667 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22251) );
  INV_X1 U12668 ( .A(n20497), .ZN(n20509) );
  INV_X1 U12669 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n22263) );
  XNOR2_X1 U12670 ( .A(n16412), .B(n13984), .ZN(n16870) );
  NAND2_X1 U12671 ( .A1(n16233), .A2(n16232), .ZN(n16412) );
  NAND2_X1 U12672 ( .A1(n16198), .A2(n16199), .ZN(n16203) );
  NAND2_X1 U12673 ( .A1(n16182), .A2(n16183), .ZN(n16190) );
  INV_X1 U12674 ( .A(n18926), .ZN(n18932) );
  OR2_X1 U12675 ( .A1(n13440), .A2(n13439), .ZN(n14921) );
  OR2_X1 U12676 ( .A1(n13381), .A2(n13380), .ZN(n14748) );
  CLKBUF_X1 U12677 ( .A(n14421), .Z(n14497) );
  AND2_X1 U12678 ( .A1(n16885), .A2(n16884), .ZN(n17366) );
  INV_X1 U12679 ( .A(n19247), .ZN(n18852) );
  INV_X1 U12680 ( .A(n20222), .ZN(n20279) );
  INV_X1 U12681 ( .A(n17664), .ZN(n14550) );
  INV_X1 U12682 ( .A(n17664), .ZN(n14574) );
  NAND2_X1 U12683 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n14209), .ZN(
        n14213) );
  INV_X1 U12684 ( .A(n13203), .ZN(n13204) );
  NAND2_X1 U12685 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n14186), .ZN(
        n14185) );
  AND2_X2 U12686 ( .A1(n12634), .A2(n12620), .ZN(n18865) );
  XNOR2_X1 U12687 ( .A(n17422), .B(n17411), .ZN(n17811) );
  NAND2_X1 U12688 ( .A1(n19153), .A2(n17448), .ZN(n17454) );
  AND2_X1 U12689 ( .A1(n15125), .A2(n13198), .ZN(n17520) );
  AND2_X1 U12690 ( .A1(n13523), .A2(n13278), .ZN(n17451) );
  AND2_X1 U12691 ( .A1(n13523), .A2(n13260), .ZN(n19160) );
  XNOR2_X1 U12692 ( .A(n14463), .B(n14462), .ZN(n19909) );
  NAND2_X1 U12693 ( .A1(n19197), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19236) );
  NOR2_X1 U12694 ( .A1(n19947), .A2(n19904), .ZN(n20378) );
  INV_X1 U12695 ( .A(n20368), .ZN(n20370) );
  OR2_X1 U12696 ( .A1(n19900), .A2(n19896), .ZN(n19894) );
  OAI21_X1 U12697 ( .B1(n19866), .B2(n19865), .A(n19864), .ZN(n20349) );
  INV_X1 U12698 ( .A(n19989), .ZN(n20343) );
  NOR2_X1 U12699 ( .A1(n19872), .A2(n19884), .ZN(n20246) );
  INV_X1 U12700 ( .A(n19984), .ZN(n20331) );
  OAI21_X1 U12701 ( .B1(n19811), .B2(n19810), .A(n19809), .ZN(n20325) );
  NOR2_X1 U12702 ( .A1(n19776), .A2(n19946), .ZN(n20313) );
  INV_X1 U12703 ( .A(n20389), .ZN(n20393) );
  INV_X1 U12704 ( .A(n20303), .ZN(n20306) );
  INV_X1 U12705 ( .A(n20166), .ZN(n20155) );
  INV_X1 U12706 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19835) );
  AND2_X1 U12707 ( .A1(n19221), .A2(n19220), .ZN(n19234) );
  NAND2_X1 U12708 ( .A1(n21872), .A2(n21839), .ZN(n20724) );
  INV_X1 U12709 ( .A(n17656), .ZN(n20720) );
  OR2_X1 U12710 ( .A1(n21152), .A2(n21151), .ZN(n21164) );
  NOR2_X1 U12711 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n21057), .ZN(n21077) );
  INV_X1 U12712 ( .A(n21185), .ZN(n21160) );
  NOR2_X1 U12713 ( .A1(n20962), .A2(n20961), .ZN(n21049) );
  NOR3_X1 U12714 ( .A1(n21081), .A2(n21535), .A3(n20920), .ZN(n21067) );
  NOR2_X1 U12715 ( .A1(n21873), .A2(n14146), .ZN(n21103) );
  NOR2_X1 U12716 ( .A1(n20720), .A2(n19610), .ZN(n14144) );
  NAND4_X1 U12717 ( .A1(n21808), .A2(n20720), .A3(n21882), .A4(n21894), .ZN(
        n21184) );
  NOR2_X2 U12718 ( .A1(n14107), .A2(n14106), .ZN(n19560) );
  NAND2_X1 U12719 ( .A1(n21316), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n21315) );
  NOR2_X1 U12720 ( .A1(n21290), .A2(n21333), .ZN(n21328) );
  NAND2_X1 U12721 ( .A1(n21350), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21340) );
  NAND4_X1 U12722 ( .A1(n21358), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n21250), .ZN(n21352) );
  NOR2_X1 U12723 ( .A1(n21365), .A2(n21247), .ZN(n21358) );
  INV_X1 U12724 ( .A(n21363), .ZN(n21372) );
  INV_X1 U12725 ( .A(n19610), .ZN(n18802) );
  NOR2_X1 U12726 ( .A1(n21650), .A2(n21641), .ZN(n21649) );
  NAND2_X1 U12727 ( .A1(n18494), .A2(n21627), .ZN(n21612) );
  INV_X1 U12728 ( .A(n18580), .ZN(n18570) );
  NOR2_X2 U12729 ( .A1(n20710), .A2(n21900), .ZN(n18700) );
  XNOR2_X1 U12730 ( .A(n15583), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18722) );
  NOR2_X1 U12731 ( .A1(n19560), .A2(n21900), .ZN(n18704) );
  AND2_X1 U12732 ( .A1(n21656), .A2(n21828), .ZN(n21657) );
  NAND2_X1 U12733 ( .A1(n18466), .A2(n18465), .ZN(n18474) );
  OAI21_X1 U12734 ( .B1(n18304), .B2(n18303), .A(n18302), .ZN(n18648) );
  NOR2_X1 U12735 ( .A1(n19560), .A2(n21727), .ZN(n21483) );
  NOR2_X2 U12736 ( .A1(n20710), .A2(n21727), .ZN(n21834) );
  NOR2_X1 U12737 ( .A1(n19518), .A2(n19333), .ZN(n18750) );
  INV_X1 U12738 ( .A(n21421), .ZN(n21887) );
  OAI21_X1 U12739 ( .B1(n21695), .B2(n18307), .A(n11241), .ZN(n21871) );
  OR2_X1 U12740 ( .A1(n20710), .A2(n18223), .ZN(n21874) );
  NAND2_X1 U12741 ( .A1(n16463), .A2(n14286), .ZN(n16451) );
  INV_X1 U12742 ( .A(n22139), .ZN(n22122) );
  NAND2_X1 U12743 ( .A1(n22095), .A2(n14897), .ZN(n22181) );
  INV_X1 U12744 ( .A(n16557), .ZN(n22202) );
  INV_X1 U12745 ( .A(n13596), .ZN(n13597) );
  NOR2_X1 U12746 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  INV_X1 U12747 ( .A(n15728), .ZN(n16612) );
  INV_X1 U12748 ( .A(n15903), .ZN(n15819) );
  INV_X1 U12749 ( .A(n20453), .ZN(n20473) );
  AOI21_X1 U12750 ( .B1(n21907), .B2(n22242), .A(n16451), .ZN(n22299) );
  OAI21_X1 U12751 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15982) );
  NAND2_X1 U12752 ( .A1(n11919), .A2(n11918), .ZN(n22017) );
  INV_X1 U12753 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17707) );
  INV_X1 U12754 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U12755 ( .A1(n22391), .A2(n22397), .B1(n22390), .B2(n22450), .ZN(
        n22658) );
  AOI22_X1 U12756 ( .A1(n22407), .A2(n22412), .B1(n22434), .B2(n22450), .ZN(
        n22664) );
  INV_X1 U12757 ( .A(n22422), .ZN(n22671) );
  AOI21_X1 U12758 ( .B1(n15012), .B2(n15011), .A(n22480), .ZN(n15053) );
  NAND2_X1 U12759 ( .A1(n14683), .A2(n14764), .ZN(n15049) );
  AOI22_X1 U12760 ( .A1(n22436), .A2(n22441), .B1(n22435), .B2(n22434), .ZN(
        n22678) );
  AOI21_X1 U12761 ( .B1(n16813), .B2(n14686), .A(n22424), .ZN(n14746) );
  NAND2_X1 U12762 ( .A1(n14790), .A2(n14764), .ZN(n22684) );
  AOI22_X1 U12763 ( .A1(n22452), .A2(n22461), .B1(n22451), .B2(n22450), .ZN(
        n22693) );
  NAND2_X1 U12764 ( .A1(n14790), .A2(n22403), .ZN(n22699) );
  INV_X1 U12765 ( .A(n22488), .ZN(n22487) );
  AOI22_X1 U12766 ( .A1(n22473), .A2(n22483), .B1(n22472), .B2(n22477), .ZN(
        n22708) );
  OR2_X1 U12767 ( .A1(n14828), .A2(n14706), .ZN(n22715) );
  OR2_X1 U12768 ( .A1(n14706), .A2(n14555), .ZN(n22725) );
  INV_X1 U12769 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17727) );
  INV_X1 U12770 ( .A(n22226), .ZN(n17683) );
  OR2_X1 U12771 ( .A1(n19193), .A2(n14229), .ZN(n14502) );
  INV_X1 U12772 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19237) );
  OR2_X1 U12773 ( .A1(n19205), .A2(n19247), .ZN(n19250) );
  NAND2_X1 U12774 ( .A1(n14574), .A2(n19218), .ZN(n19072) );
  OR2_X1 U12775 ( .A1(n15705), .A2(n15656), .ZN(n18948) );
  AND2_X1 U12776 ( .A1(n14346), .A2(n18852), .ZN(n17125) );
  NAND2_X1 U12777 ( .A1(n14382), .A2(n14385), .ZN(n20015) );
  AND2_X1 U12778 ( .A1(n13999), .A2(n13998), .ZN(n14000) );
  AND2_X2 U12779 ( .A1(n13968), .A2(n18852), .ZN(n20066) );
  NAND2_X1 U12780 ( .A1(n20066), .A2(n13243), .ZN(n20222) );
  INV_X1 U12781 ( .A(n17883), .ZN(n17881) );
  OR2_X1 U12782 ( .A1(n14502), .A2(n19096), .ZN(n17664) );
  AOI21_X1 U12783 ( .B1(n16429), .B2(n17321), .A(n16410), .ZN(n16411) );
  AOI21_X1 U12784 ( .B1(n17811), .B2(n17820), .A(n17810), .ZN(n17812) );
  NAND2_X1 U12785 ( .A1(n19250), .A2(n12958), .ZN(n17789) );
  INV_X1 U12786 ( .A(n17777), .ZN(n17827) );
  NAND2_X1 U12787 ( .A1(n13524), .A2(n19157), .ZN(n13525) );
  AOI21_X1 U12788 ( .B1(n17792), .B2(n17454), .A(n17486), .ZN(n19139) );
  INV_X1 U12789 ( .A(n19157), .ZN(n19153) );
  INV_X1 U12790 ( .A(n19160), .ZN(n19123) );
  INV_X1 U12791 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19910) );
  INV_X1 U12792 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19101) );
  INV_X1 U12793 ( .A(n20392), .ZN(n20273) );
  INV_X1 U12794 ( .A(n20262), .ZN(n20388) );
  INV_X1 U12795 ( .A(n20378), .ZN(n20375) );
  AND2_X1 U12796 ( .A1(n19894), .A2(n19893), .ZN(n20363) );
  NAND2_X1 U12797 ( .A1(n19870), .A2(n19869), .ZN(n20360) );
  INV_X1 U12798 ( .A(n20355), .ZN(n20353) );
  INV_X1 U12799 ( .A(n20350), .ZN(n20200) );
  INV_X1 U12800 ( .A(n20246), .ZN(n20346) );
  OR2_X1 U12801 ( .A1(n19821), .A2(n19946), .ZN(n20249) );
  AND2_X1 U12802 ( .A1(n19820), .A2(n19819), .ZN(n19984) );
  OR2_X1 U12803 ( .A1(n19821), .A2(n19925), .ZN(n20334) );
  OR2_X1 U12804 ( .A1(n19821), .A2(n19904), .ZN(n20240) );
  INV_X1 U12805 ( .A(n20313), .ZN(n20310) );
  OR2_X1 U12806 ( .A1(n19776), .A2(n19925), .ZN(n20303) );
  OR2_X1 U12807 ( .A1(n19776), .A2(n19904), .ZN(n20232) );
  OR2_X1 U12808 ( .A1(n19776), .A2(n19884), .ZN(n20399) );
  INV_X1 U12809 ( .A(n19234), .ZN(n19233) );
  INV_X1 U12810 ( .A(n22231), .ZN(n17660) );
  INV_X1 U12811 ( .A(n21092), .ZN(n21170) );
  NOR2_X1 U12812 ( .A1(n21076), .A2(n18138), .ZN(n18143) );
  INV_X1 U12813 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18233) );
  NOR2_X2 U12814 ( .A1(n18218), .A2(n21366), .ZN(n18219) );
  INV_X1 U12815 ( .A(n18332), .ZN(n21439) );
  NOR2_X1 U12816 ( .A1(n15607), .A2(n15606), .ZN(n21233) );
  AOI221_X2 U12817 ( .B1(n21194), .B2(n21193), .C1(n21192), .C2(n21193), .A(
        n21897), .ZN(n21375) );
  NAND2_X1 U12818 ( .A1(n20726), .A2(n17655), .ZN(n18801) );
  INV_X1 U12819 ( .A(n18586), .ZN(n18523) );
  AOI22_X1 U12820 ( .A1(n21520), .A2(n18700), .B1(n21521), .B2(n18660), .ZN(
        n18646) );
  INV_X1 U12821 ( .A(n18736), .ZN(n18726) );
  INV_X1 U12822 ( .A(n18704), .ZN(n18739) );
  NAND2_X1 U12823 ( .A1(n21668), .A2(n21688), .ZN(n21813) );
  OR2_X1 U12824 ( .A1(n21668), .A2(n21801), .ZN(n21793) );
  INV_X1 U12825 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21852) );
  INV_X1 U12826 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21885) );
  INV_X1 U12827 ( .A(n22236), .ZN(n17652) );
  OR4_X1 U12828 ( .A1(n14272), .A2(n14271), .A3(n14270), .A4(n14269), .ZN(
        P2_U2827) );
  OAI21_X1 U12829 ( .B1(n17515), .B2(n17779), .A(n13206), .ZN(P2_U3002) );
  OR4_X1 U12830 ( .A1(n14153), .A2(n14152), .A3(n14151), .A4(n14150), .ZN(
        P3_U2651) );
  AND2_X2 U12831 ( .A1(n11309), .A2(n11312), .ZN(n11516) );
  AND2_X2 U12832 ( .A1(n16828), .A2(n14304), .ZN(n12231) );
  AOI22_X1 U12833 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11308) );
  INV_X1 U12834 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11304) );
  NOR2_X4 U12835 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16829) );
  AND2_X2 U12836 ( .A1(n11313), .A2(n16828), .ZN(n11443) );
  AOI22_X1 U12837 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11443), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11307) );
  AND2_X2 U12838 ( .A1(n11309), .A2(n14474), .ZN(n11457) );
  AOI22_X1 U12839 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11306) );
  NOR2_X4 U12840 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U12841 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U12842 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U12843 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U12844 ( .A1(n11311), .A2(n11310), .ZN(n11317) );
  AOI22_X1 U12845 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U12846 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  NOR2_X1 U12847 ( .A1(n11317), .A2(n11316), .ZN(n11318) );
  AOI22_X1 U12848 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U12849 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11443), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U12850 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11319) );
  NAND4_X1 U12851 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11328) );
  AOI22_X1 U12852 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U12853 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11169), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U12854 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U12855 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U12856 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11327) );
  AOI22_X1 U12857 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U12858 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U12859 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U12860 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11329) );
  NAND4_X1 U12861 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11339) );
  AOI22_X1 U12862 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U12863 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U12864 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11335) );
  INV_X2 U12865 ( .A(n11982), .ZN(n13530) );
  AOI22_X1 U12866 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U12867 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  AOI22_X1 U12868 ( .A1(n12231), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U12869 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U12870 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11394), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U12871 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U12872 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11349) );
  AOI22_X1 U12873 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11443), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U12874 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U12875 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11216), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U12876 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11169), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U12877 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11348) );
  NAND2_X1 U12878 ( .A1(n11717), .A2(n11588), .ZN(n11617) );
  AOI22_X1 U12879 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U12880 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11169), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U12881 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11216), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U12882 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11350) );
  NAND4_X1 U12883 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11359) );
  AOI22_X1 U12884 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U12885 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U12886 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U12887 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U12888 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11358) );
  OR2_X2 U12889 ( .A1(n11359), .A2(n11358), .ZN(n11603) );
  NAND3_X1 U12890 ( .A1(n12058), .A2(n11617), .A3(n14580), .ZN(n11373) );
  INV_X1 U12891 ( .A(n11420), .ZN(n11372) );
  AOI22_X1 U12892 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U12893 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U12894 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U12895 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U12896 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11395), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U12897 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U12898 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11366) );
  NAND2_X2 U12899 ( .A1(n11370), .A2(n11297), .ZN(n11416) );
  NAND2_X1 U12900 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11377) );
  NAND2_X1 U12901 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11376) );
  NAND2_X1 U12902 ( .A1(n11169), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11375) );
  NAND2_X1 U12903 ( .A1(n11360), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11374) );
  NAND2_X1 U12904 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U12905 ( .A1(n11950), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11380) );
  NAND2_X1 U12906 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11379) );
  NAND2_X1 U12907 ( .A1(n16824), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11378) );
  NAND2_X1 U12908 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U12909 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U12910 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U12911 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U12912 ( .A1(n12231), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U12913 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U12914 ( .A1(n11395), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U12915 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11386) );
  AOI22_X1 U12916 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11394), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U12917 ( .A1(n11169), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11360), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U12918 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11395), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U12919 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11396) );
  NAND4_X1 U12920 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11405) );
  AOI22_X1 U12921 ( .A1(n12231), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U12922 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U12923 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U12924 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11404) );
  OR2_X2 U12925 ( .A1(n11405), .A2(n11404), .ZN(n11788) );
  INV_X2 U12926 ( .A(n11788), .ZN(n14587) );
  NAND2_X1 U12927 ( .A1(n11711), .A2(n14587), .ZN(n11787) );
  INV_X1 U12928 ( .A(n14898), .ZN(n11406) );
  NAND2_X1 U12929 ( .A1(n11406), .A2(n13588), .ZN(n13562) );
  OR2_X2 U12930 ( .A1(n13562), .A2(n13577), .ZN(n11786) );
  XNOR2_X1 U12931 ( .A(n22251), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n11715) );
  OAI21_X1 U12932 ( .B1(n11715), .B2(n14287), .A(n14279), .ZN(n11409) );
  AND3_X2 U12933 ( .A1(n11787), .A2(n11786), .A3(n11409), .ZN(n11436) );
  INV_X1 U12934 ( .A(n11410), .ZN(n11411) );
  OAI21_X1 U12935 ( .B1(n11414), .B2(n16332), .A(n11413), .ZN(n11799) );
  NAND2_X1 U12936 ( .A1(n11298), .A2(n11408), .ZN(n11419) );
  NAND2_X1 U12937 ( .A1(n11419), .A2(n14909), .ZN(n11417) );
  NAND2_X1 U12938 ( .A1(n11705), .A2(n14287), .ZN(n14915) );
  OAI211_X1 U12939 ( .C1(n11794), .C2(n11173), .A(n11417), .B(n14915), .ZN(
        n11418) );
  INV_X1 U12940 ( .A(n11419), .ZN(n11421) );
  NAND2_X1 U12941 ( .A1(n11421), .A2(n14622), .ZN(n11707) );
  AOI21_X1 U12942 ( .B1(n11707), .B2(n11422), .A(n16825), .ZN(n11423) );
  NAND3_X1 U12943 ( .A1(n11436), .A2(n11432), .A3(n11423), .ZN(n11424) );
  NAND2_X1 U12944 ( .A1(n11424), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11435) );
  INV_X1 U12945 ( .A(n11435), .ZN(n11506) );
  NAND2_X1 U12946 ( .A1(n11506), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11427) );
  INV_X1 U12947 ( .A(n22207), .ZN(n11425) );
  NOR2_X1 U12948 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17648) );
  NAND2_X1 U12949 ( .A1(n17648), .A2(n22210), .ZN(n12411) );
  MUX2_X1 U12950 ( .A(n11425), .B(n12411), .S(n22454), .Z(n11426) );
  NAND3_X1 U12951 ( .A1(n11707), .A2(n14287), .A3(n11422), .ZN(n11430) );
  AND2_X1 U12952 ( .A1(n14898), .A2(n11854), .ZN(n14284) );
  NAND2_X1 U12953 ( .A1(n14622), .A2(n11603), .ZN(n11428) );
  NAND2_X1 U12954 ( .A1(n17648), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20636) );
  AOI21_X1 U12955 ( .B1(n14284), .B2(n11428), .A(n20636), .ZN(n11429) );
  NAND2_X1 U12956 ( .A1(n11432), .A2(n11431), .ZN(n11475) );
  NAND2_X1 U12957 ( .A1(n11477), .A2(n11475), .ZN(n11440) );
  INV_X1 U12958 ( .A(n11440), .ZN(n11439) );
  XNOR2_X1 U12959 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22477) );
  NAND2_X1 U12960 ( .A1(n22207), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11501) );
  OAI21_X1 U12961 ( .B1(n12411), .B2(n22477), .A(n11501), .ZN(n11433) );
  INV_X1 U12962 ( .A(n11433), .ZN(n11434) );
  OAI21_X2 U12963 ( .B1(n11435), .B2(n14307), .A(n11434), .ZN(n11438) );
  INV_X1 U12964 ( .A(n11436), .ZN(n11437) );
  XNOR2_X1 U12965 ( .A(n11438), .B(n11503), .ZN(n11441) );
  INV_X1 U12966 ( .A(n11441), .ZN(n14561) );
  NAND2_X1 U12967 ( .A1(n11440), .A2(n11441), .ZN(n14701) );
  NAND2_X1 U12968 ( .A1(n11505), .A2(n14701), .ZN(n14932) );
  AOI22_X1 U12969 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U12970 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11447) );
  BUF_X1 U12971 ( .A(n11517), .Z(n11478) );
  AOI22_X1 U12972 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U12973 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11445) );
  NAND4_X1 U12974 ( .A1(n11448), .A2(n11447), .A3(n11446), .A4(n11445), .ZN(
        n11454) );
  AOI22_X1 U12975 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U12976 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U12977 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U12978 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11449) );
  NAND4_X1 U12979 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11453) );
  NAND2_X1 U12980 ( .A1(n11490), .A2(n11614), .ZN(n11455) );
  INV_X1 U12981 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11472) );
  INV_X1 U12982 ( .A(n11490), .ZN(n11498) );
  AOI22_X1 U12983 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U12984 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11461) );
  INV_X1 U12985 ( .A(n11457), .ZN(n11986) );
  AOI22_X1 U12986 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U12987 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11459) );
  NAND4_X1 U12988 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11468) );
  AOI22_X1 U12989 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U12990 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U12991 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U12992 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11444), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U12993 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11467) );
  NAND3_X1 U12994 ( .A1(n14611), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n11614), 
        .ZN(n11469) );
  OAI21_X1 U12995 ( .B1(n11498), .B2(n11681), .A(n11469), .ZN(n11470) );
  INV_X1 U12996 ( .A(n11470), .ZN(n11471) );
  OAI21_X1 U12997 ( .B1(n11736), .B2(n11472), .A(n11471), .ZN(n11473) );
  NAND2_X1 U12998 ( .A1(n11207), .A2(n11473), .ZN(n11474) );
  AND2_X2 U12999 ( .A1(n11499), .A2(n11474), .ZN(n12066) );
  INV_X1 U13000 ( .A(n11475), .ZN(n11476) );
  AOI22_X1 U13001 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U13002 ( .A1(n11955), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U13003 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U13004 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U13005 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11489) );
  AOI22_X1 U13006 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U13007 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U13008 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U13009 ( .A1(n11442), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U13010 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11488) );
  XNOR2_X1 U13011 ( .A(n11669), .B(n11610), .ZN(n11491) );
  NAND2_X1 U13012 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  INV_X1 U13013 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U13014 ( .A1(n14611), .A2(n11610), .ZN(n11494) );
  OAI211_X1 U13015 ( .C1(n11669), .C2(n11416), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n11494), .ZN(n11495) );
  INV_X1 U13016 ( .A(n11495), .ZN(n11496) );
  NAND2_X1 U13017 ( .A1(n12066), .A2(n12068), .ZN(n11500) );
  INV_X1 U13018 ( .A(n11599), .ZN(n11530) );
  NAND2_X1 U13019 ( .A1(n11501), .A2(n14307), .ZN(n11502) );
  NAND2_X1 U13020 ( .A1(n11503), .A2(n11502), .ZN(n11504) );
  NAND2_X1 U13021 ( .A1(n11507), .A2(n17687), .ZN(n11512) );
  INV_X1 U13022 ( .A(n12411), .ZN(n11533) );
  NAND2_X1 U13023 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11508) );
  NAND2_X1 U13024 ( .A1(n17707), .A2(n11508), .ZN(n11510) );
  NAND2_X1 U13025 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22437) );
  INV_X1 U13026 ( .A(n22437), .ZN(n11509) );
  NAND2_X1 U13027 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11509), .ZN(
        n14684) );
  AND2_X1 U13028 ( .A1(n11510), .A2(n14684), .ZN(n14938) );
  AOI22_X1 U13029 ( .A1(n11533), .A2(n14938), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n22207), .ZN(n11511) );
  NAND2_X2 U13030 ( .A1(n17645), .A2(n11515), .ZN(n14822) );
  AOI22_X1 U13031 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U13032 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U13033 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U13034 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11518) );
  NAND4_X1 U13035 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n11527) );
  AOI22_X1 U13036 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U13037 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U13038 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U13039 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U13040 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11526) );
  AOI22_X1 U13041 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11744), .B2(n11631), .ZN(n11528) );
  NAND2_X1 U13042 ( .A1(n11530), .A2(n11598), .ZN(n11629) );
  INV_X1 U13043 ( .A(n11629), .ZN(n11548) );
  NAND2_X1 U13044 ( .A1(n11507), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11535) );
  INV_X1 U13045 ( .A(n14684), .ZN(n11531) );
  NAND2_X1 U13046 ( .A1(n11531), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14615) );
  NAND2_X1 U13047 ( .A1(n17709), .A2(n14684), .ZN(n11532) );
  AOI22_X1 U13048 ( .A1(n22478), .A2(n11533), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n22207), .ZN(n11534) );
  AOI22_X1 U13049 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U13050 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U13051 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11537) );
  INV_X1 U13052 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U13053 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11536) );
  NAND4_X1 U13054 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11545) );
  AOI22_X1 U13055 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U13056 ( .A1(n11361), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U13057 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U13058 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U13059 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11544) );
  AOI22_X1 U13060 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11744), .B2(n11642), .ZN(n11546) );
  INV_X1 U13061 ( .A(n11641), .ZN(n11561) );
  INV_X1 U13062 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U13063 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13535), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U13064 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13536), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13065 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11180), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U13066 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11549) );
  NAND4_X1 U13067 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11558) );
  AOI22_X1 U13068 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11179), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U13069 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U13070 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U13071 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U13072 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  NAND2_X1 U13073 ( .A1(n11744), .A2(n11651), .ZN(n11559) );
  OAI21_X1 U13074 ( .B1(n11736), .B2(n11560), .A(n11559), .ZN(n11640) );
  INV_X1 U13075 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U13076 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U13077 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13078 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13079 ( .A1(n11442), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U13080 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11571) );
  AOI22_X1 U13081 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13082 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U13083 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U13084 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U13085 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  NAND2_X1 U13086 ( .A1(n11744), .A2(n11662), .ZN(n11572) );
  OAI21_X1 U13087 ( .B1(n11736), .B2(n11573), .A(n11572), .ZN(n11649) );
  INV_X1 U13088 ( .A(n11660), .ZN(n11587) );
  NAND2_X1 U13089 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11585) );
  AOI22_X1 U13090 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U13091 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U13092 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13093 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U13094 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11583) );
  AOI22_X1 U13095 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U13096 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U13097 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U13098 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11578) );
  NAND4_X1 U13099 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11582) );
  NAND2_X1 U13100 ( .A1(n11744), .A2(n11674), .ZN(n11584) );
  AND2_X1 U13101 ( .A1(n11589), .A2(n11746), .ZN(n11590) );
  INV_X1 U13102 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n22024) );
  INV_X1 U13103 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21921) );
  NAND2_X1 U13104 ( .A1(n11597), .A2(n21921), .ZN(n11591) );
  NAND2_X1 U13105 ( .A1(n15830), .A2(n11591), .ZN(n15976) );
  INV_X1 U13106 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21993) );
  NAND2_X1 U13107 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U13108 ( .A1(n11597), .A2(n11592), .ZN(n15972) );
  NAND2_X1 U13109 ( .A1(n15974), .A2(n15972), .ZN(n11593) );
  INV_X1 U13110 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U13111 ( .A1(n16794), .A2(n11870), .ZN(n11594) );
  INV_X1 U13112 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22006) );
  OR2_X1 U13113 ( .A1(n20593), .A2(n22006), .ZN(n15931) );
  NOR2_X1 U13114 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11688) );
  OR2_X1 U13115 ( .A1(n20593), .A2(n11688), .ZN(n11596) );
  NAND2_X1 U13116 ( .A1(n15931), .A2(n11596), .ZN(n20617) );
  XNOR2_X1 U13117 ( .A(n16794), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15933) );
  NAND2_X1 U13118 ( .A1(n16794), .A2(n22006), .ZN(n15932) );
  AOI21_X1 U13119 ( .B1(n16794), .B2(n22024), .A(n20615), .ZN(n11690) );
  NAND2_X1 U13120 ( .A1(n12057), .A2(n11746), .ZN(n11607) );
  NAND2_X1 U13121 ( .A1(n11610), .A2(n11614), .ZN(n11633) );
  AND2_X1 U13122 ( .A1(n14909), .A2(n11633), .ZN(n11620) );
  INV_X1 U13123 ( .A(n11620), .ZN(n11602) );
  INV_X1 U13124 ( .A(n11633), .ZN(n11600) );
  NAND2_X1 U13125 ( .A1(n14909), .A2(n11600), .ZN(n11601) );
  MUX2_X1 U13126 ( .A(n11602), .B(n11601), .S(n11631), .Z(n11605) );
  AND2_X1 U13127 ( .A1(n14611), .A2(n11603), .ZN(n11611) );
  INV_X1 U13128 ( .A(n11611), .ZN(n11604) );
  AND2_X1 U13129 ( .A1(n11605), .A2(n11604), .ZN(n11606) );
  NAND2_X1 U13130 ( .A1(n11607), .A2(n11606), .ZN(n14435) );
  INV_X1 U13131 ( .A(n11610), .ZN(n11616) );
  AOI21_X1 U13132 ( .B1(n11616), .B2(n14909), .A(n11611), .ZN(n11612) );
  OR2_X1 U13133 ( .A1(n11207), .A2(n11704), .ZN(n11622) );
  INV_X1 U13134 ( .A(n11614), .ZN(n11615) );
  NAND2_X1 U13135 ( .A1(n11616), .A2(n11615), .ZN(n11619) );
  OR2_X1 U13136 ( .A1(n11617), .A2(n14580), .ZN(n11618) );
  AOI21_X1 U13137 ( .B1(n11620), .B2(n11619), .A(n11618), .ZN(n11621) );
  NAND2_X1 U13138 ( .A1(n11622), .A2(n11621), .ZN(n11624) );
  INV_X1 U13139 ( .A(n11623), .ZN(n14291) );
  NAND2_X1 U13140 ( .A1(n14291), .A2(n11624), .ZN(n11625) );
  NAND2_X1 U13141 ( .A1(n14327), .A2(n11625), .ZN(n11627) );
  NAND2_X1 U13142 ( .A1(n11156), .A2(n11626), .ZN(n14437) );
  NAND2_X1 U13143 ( .A1(n14435), .A2(n14437), .ZN(n11628) );
  NAND2_X1 U13144 ( .A1(n11627), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14436) );
  NAND2_X2 U13145 ( .A1(n11628), .A2(n14436), .ZN(n11638) );
  INV_X1 U13146 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21940) );
  XNOR2_X2 U13147 ( .A(n11638), .B(n21940), .ZN(n14999) );
  INV_X1 U13148 ( .A(n14554), .ZN(n14629) );
  NAND2_X1 U13149 ( .A1(n11629), .A2(n14629), .ZN(n11630) );
  OR2_X1 U13150 ( .A1(n14759), .A2(n11704), .ZN(n11637) );
  INV_X1 U13151 ( .A(n11631), .ZN(n11632) );
  NAND2_X1 U13152 ( .A1(n11633), .A2(n11632), .ZN(n11643) );
  INV_X1 U13153 ( .A(n11642), .ZN(n11634) );
  XNOR2_X1 U13154 ( .A(n11643), .B(n11634), .ZN(n11635) );
  NAND2_X1 U13155 ( .A1(n11635), .A2(n14909), .ZN(n11636) );
  NAND2_X1 U13156 ( .A1(n11637), .A2(n11636), .ZN(n14998) );
  NAND2_X1 U13157 ( .A1(n11638), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U13158 ( .A1(n14997), .A2(n11639), .ZN(n20558) );
  XNOR2_X1 U13159 ( .A(n11641), .B(n11640), .ZN(n12095) );
  NAND2_X1 U13160 ( .A1(n12095), .A2(n11746), .ZN(n11646) );
  NAND2_X1 U13161 ( .A1(n11643), .A2(n11642), .ZN(n11653) );
  XNOR2_X1 U13162 ( .A(n11653), .B(n11651), .ZN(n11644) );
  NAND2_X1 U13163 ( .A1(n11644), .A2(n14909), .ZN(n11645) );
  NAND2_X1 U13164 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  INV_X1 U13165 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21933) );
  XNOR2_X1 U13166 ( .A(n11647), .B(n21933), .ZN(n20557) );
  NAND2_X1 U13167 ( .A1(n20558), .A2(n20557), .ZN(n20560) );
  NAND2_X1 U13168 ( .A1(n11647), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U13169 ( .A1(n20560), .A2(n11648), .ZN(n20568) );
  XNOR2_X1 U13170 ( .A(n11650), .B(n11649), .ZN(n12106) );
  NAND2_X1 U13171 ( .A1(n12106), .A2(n11746), .ZN(n11656) );
  INV_X1 U13172 ( .A(n11651), .ZN(n11652) );
  OR2_X1 U13173 ( .A1(n11653), .A2(n11652), .ZN(n11661) );
  XNOR2_X1 U13174 ( .A(n11661), .B(n11662), .ZN(n11654) );
  NAND2_X1 U13175 ( .A1(n11654), .A2(n14909), .ZN(n11655) );
  NAND2_X1 U13176 ( .A1(n11656), .A2(n11655), .ZN(n11657) );
  INV_X1 U13177 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21952) );
  XNOR2_X1 U13178 ( .A(n11657), .B(n21952), .ZN(n20567) );
  NAND2_X1 U13179 ( .A1(n20568), .A2(n20567), .ZN(n20565) );
  NAND2_X1 U13180 ( .A1(n11657), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11658) );
  NAND2_X1 U13181 ( .A1(n20565), .A2(n11658), .ZN(n20576) );
  NAND2_X1 U13182 ( .A1(n11660), .A2(n11659), .ZN(n12115) );
  NAND3_X1 U13183 ( .A1(n11672), .A2(n11746), .A3(n12115), .ZN(n11666) );
  INV_X1 U13184 ( .A(n11661), .ZN(n11663) );
  NAND2_X1 U13185 ( .A1(n11663), .A2(n11662), .ZN(n11673) );
  XNOR2_X1 U13186 ( .A(n11673), .B(n11674), .ZN(n11664) );
  NAND2_X1 U13187 ( .A1(n11664), .A2(n14909), .ZN(n11665) );
  NAND2_X1 U13188 ( .A1(n11666), .A2(n11665), .ZN(n11667) );
  INV_X1 U13189 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21950) );
  XNOR2_X1 U13190 ( .A(n11667), .B(n21950), .ZN(n20575) );
  NAND2_X1 U13191 ( .A1(n20576), .A2(n20575), .ZN(n20574) );
  NAND2_X1 U13192 ( .A1(n11667), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11668) );
  NAND2_X1 U13193 ( .A1(n20574), .A2(n11668), .ZN(n20585) );
  INV_X1 U13194 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11670) );
  INV_X1 U13195 ( .A(n11744), .ZN(n11740) );
  OAI22_X1 U13196 ( .A1(n11736), .A2(n11670), .B1(n11740), .B2(n11669), .ZN(
        n11671) );
  NAND2_X1 U13197 ( .A1(n12054), .A2(n11746), .ZN(n11678) );
  INV_X1 U13198 ( .A(n11673), .ZN(n11675) );
  NAND2_X1 U13199 ( .A1(n11675), .A2(n11674), .ZN(n11683) );
  XNOR2_X1 U13200 ( .A(n11683), .B(n11681), .ZN(n11676) );
  NAND2_X1 U13201 ( .A1(n11676), .A2(n14909), .ZN(n11677) );
  NAND2_X1 U13202 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  INV_X1 U13203 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21970) );
  XNOR2_X1 U13204 ( .A(n11679), .B(n21970), .ZN(n20584) );
  NAND2_X1 U13205 ( .A1(n20585), .A2(n20584), .ZN(n20583) );
  NAND2_X1 U13206 ( .A1(n11679), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11680) );
  NAND2_X1 U13207 ( .A1(n20583), .A2(n11680), .ZN(n15088) );
  NAND2_X1 U13208 ( .A1(n14909), .A2(n11681), .ZN(n11682) );
  OR2_X1 U13209 ( .A1(n11683), .A2(n11682), .ZN(n11684) );
  NAND2_X1 U13210 ( .A1(n11597), .A2(n11684), .ZN(n11685) );
  INV_X1 U13211 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15092) );
  XNOR2_X1 U13212 ( .A(n11685), .B(n15092), .ZN(n15087) );
  NAND2_X1 U13213 ( .A1(n15088), .A2(n15087), .ZN(n15086) );
  NAND2_X1 U13214 ( .A1(n11685), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11686) );
  XNOR2_X1 U13215 ( .A(n16794), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15688) );
  INV_X1 U13216 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21977) );
  NOR2_X1 U13217 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15970) );
  AND2_X1 U13218 ( .A1(n15970), .A2(n21993), .ZN(n15829) );
  AOI21_X1 U13219 ( .B1(n11688), .B2(n15829), .A(n20593), .ZN(n15929) );
  NOR2_X1 U13220 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15935) );
  AOI21_X1 U13221 ( .B1(n15935), .B2(n22024), .A(n20593), .ZN(n11689) );
  INV_X1 U13222 ( .A(n11692), .ZN(n11691) );
  AND2_X1 U13223 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16770) );
  AND2_X1 U13224 ( .A1(n16770), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n22045) );
  INV_X1 U13225 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22011) );
  INV_X1 U13226 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22043) );
  NOR2_X1 U13227 ( .A1(n16685), .A2(n22043), .ZN(n11694) );
  NOR4_X1 U13228 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11693) );
  NOR2_X1 U13229 ( .A1(n11694), .A2(n16684), .ZN(n16623) );
  NOR3_X1 U13230 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16625) );
  NAND2_X1 U13231 ( .A1(n16623), .A2(n16625), .ZN(n11698) );
  INV_X1 U13232 ( .A(n11694), .ZN(n16658) );
  INV_X1 U13233 ( .A(n16658), .ZN(n11695) );
  NAND2_X1 U13234 ( .A1(n11695), .A2(n16794), .ZN(n11696) );
  NAND2_X1 U13235 ( .A1(n11698), .A2(n11696), .ZN(n11697) );
  AND2_X1 U13236 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U13237 ( .A1(n16729), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U13238 ( .A1(n16794), .A2(n11822), .ZN(n16624) );
  INV_X1 U13239 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16734) );
  NOR2_X1 U13240 ( .A1(n11160), .A2(n11699), .ZN(n16638) );
  NOR2_X1 U13241 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16708) );
  NAND2_X1 U13242 ( .A1(n16638), .A2(n16708), .ZN(n16126) );
  NAND2_X1 U13243 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16257) );
  INV_X1 U13244 ( .A(n16257), .ZN(n11700) );
  AOI21_X1 U13245 ( .B1(n16650), .B2(n11700), .A(n11595), .ZN(n11701) );
  INV_X1 U13246 ( .A(n11701), .ZN(n16128) );
  NAND2_X1 U13247 ( .A1(n16126), .A2(n16128), .ZN(n14002) );
  INV_X1 U13248 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16125) );
  XNOR2_X1 U13249 ( .A(n16794), .B(n16125), .ZN(n16127) );
  NOR2_X1 U13250 ( .A1(n11704), .A2(n11703), .ZN(n11806) );
  INV_X1 U13251 ( .A(n16332), .ZN(n14611) );
  NOR2_X1 U13252 ( .A1(n11806), .A2(n14611), .ZN(n11706) );
  AND2_X1 U13253 ( .A1(n11707), .A2(n11706), .ZN(n11798) );
  INV_X1 U13254 ( .A(n11805), .ZN(n11795) );
  NOR2_X1 U13255 ( .A1(n11422), .A2(n11795), .ZN(n14303) );
  AND2_X1 U13256 ( .A1(n11805), .A2(n16332), .ZN(n11708) );
  OR2_X1 U13257 ( .A1(n14303), .A2(n11708), .ZN(n11710) );
  OR2_X1 U13258 ( .A1(n14622), .A2(n11416), .ZN(n11709) );
  AND2_X1 U13259 ( .A1(n11298), .A2(n11709), .ZN(n11797) );
  NAND2_X1 U13260 ( .A1(n11710), .A2(n11797), .ZN(n11784) );
  INV_X1 U13261 ( .A(n11712), .ZN(n16448) );
  OAI21_X1 U13262 ( .B1(n11798), .B2(n11784), .A(n16448), .ZN(n14319) );
  INV_X1 U13263 ( .A(n14317), .ZN(n14300) );
  NAND2_X1 U13264 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22243) );
  INV_X1 U13265 ( .A(n22243), .ZN(n22242) );
  OR2_X1 U13266 ( .A1(n14300), .A2(n22242), .ZN(n13558) );
  INV_X1 U13267 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U13268 ( .A1(n11715), .A2(n11714), .ZN(n22254) );
  NAND2_X1 U13269 ( .A1(n14587), .A2(n22254), .ZN(n14903) );
  INV_X1 U13270 ( .A(n14903), .ZN(n11716) );
  OAI211_X1 U13271 ( .C1(n13558), .C2(n11716), .A(n16332), .B(n13577), .ZN(
        n11771) );
  NAND2_X1 U13272 ( .A1(n22408), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U13273 ( .A1(n14307), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U13274 ( .A1(n11719), .A2(n11718), .ZN(n11735) );
  NAND2_X1 U13275 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n22454), .ZN(
        n11737) );
  NAND2_X1 U13276 ( .A1(n11720), .A2(n11719), .ZN(n11731) );
  MUX2_X1 U13277 ( .A(n17707), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n17687), .Z(n11729) );
  NAND2_X1 U13278 ( .A1(n11731), .A2(n11729), .ZN(n11722) );
  NAND2_X1 U13279 ( .A1(n17707), .A2(n17687), .ZN(n11721) );
  NAND2_X1 U13280 ( .A1(n11722), .A2(n11721), .ZN(n11759) );
  NAND2_X1 U13281 ( .A1(n17709), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U13282 ( .A1(n17685), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U13283 ( .A1(n11759), .A2(n11758), .ZN(n11726) );
  INV_X1 U13284 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17729) );
  NAND2_X1 U13285 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17729), .ZN(
        n11724) );
  AND2_X1 U13286 ( .A1(n11755), .A2(n11724), .ZN(n11725) );
  NAND2_X1 U13287 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  NAND2_X1 U13288 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17696), .ZN(
        n11756) );
  NAND2_X1 U13289 ( .A1(n11727), .A2(n11756), .ZN(n11777) );
  INV_X1 U13290 ( .A(n11777), .ZN(n11728) );
  NAND2_X1 U13291 ( .A1(n11744), .A2(n11728), .ZN(n11770) );
  INV_X1 U13292 ( .A(n11729), .ZN(n11730) );
  XNOR2_X1 U13293 ( .A(n11731), .B(n11730), .ZN(n11773) );
  NAND2_X1 U13294 ( .A1(n11744), .A2(n11773), .ZN(n11733) );
  INV_X1 U13295 ( .A(n11733), .ZN(n11754) );
  NAND2_X1 U13296 ( .A1(n14559), .A2(n16332), .ZN(n11732) );
  NAND2_X1 U13297 ( .A1(n11732), .A2(n14587), .ZN(n11738) );
  INV_X1 U13298 ( .A(n11738), .ZN(n11753) );
  OAI211_X1 U13299 ( .C1(n11773), .C2(n11736), .A(n11733), .B(n11738), .ZN(
        n11752) );
  INV_X1 U13300 ( .A(n11737), .ZN(n11734) );
  XNOR2_X1 U13301 ( .A(n11735), .B(n11734), .ZN(n11774) );
  OAI22_X1 U13302 ( .A1(n22210), .A2(n15726), .B1(n11736), .B2(n11774), .ZN(
        n11745) );
  NOR3_X1 U13303 ( .A1(n14287), .A2(n11774), .A3(n11745), .ZN(n11750) );
  OAI21_X1 U13304 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n22454), .A(
        n11737), .ZN(n11741) );
  INV_X1 U13305 ( .A(n11741), .ZN(n11739) );
  OAI211_X1 U13306 ( .C1(n14611), .C2(n11794), .A(n11739), .B(n11738), .ZN(
        n11743) );
  OAI21_X1 U13307 ( .B1(n11741), .B2(n11740), .A(n11761), .ZN(n11742) );
  NAND2_X1 U13308 ( .A1(n11743), .A2(n11742), .ZN(n11749) );
  NAND3_X1 U13309 ( .A1(n11744), .A2(n14287), .A3(n11774), .ZN(n11748) );
  OAI21_X1 U13310 ( .B1(n11746), .B2(n11774), .A(n11745), .ZN(n11747) );
  OAI211_X1 U13311 ( .C1(n11750), .C2(n11749), .A(n11748), .B(n11747), .ZN(
        n11751) );
  AOI22_X1 U13312 ( .A1(n11754), .A2(n11753), .B1(n11752), .B2(n11751), .ZN(
        n11764) );
  INV_X1 U13313 ( .A(n11755), .ZN(n11757) );
  OAI22_X1 U13314 ( .A1(n11759), .A2(n11758), .B1(n11757), .B2(n11756), .ZN(
        n11776) );
  INV_X1 U13315 ( .A(n11776), .ZN(n11762) );
  NOR2_X1 U13316 ( .A1(n11760), .A2(n11762), .ZN(n11763) );
  OAI22_X1 U13317 ( .A1(n11764), .A2(n11763), .B1(n11762), .B2(n11761), .ZN(
        n11765) );
  AOI21_X1 U13318 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n22210), .A(
        n11765), .ZN(n11766) );
  INV_X1 U13319 ( .A(n11766), .ZN(n11767) );
  NAND3_X1 U13320 ( .A1(n11771), .A2(n11411), .A3(n16461), .ZN(n11782) );
  INV_X1 U13321 ( .A(n11806), .ZN(n11772) );
  OR2_X1 U13322 ( .A1(n16461), .A2(n11772), .ZN(n11781) );
  NAND2_X1 U13323 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  OR2_X1 U13324 ( .A1(n11776), .A2(n11775), .ZN(n11778) );
  AND2_X1 U13325 ( .A1(n11778), .A2(n11777), .ZN(n16447) );
  NAND2_X1 U13326 ( .A1(n14287), .A2(n22254), .ZN(n11779) );
  NAND4_X1 U13327 ( .A1(n16447), .A2(n22243), .A3(n11410), .A4(n11779), .ZN(
        n11780) );
  NAND4_X1 U13328 ( .A1(n14319), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11783) );
  NOR2_X1 U13329 ( .A1(n11784), .A2(n11794), .ZN(n17690) );
  INV_X1 U13330 ( .A(n14898), .ZN(n16462) );
  NAND2_X1 U13331 ( .A1(n14303), .A2(n16462), .ZN(n13557) );
  INV_X1 U13332 ( .A(n13557), .ZN(n11785) );
  OR2_X1 U13333 ( .A1(n17690), .A2(n11785), .ZN(n16460) );
  INV_X1 U13334 ( .A(n16460), .ZN(n11792) );
  CLKBUF_X1 U13335 ( .A(n11786), .Z(n11917) );
  NAND2_X1 U13336 ( .A1(n14317), .A2(n11174), .ZN(n11789) );
  OAI211_X1 U13337 ( .C1(n11408), .C2(n11917), .A(n11192), .B(n11789), .ZN(
        n11790) );
  INV_X1 U13338 ( .A(n11790), .ZN(n11791) );
  NAND2_X1 U13339 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  INV_X1 U13340 ( .A(n16825), .ZN(n14305) );
  INV_X1 U13342 ( .A(n14915), .ZN(n14315) );
  AOI22_X1 U13343 ( .A1(n11795), .A2(n16254), .B1(n14315), .B2(n11794), .ZN(
        n11796) );
  OAI21_X1 U13344 ( .B1(n11797), .B2(n11854), .A(n11796), .ZN(n11800) );
  OR3_X1 U13345 ( .A1(n11800), .A2(n11799), .A3(n11798), .ZN(n14302) );
  INV_X1 U13346 ( .A(n14302), .ZN(n11801) );
  OAI21_X1 U13347 ( .B1(n11703), .B2(n14305), .A(n11801), .ZN(n11802) );
  NAND2_X1 U13348 ( .A1(n11919), .A2(n11802), .ZN(n15846) );
  INV_X1 U13349 ( .A(n15846), .ZN(n15848) );
  INV_X1 U13350 ( .A(n16729), .ZN(n11815) );
  NAND2_X1 U13351 ( .A1(n11919), .A2(n16834), .ZN(n15845) );
  INV_X1 U13352 ( .A(n14621), .ZN(n15727) );
  NOR2_X1 U13353 ( .A1(n15727), .A2(n11803), .ZN(n11804) );
  INV_X1 U13354 ( .A(n11822), .ZN(n11807) );
  AOI21_X1 U13355 ( .B1(n15845), .B2(n15936), .A(n11807), .ZN(n11814) );
  NAND2_X1 U13356 ( .A1(n15845), .A2(n15846), .ZN(n21981) );
  INV_X1 U13357 ( .A(n21981), .ZN(n21944) );
  AND2_X1 U13358 ( .A1(n22045), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11817) );
  OR2_X1 U13359 ( .A1(n15846), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11808) );
  OR2_X1 U13360 ( .A1(n11919), .A2(n22040), .ZN(n14329) );
  INV_X1 U13361 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n22003) );
  NOR2_X1 U13362 ( .A1(n21933), .A2(n21940), .ZN(n21927) );
  NAND3_X1 U13363 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21927), .ZN(n21965) );
  NOR2_X1 U13364 ( .A1(n21952), .A2(n21965), .ZN(n15090) );
  NOR3_X1 U13365 ( .A1(n15092), .A2(n21970), .A3(n21950), .ZN(n15872) );
  AND2_X1 U13366 ( .A1(n15090), .A2(n15872), .ZN(n15874) );
  NAND3_X1 U13367 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n15874), .ZN(n21980) );
  NOR3_X1 U13368 ( .A1(n22003), .A2(n21993), .A3(n21980), .ZN(n21916) );
  NOR2_X1 U13369 ( .A1(n11870), .A2(n21921), .ZN(n15938) );
  NAND2_X1 U13370 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22026) );
  NOR2_X1 U13371 ( .A1(n22024), .A2(n22026), .ZN(n22014) );
  NAND2_X1 U13372 ( .A1(n15938), .A2(n22014), .ZN(n22023) );
  NOR2_X1 U13373 ( .A1(n22011), .A2(n22023), .ZN(n11810) );
  NAND2_X1 U13374 ( .A1(n21916), .A2(n11810), .ZN(n11819) );
  NAND2_X1 U13375 ( .A1(n21981), .A2(n11819), .ZN(n11809) );
  NAND2_X1 U13376 ( .A1(n15873), .A2(n11809), .ZN(n16783) );
  INV_X1 U13377 ( .A(n16783), .ZN(n11813) );
  INV_X1 U13378 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16750) );
  INV_X1 U13379 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15877) );
  INV_X1 U13380 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14388) );
  INV_X1 U13381 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14444) );
  OAI21_X1 U13382 ( .B1(n14388), .B2(n14444), .A(n11626), .ZN(n21925) );
  NAND2_X1 U13383 ( .A1(n21927), .A2(n21925), .ZN(n21956) );
  NOR2_X1 U13384 ( .A1(n21952), .A2(n21956), .ZN(n15089) );
  NAND2_X1 U13385 ( .A1(n15872), .A2(n15089), .ZN(n15876) );
  NOR3_X1 U13386 ( .A1(n21977), .A2(n15877), .A3(n15876), .ZN(n15839) );
  NAND2_X1 U13387 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15839), .ZN(
        n21984) );
  NOR2_X1 U13388 ( .A1(n21993), .A2(n21984), .ZN(n15937) );
  NAND2_X1 U13389 ( .A1(n11810), .A2(n15937), .ZN(n16784) );
  INV_X1 U13390 ( .A(n16784), .ZN(n11811) );
  NAND2_X1 U13391 ( .A1(n11811), .A2(n11817), .ZN(n11820) );
  OAI21_X1 U13392 ( .B1(n16750), .B2(n11820), .A(n21985), .ZN(n11812) );
  OAI211_X1 U13393 ( .C1(n21944), .C2(n11817), .A(n11813), .B(n11812), .ZN(
        n16762) );
  AOI211_X1 U13394 ( .C1(n15848), .C2(n11815), .A(n11814), .B(n16762), .ZN(
        n16739) );
  NAND3_X1 U13395 ( .A1(n16739), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16134) );
  INV_X1 U13396 ( .A(n16134), .ZN(n11816) );
  AND2_X1 U13397 ( .A1(n15936), .A2(n15846), .ZN(n14296) );
  AND2_X1 U13398 ( .A1(n14296), .A2(n15845), .ZN(n22015) );
  NAND2_X1 U13399 ( .A1(n22015), .A2(n15873), .ZN(n16776) );
  INV_X1 U13400 ( .A(n16776), .ZN(n16260) );
  AOI21_X1 U13401 ( .B1(n11816), .B2(n11700), .A(n16260), .ZN(n16132) );
  INV_X1 U13402 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n16480) );
  NOR2_X1 U13403 ( .A1(n22016), .A2(n16480), .ZN(n12414) );
  NAND2_X1 U13404 ( .A1(n14388), .A2(n15845), .ZN(n14331) );
  NAND2_X1 U13405 ( .A1(n21981), .A2(n14331), .ZN(n15838) );
  INV_X1 U13406 ( .A(n11817), .ZN(n11818) );
  OR3_X1 U13407 ( .A1(n15838), .A2(n11819), .A3(n11818), .ZN(n16749) );
  OR2_X1 U13408 ( .A1(n15936), .A2(n11820), .ZN(n11821) );
  NOR2_X1 U13409 ( .A1(n16764), .A2(n11822), .ZN(n16735) );
  NAND2_X1 U13410 ( .A1(n16735), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16717) );
  NOR2_X1 U13411 ( .A1(n16717), .A2(n16257), .ZN(n16264) );
  INV_X1 U13412 ( .A(n16264), .ZN(n11823) );
  NOR2_X1 U13413 ( .A1(n11823), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11824) );
  AOI211_X1 U13414 ( .C1(n16132), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12414), .B(n11824), .ZN(n11825) );
  OAI22_X1 U13415 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n11229), .ZN(n13593) );
  MUX2_X1 U13416 ( .A(P1_EBX_REG_29__SCAN_IN), .B(n13593), .S(n11173), .Z(
        n11916) );
  NAND2_X1 U13417 ( .A1(n11231), .A2(n14444), .ZN(n11828) );
  INV_X1 U13418 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U13419 ( .A1(n11174), .A2(n15315), .ZN(n11827) );
  NAND3_X1 U13420 ( .A1(n11828), .A2(n11827), .A3(n11173), .ZN(n11829) );
  MUX2_X1 U13421 ( .A(n11830), .B(n11231), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14294) );
  INV_X1 U13422 ( .A(n14294), .ZN(n11831) );
  OAI21_X1 U13423 ( .B1(n14325), .B2(n11228), .A(n11832), .ZN(n14442) );
  INV_X1 U13424 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n16315) );
  NAND2_X1 U13425 ( .A1(n11899), .A2(n16315), .ZN(n11835) );
  NAND2_X1 U13426 ( .A1(n11907), .A2(n11626), .ZN(n11833) );
  OAI211_X1 U13427 ( .C1(n11228), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11833), .B(
        n11173), .ZN(n11834) );
  MUX2_X1 U13428 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11840) );
  OR2_X1 U13429 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U13430 ( .A1(n11840), .A2(n11839), .ZN(n14799) );
  NAND2_X1 U13431 ( .A1(n11907), .A2(n21933), .ZN(n11841) );
  OAI211_X1 U13432 ( .C1(P1_EBX_REG_4__SCAN_IN), .C2(n11229), .A(n11841), .B(
        n11854), .ZN(n11842) );
  OAI21_X1 U13433 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n11913), .A(n11842), .ZN(
        n14818) );
  NAND2_X1 U13434 ( .A1(n14819), .A2(n14818), .ZN(n14817) );
  INV_X1 U13435 ( .A(n14817), .ZN(n11847) );
  OR2_X1 U13436 ( .A1(n11910), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U13437 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11843) );
  OAI211_X1 U13438 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n11229), .A(n11907), .B(
        n11843), .ZN(n11844) );
  NAND2_X1 U13439 ( .A1(n11845), .A2(n11844), .ZN(n14990) );
  NAND2_X1 U13440 ( .A1(n11847), .A2(n11846), .ZN(n14960) );
  INV_X1 U13441 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14963) );
  NAND2_X1 U13442 ( .A1(n11899), .A2(n14963), .ZN(n11850) );
  NAND2_X1 U13443 ( .A1(n11907), .A2(n21950), .ZN(n11848) );
  OAI211_X1 U13444 ( .C1(P1_EBX_REG_6__SCAN_IN), .C2(n11229), .A(n11848), .B(
        n11854), .ZN(n11849) );
  OR2_X2 U13445 ( .A1(n14960), .A2(n14961), .ZN(n15120) );
  OR2_X1 U13446 ( .A1(n11910), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11853) );
  NAND2_X1 U13447 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11851) );
  OAI211_X1 U13448 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n11229), .A(n11907), .B(
        n11851), .ZN(n11852) );
  NAND2_X1 U13449 ( .A1(n11853), .A2(n11852), .ZN(n15119) );
  NAND2_X1 U13450 ( .A1(n11907), .A2(n15092), .ZN(n11855) );
  OAI211_X1 U13451 ( .C1(P1_EBX_REG_8__SCAN_IN), .C2(n11229), .A(n11855), .B(
        n11854), .ZN(n11856) );
  OAI21_X1 U13452 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n11913), .A(n11856), .ZN(
        n15094) );
  MUX2_X1 U13453 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11858) );
  OR2_X1 U13454 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U13455 ( .A1(n11858), .A2(n11857), .ZN(n15713) );
  INV_X1 U13456 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15484) );
  NAND2_X1 U13457 ( .A1(n11899), .A2(n15484), .ZN(n11861) );
  NAND2_X1 U13458 ( .A1(n11907), .A2(n15877), .ZN(n11859) );
  OAI211_X1 U13459 ( .C1(P1_EBX_REG_10__SCAN_IN), .C2(n11228), .A(n11859), .B(
        n11854), .ZN(n11860) );
  OR2_X1 U13460 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11863) );
  MUX2_X1 U13461 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11862) );
  AND2_X1 U13462 ( .A1(n11863), .A2(n11862), .ZN(n15698) );
  NAND2_X1 U13463 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U13464 ( .A1(n11907), .A2(n11864), .ZN(n11866) );
  OR2_X1 U13465 ( .A1(n11229), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U13466 ( .A1(n11866), .A2(n11865), .ZN(n11867) );
  OAI21_X1 U13467 ( .B1(n11913), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11867), .ZN(
        n15906) );
  MUX2_X1 U13468 ( .A(n11910), .B(n11854), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11869) );
  OR2_X1 U13469 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U13470 ( .A1(n11869), .A2(n11868), .ZN(n15895) );
  INV_X1 U13471 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n22104) );
  NAND2_X1 U13472 ( .A1(n11899), .A2(n22104), .ZN(n11873) );
  NAND2_X1 U13473 ( .A1(n11907), .A2(n11870), .ZN(n11871) );
  OAI211_X1 U13474 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n11229), .A(n11871), .B(
        n11854), .ZN(n11872) );
  NAND2_X1 U13475 ( .A1(n11185), .A2(n11874), .ZN(n11875) );
  MUX2_X1 U13476 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11877) );
  OR2_X1 U13477 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11876) );
  INV_X1 U13478 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20614) );
  NAND2_X1 U13479 ( .A1(n11907), .A2(n20614), .ZN(n11878) );
  OAI211_X1 U13480 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n11229), .A(n11878), .B(
        n11173), .ZN(n11879) );
  OAI21_X1 U13481 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(n11913), .A(n11879), .ZN(
        n15785) );
  NAND2_X1 U13482 ( .A1(n15798), .A2(n15785), .ZN(n15750) );
  MUX2_X1 U13483 ( .A(n11910), .B(n11854), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11881) );
  OR2_X1 U13484 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U13485 ( .A1(n11881), .A2(n11880), .ZN(n15751) );
  INV_X1 U13486 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n22127) );
  NAND2_X1 U13487 ( .A1(n11899), .A2(n22127), .ZN(n11884) );
  NAND2_X1 U13488 ( .A1(n11907), .A2(n22011), .ZN(n11882) );
  OAI211_X1 U13489 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n11228), .A(n11882), .B(
        n11173), .ZN(n11883) );
  AND2_X1 U13490 ( .A1(n11884), .A2(n11883), .ZN(n15863) );
  MUX2_X1 U13491 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11886) );
  OAI21_X1 U13492 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16254), .A(
        n11886), .ZN(n15983) );
  INV_X1 U13493 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16785) );
  NAND2_X1 U13494 ( .A1(n11907), .A2(n16785), .ZN(n11888) );
  INV_X1 U13495 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15993) );
  NAND2_X1 U13496 ( .A1(n11174), .A2(n15993), .ZN(n11887) );
  NAND3_X1 U13497 ( .A1(n11888), .A2(n11887), .A3(n11173), .ZN(n11889) );
  OAI21_X1 U13498 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n11913), .A(n11889), .ZN(
        n15990) );
  MUX2_X1 U13499 ( .A(n11910), .B(n11854), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11891) );
  OR2_X1 U13500 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11890) );
  AND2_X1 U13501 ( .A1(n11891), .A2(n11890), .ZN(n16773) );
  NAND2_X1 U13502 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U13503 ( .A1(n11907), .A2(n11892), .ZN(n11894) );
  OR2_X1 U13504 ( .A1(n11229), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U13505 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  OAI21_X1 U13506 ( .B1(n11913), .B2(P1_EBX_REG_22__SCAN_IN), .A(n11895), .ZN(
        n16547) );
  MUX2_X1 U13507 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11897) );
  OR2_X1 U13508 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11896) );
  NAND2_X1 U13509 ( .A1(n11897), .A2(n11896), .ZN(n16758) );
  INV_X1 U13510 ( .A(n11898), .ZN(n16760) );
  INV_X1 U13511 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n22190) );
  NAND2_X1 U13512 ( .A1(n11899), .A2(n22190), .ZN(n11903) );
  NAND2_X1 U13513 ( .A1(n11854), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U13514 ( .A1(n11907), .A2(n11900), .ZN(n11901) );
  OAI21_X1 U13515 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n11229), .A(n11901), .ZN(
        n11902) );
  AND2_X1 U13516 ( .A1(n11903), .A2(n11902), .ZN(n16566) );
  OR2_X1 U13517 ( .A1(n11910), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U13518 ( .A1(n11173), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11904) );
  OAI211_X1 U13519 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n11229), .A(n11907), .B(
        n11904), .ZN(n11905) );
  AND2_X1 U13520 ( .A1(n11906), .A2(n11905), .ZN(n16528) );
  AND2_X2 U13521 ( .A1(n16527), .A2(n16528), .ZN(n16530) );
  INV_X1 U13522 ( .A(n11907), .ZN(n11912) );
  AOI21_X1 U13523 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n11854), .A(
        n11912), .ZN(n11909) );
  NOR2_X1 U13524 ( .A1(n11229), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n11908) );
  OAI22_X1 U13525 ( .A1(n11909), .A2(n11908), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n11913), .ZN(n16522) );
  MUX2_X1 U13526 ( .A(n11910), .B(n11173), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11911) );
  OAI21_X1 U13527 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16254), .A(
        n11911), .ZN(n16511) );
  AOI21_X1 U13528 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11173), .A(
        n11912), .ZN(n11915) );
  NOR2_X1 U13529 ( .A1(n11228), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n11914) );
  OAI22_X1 U13530 ( .A1(n11915), .A2(n11914), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n11913), .ZN(n16498) );
  NOR2_X4 U13531 ( .A1(n13592), .A2(n11916), .ZN(n16251) );
  AOI21_X1 U13532 ( .B1(n11916), .B2(n16497), .A(n16251), .ZN(n16559) );
  NAND2_X1 U13533 ( .A1(n14317), .A2(n14909), .ZN(n17718) );
  OAI21_X1 U13534 ( .B1(n11917), .B2(n11416), .A(n17718), .ZN(n11918) );
  OAI21_X1 U13535 ( .B1(n12418), .B2(n22033), .A(n11921), .ZN(P1_U3002) );
  INV_X1 U13536 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15753) );
  INV_X1 U13537 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16551) );
  INV_X1 U13538 ( .A(n12368), .ZN(n11924) );
  INV_X1 U13539 ( .A(n12382), .ZN(n11925) );
  INV_X1 U13540 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11926) );
  INV_X1 U13541 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U13542 ( .A1(n11928), .A2(n11927), .ZN(n11929) );
  NAND2_X1 U13543 ( .A1(n14015), .A2(n11929), .ZN(n16484) );
  AOI22_X1 U13544 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11443), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13545 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U13546 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U13547 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11930) );
  NAND4_X1 U13548 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11939) );
  AOI22_X1 U13549 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12333), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U13550 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U13551 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U13552 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11934) );
  NAND4_X1 U13553 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11938) );
  NOR2_X1 U13554 ( .A1(n11939), .A2(n11938), .ZN(n12393) );
  AOI22_X1 U13555 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U13556 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U13557 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U13558 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U13559 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11949) );
  AOI22_X1 U13560 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U13561 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13536), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U13562 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13563 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U13564 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11948) );
  NOR2_X1 U13565 ( .A1(n11949), .A2(n11948), .ZN(n12377) );
  AOI22_X1 U13566 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U13567 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U13568 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U13569 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U13570 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11961) );
  AOI22_X1 U13571 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U13572 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13573 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13574 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U13575 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  NOR2_X1 U13576 ( .A1(n11961), .A2(n11960), .ZN(n12352) );
  AOI22_X1 U13577 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13536), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U13578 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U13579 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U13580 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11962) );
  NAND4_X1 U13581 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n11971) );
  AOI22_X1 U13582 ( .A1(n11442), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U13583 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13584 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13585 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U13586 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  NOR2_X1 U13587 ( .A1(n11971), .A2(n11970), .ZN(n12351) );
  NOR2_X1 U13588 ( .A1(n12352), .A2(n12351), .ZN(n12364) );
  AOI22_X1 U13589 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U13590 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U13591 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13592 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11972) );
  NAND4_X1 U13593 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n11981) );
  AOI22_X1 U13594 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U13595 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U13596 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U13597 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U13598 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11980) );
  OR2_X1 U13599 ( .A1(n11981), .A2(n11980), .ZN(n12362) );
  NAND2_X1 U13600 ( .A1(n12364), .A2(n12362), .ZN(n12376) );
  NOR2_X1 U13601 ( .A1(n12377), .A2(n12376), .ZN(n12383) );
  INV_X1 U13602 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15018) );
  NOR2_X1 U13603 ( .A1(n11982), .A2(n15018), .ZN(n11988) );
  INV_X1 U13604 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11985) );
  OAI22_X1 U13605 ( .A1(n11986), .A2(n11985), .B1(n11230), .B2(n11983), .ZN(
        n11987) );
  AOI211_X1 U13606 ( .C1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .C2(n11517), .A(
        n11988), .B(n11987), .ZN(n11996) );
  AOI22_X1 U13607 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U13608 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U13609 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U13610 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11989) );
  AND4_X1 U13611 ( .A1(n11992), .A2(n11991), .A3(n11990), .A4(n11989), .ZN(
        n11995) );
  AOI22_X1 U13612 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U13613 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U13614 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12384) );
  NAND2_X1 U13615 ( .A1(n12383), .A2(n12384), .ZN(n12394) );
  NOR2_X1 U13616 ( .A1(n12393), .A2(n12394), .ZN(n12402) );
  AOI22_X1 U13617 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U13618 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U13619 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U13620 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U13621 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12006) );
  AOI22_X1 U13622 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U13623 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U13624 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U13625 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12001) );
  NAND4_X1 U13626 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  OR2_X1 U13627 ( .A1(n12006), .A2(n12005), .ZN(n12403) );
  NAND2_X1 U13628 ( .A1(n12402), .A2(n12403), .ZN(n13526) );
  AOI22_X1 U13629 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U13630 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U13631 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U13632 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12007) );
  NAND4_X1 U13633 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12016) );
  AOI22_X1 U13634 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13536), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U13635 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U13636 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U13637 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12011) );
  NAND4_X1 U13638 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12015) );
  NOR2_X1 U13639 ( .A1(n12016), .A2(n12015), .ZN(n13527) );
  XNOR2_X1 U13640 ( .A(n13526), .B(n13527), .ZN(n12019) );
  AOI21_X1 U13641 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22476), .A(
        n13548), .ZN(n12018) );
  NAND2_X1 U13642 ( .A1(n13553), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12017) );
  OAI211_X1 U13643 ( .C1(n12019), .C2(n12397), .A(n12018), .B(n12017), .ZN(
        n12020) );
  OAI21_X1 U13644 ( .B1(n12400), .B2(n16484), .A(n12020), .ZN(n12410) );
  XOR2_X1 U13645 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12021), .Z(n22084) );
  INV_X1 U13646 ( .A(n22084), .ZN(n12036) );
  INV_X1 U13647 ( .A(n12239), .ZN(n12256) );
  AOI22_X1 U13648 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U13649 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U13650 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U13651 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12022) );
  NAND4_X1 U13652 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n12031) );
  AOI22_X1 U13653 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U13654 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U13655 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U13656 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U13657 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12030) );
  NOR2_X1 U13658 ( .A1(n12031), .A2(n12030), .ZN(n12034) );
  NAND2_X1 U13659 ( .A1(n13553), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U13660 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12032) );
  OAI211_X1 U13661 ( .C1(n12256), .C2(n12034), .A(n12033), .B(n12032), .ZN(
        n12035) );
  AOI21_X1 U13662 ( .B1(n12036), .B2(n12312), .A(n12035), .ZN(n15686) );
  XNOR2_X1 U13663 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12050), .ZN(
        n15644) );
  INV_X1 U13664 ( .A(n13552), .ZN(n12129) );
  OAI22_X1 U13665 ( .A1(n12400), .A2(n15644), .B1(n12129), .B2(n15647), .ZN(
        n12037) );
  AOI21_X1 U13666 ( .B1(n13553), .B2(P1_EAX_REG_8__SCAN_IN), .A(n12037), .ZN(
        n12049) );
  AOI22_X1 U13667 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U13668 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U13669 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U13670 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U13671 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12047) );
  AOI22_X1 U13672 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U13673 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U13674 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U13675 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12042) );
  NAND4_X1 U13676 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n12046) );
  OAI21_X1 U13677 ( .B1(n12047), .B2(n12046), .A(n12239), .ZN(n12048) );
  NOR2_X1 U13678 ( .A1(n15686), .A2(n15633), .ZN(n12056) );
  INV_X1 U13679 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12052) );
  OAI21_X1 U13680 ( .B1(n12116), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12050), .ZN(n22079) );
  AOI22_X1 U13681 ( .A1(n22079), .A2(n12312), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12051) );
  OAI21_X1 U13682 ( .B1(n12405), .B2(n12052), .A(n12051), .ZN(n12053) );
  INV_X1 U13683 ( .A(n15117), .ZN(n12055) );
  NAND2_X1 U13684 ( .A1(n12056), .A2(n12055), .ZN(n12126) );
  NAND2_X1 U13685 ( .A1(n12057), .A2(n12239), .ZN(n12065) );
  NAND2_X1 U13686 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12085) );
  INV_X1 U13687 ( .A(n12085), .ZN(n12063) );
  AND2_X1 U13688 ( .A1(n12058), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12092) );
  INV_X1 U13689 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12060) );
  XNOR2_X1 U13690 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16318) );
  AOI21_X1 U13691 ( .B1(n13548), .B2(n16318), .A(n13552), .ZN(n12059) );
  OAI21_X1 U13692 ( .B1(n12405), .B2(n12060), .A(n12059), .ZN(n12061) );
  AOI21_X1 U13693 ( .B1(n12092), .B2(n17687), .A(n12061), .ZN(n12062) );
  OR2_X1 U13694 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U13696 ( .A1(n14479), .A2(n12239), .ZN(n12073) );
  INV_X1 U13697 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12070) );
  INV_X1 U13698 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12069) );
  OAI22_X1 U13699 ( .A1(n12405), .A2(n12070), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12069), .ZN(n12071) );
  AOI21_X1 U13700 ( .B1(n12092), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12071), .ZN(n12072) );
  NAND2_X1 U13701 ( .A1(n12073), .A2(n12072), .ZN(n14619) );
  NAND2_X1 U13702 ( .A1(n12075), .A2(n12076), .ZN(n12077) );
  NAND2_X1 U13703 ( .A1(n12077), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14451) );
  INV_X1 U13704 ( .A(n12092), .ZN(n12102) );
  INV_X1 U13705 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14391) );
  NAND2_X1 U13706 ( .A1(n13553), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U13707 ( .A1(n22476), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12079) );
  OAI211_X1 U13708 ( .C1(n12102), .C2(n14391), .A(n12080), .B(n12079), .ZN(
        n12081) );
  AOI21_X1 U13709 ( .B1(n16804), .B2(n12239), .A(n12081), .ZN(n12082) );
  OR2_X1 U13710 ( .A1(n14451), .A2(n12082), .ZN(n14452) );
  INV_X1 U13711 ( .A(n12082), .ZN(n14453) );
  OR2_X1 U13712 ( .A1(n14453), .A2(n12400), .ZN(n12083) );
  NAND2_X1 U13713 ( .A1(n14452), .A2(n12083), .ZN(n14620) );
  NAND2_X1 U13714 ( .A1(n14619), .A2(n14620), .ZN(n14627) );
  OR2_X1 U13715 ( .A1(n14759), .A2(n12256), .ZN(n12094) );
  INV_X1 U13716 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12090) );
  INV_X1 U13717 ( .A(n12086), .ZN(n12088) );
  INV_X1 U13718 ( .A(n12087), .ZN(n12097) );
  OAI21_X1 U13719 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12088), .A(
        n12097), .ZN(n15002) );
  AOI22_X1 U13720 ( .A1(n13548), .A2(n15002), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12089) );
  OAI21_X1 U13721 ( .B1(n12405), .B2(n12090), .A(n12089), .ZN(n12091) );
  AOI21_X1 U13722 ( .B1(n12092), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12091), .ZN(n12093) );
  NAND2_X1 U13723 ( .A1(n14797), .A2(n14798), .ZN(n14757) );
  NAND2_X1 U13724 ( .A1(n12095), .A2(n12239), .ZN(n12105) );
  INV_X1 U13725 ( .A(n12096), .ZN(n12109) );
  INV_X1 U13726 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U13727 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND2_X1 U13728 ( .A1(n12109), .A2(n12099), .ZN(n22067) );
  INV_X1 U13729 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22223) );
  OAI21_X1 U13730 ( .B1(n22223), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22476), .ZN(n12101) );
  NAND2_X1 U13731 ( .A1(n13553), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12100) );
  OAI211_X1 U13732 ( .C1(n12102), .C2(n17696), .A(n12101), .B(n12100), .ZN(
        n12103) );
  OAI21_X1 U13733 ( .B1(n12400), .B2(n22067), .A(n12103), .ZN(n12104) );
  NAND2_X1 U13734 ( .A1(n12106), .A2(n12239), .ZN(n12114) );
  INV_X1 U13735 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14869) );
  INV_X1 U13736 ( .A(n12107), .ZN(n12118) );
  INV_X1 U13737 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U13738 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  NAND2_X1 U13739 ( .A1(n12118), .A2(n12110), .ZN(n20573) );
  AOI22_X1 U13740 ( .A1(n20573), .A2(n13548), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12111) );
  OAI21_X1 U13741 ( .B1(n12405), .B2(n14869), .A(n12111), .ZN(n12112) );
  INV_X1 U13742 ( .A(n12112), .ZN(n12113) );
  NAND2_X1 U13743 ( .A1(n12114), .A2(n12113), .ZN(n14867) );
  NAND2_X1 U13744 ( .A1(n12115), .A2(n12239), .ZN(n12125) );
  INV_X1 U13745 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12122) );
  INV_X1 U13746 ( .A(n12116), .ZN(n12120) );
  INV_X1 U13747 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U13748 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U13749 ( .A1(n12120), .A2(n12119), .ZN(n20582) );
  AOI22_X1 U13750 ( .A1(n20582), .A2(n12312), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12121) );
  OAI21_X1 U13751 ( .B1(n12405), .B2(n12122), .A(n12121), .ZN(n12123) );
  INV_X1 U13752 ( .A(n12123), .ZN(n12124) );
  NAND2_X1 U13753 ( .A1(n12125), .A2(n12124), .ZN(n14931) );
  XNOR2_X1 U13754 ( .A(n12127), .B(n12128), .ZN(n15885) );
  NAND2_X1 U13755 ( .A1(n15885), .A2(n12312), .ZN(n12145) );
  INV_X1 U13756 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15134) );
  OAI22_X1 U13757 ( .A1(n12405), .A2(n15134), .B1(n12129), .B2(n12128), .ZN(
        n12130) );
  INV_X1 U13758 ( .A(n12130), .ZN(n12143) );
  AOI22_X1 U13759 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U13760 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13761 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U13762 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U13763 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12141) );
  AOI22_X1 U13764 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U13765 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U13766 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U13767 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U13768 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  OAI21_X1 U13769 ( .B1(n12141), .B2(n12140), .A(n12239), .ZN(n12142) );
  AND2_X1 U13770 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  NAND2_X1 U13771 ( .A1(n12145), .A2(n12144), .ZN(n15103) );
  INV_X1 U13772 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15696) );
  OAI21_X1 U13773 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12147), .A(
        n12146), .ZN(n20595) );
  AOI22_X1 U13774 ( .A1(n13548), .A2(n20595), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12148) );
  OAI21_X1 U13775 ( .B1(n12405), .B2(n15696), .A(n12148), .ZN(n15695) );
  AOI22_X1 U13776 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13777 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U13778 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U13779 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12149) );
  NAND4_X1 U13780 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12158) );
  AOI22_X1 U13781 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U13782 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U13783 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13784 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U13785 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  OR2_X1 U13786 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  NAND2_X1 U13787 ( .A1(n12239), .A2(n12159), .ZN(n15856) );
  NAND2_X1 U13788 ( .A1(n15100), .A2(n12160), .ZN(n12161) );
  XOR2_X1 U13789 ( .A(n15753), .B(n12162), .Z(n20622) );
  INV_X1 U13790 ( .A(n20622), .ZN(n12177) );
  AOI22_X1 U13791 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U13792 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U13793 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U13794 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U13795 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12172) );
  AOI22_X1 U13796 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U13797 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U13798 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U13799 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U13800 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  NOR2_X1 U13801 ( .A1(n12172), .A2(n12171), .ZN(n12175) );
  NAND2_X1 U13802 ( .A1(n13553), .A2(P1_EAX_REG_17__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U13803 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12173) );
  OAI211_X1 U13804 ( .C1(n12397), .C2(n12175), .A(n12174), .B(n12173), .ZN(
        n12176) );
  AOI21_X1 U13805 ( .B1(n12177), .B2(n12312), .A(n12176), .ZN(n15740) );
  INV_X1 U13806 ( .A(n15740), .ZN(n12261) );
  INV_X1 U13807 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12178) );
  XNOR2_X1 U13808 ( .A(n12179), .B(n12178), .ZN(n22117) );
  AOI22_X1 U13809 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U13810 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U13811 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U13812 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U13813 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12189) );
  AOI22_X1 U13814 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13815 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U13816 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U13817 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12184) );
  NAND4_X1 U13818 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12188) );
  OR2_X1 U13819 ( .A1(n12189), .A2(n12188), .ZN(n12193) );
  INV_X1 U13820 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12191) );
  OAI21_X1 U13821 ( .B1(n22223), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n22476), .ZN(n12190) );
  OAI21_X1 U13822 ( .B1(n12405), .B2(n12191), .A(n12190), .ZN(n12192) );
  AOI21_X1 U13823 ( .B1(n13545), .B2(n12193), .A(n12192), .ZN(n12194) );
  AOI21_X1 U13824 ( .B1(n22117), .B2(n12312), .A(n12194), .ZN(n15724) );
  XOR2_X1 U13825 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12195), .Z(
        n20610) );
  INV_X1 U13826 ( .A(n20610), .ZN(n15800) );
  AOI22_X1 U13827 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U13828 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U13829 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U13830 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U13831 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12205) );
  AOI22_X1 U13832 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U13833 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U13834 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13835 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U13836 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12204) );
  NOR2_X1 U13837 ( .A1(n12205), .A2(n12204), .ZN(n12208) );
  NAND2_X1 U13838 ( .A1(n13553), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U13839 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12206) );
  OAI211_X1 U13840 ( .C1(n12256), .C2(n12208), .A(n12207), .B(n12206), .ZN(
        n12209) );
  AOI21_X1 U13841 ( .B1(n15800), .B2(n12312), .A(n12209), .ZN(n15796) );
  INV_X1 U13842 ( .A(n15796), .ZN(n12260) );
  XNOR2_X1 U13843 ( .A(n12210), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n22108) );
  AOI22_X1 U13844 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U13845 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U13846 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U13847 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U13848 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12220) );
  AOI22_X1 U13849 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U13850 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U13851 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U13852 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U13853 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  NOR2_X1 U13854 ( .A1(n12220), .A2(n12219), .ZN(n12223) );
  NAND2_X1 U13855 ( .A1(n13553), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U13856 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12221) );
  OAI211_X1 U13857 ( .C1(n12256), .C2(n12223), .A(n12222), .B(n12221), .ZN(
        n12224) );
  AOI21_X1 U13858 ( .B1(n22108), .B2(n12312), .A(n12224), .ZN(n15792) );
  INV_X1 U13859 ( .A(n15792), .ZN(n12259) );
  XOR2_X1 U13860 ( .A(n12226), .B(n12225), .Z(n15979) );
  AOI22_X1 U13861 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U13862 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U13863 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U13864 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U13865 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12237) );
  AOI22_X1 U13866 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12231), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U13867 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U13868 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U13869 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U13870 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12236) );
  OR2_X1 U13871 ( .A1(n12237), .A2(n12236), .ZN(n12238) );
  AOI22_X1 U13872 ( .A1(n12239), .A2(n12238), .B1(n13552), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U13873 ( .A1(n13553), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12240) );
  OAI211_X1 U13874 ( .C1(n15979), .C2(n12400), .A(n12241), .B(n12240), .ZN(
        n15892) );
  XOR2_X1 U13875 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12242), .Z(
        n22099) );
  AOI22_X1 U13876 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U13877 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U13878 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U13879 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11478), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U13880 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12252) );
  AOI22_X1 U13881 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12333), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13882 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11180), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U13883 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U13884 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12247) );
  NAND4_X1 U13885 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12251) );
  NOR2_X1 U13886 ( .A1(n12252), .A2(n12251), .ZN(n12255) );
  NAND2_X1 U13887 ( .A1(n13553), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U13888 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12253) );
  OAI211_X1 U13889 ( .C1(n12256), .C2(n12255), .A(n12254), .B(n12253), .ZN(
        n12257) );
  INV_X1 U13890 ( .A(n12257), .ZN(n12258) );
  OAI21_X1 U13891 ( .B1(n22099), .B2(n12400), .A(n12258), .ZN(n15858) );
  AND2_X1 U13892 ( .A1(n15892), .A2(n15858), .ZN(n15788) );
  AND2_X1 U13893 ( .A1(n12259), .A2(n15788), .ZN(n15789) );
  NAND2_X1 U13894 ( .A1(n15721), .A2(n12262), .ZN(n15739) );
  INV_X1 U13895 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15996) );
  XNOR2_X1 U13896 ( .A(n12263), .B(n15996), .ZN(n22129) );
  NAND2_X1 U13897 ( .A1(n22129), .A2(n12312), .ZN(n12278) );
  AOI22_X1 U13898 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U13899 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U13900 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U13901 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U13902 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12273) );
  AOI22_X1 U13903 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U13904 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U13905 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U13906 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12268) );
  NAND4_X1 U13907 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  NOR2_X1 U13908 ( .A1(n12273), .A2(n12272), .ZN(n12276) );
  AOI21_X1 U13909 ( .B1(n15996), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12274) );
  AOI21_X1 U13910 ( .B1(n13553), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12274), .ZN(
        n12275) );
  OAI21_X1 U13911 ( .B1(n12397), .B2(n12276), .A(n12275), .ZN(n12277) );
  NAND2_X1 U13912 ( .A1(n12278), .A2(n12277), .ZN(n15821) );
  AOI22_X1 U13913 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U13914 ( .A1(n11443), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U13915 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13528), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U13916 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12280) );
  NAND4_X1 U13917 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12289) );
  AOI22_X1 U13918 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U13919 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U13920 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U13921 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U13922 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  NOR2_X1 U13923 ( .A1(n12289), .A2(n12288), .ZN(n12293) );
  INV_X1 U13924 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n22316) );
  OAI21_X1 U13925 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n22223), .A(
        n22476), .ZN(n12290) );
  OAI21_X1 U13926 ( .B1(n12405), .B2(n22316), .A(n12290), .ZN(n12291) );
  INV_X1 U13927 ( .A(n12291), .ZN(n12292) );
  OAI21_X1 U13928 ( .B1(n12397), .B2(n12293), .A(n12292), .ZN(n12296) );
  OAI21_X1 U13929 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12294), .A(
        n12311), .ZN(n22142) );
  OR2_X1 U13930 ( .A1(n12400), .A2(n22142), .ZN(n12295) );
  AOI22_X1 U13931 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11443), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U13932 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11516), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U13933 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U13934 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U13935 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12306) );
  AOI22_X1 U13936 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13536), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U13937 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U13938 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U13939 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U13940 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12305) );
  NOR2_X1 U13941 ( .A1(n12306), .A2(n12305), .ZN(n12310) );
  INV_X1 U13942 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n22321) );
  NAND2_X1 U13943 ( .A1(n22476), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12307) );
  OAI211_X1 U13944 ( .C1(n12405), .C2(n22321), .A(n12400), .B(n12307), .ZN(
        n12308) );
  INV_X1 U13945 ( .A(n12308), .ZN(n12309) );
  OAI21_X1 U13946 ( .B1(n12397), .B2(n12310), .A(n12309), .ZN(n12314) );
  XNOR2_X1 U13947 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12311), .ZN(
        n22161) );
  NAND2_X1 U13948 ( .A1(n22161), .A2(n12312), .ZN(n12313) );
  NAND2_X1 U13949 ( .A1(n15920), .A2(n15924), .ZN(n15922) );
  AOI22_X1 U13950 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U13951 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U13952 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U13953 ( .A1(n11457), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12315) );
  NAND4_X1 U13954 ( .A1(n12318), .A2(n12317), .A3(n12316), .A4(n12315), .ZN(
        n12324) );
  AOI22_X1 U13955 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U13956 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U13957 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U13958 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U13959 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12323) );
  NOR2_X1 U13960 ( .A1(n12324), .A2(n12323), .ZN(n12328) );
  INV_X1 U13961 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n22327) );
  NAND2_X1 U13962 ( .A1(n22476), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12325) );
  OAI211_X1 U13963 ( .C1(n12405), .C2(n22327), .A(n12400), .B(n12325), .ZN(
        n12326) );
  INV_X1 U13964 ( .A(n12326), .ZN(n12327) );
  OAI21_X1 U13965 ( .B1(n12397), .B2(n12328), .A(n12327), .ZN(n12331) );
  OAI21_X1 U13966 ( .B1(n12329), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n12348), .ZN(n22174) );
  OR2_X1 U13967 ( .A1(n22174), .A2(n12400), .ZN(n12330) );
  NAND2_X1 U13968 ( .A1(n12331), .A2(n12330), .ZN(n16002) );
  AOI22_X1 U13969 ( .A1(n13535), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11442), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U13970 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U13971 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U13972 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12335) );
  NAND4_X1 U13973 ( .A1(n12338), .A2(n12337), .A3(n12336), .A4(n12335), .ZN(
        n12344) );
  AOI22_X1 U13974 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U13975 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13530), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U13976 ( .A1(n13528), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U13977 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16824), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12339) );
  NAND4_X1 U13978 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12343) );
  NOR2_X1 U13979 ( .A1(n12344), .A2(n12343), .ZN(n12347) );
  OAI21_X1 U13980 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n16551), .A(n12400), 
        .ZN(n12345) );
  AOI21_X1 U13981 ( .B1(n13553), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12345), .ZN(
        n12346) );
  OAI21_X1 U13982 ( .B1(n12397), .B2(n12347), .A(n12346), .ZN(n12350) );
  XNOR2_X1 U13983 ( .A(n12348), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16550) );
  NAND2_X1 U13984 ( .A1(n16550), .A2(n13548), .ZN(n12349) );
  NAND2_X1 U13985 ( .A1(n12350), .A2(n12349), .ZN(n16544) );
  XNOR2_X1 U13986 ( .A(n12352), .B(n12351), .ZN(n12356) );
  INV_X1 U13987 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n22337) );
  OAI21_X1 U13988 ( .B1(n22223), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n22476), .ZN(n12353) );
  OAI21_X1 U13989 ( .B1(n12405), .B2(n22337), .A(n12353), .ZN(n12354) );
  INV_X1 U13990 ( .A(n12354), .ZN(n12355) );
  OAI21_X1 U13991 ( .B1(n12397), .B2(n12356), .A(n12355), .ZN(n12361) );
  INV_X1 U13992 ( .A(n12357), .ZN(n12358) );
  INV_X1 U13993 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n22176) );
  NAND2_X1 U13994 ( .A1(n12358), .A2(n22176), .ZN(n12359) );
  NAND2_X1 U13995 ( .A1(n12368), .A2(n12359), .ZN(n22187) );
  INV_X1 U13996 ( .A(n12362), .ZN(n12363) );
  XNOR2_X1 U13997 ( .A(n12364), .B(n12363), .ZN(n12365) );
  NAND2_X1 U13998 ( .A1(n12365), .A2(n13545), .ZN(n12371) );
  INV_X1 U13999 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n22343) );
  NAND2_X1 U14000 ( .A1(n22476), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12366) );
  OAI211_X1 U14001 ( .C1(n12405), .C2(n22343), .A(n12400), .B(n12366), .ZN(
        n12367) );
  INV_X1 U14002 ( .A(n12367), .ZN(n12370) );
  XNOR2_X1 U14003 ( .A(n12368), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n22196) );
  AOI21_X1 U14004 ( .B1(n12371), .B2(n12370), .A(n12369), .ZN(n16569) );
  INV_X1 U14005 ( .A(n12372), .ZN(n12374) );
  INV_X1 U14006 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U14007 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  NAND2_X1 U14008 ( .A1(n12382), .A2(n12375), .ZN(n16664) );
  XNOR2_X1 U14009 ( .A(n12377), .B(n12376), .ZN(n12380) );
  AOI21_X1 U14010 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n22476), .A(
        n13548), .ZN(n12379) );
  NAND2_X1 U14011 ( .A1(n13553), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12378) );
  OAI211_X1 U14012 ( .C1(n12380), .C2(n12397), .A(n12379), .B(n12378), .ZN(
        n12381) );
  OAI21_X1 U14013 ( .B1(n12400), .B2(n16664), .A(n12381), .ZN(n16532) );
  NOR2_X2 U14014 ( .A1(n16531), .A2(n16532), .ZN(n16514) );
  XNOR2_X1 U14015 ( .A(n12382), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16653) );
  XOR2_X1 U14016 ( .A(n12384), .B(n12383), .Z(n12387) );
  INV_X1 U14017 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n22356) );
  AOI21_X1 U14018 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n22476), .A(
        n13548), .ZN(n12385) );
  OAI21_X1 U14019 ( .B1(n12405), .B2(n22356), .A(n12385), .ZN(n12386) );
  AOI21_X1 U14020 ( .B1(n12387), .B2(n13545), .A(n12386), .ZN(n12388) );
  AOI21_X1 U14021 ( .B1(n13548), .B2(n16653), .A(n12388), .ZN(n16516) );
  NAND2_X1 U14022 ( .A1(n16514), .A2(n16516), .ZN(n16503) );
  INV_X1 U14023 ( .A(n12389), .ZN(n12391) );
  INV_X1 U14024 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12390) );
  NAND2_X1 U14025 ( .A1(n12391), .A2(n12390), .ZN(n12392) );
  NAND2_X1 U14026 ( .A1(n12401), .A2(n12392), .ZN(n16643) );
  XNOR2_X1 U14027 ( .A(n12394), .B(n12393), .ZN(n12398) );
  AOI21_X1 U14028 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22476), .A(
        n13548), .ZN(n12396) );
  NAND2_X1 U14029 ( .A1(n13553), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12395) );
  OAI211_X1 U14030 ( .C1(n12398), .C2(n12397), .A(n12396), .B(n12395), .ZN(
        n12399) );
  OAI21_X1 U14031 ( .B1(n12400), .B2(n16643), .A(n12399), .ZN(n16505) );
  NOR2_X2 U14032 ( .A1(n16503), .A2(n16505), .ZN(n16488) );
  XNOR2_X1 U14033 ( .A(n12401), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16492) );
  XOR2_X1 U14034 ( .A(n12403), .B(n12402), .Z(n12407) );
  INV_X1 U14035 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n22368) );
  AOI21_X1 U14036 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n22476), .A(
        n13548), .ZN(n12404) );
  OAI21_X1 U14037 ( .B1(n12405), .B2(n22368), .A(n12404), .ZN(n12406) );
  AOI21_X1 U14038 ( .B1(n12407), .B2(n13545), .A(n12406), .ZN(n12408) );
  AOI21_X1 U14039 ( .B1(n13548), .B2(n16492), .A(n12408), .ZN(n16491) );
  NAND2_X1 U14040 ( .A1(n16488), .A2(n16491), .ZN(n12409) );
  AOI21_X1 U14041 ( .B1(n12410), .B2(n16490), .A(n13585), .ZN(n16479) );
  NAND3_X1 U14042 ( .A1(n22210), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17723) );
  INV_X1 U14043 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22211) );
  NAND2_X1 U14044 ( .A1(n12411), .A2(n22465), .ZN(n21904) );
  NAND2_X1 U14045 ( .A1(n21904), .A2(n22210), .ZN(n12412) );
  NAND2_X1 U14046 ( .A1(n22210), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17720) );
  NAND2_X1 U14047 ( .A1(n22223), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12413) );
  AND2_X1 U14048 ( .A1(n17720), .A2(n12413), .ZN(n14456) );
  AOI21_X1 U14049 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12414), .ZN(n12415) );
  OAI21_X1 U14050 ( .B1(n20633), .B2(n16484), .A(n12415), .ZN(n12416) );
  AOI21_X1 U14051 ( .B1(n16479), .B2(n20628), .A(n12416), .ZN(n12417) );
  OAI21_X1 U14052 ( .B1(n12418), .B2(n22203), .A(n12417), .ZN(P1_U2970) );
  INV_X1 U14053 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12667) );
  NAND2_X2 U14054 ( .A1(n12663), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13707) );
  AOI22_X1 U14055 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12425) );
  AND2_X4 U14056 ( .A1(n12664), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12673) );
  INV_X2 U14057 ( .A(n13705), .ZN(n13945) );
  AOI22_X1 U14058 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12673), .B1(
        n13945), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12424) );
  AND2_X4 U14059 ( .A1(n12664), .A2(n17630), .ZN(n13615) );
  NAND2_X2 U14060 ( .A1(n12660), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12459) );
  INV_X2 U14061 ( .A(n12459), .ZN(n12503) );
  AOI22_X1 U14062 ( .A1(n13615), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12423) );
  NAND2_X2 U14063 ( .A1(n12659), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13715) );
  INV_X4 U14064 ( .A(n13715), .ZN(n13672) );
  NOR2_X2 U14065 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12421) );
  AND2_X4 U14066 ( .A1(n12421), .A2(n12945), .ZN(n13952) );
  AOI22_X1 U14067 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12422) );
  NAND4_X1 U14068 ( .A1(n12425), .A2(n12424), .A3(n12423), .A4(n12422), .ZN(
        n12426) );
  INV_X2 U14069 ( .A(n13713), .ZN(n12514) );
  AOI22_X1 U14070 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12427) );
  NAND3_X1 U14071 ( .A1(n12429), .A2(n12428), .A3(n12427), .ZN(n12432) );
  INV_X2 U14072 ( .A(n13707), .ZN(n12521) );
  INV_X1 U14073 ( .A(n12430), .ZN(n12431) );
  OAI21_X2 U14074 ( .B1(n12432), .B2(n12431), .A(n12519), .ZN(n12433) );
  AOI22_X1 U14075 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U14076 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U14077 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U14078 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  AOI22_X1 U14079 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U14080 ( .A1(n13615), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12440) );
  NAND4_X1 U14081 ( .A1(n12443), .A2(n12442), .A3(n12441), .A4(n12440), .ZN(
        n12444) );
  NAND2_X2 U14082 ( .A1(n12446), .A2(n12445), .ZN(n12564) );
  AOI22_X1 U14083 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U14084 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U14085 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U14086 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U14087 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12451) );
  NAND2_X1 U14088 ( .A1(n12451), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12458) );
  AOI22_X1 U14089 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U14090 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U14091 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U14092 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U14093 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12456) );
  AOI22_X1 U14094 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12461) );
  INV_X2 U14095 ( .A(n13715), .ZN(n13951) );
  AOI22_X1 U14096 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12460) );
  NAND3_X1 U14097 ( .A1(n12462), .A2(n12461), .A3(n12460), .ZN(n12465) );
  AOI22_X1 U14098 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12463) );
  INV_X1 U14099 ( .A(n12463), .ZN(n12464) );
  AOI22_X1 U14100 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14101 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U14102 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U14103 ( .A1(n13953), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U14104 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12470) );
  NAND2_X1 U14105 ( .A1(n12470), .A2(n12519), .ZN(n12471) );
  AOI22_X1 U14106 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U14107 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U14108 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U14109 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U14110 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12478) );
  NAND2_X1 U14111 ( .A1(n12478), .A2(n12519), .ZN(n12485) );
  AOI22_X1 U14112 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U14113 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U14114 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U14115 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12479) );
  NAND4_X1 U14116 ( .A1(n12482), .A2(n12481), .A3(n12480), .A4(n12479), .ZN(
        n12483) );
  NAND2_X1 U14117 ( .A1(n12483), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12484) );
  NAND2_X2 U14118 ( .A1(n12485), .A2(n12484), .ZN(n12569) );
  AOI22_X1 U14119 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U14120 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U14121 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U14122 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U14123 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  NAND2_X1 U14124 ( .A1(n12490), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12497) );
  AOI22_X1 U14125 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U14126 ( .A1(n11217), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U14127 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U14128 ( .A1(n13941), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U14129 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  NAND2_X1 U14130 ( .A1(n12495), .A2(n12519), .ZN(n12496) );
  AOI22_X1 U14131 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U14132 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U14133 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U14134 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12498) );
  NAND4_X1 U14135 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n12502) );
  AOI22_X1 U14136 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U14137 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14138 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U14139 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12504) );
  NAND4_X1 U14140 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12508) );
  NAND2_X1 U14141 ( .A1(n20179), .A2(n13300), .ZN(n12513) );
  INV_X1 U14142 ( .A(n12543), .ZN(n12512) );
  OAI21_X1 U14143 ( .B1(n12955), .B2(n12513), .A(n13250), .ZN(n13295) );
  AOI22_X1 U14144 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U14145 ( .A1(n13941), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U14146 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U14147 ( .A1(n13953), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12503), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12515) );
  NAND4_X1 U14148 ( .A1(n12518), .A2(n12517), .A3(n12516), .A4(n12515), .ZN(
        n12520) );
  AOI22_X1 U14149 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U14150 ( .A1(n12673), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13615), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U14151 ( .A1(n13941), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U14152 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12526) );
  NAND2_X1 U14153 ( .A1(n13230), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18853) );
  INV_X1 U14154 ( .A(n12564), .ZN(n12531) );
  NAND2_X1 U14155 ( .A1(n20081), .A2(n12533), .ZN(n12560) );
  OAI21_X1 U14156 ( .B1(n12534), .B2(n13232), .A(n12560), .ZN(n12535) );
  NAND2_X1 U14157 ( .A1(n12562), .A2(n12535), .ZN(n12536) );
  INV_X2 U14158 ( .A(n12565), .ZN(n20289) );
  NAND2_X1 U14159 ( .A1(n12536), .A2(n20289), .ZN(n13274) );
  INV_X1 U14160 ( .A(n13243), .ZN(n12537) );
  NAND2_X1 U14161 ( .A1(n12581), .A2(n20289), .ZN(n12538) );
  NAND2_X1 U14162 ( .A1(n13274), .A2(n12538), .ZN(n12539) );
  NAND2_X1 U14163 ( .A1(n12539), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12540) );
  AND2_X2 U14164 ( .A1(n12541), .A2(n12540), .ZN(n12577) );
  NAND2_X1 U14165 ( .A1(n12543), .A2(n12542), .ZN(n13236) );
  NAND2_X1 U14166 ( .A1(n12544), .A2(n14347), .ZN(n13262) );
  NAND2_X2 U14167 ( .A1(n13300), .A2(n12565), .ZN(n19189) );
  NAND2_X1 U14168 ( .A1(n12580), .A2(n12546), .ZN(n12545) );
  NAND2_X2 U14169 ( .A1(n12577), .A2(n12545), .ZN(n12608) );
  INV_X1 U14170 ( .A(n12546), .ZN(n12548) );
  NOR2_X2 U14171 ( .A1(n13232), .A2(n12564), .ZN(n13267) );
  INV_X1 U14172 ( .A(n13267), .ZN(n12547) );
  NOR2_X1 U14173 ( .A1(n12548), .A2(n12547), .ZN(n12550) );
  NAND3_X2 U14174 ( .A1(n12549), .A2(n13267), .A3(n14261), .ZN(n13277) );
  INV_X1 U14175 ( .A(n12567), .ZN(n13736) );
  NAND2_X1 U14176 ( .A1(n13301), .A2(n20289), .ZN(n12553) );
  INV_X1 U14177 ( .A(n12554), .ZN(n12555) );
  NOR2_X1 U14178 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U14179 ( .A1(n17629), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19222), .ZN(n12558) );
  NAND2_X1 U14180 ( .A1(n12559), .A2(n12558), .ZN(n12616) );
  NOR2_X1 U14181 ( .A1(n12560), .A2(n13230), .ZN(n12561) );
  NOR2_X1 U14182 ( .A1(n13300), .A2(n12563), .ZN(n13253) );
  NOR2_X1 U14183 ( .A1(n12565), .A2(n12564), .ZN(n12566) );
  NAND2_X1 U14184 ( .A1(n13253), .A2(n12566), .ZN(n13270) );
  NAND2_X1 U14185 ( .A1(n12567), .A2(n12568), .ZN(n13996) );
  INV_X1 U14186 ( .A(n12570), .ZN(n12571) );
  NAND2_X1 U14187 ( .A1(n14228), .A2(n13301), .ZN(n19217) );
  NAND3_X1 U14188 ( .A1(n12572), .A2(n12585), .A3(n19217), .ZN(n12573) );
  AND2_X2 U14189 ( .A1(n12573), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U14190 ( .A1(n12603), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12584) );
  INV_X1 U14191 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18862) );
  AND2_X1 U14192 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12574) );
  NOR2_X1 U14193 ( .A1(n19222), .A2(n12574), .ZN(n12576) );
  NAND2_X1 U14194 ( .A1(n12604), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12575) );
  OAI211_X1 U14195 ( .C1(n12605), .C2(n18862), .A(n12576), .B(n12575), .ZN(
        n12579) );
  INV_X1 U14196 ( .A(n12577), .ZN(n12578) );
  NOR2_X1 U14197 ( .A1(n12579), .A2(n12578), .ZN(n12583) );
  NAND3_X1 U14198 ( .A1(n12584), .A2(n12583), .A3(n12582), .ZN(n12617) );
  NAND2_X1 U14199 ( .A1(n12608), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12587) );
  NAND2_X2 U14200 ( .A1(n12585), .A2(n13294), .ZN(n19082) );
  AOI22_X2 U14201 ( .A1(n19082), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19222), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12586) );
  NAND2_X2 U14202 ( .A1(n12587), .A2(n12586), .ZN(n12621) );
  NAND2_X1 U14203 ( .A1(n12603), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12591) );
  NAND2_X1 U14204 ( .A1(n12971), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U14205 ( .A1(n12604), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12588) );
  NOR2_X2 U14206 ( .A1(n12621), .A2(n12592), .ZN(n12594) );
  INV_X1 U14207 ( .A(n12621), .ZN(n12593) );
  OAI22_X2 U14208 ( .A1(n12615), .A2(n12594), .B1(n12622), .B2(n12593), .ZN(
        n12611) );
  OAI21_X1 U14209 ( .B1(n19906), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17661), 
        .ZN(n12595) );
  INV_X1 U14210 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U14211 ( .A1(n12604), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U14212 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U14213 ( .A1(n12600), .A2(n12599), .ZN(n12602) );
  NAND2_X1 U14214 ( .A1(n12602), .A2(n12601), .ZN(n12612) );
  OR2_X2 U14215 ( .A1(n12611), .A2(n12612), .ZN(n12614) );
  NAND2_X2 U14216 ( .A1(n12614), .A2(n12602), .ZN(n12964) );
  INV_X1 U14217 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U14218 ( .A1(n16360), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12607) );
  NAND2_X1 U14219 ( .A1(n13028), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U14220 ( .A1(n11155), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12610) );
  NAND2_X1 U14221 ( .A1(n19222), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12609) );
  XNOR2_X2 U14222 ( .A(n12964), .B(n12962), .ZN(n13729) );
  INV_X2 U14223 ( .A(n13729), .ZN(n12643) );
  NAND2_X1 U14224 ( .A1(n12611), .A2(n12612), .ZN(n12613) );
  INV_X1 U14225 ( .A(n12616), .ZN(n12619) );
  INV_X1 U14226 ( .A(n12617), .ZN(n12618) );
  NAND2_X1 U14227 ( .A1(n12619), .A2(n12618), .ZN(n12620) );
  XNOR2_X1 U14228 ( .A(n12622), .B(n12621), .ZN(n12624) );
  INV_X1 U14229 ( .A(n12624), .ZN(n12635) );
  AND2_X1 U14230 ( .A1(n18865), .A2(n12635), .ZN(n12649) );
  INV_X1 U14231 ( .A(n12649), .ZN(n12646) );
  NOR2_X1 U14232 ( .A1(n17054), .A2(n12646), .ZN(n12623) );
  INV_X1 U14233 ( .A(n12638), .ZN(n12625) );
  NOR2_X1 U14234 ( .A1(n17054), .A2(n12625), .ZN(n12626) );
  NAND2_X2 U14235 ( .A1(n12643), .A2(n12626), .ZN(n19794) );
  INV_X1 U14236 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12627) );
  OAI22_X1 U14237 ( .A1(n12667), .A2(n12814), .B1(n19794), .B2(n12627), .ZN(
        n12633) );
  INV_X1 U14238 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12631) );
  AND2_X1 U14239 ( .A1(n17054), .A2(n12649), .ZN(n12628) );
  NAND2_X2 U14240 ( .A1(n12643), .A2(n12628), .ZN(n19772) );
  AND2_X1 U14241 ( .A1(n17054), .A2(n12638), .ZN(n12629) );
  NAND2_X1 U14242 ( .A1(n12643), .A2(n12629), .ZN(n12816) );
  INV_X1 U14243 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12630) );
  OAI22_X1 U14244 ( .A1(n12631), .A2(n19772), .B1(n12816), .B2(n12630), .ZN(
        n12632) );
  AND2_X2 U14245 ( .A1(n13729), .A2(n14411), .ZN(n12647) );
  XNOR2_X2 U14246 ( .A(n12635), .B(n12634), .ZN(n13741) );
  AND2_X2 U14247 ( .A1(n13729), .A2(n17054), .ZN(n12651) );
  AND2_X2 U14248 ( .A1(n12651), .A2(n12638), .ZN(n19850) );
  AOI22_X1 U14249 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19927), .B1(
        n19850), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12641) );
  INV_X1 U14250 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12636) );
  INV_X1 U14251 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13678) );
  INV_X1 U14252 ( .A(n12637), .ZN(n12640) );
  AND2_X2 U14253 ( .A1(n12647), .A2(n12638), .ZN(n19915) );
  AND2_X1 U14254 ( .A1(n13741), .A2(n14399), .ZN(n12645) );
  AND2_X2 U14255 ( .A1(n12647), .A2(n12645), .ZN(n19962) );
  AOI22_X1 U14256 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19915), .B1(
        n19962), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12639) );
  NOR2_X1 U14257 ( .A1(n12654), .A2(n17595), .ZN(n12827) );
  NAND2_X1 U14258 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12658) );
  INV_X1 U14259 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20152) );
  NAND2_X2 U14260 ( .A1(n12647), .A2(n12649), .ZN(n19941) );
  INV_X1 U14261 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12661) );
  OAI22_X1 U14262 ( .A1(n20152), .A2(n19892), .B1(n19941), .B2(n12661), .ZN(
        n12648) );
  INV_X1 U14263 ( .A(n12648), .ZN(n12657) );
  NAND2_X1 U14264 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19877), .ZN(
        n12653) );
  NAND2_X1 U14265 ( .A1(n12813), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12652) );
  AND2_X1 U14266 ( .A1(n12653), .A2(n12652), .ZN(n12656) );
  NOR2_X1 U14267 ( .A1(n12654), .A2(n17621), .ZN(n12826) );
  NAND2_X1 U14268 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12655) );
  AND2_X4 U14269 ( .A1(n13940), .A2(n12519), .ZN(n13878) );
  NAND2_X1 U14270 ( .A1(n13616), .A2(n12659), .ZN(n13876) );
  OAI22_X1 U14271 ( .A1(n13876), .A2(n12661), .B1(n13874), .B2(n20152), .ZN(
        n12662) );
  AOI21_X1 U14272 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n12662), .ZN(n12672) );
  AND2_X2 U14273 ( .A1(n13941), .A2(n12519), .ZN(n13879) );
  AND2_X2 U14274 ( .A1(n13941), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12727) );
  AOI22_X1 U14275 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12671) );
  OR2_X2 U14276 ( .A1(n13720), .A2(n12519), .ZN(n13473) );
  NAND2_X1 U14277 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12666) );
  AND2_X2 U14278 ( .A1(n12664), .A2(n13616), .ZN(n13884) );
  NAND2_X1 U14279 ( .A1(n13884), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12665) );
  OAI211_X1 U14280 ( .C1(n12667), .C2(n13473), .A(n12666), .B(n12665), .ZN(
        n12668) );
  INV_X1 U14281 ( .A(n12668), .ZN(n12670) );
  NAND2_X1 U14282 ( .A1(n13462), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12669) );
  NAND4_X1 U14283 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12679) );
  AOI22_X1 U14284 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12677) );
  AND2_X2 U14285 ( .A1(n13945), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13847) );
  AOI22_X1 U14286 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12676) );
  BUF_X4 U14287 ( .A(n12673), .Z(n13955) );
  AOI22_X1 U14288 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12675) );
  NAND3_X1 U14289 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12925) );
  NOR2_X1 U14290 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12925), .ZN(
        n12805) );
  NAND2_X1 U14291 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12674) );
  NAND4_X1 U14292 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  INV_X1 U14293 ( .A(n13327), .ZN(n12680) );
  NAND2_X1 U14294 ( .A1(n12680), .A2(n20227), .ZN(n12681) );
  AOI22_X1 U14295 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19915), .B1(
        n12825), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U14296 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19877), .B1(
        n12813), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12682) );
  INV_X1 U14297 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12730) );
  NOR2_X1 U14298 ( .A1(n19762), .A2(n12730), .ZN(n12686) );
  INV_X1 U14299 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12684) );
  INV_X1 U14300 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U14301 ( .A1(n12684), .A2(n19772), .B1(n12816), .B2(n13370), .ZN(
        n12685) );
  NOR2_X1 U14302 ( .A1(n12686), .A2(n12685), .ZN(n12690) );
  INV_X1 U14303 ( .A(n19787), .ZN(n19783) );
  INV_X1 U14304 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12687) );
  INV_X1 U14305 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12692) );
  OR2_X1 U14306 ( .A1(n12814), .A2(n12692), .ZN(n12697) );
  INV_X1 U14307 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12693) );
  INV_X1 U14308 ( .A(n12694), .ZN(n12696) );
  NAND2_X1 U14309 ( .A1(n19850), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12695) );
  NAND2_X1 U14310 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12700) );
  NAND2_X1 U14311 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12699) );
  AOI22_X1 U14312 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U14313 ( .A1(n13470), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U14314 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12703) );
  INV_X4 U14315 ( .A(n13473), .ZN(n13885) );
  NAND2_X1 U14316 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12702) );
  NAND4_X1 U14317 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12710) );
  NAND2_X1 U14318 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12708) );
  NAND2_X1 U14319 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12707) );
  NAND2_X1 U14320 ( .A1(n13445), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12706) );
  NAND3_X1 U14321 ( .A1(n12708), .A2(n12707), .A3(n12706), .ZN(n12709) );
  NOR2_X1 U14322 ( .A1(n12710), .A2(n12709), .ZN(n12724) );
  NAND2_X1 U14323 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12716) );
  NAND2_X1 U14324 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12715) );
  NAND2_X1 U14325 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12714) );
  NAND2_X1 U14326 ( .A1(n12712), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12713) );
  NAND4_X1 U14327 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12722) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U14329 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12719) );
  INV_X1 U14330 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U14331 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12718) );
  OAI211_X1 U14332 ( .C1(n13882), .C2(n12720), .A(n12719), .B(n12718), .ZN(
        n12721) );
  NOR2_X1 U14333 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  INV_X1 U14334 ( .A(n13303), .ZN(n12762) );
  NOR2_X1 U14335 ( .A1(n12762), .A2(n19096), .ZN(n14338) );
  INV_X1 U14336 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12725) );
  OAI22_X1 U14337 ( .A1(n13876), .A2(n12725), .B1(n13874), .B2(n12687), .ZN(
        n12726) );
  AOI21_X1 U14338 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n12726), .ZN(n12735) );
  NAND2_X1 U14339 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12729) );
  NAND2_X1 U14340 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12728) );
  OAI211_X1 U14341 ( .C1(n13882), .C2(n12730), .A(n12729), .B(n12728), .ZN(
        n12731) );
  INV_X1 U14342 ( .A(n12731), .ZN(n12734) );
  AOI22_X1 U14343 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U14344 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12732) );
  NAND4_X1 U14345 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12742) );
  AOI22_X1 U14346 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14347 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U14348 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12738) );
  NAND2_X1 U14349 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12737) );
  NAND4_X1 U14350 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12737), .ZN(
        n12741) );
  NAND2_X1 U14351 ( .A1(n14338), .A2(n13315), .ZN(n12765) );
  INV_X1 U14352 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12743) );
  INV_X1 U14353 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13655) );
  OAI22_X1 U14354 ( .A1(n13876), .A2(n12743), .B1(n13874), .B2(n13655), .ZN(
        n12744) );
  AOI21_X1 U14355 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n12744), .ZN(n12752) );
  INV_X1 U14356 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U14357 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12746) );
  NAND2_X1 U14358 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12745) );
  OAI211_X1 U14359 ( .C1(n13882), .C2(n12747), .A(n12746), .B(n12745), .ZN(
        n12748) );
  INV_X1 U14360 ( .A(n12748), .ZN(n12751) );
  AOI22_X1 U14361 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U14362 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12749) );
  NAND4_X1 U14363 ( .A1(n12752), .A2(n12751), .A3(n12750), .A4(n12749), .ZN(
        n12759) );
  AOI22_X1 U14364 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U14365 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U14366 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U14367 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12754) );
  NAND4_X1 U14368 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12758) );
  OR2_X2 U14369 ( .A1(n12759), .A2(n12758), .ZN(n13042) );
  INV_X1 U14370 ( .A(n13042), .ZN(n12760) );
  NAND2_X1 U14371 ( .A1(n12765), .A2(n12760), .ZN(n12761) );
  INV_X1 U14372 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14408) );
  XNOR2_X1 U14373 ( .A(n12762), .B(n13315), .ZN(n12763) );
  INV_X1 U14374 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14339) );
  NAND2_X1 U14375 ( .A1(n12763), .A2(n11280), .ZN(n12764) );
  XOR2_X1 U14376 ( .A(n12763), .B(n11280), .Z(n14358) );
  NAND2_X1 U14377 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14358), .ZN(
        n14357) );
  NAND2_X1 U14378 ( .A1(n12764), .A2(n14357), .ZN(n12766) );
  XNOR2_X1 U14379 ( .A(n14408), .B(n12766), .ZN(n14368) );
  XOR2_X1 U14380 ( .A(n13042), .B(n12765), .Z(n14367) );
  NAND2_X1 U14381 ( .A1(n14368), .A2(n14367), .ZN(n14366) );
  NAND2_X1 U14382 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12766), .ZN(
        n12767) );
  NAND2_X1 U14383 ( .A1(n14366), .A2(n12767), .ZN(n12768) );
  XNOR2_X1 U14384 ( .A(n12768), .B(n15058), .ZN(n14873) );
  NAND2_X1 U14385 ( .A1(n14872), .A2(n14873), .ZN(n12770) );
  NAND2_X1 U14386 ( .A1(n12768), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12769) );
  INV_X1 U14387 ( .A(n12771), .ZN(n12773) );
  NAND2_X1 U14388 ( .A1(n12773), .A2(n12772), .ZN(n12795) );
  INV_X1 U14389 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12774) );
  INV_X1 U14390 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U14391 ( .A1(n13876), .A2(n12774), .B1(n13874), .B2(n13688), .ZN(
        n12775) );
  AOI21_X1 U14392 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n12775), .ZN(n12783) );
  AOI22_X1 U14393 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12782) );
  INV_X1 U14394 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12778) );
  NAND2_X1 U14395 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12777) );
  NAND2_X1 U14396 ( .A1(n13884), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12776) );
  OAI211_X1 U14397 ( .C1(n12778), .C2(n13473), .A(n12777), .B(n12776), .ZN(
        n12779) );
  INV_X1 U14398 ( .A(n12779), .ZN(n12781) );
  NAND2_X1 U14399 ( .A1(n13462), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12780) );
  NAND4_X1 U14400 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n12789) );
  AOI22_X1 U14401 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U14402 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U14403 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U14404 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12784) );
  NAND4_X1 U14405 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12788) );
  INV_X1 U14406 ( .A(n13330), .ZN(n12790) );
  XNOR2_X1 U14407 ( .A(n12795), .B(n12790), .ZN(n12792) );
  INV_X1 U14408 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15672) );
  INV_X1 U14409 ( .A(n12791), .ZN(n12793) );
  NAND2_X1 U14410 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  INV_X1 U14411 ( .A(n12795), .ZN(n12796) );
  AOI22_X1 U14412 ( .A1(n13470), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U14413 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U14414 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U14415 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12797) );
  NAND4_X1 U14416 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12804) );
  INV_X1 U14417 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13710) );
  NAND2_X1 U14418 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12802) );
  NAND2_X1 U14419 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12801) );
  OAI211_X1 U14420 ( .C1(n13882), .C2(n13710), .A(n12802), .B(n12801), .ZN(
        n12803) );
  NOR2_X1 U14421 ( .A1(n12804), .A2(n12803), .ZN(n12812) );
  AOI22_X1 U14422 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U14423 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13847), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12810) );
  INV_X1 U14424 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13712) );
  INV_X1 U14425 ( .A(n12805), .ZN(n13398) );
  NAND2_X1 U14426 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12807) );
  NAND2_X1 U14427 ( .A1(n12712), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12806) );
  OAI211_X1 U14428 ( .C1(n13712), .C2(n13398), .A(n12807), .B(n12806), .ZN(
        n12808) );
  INV_X1 U14429 ( .A(n12808), .ZN(n12809) );
  NAND4_X1 U14430 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12809), .ZN(
        n13335) );
  AOI22_X1 U14431 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19850), .B1(
        n19927), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U14432 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11191), .B1(
        n19860), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12823) );
  INV_X1 U14433 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12815) );
  INV_X1 U14434 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13706) );
  OAI22_X1 U14435 ( .A1(n12815), .A2(n19798), .B1(n19824), .B2(n13706), .ZN(
        n12818) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13704) );
  OAI22_X1 U14437 ( .A1(n13704), .A2(n19772), .B1(n19746), .B2(n13712), .ZN(
        n12817) );
  INV_X1 U14438 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12819) );
  OAI22_X1 U14439 ( .A1(n12819), .A2(n19787), .B1(n19762), .B2(n13710), .ZN(
        n12820) );
  INV_X1 U14440 ( .A(n12820), .ZN(n12821) );
  NAND4_X1 U14441 ( .A1(n12822), .A2(n12823), .A3(n12824), .A4(n12821), .ZN(
        n12833) );
  AOI22_X1 U14442 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19962), .B1(
        n19915), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19897), .B1(
        n12825), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U14444 ( .A1(n19808), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12829) );
  NAND2_X1 U14445 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12828) );
  NAND4_X1 U14446 ( .A1(n12831), .A2(n12830), .A3(n12829), .A4(n12828), .ZN(
        n12832) );
  OAI21_X1 U14447 ( .B1(n19096), .B2(n13335), .A(n12834), .ZN(n12835) );
  INV_X1 U14448 ( .A(n12835), .ZN(n12838) );
  INV_X1 U14449 ( .A(n12836), .ZN(n12877) );
  NAND2_X1 U14450 ( .A1(n12887), .A2(n11182), .ZN(n12876) );
  INV_X1 U14451 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11191), .B1(
        n19860), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U14453 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19927), .B1(
        n19897), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12848) );
  INV_X1 U14454 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12839) );
  INV_X1 U14455 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13929) );
  OAI22_X1 U14456 ( .A1(n12839), .A2(n19824), .B1(n19798), .B2(n13929), .ZN(
        n12843) );
  INV_X1 U14457 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12841) );
  INV_X1 U14458 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12840) );
  OAI22_X1 U14459 ( .A1(n12841), .A2(n19772), .B1(n19746), .B2(n12840), .ZN(
        n12842) );
  NOR2_X1 U14460 ( .A1(n12843), .A2(n12842), .ZN(n12847) );
  INV_X1 U14461 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12861) );
  INV_X1 U14462 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12844) );
  OAI22_X1 U14463 ( .A1(n12861), .A2(n19762), .B1(n19787), .B2(n12844), .ZN(
        n12845) );
  INV_X1 U14464 ( .A(n12845), .ZN(n12846) );
  NAND4_X1 U14465 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n12846), .ZN(
        n12855) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19962), .B1(
        n19850), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U14467 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19915), .B1(
        n12825), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U14468 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U14469 ( .A1(n19808), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12850) );
  NAND4_X1 U14470 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12854) );
  INV_X1 U14471 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12857) );
  INV_X1 U14472 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12856) );
  OAI22_X1 U14473 ( .A1(n13876), .A2(n12857), .B1(n13874), .B2(n12856), .ZN(
        n12858) );
  AOI21_X1 U14474 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n12858), .ZN(n12866) );
  NAND2_X1 U14475 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U14476 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12859) );
  OAI211_X1 U14477 ( .C1(n13882), .C2(n12861), .A(n12860), .B(n12859), .ZN(
        n12862) );
  INV_X1 U14478 ( .A(n12862), .ZN(n12865) );
  AOI22_X1 U14479 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U14480 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12863) );
  NAND4_X1 U14481 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12872) );
  AOI22_X1 U14482 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U14483 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U14484 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U14485 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12867) );
  NAND4_X1 U14486 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n12867), .ZN(
        n12871) );
  NAND2_X1 U14487 ( .A1(n13084), .A2(n20227), .ZN(n12873) );
  NAND2_X1 U14489 ( .A1(n12876), .A2(n12875), .ZN(n12883) );
  AND2_X1 U14490 ( .A1(n12877), .A2(n15664), .ZN(n12878) );
  OR2_X1 U14491 ( .A1(n11182), .A2(n12878), .ZN(n12881) );
  NAND2_X1 U14492 ( .A1(n12883), .A2(n12882), .ZN(n12886) );
  INV_X1 U14493 ( .A(n12894), .ZN(n12884) );
  NAND3_X1 U14494 ( .A1(n12836), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n12884), .ZN(n12885) );
  NAND2_X1 U14495 ( .A1(n15761), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12892) );
  BUF_X1 U14496 ( .A(n12887), .Z(n15665) );
  OAI21_X1 U14497 ( .B1(n15665), .B2(n15664), .A(n12888), .ZN(n12890) );
  NAND2_X1 U14498 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  NAND2_X1 U14499 ( .A1(n12892), .A2(n12891), .ZN(n17340) );
  AOI22_X1 U14500 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13470), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13467), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12898) );
  NAND2_X1 U14502 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U14503 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12896) );
  NAND2_X1 U14504 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12903) );
  NAND2_X1 U14505 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12902) );
  NAND2_X1 U14506 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12901) );
  NAND2_X1 U14507 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12900) );
  INV_X1 U14508 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U14509 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12905) );
  NAND2_X1 U14510 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12904) );
  OAI211_X1 U14511 ( .C1(n13882), .C2(n12906), .A(n12905), .B(n12904), .ZN(
        n12907) );
  INV_X1 U14512 ( .A(n12907), .ZN(n12912) );
  NAND2_X1 U14513 ( .A1(n13890), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12910) );
  NAND2_X1 U14514 ( .A1(n12712), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12909) );
  NAND2_X1 U14515 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12908) );
  AND3_X1 U14516 ( .A1(n12910), .A2(n12909), .A3(n12908), .ZN(n12911) );
  NAND2_X1 U14517 ( .A1(n12914), .A2(n13093), .ZN(n12915) );
  INV_X1 U14518 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17581) );
  NOR2_X1 U14519 ( .A1(n17341), .A2(n17581), .ZN(n12916) );
  NAND2_X1 U14520 ( .A1(n17341), .A2(n17581), .ZN(n12917) );
  OAI21_X1 U14521 ( .B1(n17340), .B2(n12916), .A(n12917), .ZN(n12918) );
  NAND2_X1 U14522 ( .A1(n17747), .A2(n17746), .ZN(n17745) );
  INV_X1 U14523 ( .A(n12919), .ZN(n12920) );
  NAND2_X1 U14524 ( .A1(n12920), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12921) );
  INV_X1 U14525 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17533) );
  INV_X1 U14526 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17573) );
  INV_X1 U14527 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17546) );
  NOR3_X1 U14528 ( .A1(n17533), .A2(n17573), .A3(n17546), .ZN(n17498) );
  NAND4_X1 U14529 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n17498), .ZN(n13292) );
  INV_X1 U14530 ( .A(n13292), .ZN(n13514) );
  INV_X1 U14531 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17473) );
  NAND2_X1 U14532 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12922) );
  NAND2_X2 U14533 ( .A1(n17797), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17796) );
  INV_X1 U14534 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17437) );
  NOR2_X2 U14535 ( .A1(n17796), .A2(n17437), .ZN(n17296) );
  OR2_X1 U14536 ( .A1(n17296), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12924) );
  INV_X1 U14537 ( .A(n17472), .ZN(n12923) );
  AND2_X1 U14538 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16226) );
  NOR2_X1 U14539 ( .A1(n17473), .A2(n12922), .ZN(n13293) );
  AND2_X1 U14540 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n13293), .ZN(
        n13513) );
  AND2_X2 U14541 ( .A1(n12924), .A2(n17285), .ZN(n13524) );
  AND2_X1 U14542 ( .A1(n12925), .A2(n19101), .ZN(n19095) );
  NAND2_X1 U14543 ( .A1(n13882), .A2(n19095), .ZN(n12927) );
  INV_X1 U14544 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12926) );
  NAND2_X1 U14545 ( .A1(n12927), .A2(n12926), .ZN(n17829) );
  XNOR2_X1 U14546 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U14547 ( .A1(n12951), .A2(n12940), .ZN(n12942) );
  NAND2_X1 U14548 ( .A1(n19910), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U14549 ( .A1(n12942), .A2(n12928), .ZN(n12939) );
  XNOR2_X1 U14550 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U14551 ( .A1(n12939), .A2(n12937), .ZN(n12930) );
  NAND2_X1 U14552 ( .A1(n19906), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12929) );
  NOR2_X1 U14553 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19181), .ZN(
        n12933) );
  NAND3_X1 U14554 ( .A1(n12934), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n19101), .ZN(n13207) );
  XNOR2_X1 U14555 ( .A(n12936), .B(n12935), .ZN(n13222) );
  INV_X1 U14556 ( .A(n12937), .ZN(n12938) );
  XNOR2_X1 U14557 ( .A(n12939), .B(n12938), .ZN(n13210) );
  AND2_X1 U14558 ( .A1(n13222), .A2(n13210), .ZN(n12948) );
  INV_X1 U14559 ( .A(n12951), .ZN(n12941) );
  INV_X1 U14560 ( .A(n12940), .ZN(n12947) );
  NAND2_X1 U14561 ( .A1(n12941), .A2(n12947), .ZN(n12943) );
  AND2_X1 U14562 ( .A1(n12943), .A2(n12942), .ZN(n13211) );
  AND3_X1 U14563 ( .A1(n13207), .A2(n12948), .A3(n13211), .ZN(n12944) );
  OR2_X1 U14564 ( .A1(n13228), .A2(n12944), .ZN(n19193) );
  NAND2_X1 U14565 ( .A1(n12945), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12946) );
  AND3_X1 U14566 ( .A1(n13207), .A2(n13212), .A3(n12948), .ZN(n12949) );
  NOR2_X1 U14567 ( .A1(n19193), .A2(n12949), .ZN(n12950) );
  MUX2_X1 U14568 ( .A(n17829), .B(n12950), .S(n17661), .Z(n19242) );
  NAND2_X1 U14569 ( .A1(n19242), .A2(n14261), .ZN(n12954) );
  MUX2_X1 U14570 ( .A(n13207), .B(n13330), .S(n14261), .Z(n13064) );
  MUX2_X1 U14571 ( .A(n13327), .B(n13222), .S(n19189), .Z(n13049) );
  NAND2_X1 U14572 ( .A1(n13064), .A2(n13049), .ZN(n13224) );
  NAND2_X1 U14573 ( .A1(n19189), .A2(n13210), .ZN(n13209) );
  NAND2_X1 U14574 ( .A1(n13212), .A2(n12951), .ZN(n13216) );
  AND2_X1 U14575 ( .A1(n13209), .A2(n13216), .ZN(n12952) );
  NOR2_X1 U14576 ( .A1(n13224), .A2(n12952), .ZN(n12953) );
  NOR2_X1 U14577 ( .A1(n12953), .A2(n13228), .ZN(n19188) );
  AND2_X1 U14578 ( .A1(n20227), .A2(n13230), .ZN(n19186) );
  NAND2_X1 U14579 ( .A1(n19188), .A2(n19186), .ZN(n13233) );
  NAND2_X1 U14580 ( .A1(n12954), .A2(n13233), .ZN(n12956) );
  NAND2_X1 U14581 ( .A1(n12956), .A2(n19190), .ZN(n19205) );
  NAND3_X1 U14582 ( .A1(n17661), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19247) );
  NAND2_X1 U14583 ( .A1(n13524), .A2(n17820), .ZN(n13041) );
  NAND2_X1 U14584 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17668) );
  INV_X1 U14585 ( .A(n17668), .ZN(n12957) );
  NOR2_X1 U14586 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n12957), .ZN(n17828) );
  NAND2_X1 U14587 ( .A1(n17828), .A2(n19237), .ZN(n12958) );
  AND2_X1 U14588 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12959) );
  INV_X1 U14589 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U14590 ( .A1(n11221), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12961) );
  NAND2_X1 U14591 ( .A1(n13028), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12960) );
  OAI211_X1 U14592 ( .C1(n12985), .C2(n13515), .A(n12961), .B(n12960), .ZN(
        n13033) );
  INV_X1 U14593 ( .A(n13033), .ZN(n13036) );
  INV_X1 U14594 ( .A(n12962), .ZN(n12963) );
  NAND2_X1 U14595 ( .A1(n12964), .A2(n12963), .ZN(n12970) );
  INV_X1 U14596 ( .A(n12965), .ZN(n12968) );
  INV_X1 U14597 ( .A(n12966), .ZN(n12967) );
  NAND2_X1 U14598 ( .A1(n12968), .A2(n12967), .ZN(n12969) );
  NAND2_X1 U14599 ( .A1(n12970), .A2(n12969), .ZN(n14430) );
  INV_X1 U14600 ( .A(n12985), .ZN(n12975) );
  INV_X1 U14601 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n13333) );
  NAND2_X1 U14602 ( .A1(n11221), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12973) );
  NAND2_X1 U14603 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12972) );
  OAI211_X1 U14604 ( .C1(n16236), .C2(n13333), .A(n12973), .B(n12972), .ZN(
        n12974) );
  AOI21_X1 U14605 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12974), .ZN(n14429) );
  INV_X1 U14606 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U14607 ( .A1(n16401), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U14608 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12978) );
  OAI211_X1 U14609 ( .C1(n16236), .C2(n12980), .A(n12979), .B(n12978), .ZN(
        n12981) );
  AOI21_X1 U14610 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12981), .ZN(n14422) );
  NOR2_X2 U14611 ( .A1(n14432), .A2(n14422), .ZN(n14494) );
  INV_X1 U14612 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U14613 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12983) );
  AOI22_X1 U14614 ( .A1(n16401), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12982) );
  OAI211_X1 U14615 ( .C1(n16236), .C2(n12984), .A(n12983), .B(n12982), .ZN(
        n14493) );
  NAND2_X1 U14616 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  INV_X1 U14617 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17347) );
  NAND2_X1 U14618 ( .A1(n16401), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U14619 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12986) );
  OAI211_X1 U14620 ( .C1(n16236), .C2(n17347), .A(n12987), .B(n12986), .ZN(
        n12988) );
  AOI21_X1 U14621 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12988), .ZN(n14466) );
  NOR2_X2 U14622 ( .A1(n14495), .A2(n14466), .ZN(n14467) );
  NAND2_X1 U14623 ( .A1(n12975), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12993) );
  INV_X1 U14624 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13363) );
  NAND2_X1 U14625 ( .A1(n16401), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U14626 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12989) );
  OAI211_X1 U14627 ( .C1(n16236), .C2(n13363), .A(n12990), .B(n12989), .ZN(
        n12991) );
  INV_X1 U14628 ( .A(n12991), .ZN(n12992) );
  NAND2_X1 U14629 ( .A1(n12993), .A2(n12992), .ZN(n14601) );
  NAND2_X1 U14630 ( .A1(n14467), .A2(n14601), .ZN(n14750) );
  INV_X1 U14631 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U14632 ( .A1(n16401), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12995) );
  NAND2_X1 U14633 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12994) );
  OAI211_X1 U14634 ( .C1(n16236), .C2(n13384), .A(n12995), .B(n12994), .ZN(
        n12996) );
  AOI21_X1 U14635 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12996), .ZN(n14751) );
  INV_X1 U14636 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U14637 ( .A1(n11221), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U14638 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12999) );
  OAI211_X1 U14639 ( .C1(n16236), .C2(n13405), .A(n13000), .B(n12999), .ZN(
        n13001) );
  AOI21_X1 U14640 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n13001), .ZN(n14855) );
  INV_X1 U14641 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17322) );
  NAND2_X1 U14642 ( .A1(n12975), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13003) );
  AOI22_X1 U14643 ( .A1(n11221), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n13002) );
  OAI211_X1 U14644 ( .C1(n16236), .C2(n17322), .A(n13003), .B(n13002), .ZN(
        n14925) );
  INV_X1 U14645 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n13505) );
  NAND2_X1 U14646 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13005) );
  AOI22_X1 U14647 ( .A1(n16401), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n13004) );
  OAI211_X1 U14648 ( .C1(n16236), .C2(n13505), .A(n13005), .B(n13004), .ZN(
        n15706) );
  INV_X1 U14649 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U14650 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13007) );
  AOI22_X1 U14651 ( .A1(n16401), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n13006) );
  OAI211_X1 U14652 ( .C1(n16236), .C2(n13484), .A(n13007), .B(n13006), .ZN(
        n15654) );
  INV_X1 U14653 ( .A(n15654), .ZN(n13014) );
  INV_X1 U14654 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U14655 ( .A1(n16401), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U14656 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13008) );
  OAI211_X1 U14657 ( .C1(n16236), .C2(n13461), .A(n13009), .B(n13008), .ZN(
        n13010) );
  AOI21_X1 U14658 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n13010), .ZN(n15124) );
  INV_X1 U14659 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U14660 ( .A1(n16401), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U14661 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13011) );
  OAI211_X1 U14662 ( .C1(n16236), .C2(n13443), .A(n13012), .B(n13011), .ZN(
        n13013) );
  AOI21_X1 U14663 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n13013), .ZN(n13197) );
  OR2_X1 U14664 ( .A1(n15124), .A2(n13197), .ZN(n15126) );
  NOR2_X1 U14665 ( .A1(n13014), .A2(n15126), .ZN(n15652) );
  NAND2_X1 U14666 ( .A1(n15653), .A2(n13015), .ZN(n15704) );
  INV_X1 U14667 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n13018) );
  NAND2_X1 U14668 ( .A1(n11221), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U14669 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13016) );
  OAI211_X1 U14670 ( .C1(n16236), .C2(n13018), .A(n13017), .B(n13016), .ZN(
        n13019) );
  AOI21_X1 U14671 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n13019), .ZN(n15717) );
  INV_X1 U14672 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17457) );
  NAND2_X1 U14673 ( .A1(n16401), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13023) );
  NAND2_X1 U14674 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13022) );
  OAI211_X1 U14675 ( .C1(n16236), .C2(n17457), .A(n13023), .B(n13022), .ZN(
        n13024) );
  AOI21_X1 U14676 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13024), .ZN(n17129) );
  NOR2_X2 U14677 ( .A1(n15716), .A2(n17129), .ZN(n17131) );
  INV_X1 U14678 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U14679 ( .A1(n12975), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13026) );
  AOI22_X1 U14680 ( .A1(n11221), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n13025) );
  OAI211_X1 U14681 ( .C1(n16236), .C2(n13027), .A(n13026), .B(n13025), .ZN(
        n17121) );
  AND2_X2 U14682 ( .A1(n17131), .A2(n17121), .ZN(n17122) );
  NAND2_X1 U14683 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13032) );
  NAND2_X1 U14684 ( .A1(n13028), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14685 ( .A1(n16401), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n13029) );
  AND2_X1 U14686 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  NAND2_X1 U14687 ( .A1(n13032), .A2(n13031), .ZN(n17111) );
  INV_X1 U14688 ( .A(n13034), .ZN(n13035) );
  AND2_X2 U14689 ( .A1(n13034), .A2(n13033), .ZN(n14244) );
  AOI21_X1 U14690 ( .B1(n13036), .B2(n13035), .A(n14244), .ZN(n17103) );
  AND2_X1 U14691 ( .A1(n17807), .A2(n17103), .ZN(n13040) );
  NAND2_X1 U14692 ( .A1(n19237), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19215) );
  INV_X1 U14693 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22228) );
  NAND2_X1 U14694 ( .A1(n22228), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U14695 ( .A1(n19215), .A2(n13037), .ZN(n14341) );
  INV_X1 U14696 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17297) );
  INV_X1 U14697 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14203) );
  INV_X1 U14698 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17784) );
  OAI21_X1 U14699 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14204), .A(
        n14207), .ZN(n14179) );
  NAND2_X1 U14700 ( .A1(n17661), .A2(n19834), .ZN(n19224) );
  INV_X1 U14701 ( .A(n19224), .ZN(n17625) );
  NAND2_X1 U14702 ( .A1(n17625), .A2(n19835), .ZN(n17732) );
  INV_X1 U14703 ( .A(n17732), .ZN(n14275) );
  NAND2_X1 U14704 ( .A1(n19237), .A2(n14275), .ZN(n18958) );
  INV_X2 U14705 ( .A(n18958), .ZN(n19142) );
  AOI22_X1 U14706 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19142), .ZN(n13038) );
  OAI21_X1 U14707 ( .B1(n17827), .B2(n14179), .A(n13038), .ZN(n13039) );
  NAND2_X1 U14708 ( .A1(n14872), .A2(n13093), .ZN(n13052) );
  NAND2_X1 U14709 ( .A1(n14261), .A2(n13042), .ZN(n13043) );
  NAND2_X1 U14710 ( .A1(n13043), .A2(n13209), .ZN(n13045) );
  INV_X1 U14711 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13044) );
  MUX2_X2 U14712 ( .A(n13045), .B(n13044), .S(n20026), .Z(n13059) );
  INV_X1 U14713 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14351) );
  INV_X1 U14714 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13046) );
  AND2_X1 U14715 ( .A1(n14351), .A2(n13046), .ZN(n13047) );
  MUX2_X1 U14716 ( .A(n13047), .B(n13315), .S(n16391), .Z(n13058) );
  NAND2_X1 U14717 ( .A1(n13059), .A2(n13058), .ZN(n13057) );
  INV_X1 U14718 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13048) );
  MUX2_X1 U14719 ( .A(n13049), .B(n13048), .S(n20026), .Z(n13050) );
  OAI21_X1 U14720 ( .B1(n13051), .B2(n13050), .A(n13067), .ZN(n17041) );
  NAND2_X1 U14721 ( .A1(n13052), .A2(n17041), .ZN(n13061) );
  MUX2_X1 U14722 ( .A(n13212), .B(n13303), .S(n14261), .Z(n13053) );
  MUX2_X1 U14723 ( .A(n13053), .B(P2_EBX_REG_0__SCAN_IN), .S(n20026), .Z(
        n18864) );
  INV_X1 U14724 ( .A(n18864), .ZN(n13054) );
  NOR2_X1 U14725 ( .A1(n13054), .A2(n14339), .ZN(n13056) );
  AND2_X1 U14726 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n13055) );
  AOI21_X1 U14727 ( .B1(n20026), .B2(n13055), .A(n13058), .ZN(n17064) );
  NOR2_X1 U14728 ( .A1(n13056), .A2(n17064), .ZN(n14356) );
  AND2_X1 U14729 ( .A1(n13056), .A2(n17064), .ZN(n14355) );
  NOR2_X1 U14730 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14355), .ZN(
        n14354) );
  NOR2_X1 U14731 ( .A1(n14356), .A2(n14354), .ZN(n14365) );
  OAI21_X1 U14732 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n17052) );
  XNOR2_X1 U14733 ( .A(n17052), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14364) );
  NOR2_X1 U14734 ( .A1(n17052), .A2(n14408), .ZN(n13060) );
  AOI21_X1 U14735 ( .B1(n14365), .B2(n14364), .A(n13060), .ZN(n14870) );
  NAND2_X1 U14736 ( .A1(n13061), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13062) );
  INV_X1 U14737 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13063) );
  MUX2_X1 U14738 ( .A(n13064), .B(n13063), .S(n20026), .Z(n13065) );
  NAND2_X1 U14739 ( .A1(n13066), .A2(n13067), .ZN(n13068) );
  NOR2_X2 U14740 ( .A1(n13067), .A2(n13066), .ZN(n13074) );
  INV_X1 U14741 ( .A(n13074), .ZN(n13077) );
  NAND2_X1 U14742 ( .A1(n13068), .A2(n13077), .ZN(n17030) );
  XNOR2_X1 U14743 ( .A(n17030), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15055) );
  NAND2_X1 U14744 ( .A1(n15054), .A2(n15055), .ZN(n13071) );
  INV_X1 U14745 ( .A(n17030), .ZN(n13069) );
  NAND2_X1 U14746 ( .A1(n13069), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13070) );
  NAND2_X1 U14747 ( .A1(n13071), .A2(n13070), .ZN(n15667) );
  NAND2_X1 U14748 ( .A1(n13072), .A2(n13093), .ZN(n13079) );
  INV_X1 U14749 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13073) );
  MUX2_X1 U14750 ( .A(n13073), .B(n13335), .S(n16391), .Z(n13075) );
  NAND2_X1 U14751 ( .A1(n13074), .A2(n13075), .ZN(n13085) );
  INV_X1 U14752 ( .A(n13075), .ZN(n13076) );
  NAND2_X1 U14753 ( .A1(n13077), .A2(n13076), .ZN(n13078) );
  NAND2_X1 U14754 ( .A1(n13085), .A2(n13078), .ZN(n17016) );
  NAND2_X1 U14755 ( .A1(n15667), .A2(n15666), .ZN(n13082) );
  NAND2_X1 U14756 ( .A1(n13080), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13081) );
  NAND2_X1 U14757 ( .A1(n13082), .A2(n13081), .ZN(n15763) );
  NAND2_X1 U14758 ( .A1(n13083), .A2(n13093), .ZN(n13088) );
  MUX2_X1 U14759 ( .A(n13084), .B(P2_EBX_REG_6__SCAN_IN), .S(n20026), .Z(
        n13086) );
  NOR2_X2 U14760 ( .A1(n13085), .A2(n13086), .ZN(n13099) );
  INV_X1 U14761 ( .A(n13099), .ZN(n13096) );
  NAND2_X1 U14762 ( .A1(n13085), .A2(n13086), .ZN(n13087) );
  NAND2_X1 U14763 ( .A1(n13096), .A2(n13087), .ZN(n18875) );
  INV_X1 U14764 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13089) );
  NAND2_X1 U14765 ( .A1(n15763), .A2(n15762), .ZN(n13092) );
  NAND2_X1 U14766 ( .A1(n13090), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13091) );
  NAND2_X1 U14767 ( .A1(n13092), .A2(n13091), .ZN(n17343) );
  INV_X1 U14768 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U14769 ( .A(n13094), .B(n16393), .S(n16391), .Z(n13098) );
  INV_X1 U14770 ( .A(n13098), .ZN(n13095) );
  XNOR2_X1 U14771 ( .A(n13096), .B(n13095), .ZN(n18894) );
  XNOR2_X1 U14772 ( .A(n18894), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17345) );
  NAND2_X1 U14773 ( .A1(n17343), .A2(n17345), .ZN(n16155) );
  INV_X1 U14774 ( .A(n18894), .ZN(n13097) );
  NAND2_X1 U14775 ( .A1(n13097), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16153) );
  NAND2_X1 U14776 ( .A1(n16155), .A2(n16153), .ZN(n13188) );
  NAND2_X1 U14777 ( .A1(n13099), .A2(n13098), .ZN(n13103) );
  INV_X1 U14778 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n17006) );
  XNOR2_X1 U14779 ( .A(n13103), .B(n11244), .ZN(n17007) );
  NAND2_X1 U14780 ( .A1(n17007), .A2(n16393), .ZN(n13101) );
  INV_X1 U14781 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U14782 ( .A1(n13101), .A2(n13100), .ZN(n17741) );
  NAND2_X1 U14783 ( .A1(n13188), .A2(n17741), .ZN(n13102) );
  OR2_X1 U14784 ( .A1(n13101), .A2(n13100), .ZN(n17742) );
  NAND2_X1 U14785 ( .A1(n13102), .A2(n17742), .ZN(n17327) );
  INV_X1 U14786 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13105) );
  NOR2_X1 U14787 ( .A1(n16391), .A2(n13105), .ZN(n13108) );
  INV_X1 U14788 ( .A(n13108), .ZN(n13106) );
  XNOR2_X1 U14789 ( .A(n13109), .B(n13106), .ZN(n16988) );
  NAND2_X1 U14790 ( .A1(n16988), .A2(n16393), .ZN(n13107) );
  NAND2_X1 U14791 ( .A1(n13107), .A2(n17573), .ZN(n17328) );
  NOR2_X2 U14792 ( .A1(n13109), .A2(n13108), .ZN(n13113) );
  INV_X1 U14793 ( .A(n13113), .ZN(n13110) );
  NAND2_X1 U14794 ( .A1(n20026), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13112) );
  XNOR2_X1 U14795 ( .A(n13110), .B(n13112), .ZN(n18908) );
  AOI21_X1 U14796 ( .B1(n18908), .B2(n16393), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17557) );
  INV_X1 U14797 ( .A(n17557), .ZN(n13111) );
  AND2_X1 U14798 ( .A1(n17328), .A2(n13111), .ZN(n13189) );
  AND2_X2 U14799 ( .A1(n13113), .A2(n13112), .ZN(n13128) );
  NAND2_X1 U14800 ( .A1(n20026), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U14801 ( .A1(n13128), .A2(n13129), .ZN(n13122) );
  INV_X1 U14802 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13114) );
  NOR2_X1 U14803 ( .A1(n16391), .A2(n13114), .ZN(n13123) );
  INV_X1 U14804 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13115) );
  NOR2_X1 U14805 ( .A1(n16391), .A2(n13115), .ZN(n13118) );
  NAND2_X1 U14806 ( .A1(n20026), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U14807 ( .A1(n20026), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13150) );
  XNOR2_X1 U14808 ( .A(n13149), .B(n13150), .ZN(n18963) );
  NAND2_X1 U14809 ( .A1(n18963), .A2(n16393), .ZN(n13137) );
  AND2_X1 U14810 ( .A1(n13137), .A2(n17473), .ZN(n17469) );
  INV_X1 U14811 ( .A(n13116), .ZN(n13117) );
  XNOR2_X1 U14812 ( .A(n13119), .B(n13117), .ZN(n18945) );
  NAND2_X1 U14813 ( .A1(n18945), .A2(n16393), .ZN(n13138) );
  INV_X1 U14814 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17511) );
  AND2_X1 U14815 ( .A1(n13125), .A2(n13118), .ZN(n13120) );
  OR2_X1 U14816 ( .A1(n13120), .A2(n13119), .ZN(n13135) );
  INV_X1 U14817 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U14818 ( .B1(n13135), .B2(n13093), .A(n13121), .ZN(n17759) );
  NAND2_X1 U14819 ( .A1(n13122), .A2(n13123), .ZN(n13124) );
  NAND2_X1 U14820 ( .A1(n13125), .A2(n13124), .ZN(n16984) );
  OR2_X1 U14821 ( .A1(n16984), .A2(n13093), .ZN(n13126) );
  INV_X1 U14822 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19129) );
  NAND2_X1 U14823 ( .A1(n13126), .A2(n19129), .ZN(n17465) );
  NAND2_X1 U14824 ( .A1(n17759), .A2(n17465), .ZN(n13127) );
  INV_X1 U14825 ( .A(n13128), .ZN(n13131) );
  INV_X1 U14826 ( .A(n13129), .ZN(n13130) );
  NAND2_X1 U14827 ( .A1(n13131), .A2(n13130), .ZN(n13132) );
  NAND2_X1 U14828 ( .A1(n13122), .A2(n13132), .ZN(n18911) );
  NAND2_X1 U14829 ( .A1(n13140), .A2(n17533), .ZN(n17318) );
  NAND2_X1 U14830 ( .A1(n17316), .A2(n13134), .ZN(n13148) );
  INV_X1 U14831 ( .A(n13135), .ZN(n18936) );
  AND2_X1 U14832 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13136) );
  NAND2_X1 U14833 ( .A1(n18936), .A2(n13136), .ZN(n17758) );
  NOR2_X1 U14834 ( .A1(n17473), .A2(n13137), .ZN(n17468) );
  NOR2_X1 U14835 ( .A1(n17511), .A2(n13138), .ZN(n17492) );
  NOR2_X1 U14836 ( .A1(n17468), .A2(n17492), .ZN(n13139) );
  NAND2_X1 U14837 ( .A1(n17758), .A2(n13139), .ZN(n16173) );
  INV_X1 U14838 ( .A(n13140), .ZN(n13141) );
  NAND2_X1 U14839 ( .A1(n13141), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17317) );
  AND2_X1 U14840 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13142) );
  AND2_X1 U14841 ( .A1(n16988), .A2(n13142), .ZN(n17331) );
  AND2_X1 U14842 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13143) );
  AND2_X1 U14843 ( .A1(n18908), .A2(n13143), .ZN(n17556) );
  NOR2_X1 U14844 ( .A1(n17331), .A2(n17556), .ZN(n13144) );
  NAND2_X1 U14845 ( .A1(n17317), .A2(n13144), .ZN(n13191) );
  NAND2_X1 U14846 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13145) );
  NOR2_X1 U14847 ( .A1(n16984), .A2(n13145), .ZN(n16150) );
  OR2_X1 U14848 ( .A1(n13191), .A2(n16150), .ZN(n13146) );
  NOR2_X1 U14849 ( .A1(n16173), .A2(n13146), .ZN(n13147) );
  NAND2_X1 U14850 ( .A1(n13151), .A2(n13150), .ZN(n13154) );
  INV_X1 U14851 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13152) );
  NOR2_X1 U14852 ( .A1(n16391), .A2(n13152), .ZN(n13153) );
  OR2_X2 U14853 ( .A1(n13154), .A2(n13153), .ZN(n13162) );
  NAND2_X1 U14854 ( .A1(n13154), .A2(n13153), .ZN(n13155) );
  NAND2_X1 U14855 ( .A1(n13162), .A2(n13155), .ZN(n16968) );
  INV_X1 U14856 ( .A(n16968), .ZN(n13157) );
  AND2_X1 U14857 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13156) );
  NAND2_X1 U14858 ( .A1(n13157), .A2(n13156), .ZN(n17305) );
  INV_X1 U14859 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U14860 ( .B1(n16968), .B2(n13093), .A(n19140), .ZN(n13158) );
  NAND2_X1 U14861 ( .A1(n17785), .A2(n17786), .ZN(n17306) );
  NAND2_X1 U14862 ( .A1(n20026), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13160) );
  XNOR2_X1 U14863 ( .A(n13162), .B(n13160), .ZN(n18969) );
  AND2_X1 U14864 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13159) );
  NAND2_X1 U14865 ( .A1(n18969), .A2(n13159), .ZN(n17303) );
  AND2_X1 U14866 ( .A1(n17303), .A2(n17305), .ZN(n16175) );
  AOI21_X1 U14867 ( .B1(n18969), .B2(n16393), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16159) );
  AOI21_X2 U14868 ( .B1(n17306), .B2(n16175), .A(n16159), .ZN(n17798) );
  INV_X1 U14869 ( .A(n13160), .ZN(n13161) );
  NAND2_X1 U14870 ( .A1(n20026), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13164) );
  INV_X1 U14871 ( .A(n13163), .ZN(n13166) );
  INV_X1 U14872 ( .A(n13164), .ZN(n13165) );
  NAND2_X1 U14873 ( .A1(n13166), .A2(n13165), .ZN(n13167) );
  NAND2_X1 U14874 ( .A1(n13171), .A2(n13167), .ZN(n18982) );
  NAND2_X1 U14875 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13168) );
  NOR2_X1 U14876 ( .A1(n18982), .A2(n13168), .ZN(n16172) );
  INV_X1 U14877 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n13169) );
  NOR2_X1 U14878 ( .A1(n16391), .A2(n13169), .ZN(n13170) );
  NAND2_X1 U14879 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  NAND2_X1 U14880 ( .A1(n13180), .A2(n13172), .ZN(n18997) );
  INV_X1 U14881 ( .A(n18997), .ZN(n13174) );
  AND2_X1 U14882 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U14883 ( .A1(n13174), .A2(n13173), .ZN(n17290) );
  OAI21_X1 U14884 ( .B1(n18997), .B2(n13093), .A(n17437), .ZN(n17291) );
  OR2_X1 U14885 ( .A1(n18982), .A2(n13093), .ZN(n13176) );
  INV_X1 U14886 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U14887 ( .A1(n13176), .A2(n13175), .ZN(n17799) );
  NAND2_X1 U14888 ( .A1(n17291), .A2(n17799), .ZN(n16163) );
  NAND2_X1 U14889 ( .A1(n20026), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U14890 ( .A1(n13177), .A2(n13178), .ZN(n16157) );
  INV_X1 U14891 ( .A(n13178), .ZN(n13179) );
  NAND2_X1 U14892 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  AND2_X1 U14893 ( .A1(n16157), .A2(n13181), .ZN(n16947) );
  OAI21_X1 U14894 ( .B1(n13182), .B2(n16177), .A(n17277), .ZN(n13183) );
  NOR2_X2 U14895 ( .A1(n19250), .A2(n20227), .ZN(n17818) );
  NAND2_X1 U14896 ( .A1(n11236), .A2(n11294), .ZN(P2_U2994) );
  INV_X1 U14897 ( .A(n13185), .ZN(n17333) );
  NOR2_X2 U14898 ( .A1(n17333), .A2(n17573), .ZN(n17332) );
  NAND2_X1 U14899 ( .A1(n17332), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17544) );
  NOR2_X2 U14900 ( .A1(n17544), .A2(n17533), .ZN(n17510) );
  INV_X1 U14901 ( .A(n17510), .ZN(n13186) );
  NOR2_X1 U14902 ( .A1(n17510), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13187) );
  AND2_X1 U14903 ( .A1(n17318), .A2(n13189), .ZN(n13190) );
  AND2_X1 U14904 ( .A1(n17741), .A2(n13190), .ZN(n16166) );
  NAND2_X1 U14905 ( .A1(n17744), .A2(n16166), .ZN(n17464) );
  INV_X1 U14906 ( .A(n13191), .ZN(n13192) );
  AND2_X1 U14907 ( .A1(n17742), .A2(n13192), .ZN(n16151) );
  AND2_X1 U14908 ( .A1(n17464), .A2(n16151), .ZN(n13195) );
  INV_X1 U14909 ( .A(n17465), .ZN(n13193) );
  NOR2_X1 U14910 ( .A1(n13193), .A2(n16150), .ZN(n13194) );
  XNOR2_X1 U14911 ( .A(n13195), .B(n13194), .ZN(n17522) );
  INV_X1 U14912 ( .A(n17818), .ZN(n13196) );
  INV_X1 U14913 ( .A(n15653), .ZN(n15127) );
  OR2_X1 U14914 ( .A1(n15127), .A2(n13197), .ZN(n15125) );
  NAND2_X1 U14915 ( .A1(n15127), .A2(n13197), .ZN(n13198) );
  INV_X1 U14916 ( .A(n17520), .ZN(n13200) );
  INV_X1 U14917 ( .A(n17807), .ZN(n13199) );
  OAI21_X1 U14918 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14192), .A(
        n14197), .ZN(n16973) );
  AOI22_X1 U14919 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19142), .ZN(n13202) );
  OAI21_X1 U14920 ( .B1(n17827), .B2(n16973), .A(n13202), .ZN(n13203) );
  NOR2_X1 U14921 ( .A1(n13207), .A2(n19189), .ZN(n13208) );
  OR2_X1 U14922 ( .A1(n13228), .A2(n13208), .ZN(n13226) );
  INV_X1 U14923 ( .A(n13209), .ZN(n13221) );
  AOI21_X1 U14924 ( .B1(n18853), .B2(n19096), .A(n13210), .ZN(n13220) );
  INV_X1 U14925 ( .A(n13210), .ZN(n13214) );
  OAI21_X1 U14926 ( .B1(n19096), .B2(n13212), .A(n13211), .ZN(n13213) );
  OAI21_X1 U14927 ( .B1(n13214), .B2(n19096), .A(n13213), .ZN(n13215) );
  NAND2_X1 U14928 ( .A1(n13215), .A2(n20289), .ZN(n13218) );
  NAND2_X1 U14929 ( .A1(n14261), .A2(n13216), .ZN(n13217) );
  NAND2_X1 U14930 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  OAI21_X1 U14931 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n13223) );
  AOI22_X1 U14932 ( .A1(n13224), .A2(n19189), .B1(n13223), .B2(n13222), .ZN(
        n13225) );
  NOR2_X1 U14933 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  MUX2_X1 U14934 ( .A(n19101), .B(n13227), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n13231) );
  INV_X1 U14935 ( .A(n18853), .ZN(n17882) );
  NAND2_X1 U14936 ( .A1(n19197), .A2(n19096), .ZN(n17666) );
  OAI211_X1 U14937 ( .C1(n13231), .C2(n13230), .A(n17666), .B(n13238), .ZN(
        n13258) );
  INV_X1 U14938 ( .A(n17666), .ZN(n17612) );
  NAND2_X1 U14939 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n22264) );
  INV_X1 U14940 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22270) );
  INV_X1 U14941 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n22282) );
  NAND2_X1 U14942 ( .A1(n22263), .A2(n22282), .ZN(n22266) );
  NOR2_X1 U14943 ( .A1(n22263), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n17855) );
  OAI21_X1 U14944 ( .B1(n22270), .B2(n22266), .A(n17939), .ZN(n22272) );
  NAND2_X1 U14945 ( .A1(n22264), .A2(n22272), .ZN(n14266) );
  INV_X1 U14946 ( .A(n14266), .ZN(n19201) );
  NAND3_X1 U14947 ( .A1(n17612), .A2(n19201), .A3(n13232), .ZN(n13257) );
  INV_X1 U14948 ( .A(n13233), .ZN(n13249) );
  NAND2_X1 U14949 ( .A1(n13234), .A2(n19201), .ZN(n13235) );
  OR2_X1 U14950 ( .A1(n19193), .A2(n13235), .ZN(n13248) );
  CLKBUF_X1 U14951 ( .A(n13236), .Z(n13237) );
  INV_X1 U14952 ( .A(n13237), .ZN(n13242) );
  NAND2_X1 U14953 ( .A1(n20227), .A2(n13238), .ZN(n13279) );
  NAND2_X1 U14954 ( .A1(n13279), .A2(n20289), .ZN(n13240) );
  NAND2_X1 U14955 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  AOI22_X1 U14956 ( .A1(n13242), .A2(n20081), .B1(n20179), .B2(n13241), .ZN(
        n13247) );
  OAI21_X1 U14957 ( .B1(n13243), .B2(n20081), .A(n20179), .ZN(n13244) );
  NAND2_X1 U14958 ( .A1(n14230), .A2(n13244), .ZN(n13246) );
  NAND2_X1 U14959 ( .A1(n13237), .A2(n14347), .ZN(n13245) );
  NAND2_X1 U14960 ( .A1(n13245), .A2(n19186), .ZN(n13263) );
  NAND2_X1 U14961 ( .A1(n13248), .A2(n13281), .ZN(n17608) );
  AOI21_X1 U14962 ( .B1(n13249), .B2(n19190), .A(n17608), .ZN(n13256) );
  INV_X1 U14963 ( .A(n19193), .ZN(n13252) );
  INV_X1 U14964 ( .A(n22264), .ZN(n22275) );
  AOI21_X1 U14965 ( .B1(n13250), .B2(n19096), .A(n22275), .ZN(n13251) );
  AOI22_X1 U14966 ( .A1(n19242), .A2(n19190), .B1(n13252), .B2(n13251), .ZN(
        n13254) );
  OR2_X1 U14967 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  NAND4_X1 U14968 ( .A1(n13258), .A2(n13257), .A3(n13256), .A4(n13255), .ZN(
        n13259) );
  AND2_X1 U14969 ( .A1(n19190), .A2(n14261), .ZN(n13260) );
  NAND2_X1 U14970 ( .A1(n13262), .A2(n19096), .ZN(n17604) );
  NAND2_X1 U14971 ( .A1(n17604), .A2(n13263), .ZN(n13264) );
  NAND2_X1 U14972 ( .A1(n13264), .A2(n12564), .ZN(n13276) );
  OAI21_X1 U14973 ( .B1(n12549), .B2(n13266), .A(n14274), .ZN(n13268) );
  NAND2_X1 U14974 ( .A1(n13268), .A2(n13267), .ZN(n13273) );
  OAI22_X1 U14975 ( .A1(n14274), .A2(n20081), .B1(n20289), .B2(n20179), .ZN(
        n13269) );
  INV_X1 U14976 ( .A(n13269), .ZN(n13272) );
  OR2_X1 U14977 ( .A1(n13271), .A2(n13270), .ZN(n13967) );
  AND4_X1 U14978 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13967), .ZN(
        n13275) );
  NAND2_X1 U14979 ( .A1(n19074), .A2(n13277), .ZN(n13278) );
  INV_X1 U14980 ( .A(n17451), .ZN(n13282) );
  NAND2_X1 U14981 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17597) );
  NOR2_X1 U14982 ( .A1(n14408), .A2(n17597), .ZN(n14878) );
  NAND2_X1 U14983 ( .A1(n14408), .A2(n17597), .ZN(n14879) );
  INV_X1 U14984 ( .A(n14879), .ZN(n14410) );
  NOR4_X1 U14985 ( .A1(n13089), .A2(n15058), .A3(n15664), .A4(n15672), .ZN(
        n15773) );
  INV_X1 U14986 ( .A(n15773), .ZN(n13290) );
  NAND2_X1 U14987 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19162) );
  NOR3_X1 U14988 ( .A1(n14410), .A2(n13290), .A3(n19162), .ZN(n13283) );
  NAND2_X1 U14989 ( .A1(n14878), .A2(n13283), .ZN(n16223) );
  NOR2_X1 U14990 ( .A1(n13292), .A2(n16223), .ZN(n17449) );
  OAI21_X1 U14991 ( .B1(n13282), .B2(n17449), .A(n13293), .ZN(n13289) );
  INV_X1 U14992 ( .A(n13279), .ZN(n13280) );
  NAND2_X1 U14993 ( .A1(n17448), .A2(n13282), .ZN(n17598) );
  INV_X1 U14994 ( .A(n13283), .ZN(n13284) );
  NAND2_X1 U14995 ( .A1(n17447), .A2(n13284), .ZN(n13286) );
  INV_X1 U14996 ( .A(n13523), .ZN(n13285) );
  NAND2_X1 U14997 ( .A1(n13285), .A2(n17323), .ZN(n14409) );
  AND2_X1 U14998 ( .A1(n13286), .A2(n14409), .ZN(n16225) );
  NAND2_X1 U14999 ( .A1(n17447), .A2(n13292), .ZN(n13287) );
  AND2_X1 U15000 ( .A1(n16225), .A2(n13287), .ZN(n17453) );
  INV_X1 U15001 ( .A(n17453), .ZN(n13288) );
  AOI21_X1 U15002 ( .B1(n13289), .B2(n17598), .A(n13288), .ZN(n19145) );
  AOI22_X1 U15003 ( .A1(n17447), .A2(n14879), .B1(n17451), .B2(n14878), .ZN(
        n15771) );
  NOR2_X1 U15004 ( .A1(n15771), .A2(n13290), .ZN(n19163) );
  INV_X1 U15005 ( .A(n19162), .ZN(n13291) );
  NAND2_X1 U15006 ( .A1(n19163), .A2(n13291), .ZN(n17566) );
  NOR2_X1 U15007 ( .A1(n13292), .A2(n17566), .ZN(n17480) );
  NAND3_X1 U15008 ( .A1(n13293), .A2(n17480), .A3(n13175), .ZN(n19144) );
  NAND2_X1 U15009 ( .A1(n19145), .A2(n19144), .ZN(n17442) );
  NAND2_X1 U15010 ( .A1(n13294), .A2(n14230), .ZN(n19192) );
  NAND2_X1 U15011 ( .A1(n19192), .A2(n19096), .ZN(n13296) );
  NAND2_X1 U15012 ( .A1(n13295), .A2(n17602), .ZN(n14344) );
  NAND2_X1 U15013 ( .A1(n13296), .A2(n14344), .ZN(n13297) );
  INV_X1 U15014 ( .A(n13298), .ZN(n13299) );
  NOR2_X1 U15015 ( .A1(n14347), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13310) );
  AND2_X1 U15016 ( .A1(n13300), .A2(n19834), .ZN(n13345) );
  AOI222_X1 U15017 ( .A1(n16415), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n16414), 
        .B2(P2_EAX_REG_20__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), 
        .C2(n13343), .ZN(n13512) );
  NAND2_X1 U15018 ( .A1(n13243), .A2(n13345), .ZN(n13320) );
  NAND2_X1 U15019 ( .A1(n13502), .A2(n13303), .ZN(n13305) );
  MUX2_X1 U15020 ( .A(n14347), .B(n19856), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13304) );
  NAND3_X1 U15021 ( .A1(n13320), .A2(n13305), .A3(n13304), .ZN(n14396) );
  INV_X1 U15022 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U15023 ( .A1(n13300), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13306) );
  OAI211_X1 U15024 ( .C1(n14347), .C2(n13307), .A(n13306), .B(n19834), .ZN(
        n13308) );
  INV_X1 U15025 ( .A(n13308), .ZN(n13309) );
  INV_X1 U15026 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U15027 ( .A1(n13310), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13345), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13311) );
  OAI21_X1 U15028 ( .B1(n13983), .B2(n17918), .A(n13311), .ZN(n13318) );
  INV_X1 U15029 ( .A(n13318), .ZN(n13312) );
  NOR2_X1 U15030 ( .A1(n13243), .A2(n13313), .ZN(n13314) );
  MUX2_X1 U15031 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n13314), .S(
        n19834), .Z(n13317) );
  AND2_X1 U15032 ( .A1(n11147), .A2(n13315), .ZN(n13316) );
  NOR2_X1 U15033 ( .A1(n13317), .A2(n13316), .ZN(n14484) );
  NAND2_X1 U15034 ( .A1(n14483), .A2(n14484), .ZN(n14488) );
  OR2_X1 U15035 ( .A1(n14398), .A2(n13318), .ZN(n13322) );
  NAND2_X1 U15036 ( .A1(n11147), .A2(n13042), .ZN(n13319) );
  OAI211_X1 U15037 ( .C1(n19834), .C2(n19906), .A(n13320), .B(n13319), .ZN(
        n13321) );
  AND3_X1 U15038 ( .A1(n14488), .A2(n13322), .A3(n13321), .ZN(n13323) );
  AOI22_X1 U15039 ( .A1(n16414), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U15040 ( .B1(n13980), .B2(n14369), .A(n13324), .ZN(n14406) );
  NOR2_X1 U15041 ( .A1(n14407), .A2(n14406), .ZN(n13325) );
  INV_X1 U15042 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U15043 ( .A1(n11147), .A2(n13327), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U15044 ( .A1(n16414), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13328) );
  OAI211_X1 U15045 ( .C1(n13980), .C2(n14886), .A(n13329), .B(n13328), .ZN(
        n14874) );
  NAND2_X1 U15046 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  AOI22_X1 U15047 ( .A1(n16414), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U15048 ( .A1(n11147), .A2(n13330), .ZN(n13331) );
  OAI211_X1 U15049 ( .C1(n13980), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        n15062) );
  INV_X1 U15050 ( .A(n15062), .ZN(n13334) );
  AOI22_X1 U15051 ( .A1(n16415), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11147), 
        .B2(n13335), .ZN(n13337) );
  AOI22_X1 U15052 ( .A1(n16414), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13336) );
  NAND2_X1 U15053 ( .A1(n13337), .A2(n13336), .ZN(n15670) );
  NAND2_X1 U15054 ( .A1(n15063), .A2(n15670), .ZN(n15669) );
  NAND2_X1 U15055 ( .A1(n11147), .A2(n13338), .ZN(n15777) );
  NAND2_X1 U15056 ( .A1(n11147), .A2(n16393), .ZN(n13339) );
  AND2_X1 U15057 ( .A1(n15777), .A2(n13339), .ZN(n13342) );
  INV_X1 U15058 ( .A(n13339), .ZN(n13341) );
  AOI22_X1 U15059 ( .A1(n16414), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13340) );
  OAI21_X1 U15060 ( .B1(n13980), .B2(n12984), .A(n13340), .ZN(n15778) );
  AOI22_X1 U15061 ( .A1(n16414), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13344) );
  OAI21_X1 U15062 ( .B1(n13980), .B2(n17347), .A(n13344), .ZN(n17578) );
  NAND2_X1 U15063 ( .A1(n17579), .A2(n17578), .ZN(n16999) );
  AOI22_X1 U15064 ( .A1(n16414), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U15065 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13847), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U15066 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U15067 ( .A1(n13890), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U15068 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13346) );
  NAND4_X1 U15069 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13360) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13351) );
  INV_X1 U15071 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13350) );
  OAI22_X1 U15072 ( .A1(n13876), .A2(n13351), .B1(n13874), .B2(n13350), .ZN(
        n13352) );
  AOI21_X1 U15073 ( .B1(n13462), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13352), .ZN(n13358) );
  AOI22_X1 U15074 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U15075 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13353) );
  AND2_X1 U15076 ( .A1(n13354), .A2(n13353), .ZN(n13357) );
  AOI22_X1 U15077 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13885), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U15078 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13355) );
  NAND4_X1 U15079 ( .A1(n13358), .A2(n13357), .A3(n13356), .A4(n13355), .ZN(
        n13359) );
  NAND2_X1 U15080 ( .A1(n11147), .A2(n14604), .ZN(n13361) );
  OAI211_X1 U15081 ( .C1(n13980), .C2(n13363), .A(n13362), .B(n13361), .ZN(
        n17001) );
  INV_X1 U15082 ( .A(n17001), .ZN(n13364) );
  AOI22_X1 U15083 ( .A1(n16414), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13343), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13383) );
  INV_X1 U15084 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13366) );
  INV_X1 U15085 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13365) );
  OAI22_X1 U15086 ( .A1(n13876), .A2(n13366), .B1(n13874), .B2(n13365), .ZN(
        n13367) );
  AOI21_X1 U15087 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n13367), .ZN(n13375) );
  NAND2_X1 U15088 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13369) );
  NAND2_X1 U15089 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13368) );
  OAI211_X1 U15090 ( .C1(n13882), .C2(n13370), .A(n13369), .B(n13368), .ZN(
        n13371) );
  INV_X1 U15091 ( .A(n13371), .ZN(n13374) );
  AOI22_X1 U15092 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13373) );
  NAND2_X1 U15093 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13372) );
  NAND4_X1 U15094 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13381) );
  AOI22_X1 U15095 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U15096 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U15097 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U15098 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13376) );
  NAND4_X1 U15099 ( .A1(n13379), .A2(n13378), .A3(n13377), .A4(n13376), .ZN(
        n13380) );
  NAND2_X1 U15100 ( .A1(n11147), .A2(n14748), .ZN(n13382) );
  OAI211_X1 U15101 ( .C1(n13980), .C2(n13384), .A(n13383), .B(n13382), .ZN(
        n16991) );
  AOI22_X1 U15102 ( .A1(n16414), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U15103 ( .A1(n13470), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U15104 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U15105 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13386) );
  NAND2_X1 U15106 ( .A1(n12712), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13385) );
  NAND4_X1 U15107 ( .A1(n13388), .A2(n13387), .A3(n13386), .A4(n13385), .ZN(
        n13393) );
  INV_X1 U15108 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13391) );
  NAND2_X1 U15109 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13390) );
  NAND2_X1 U15110 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13389) );
  OAI211_X1 U15111 ( .C1(n13882), .C2(n13391), .A(n13390), .B(n13389), .ZN(
        n13392) );
  NOR2_X1 U15112 ( .A1(n13393), .A2(n13392), .ZN(n13402) );
  AOI22_X1 U15113 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U15114 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13394) );
  AND2_X1 U15115 ( .A1(n13395), .A2(n13394), .ZN(n13401) );
  INV_X1 U15116 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U15117 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13397) );
  NAND2_X1 U15118 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13396) );
  OAI211_X1 U15119 ( .C1(n13841), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        n13399) );
  INV_X1 U15120 ( .A(n13399), .ZN(n13400) );
  INV_X1 U15121 ( .A(n13766), .ZN(n14861) );
  NAND2_X1 U15122 ( .A1(n11147), .A2(n14861), .ZN(n13403) );
  OAI211_X1 U15123 ( .C1(n13980), .C2(n13405), .A(n13404), .B(n13403), .ZN(
        n17552) );
  INV_X1 U15124 ( .A(n17552), .ZN(n13406) );
  AOI22_X1 U15125 ( .A1(n16414), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U15126 ( .A1(n13462), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13865), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U15127 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U15128 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U15129 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13407) );
  NAND4_X1 U15130 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13421) );
  INV_X1 U15131 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13412) );
  INV_X1 U15132 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13411) );
  OAI22_X1 U15133 ( .A1(n13876), .A2(n13412), .B1(n13874), .B2(n13411), .ZN(
        n13413) );
  AOI21_X1 U15134 ( .B1(n11219), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n13413), .ZN(n13419) );
  AOI22_X1 U15135 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U15136 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13414) );
  AND2_X1 U15137 ( .A1(n13415), .A2(n13414), .ZN(n13418) );
  AOI22_X1 U15138 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13885), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U15139 ( .A1(n13890), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13416) );
  NAND4_X1 U15140 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        n13420) );
  NAND2_X1 U15141 ( .A1(n11147), .A2(n14927), .ZN(n13422) );
  OAI211_X1 U15142 ( .C1(n13980), .C2(n17322), .A(n13423), .B(n13422), .ZN(
        n17529) );
  NAND2_X1 U15143 ( .A1(n17528), .A2(n17529), .ZN(n16975) );
  AOI22_X1 U15144 ( .A1(n16414), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13442) );
  INV_X1 U15145 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13425) );
  INV_X1 U15146 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13424) );
  OAI22_X1 U15147 ( .A1(n13876), .A2(n13425), .B1(n13874), .B2(n13424), .ZN(
        n13426) );
  AOI21_X1 U15148 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n13426), .ZN(n13434) );
  INV_X1 U15149 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13429) );
  NAND2_X1 U15150 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13428) );
  NAND2_X1 U15151 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13427) );
  OAI211_X1 U15152 ( .C1(n13882), .C2(n13429), .A(n13428), .B(n13427), .ZN(
        n13430) );
  INV_X1 U15153 ( .A(n13430), .ZN(n13433) );
  AOI22_X1 U15154 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U15155 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13431) );
  NAND4_X1 U15156 ( .A1(n13434), .A2(n13433), .A3(n13432), .A4(n13431), .ZN(
        n13440) );
  AOI22_X1 U15157 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15158 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U15159 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U15160 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13435) );
  NAND4_X1 U15161 ( .A1(n13438), .A2(n13437), .A3(n13436), .A4(n13435), .ZN(
        n13439) );
  NAND2_X1 U15162 ( .A1(n11147), .A2(n14921), .ZN(n13441) );
  OAI211_X1 U15163 ( .C1(n13980), .C2(n13443), .A(n13442), .B(n13441), .ZN(
        n16977) );
  INV_X1 U15164 ( .A(n16977), .ZN(n13444) );
  NOR2_X2 U15165 ( .A1(n16975), .A2(n13444), .ZN(n18927) );
  AOI22_X1 U15166 ( .A1(n16414), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13460) );
  INV_X1 U15167 ( .A(n13445), .ZN(n13452) );
  AOI22_X1 U15168 ( .A1(n13470), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U15169 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U15170 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13447) );
  NAND2_X1 U15171 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13446) );
  AND4_X1 U15172 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        n13451) );
  AOI22_X1 U15173 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13450) );
  OAI211_X1 U15174 ( .C1(n13452), .C2(n13704), .A(n13451), .B(n13450), .ZN(
        n13458) );
  AOI22_X1 U15175 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U15176 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13847), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15177 ( .A1(n13462), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U15178 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13453) );
  NAND4_X1 U15179 ( .A1(n13456), .A2(n13455), .A3(n13454), .A4(n13453), .ZN(
        n13457) );
  NAND2_X1 U15180 ( .A1(n11147), .A2(n15130), .ZN(n13459) );
  OAI211_X1 U15181 ( .C1(n13980), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        n18928) );
  NAND2_X1 U15182 ( .A1(n18927), .A2(n18928), .ZN(n17502) );
  AOI22_X1 U15183 ( .A1(n16414), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15184 ( .A1(n13462), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13878), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U15185 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U15186 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13464) );
  NAND2_X1 U15187 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13463) );
  NAND4_X1 U15188 ( .A1(n13466), .A2(n13465), .A3(n13464), .A4(n13463), .ZN(
        n13481) );
  AOI22_X1 U15189 ( .A1(n13467), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U15190 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13468) );
  AND2_X1 U15191 ( .A1(n13469), .A2(n13468), .ZN(n13479) );
  AOI22_X1 U15192 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13478) );
  INV_X1 U15193 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U15194 ( .A1(n13470), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13472) );
  NAND2_X1 U15195 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13471) );
  OAI211_X1 U15196 ( .C1(n13474), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        n13475) );
  INV_X1 U15197 ( .A(n13475), .ZN(n13477) );
  NAND2_X1 U15198 ( .A1(n13890), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13476) );
  NAND4_X1 U15199 ( .A1(n13479), .A2(n13478), .A3(n13477), .A4(n13476), .ZN(
        n13480) );
  NOR2_X1 U15200 ( .A1(n13481), .A2(n13480), .ZN(n13767) );
  INV_X1 U15201 ( .A(n13767), .ZN(n15660) );
  NAND2_X1 U15202 ( .A1(n11147), .A2(n15660), .ZN(n13482) );
  OAI211_X1 U15203 ( .C1(n13980), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        n17504) );
  AOI22_X1 U15204 ( .A1(n16414), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13504) );
  INV_X1 U15205 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13486) );
  INV_X1 U15206 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13485) );
  OAI22_X1 U15207 ( .A1(n13486), .A2(n13876), .B1(n13874), .B2(n13485), .ZN(
        n13487) );
  AOI21_X1 U15208 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n13487), .ZN(n13495) );
  INV_X1 U15209 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U15210 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13489) );
  NAND2_X1 U15211 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13488) );
  OAI211_X1 U15212 ( .C1(n13882), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        n13491) );
  INV_X1 U15213 ( .A(n13491), .ZN(n13494) );
  AOI22_X1 U15214 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13884), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U15215 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13492) );
  NAND4_X1 U15216 ( .A1(n13495), .A2(n13494), .A3(n13493), .A4(n13492), .ZN(
        n13501) );
  AOI22_X1 U15217 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U15218 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15219 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U15220 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13496) );
  NAND4_X1 U15221 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        n13500) );
  OR2_X1 U15222 ( .A1(n13501), .A2(n13500), .ZN(n15703) );
  NAND2_X1 U15223 ( .A1(n11147), .A2(n15703), .ZN(n13503) );
  OAI211_X1 U15224 ( .C1(n13980), .C2(n13505), .A(n13504), .B(n13503), .ZN(
        n17478) );
  NAND2_X1 U15225 ( .A1(n17476), .A2(n17478), .ZN(n15732) );
  NAND2_X1 U15226 ( .A1(n16415), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U15227 ( .A1(n16414), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U15228 ( .A1(n16414), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13508) );
  OAI21_X1 U15229 ( .B1(n13980), .B2(n17457), .A(n13508), .ZN(n17198) );
  NAND2_X1 U15230 ( .A1(n17196), .A2(n17198), .ZN(n18984) );
  NAND2_X1 U15231 ( .A1(n16415), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U15232 ( .A1(n16414), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13509) );
  NOR2_X2 U15233 ( .A1(n18984), .A2(n18985), .ZN(n17186) );
  INV_X1 U15234 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U15235 ( .A1(n16414), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13511) );
  OAI21_X1 U15236 ( .B1(n13980), .B2(n17929), .A(n13511), .ZN(n17187) );
  NOR2_X2 U15237 ( .A1(n17188), .A2(n13512), .ZN(n13970) );
  AOI21_X1 U15238 ( .B1(n13512), .B2(n17188), .A(n13970), .ZN(n20069) );
  AOI22_X1 U15239 ( .A1(n17442), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19154), .B2(n20069), .ZN(n13518) );
  NAND2_X1 U15240 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19142), .ZN(n13517) );
  NAND2_X1 U15241 ( .A1(n13514), .A2(n13513), .ZN(n16228) );
  NOR2_X1 U15242 ( .A1(n16228), .A2(n17566), .ZN(n17438) );
  OAI221_X1 U15243 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C1(n13515), .C2(n17437), .A(
        n17438), .ZN(n13516) );
  AND3_X1 U15244 ( .A1(n13518), .A2(n13517), .A3(n13516), .ZN(n13521) );
  NAND2_X1 U15245 ( .A1(n19082), .A2(n20227), .ZN(n13519) );
  NAND2_X1 U15246 ( .A1(n12572), .A2(n13519), .ZN(n13520) );
  AND2_X1 U15247 ( .A1(n19190), .A2(n19186), .ZN(n13522) );
  NAND3_X1 U15248 ( .A1(n11296), .A2(n11271), .A3(n13525), .ZN(P2_U3026) );
  NOR2_X1 U15249 ( .A1(n13527), .A2(n13526), .ZN(n13544) );
  AOI22_X1 U15250 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U15251 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U15252 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U15253 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11984), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13531) );
  NAND4_X1 U15254 ( .A1(n13534), .A2(n13533), .A3(n13532), .A4(n13531), .ZN(
        n13542) );
  AOI22_X1 U15255 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13535), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15256 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13539) );
  AOI22_X1 U15257 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U15258 ( .A1(n13536), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13537) );
  NAND4_X1 U15259 ( .A1(n13540), .A2(n13539), .A3(n13538), .A4(n13537), .ZN(
        n13541) );
  NOR2_X1 U15260 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  XNOR2_X1 U15261 ( .A(n13544), .B(n13543), .ZN(n13546) );
  NAND2_X1 U15262 ( .A1(n13546), .A2(n13545), .ZN(n13551) );
  INV_X1 U15263 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16469) );
  AOI21_X1 U15264 ( .B1(n16469), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13547) );
  AOI21_X1 U15265 ( .B1(n13553), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13547), .ZN(
        n13550) );
  XNOR2_X1 U15266 ( .A(n14015), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16141) );
  AOI21_X1 U15267 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n13583) );
  NAND2_X1 U15268 ( .A1(n13585), .A2(n13583), .ZN(n13556) );
  AOI22_X1 U15269 ( .A1(n13553), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13552), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13554) );
  INV_X1 U15270 ( .A(n13554), .ZN(n13555) );
  INV_X1 U15271 ( .A(n11192), .ZN(n17688) );
  NAND3_X1 U15272 ( .A1(n17688), .A2(n22243), .A3(n16447), .ZN(n13561) );
  OAI21_X1 U15273 ( .B1(n13558), .B2(n11229), .A(n13557), .ZN(n13559) );
  NAND2_X1 U15274 ( .A1(n13559), .A2(n16461), .ZN(n13560) );
  NAND2_X1 U15275 ( .A1(n13561), .A2(n13560), .ZN(n14314) );
  NAND4_X1 U15276 ( .A1(n15727), .A2(n11408), .A3(n14278), .A4(n11703), .ZN(
        n13586) );
  OR2_X1 U15277 ( .A1(n14299), .A2(n13586), .ZN(n13563) );
  AND2_X1 U15278 ( .A1(n16612), .A2(n15727), .ZN(n13565) );
  NAND2_X1 U15279 ( .A1(n11208), .A2(n13565), .ZN(n13582) );
  NOR4_X1 U15280 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13569) );
  NOR4_X1 U15281 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13568) );
  NOR4_X1 U15282 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13567) );
  NOR4_X1 U15283 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13566) );
  AND4_X1 U15284 ( .A1(n13569), .A2(n13568), .A3(n13567), .A4(n13566), .ZN(
        n13574) );
  NOR4_X1 U15285 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13572) );
  NOR4_X1 U15286 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13571) );
  NOR4_X1 U15287 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13570) );
  INV_X1 U15288 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20475) );
  AND4_X1 U15289 ( .A1(n13572), .A2(n13571), .A3(n13570), .A4(n20475), .ZN(
        n13573) );
  NAND2_X1 U15290 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  NOR2_X1 U15291 ( .A1(n13577), .A2(n15902), .ZN(n13576) );
  INV_X1 U15292 ( .A(DATAI_31_), .ZN(n15149) );
  INV_X1 U15293 ( .A(n15902), .ZN(n14671) );
  NOR3_X4 U15294 ( .A1(n15728), .A2(n13577), .A3(n14671), .ZN(n16616) );
  AOI22_X1 U15295 ( .A1(n16616), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15728), .ZN(n13578) );
  INV_X1 U15296 ( .A(n13578), .ZN(n13579) );
  NAND2_X1 U15297 ( .A1(n13582), .A2(n13581), .ZN(P1_U2873) );
  NAND3_X1 U15298 ( .A1(n16459), .A2(n14278), .A3(n16454), .ZN(n13590) );
  NOR2_X1 U15299 ( .A1(n13586), .A2(n11228), .ZN(n13587) );
  NAND2_X1 U15300 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  OAI22_X1 U15301 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n11229), .ZN(n16250) );
  OAI22_X1 U15302 ( .A1(n16251), .A2(n11854), .B1(n13593), .B2(n13592), .ZN(
        n13594) );
  XOR2_X1 U15303 ( .A(n16250), .B(n13594), .Z(n16478) );
  NAND2_X2 U15304 ( .A1(n20556), .A2(n15727), .ZN(n20551) );
  INV_X1 U15305 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13595) );
  OAI22_X1 U15306 ( .A1(n16478), .A2(n20551), .B1(n13595), .B2(n20556), .ZN(
        n13596) );
  NAND2_X1 U15307 ( .A1(n13598), .A2(n13597), .ZN(P1_U2842) );
  INV_X1 U15308 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13600) );
  INV_X1 U15309 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13599) );
  OAI22_X1 U15310 ( .A1(n13876), .A2(n13600), .B1(n13874), .B2(n13599), .ZN(
        n13601) );
  AOI21_X1 U15311 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13601), .ZN(n13608) );
  INV_X1 U15312 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U15313 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13603) );
  NAND2_X1 U15314 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13602) );
  OAI211_X1 U15315 ( .C1(n13882), .C2(n13764), .A(n13603), .B(n13602), .ZN(
        n13604) );
  INV_X1 U15316 ( .A(n13604), .ZN(n13607) );
  AOI22_X1 U15317 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13884), .B1(
        n12701), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U15318 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13605) );
  NAND4_X1 U15319 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13614) );
  AOI22_X1 U15320 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15321 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15322 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U15323 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13609) );
  NAND4_X1 U15324 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13613) );
  NOR2_X1 U15325 ( .A1(n13614), .A2(n13613), .ZN(n13903) );
  INV_X1 U15326 ( .A(n13903), .ZN(n13637) );
  INV_X1 U15327 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13619) );
  INV_X1 U15328 ( .A(n13615), .ZN(n13711) );
  INV_X1 U15329 ( .A(n13711), .ZN(n13626) );
  NAND2_X1 U15330 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13618) );
  AND2_X1 U15331 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13617) );
  OR2_X1 U15332 ( .A1(n13617), .A2(n13616), .ZN(n13950) );
  OAI211_X1 U15333 ( .C1(n13720), .C2(n13619), .A(n13618), .B(n13950), .ZN(
        n13620) );
  INV_X1 U15334 ( .A(n13620), .ZN(n13625) );
  AOI22_X1 U15335 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11217), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13624) );
  CLKBUF_X1 U15336 ( .A(n13621), .Z(n13954) );
  AOI22_X1 U15337 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U15338 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13622) );
  NAND4_X1 U15339 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13635) );
  INV_X1 U15340 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13628) );
  NAND2_X1 U15341 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13627) );
  INV_X1 U15342 ( .A(n13950), .ZN(n13694) );
  OAI211_X1 U15343 ( .C1(n13720), .C2(n13628), .A(n13627), .B(n13694), .ZN(
        n13629) );
  INV_X1 U15344 ( .A(n13629), .ZN(n13633) );
  AOI22_X1 U15345 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13945), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U15346 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U15347 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13630) );
  NAND4_X1 U15348 ( .A1(n13633), .A2(n13632), .A3(n13631), .A4(n13630), .ZN(
        n13634) );
  NAND2_X1 U15349 ( .A1(n13635), .A2(n13634), .ZN(n13902) );
  INV_X1 U15350 ( .A(n13902), .ZN(n13636) );
  NAND2_X1 U15351 ( .A1(n13637), .A2(n13636), .ZN(n13906) );
  INV_X1 U15352 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13639) );
  NAND2_X1 U15353 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13638) );
  OAI211_X1 U15354 ( .C1(n13720), .C2(n13639), .A(n13638), .B(n13694), .ZN(
        n13640) );
  INV_X1 U15355 ( .A(n13640), .ZN(n13644) );
  AOI22_X1 U15356 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13955), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13643) );
  AOI22_X1 U15357 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13941), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U15358 ( .A1(n19079), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13641) );
  NAND4_X1 U15359 ( .A1(n13644), .A2(n13643), .A3(n13642), .A4(n13641), .ZN(
        n13653) );
  NAND2_X1 U15360 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13645) );
  OAI211_X1 U15361 ( .C1(n13720), .C2(n12687), .A(n13645), .B(n13950), .ZN(
        n13646) );
  INV_X1 U15362 ( .A(n13646), .ZN(n13651) );
  AOI22_X1 U15363 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13941), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13650) );
  AOI22_X1 U15364 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U15365 ( .A1(n13945), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13648) );
  NAND4_X1 U15366 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13652) );
  NAND2_X1 U15367 ( .A1(n13653), .A2(n13652), .ZN(n13907) );
  NOR2_X1 U15368 ( .A1(n13906), .A2(n13907), .ZN(n13909) );
  NAND2_X1 U15369 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13654) );
  OAI211_X1 U15370 ( .C1(n13720), .C2(n13655), .A(n13654), .B(n13950), .ZN(
        n13656) );
  INV_X1 U15371 ( .A(n13656), .ZN(n13660) );
  AOI22_X1 U15372 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U15373 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15374 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U15375 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13669) );
  INV_X1 U15376 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U15377 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13661) );
  OAI211_X1 U15378 ( .C1(n13720), .C2(n13662), .A(n13661), .B(n13694), .ZN(
        n13663) );
  INV_X1 U15379 ( .A(n13663), .ZN(n13667) );
  AOI22_X1 U15380 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U15381 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U15382 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13664) );
  NAND4_X1 U15383 ( .A1(n13667), .A2(n13666), .A3(n13665), .A4(n13664), .ZN(
        n13668) );
  AND2_X1 U15384 ( .A1(n13669), .A2(n13668), .ZN(n13911) );
  NAND2_X1 U15385 ( .A1(n13909), .A2(n13911), .ZN(n13914) );
  NAND2_X1 U15386 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13670) );
  OAI211_X1 U15387 ( .C1(n13720), .C2(n20152), .A(n13670), .B(n13950), .ZN(
        n13671) );
  INV_X1 U15388 ( .A(n13671), .ZN(n13676) );
  AOI22_X1 U15389 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13675) );
  AOI22_X1 U15390 ( .A1(n13672), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15391 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13673) );
  NAND4_X1 U15392 ( .A1(n13676), .A2(n13675), .A3(n13674), .A4(n13673), .ZN(
        n13685) );
  NAND2_X1 U15393 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13677) );
  OAI211_X1 U15394 ( .C1(n13720), .C2(n13678), .A(n13677), .B(n13694), .ZN(
        n13679) );
  INV_X1 U15395 ( .A(n13679), .ZN(n13683) );
  AOI22_X1 U15396 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13682) );
  AOI22_X1 U15397 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U15398 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13680) );
  NAND4_X1 U15399 ( .A1(n13683), .A2(n13682), .A3(n13681), .A4(n13680), .ZN(
        n13684) );
  AND2_X1 U15400 ( .A1(n13685), .A2(n13684), .ZN(n13916) );
  INV_X1 U15401 ( .A(n13916), .ZN(n13686) );
  NOR2_X1 U15402 ( .A1(n13914), .A2(n13686), .ZN(n13919) );
  NAND2_X1 U15403 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13687) );
  OAI211_X1 U15404 ( .C1(n13720), .C2(n13688), .A(n13687), .B(n13950), .ZN(
        n13689) );
  INV_X1 U15405 ( .A(n13689), .ZN(n13693) );
  AOI22_X1 U15406 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13692) );
  AOI22_X1 U15407 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13691) );
  AOI22_X1 U15408 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13690) );
  NAND4_X1 U15409 ( .A1(n13693), .A2(n13692), .A3(n13691), .A4(n13690), .ZN(
        n13703) );
  INV_X1 U15410 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U15411 ( .A1(n13626), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13695) );
  OAI211_X1 U15412 ( .C1(n13720), .C2(n13696), .A(n13695), .B(n13694), .ZN(
        n13697) );
  INV_X1 U15413 ( .A(n13697), .ZN(n13701) );
  AOI22_X1 U15414 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15415 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U15416 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13698) );
  NAND4_X1 U15417 ( .A1(n13701), .A2(n13700), .A3(n13699), .A4(n13698), .ZN(
        n13702) );
  AND2_X1 U15418 ( .A1(n13703), .A2(n13702), .ZN(n13920) );
  NAND2_X1 U15419 ( .A1(n13919), .A2(n13920), .ZN(n17070) );
  OAI22_X1 U15420 ( .A1(n13707), .A2(n13706), .B1(n11218), .B2(n13704), .ZN(
        n13718) );
  AOI22_X1 U15421 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13709) );
  AOI21_X1 U15422 ( .B1(n13952), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n13950), .ZN(n13708) );
  OAI211_X1 U15423 ( .C1(n13711), .C2(n13710), .A(n13709), .B(n13708), .ZN(
        n13717) );
  INV_X1 U15424 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13714) );
  OAI22_X1 U15425 ( .A1(n13715), .A2(n13714), .B1(n13713), .B2(n13712), .ZN(
        n13716) );
  NOR3_X1 U15426 ( .A1(n13718), .A2(n13717), .A3(n13716), .ZN(n13727) );
  INV_X1 U15427 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13719) );
  OAI21_X1 U15428 ( .B1(n13720), .B2(n13719), .A(n13950), .ZN(n13721) );
  AOI21_X1 U15429 ( .B1(n13626), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n13721), .ZN(n13725) );
  AOI22_X1 U15430 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13724) );
  AOI22_X1 U15431 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U15432 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n19079), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13722) );
  AND4_X1 U15433 ( .A1(n13725), .A2(n13724), .A3(n13723), .A4(n13722), .ZN(
        n13726) );
  NOR2_X1 U15434 ( .A1(n13727), .A2(n13726), .ZN(n17071) );
  INV_X1 U15435 ( .A(n17071), .ZN(n13728) );
  NOR3_X1 U15436 ( .A1(n17070), .A2(n20227), .A3(n13728), .ZN(n16435) );
  NOR2_X1 U15437 ( .A1(n13729), .A2(n19215), .ZN(n13735) );
  NAND2_X1 U15438 ( .A1(n12567), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13730) );
  AND2_X1 U15439 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19833) );
  NAND2_X1 U15440 ( .A1(n19833), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13750) );
  AOI21_X1 U15441 ( .B1(n13750), .B2(n19905), .A(n19953), .ZN(n13732) );
  INV_X1 U15442 ( .A(n13750), .ZN(n13731) );
  NAND2_X1 U15443 ( .A1(n13731), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19958) );
  AND2_X1 U15444 ( .A1(n13732), .A2(n19958), .ZN(n19781) );
  AOI21_X1 U15445 ( .B1(n13752), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19781), .ZN(n13733) );
  INV_X1 U15446 ( .A(n13733), .ZN(n13734) );
  NOR2_X2 U15447 ( .A1(n13735), .A2(n13734), .ZN(n13738) );
  NAND2_X1 U15448 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13737) );
  NAND2_X1 U15449 ( .A1(n13738), .A2(n13737), .ZN(n13739) );
  INV_X1 U15450 ( .A(n19833), .ZN(n19907) );
  OAI21_X1 U15451 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19907), .ZN(n19863) );
  NOR2_X1 U15452 ( .A1(n19863), .A2(n19953), .ZN(n19923) );
  AOI21_X1 U15453 ( .B1(n13752), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19923), .ZN(n13740) );
  OAI21_X1 U15454 ( .B1(n13741), .B2(n19215), .A(n13740), .ZN(n13742) );
  INV_X1 U15455 ( .A(n13742), .ZN(n14377) );
  INV_X1 U15456 ( .A(n19215), .ZN(n13743) );
  AOI22_X1 U15457 ( .A1(n13752), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19939), .B2(n19856), .ZN(n13744) );
  NAND2_X1 U15458 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13747) );
  NAND2_X1 U15459 ( .A1(n14350), .A2(n13747), .ZN(n13748) );
  NAND2_X1 U15460 ( .A1(n19907), .A2(n19906), .ZN(n13749) );
  NAND2_X1 U15461 ( .A1(n13750), .A2(n13749), .ZN(n19779) );
  NOR2_X1 U15462 ( .A1(n19779), .A2(n19953), .ZN(n13751) );
  AOI21_X1 U15463 ( .B1(n13752), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13751), .ZN(n13753) );
  NAND2_X1 U15464 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13754) );
  INV_X1 U15465 ( .A(n13754), .ZN(n13755) );
  NAND2_X1 U15466 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  NAND2_X1 U15467 ( .A1(n14461), .A2(n14462), .ZN(n13761) );
  NAND2_X1 U15468 ( .A1(n12567), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13758) );
  INV_X1 U15469 ( .A(n13918), .ZN(n13762) );
  INV_X1 U15470 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13807) );
  NOR2_X1 U15471 ( .A1(n13762), .A2(n13807), .ZN(n14426) );
  NAND2_X1 U15472 ( .A1(n14427), .A2(n14426), .ZN(n14421) );
  NAND2_X1 U15473 ( .A1(n13763), .A2(n11290), .ZN(n14465) );
  NOR2_X2 U15474 ( .A1(n14465), .A2(n13764), .ZN(n14605) );
  NAND2_X1 U15475 ( .A1(n14605), .A2(n14604), .ZN(n14603) );
  NAND2_X1 U15476 ( .A1(n13765), .A2(n14748), .ZN(n14858) );
  NOR2_X2 U15477 ( .A1(n14858), .A2(n13766), .ZN(n14859) );
  NAND2_X1 U15478 ( .A1(n11243), .A2(n15130), .ZN(n15129) );
  INV_X1 U15479 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13769) );
  INV_X1 U15480 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13768) );
  OAI22_X1 U15481 ( .A1(n13876), .A2(n13769), .B1(n13874), .B2(n13768), .ZN(
        n13770) );
  AOI21_X1 U15482 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n13770), .ZN(n13778) );
  INV_X1 U15483 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U15484 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13772) );
  NAND2_X1 U15485 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13771) );
  OAI211_X1 U15486 ( .C1(n13882), .C2(n13773), .A(n13772), .B(n13771), .ZN(
        n13774) );
  INV_X1 U15487 ( .A(n13774), .ZN(n13777) );
  AOI22_X1 U15488 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13776) );
  NAND2_X1 U15489 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13775) );
  NAND4_X1 U15490 ( .A1(n13778), .A2(n13777), .A3(n13776), .A4(n13775), .ZN(
        n13784) );
  AOI22_X1 U15491 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U15492 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U15493 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13780) );
  NAND2_X1 U15494 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13779) );
  NAND4_X1 U15495 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        n13783) );
  OR2_X1 U15496 ( .A1(n13784), .A2(n13783), .ZN(n15812) );
  INV_X1 U15497 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13786) );
  INV_X1 U15498 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13785) );
  OAI22_X1 U15499 ( .A1(n13876), .A2(n13786), .B1(n13874), .B2(n13785), .ZN(
        n13787) );
  AOI21_X1 U15500 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13787), .ZN(n13795) );
  INV_X1 U15501 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13790) );
  NAND2_X1 U15502 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13789) );
  NAND2_X1 U15503 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13788) );
  OAI211_X1 U15504 ( .C1(n13882), .C2(n13790), .A(n13789), .B(n13788), .ZN(
        n13791) );
  INV_X1 U15505 ( .A(n13791), .ZN(n13794) );
  AOI22_X1 U15506 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U15507 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13792) );
  NAND4_X1 U15508 ( .A1(n13795), .A2(n13794), .A3(n13793), .A4(n13792), .ZN(
        n13801) );
  AOI22_X1 U15509 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U15510 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U15511 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U15512 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13796) );
  NAND4_X1 U15513 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        n13800) );
  OR2_X1 U15514 ( .A1(n13801), .A2(n13800), .ZN(n15914) );
  INV_X1 U15515 ( .A(n15914), .ZN(n13872) );
  INV_X1 U15516 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13803) );
  INV_X1 U15517 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13802) );
  OAI22_X1 U15518 ( .A1(n13876), .A2(n13803), .B1(n13874), .B2(n13802), .ZN(
        n13804) );
  AOI21_X1 U15519 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n13804), .ZN(n13812) );
  NAND2_X1 U15520 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13806) );
  NAND2_X1 U15521 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13805) );
  OAI211_X1 U15522 ( .C1(n13882), .C2(n13807), .A(n13806), .B(n13805), .ZN(
        n13808) );
  INV_X1 U15523 ( .A(n13808), .ZN(n13811) );
  AOI22_X1 U15524 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U15525 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13809) );
  NAND4_X1 U15526 ( .A1(n13812), .A2(n13811), .A3(n13810), .A4(n13809), .ZN(
        n13818) );
  AOI22_X1 U15527 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U15528 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U15529 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U15530 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13813) );
  NAND4_X1 U15531 ( .A1(n13816), .A2(n13815), .A3(n13814), .A4(n13813), .ZN(
        n13817) );
  NOR2_X1 U15532 ( .A1(n13818), .A2(n13817), .ZN(n17107) );
  INV_X1 U15533 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13820) );
  INV_X1 U15534 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13819) );
  OAI22_X1 U15535 ( .A1(n13876), .A2(n13820), .B1(n13874), .B2(n13819), .ZN(
        n13821) );
  AOI21_X1 U15536 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n13821), .ZN(n13829) );
  INV_X1 U15537 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13824) );
  NAND2_X1 U15538 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13823) );
  NAND2_X1 U15539 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13822) );
  OAI211_X1 U15540 ( .C1(n13882), .C2(n13824), .A(n13823), .B(n13822), .ZN(
        n13825) );
  INV_X1 U15541 ( .A(n13825), .ZN(n13828) );
  AOI22_X1 U15542 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13827) );
  NAND2_X1 U15543 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13826) );
  NAND4_X1 U15544 ( .A1(n13829), .A2(n13828), .A3(n13827), .A4(n13826), .ZN(
        n13835) );
  AOI22_X1 U15545 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U15546 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U15547 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U15548 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13830) );
  NAND4_X1 U15549 ( .A1(n13833), .A2(n13832), .A3(n13831), .A4(n13830), .ZN(
        n13834) );
  NOR2_X1 U15550 ( .A1(n13835), .A2(n13834), .ZN(n17115) );
  INV_X1 U15551 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13837) );
  INV_X1 U15552 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13836) );
  OAI22_X1 U15553 ( .A1(n13876), .A2(n13837), .B1(n13874), .B2(n13836), .ZN(
        n13838) );
  AOI21_X1 U15554 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n13838), .ZN(n13846) );
  NAND2_X1 U15555 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13840) );
  NAND2_X1 U15556 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13839) );
  OAI211_X1 U15557 ( .C1(n13882), .C2(n13841), .A(n13840), .B(n13839), .ZN(
        n13842) );
  INV_X1 U15558 ( .A(n13842), .ZN(n13845) );
  AOI22_X1 U15559 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U15560 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13843) );
  NAND4_X1 U15561 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13843), .ZN(
        n13853) );
  AOI22_X1 U15562 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U15563 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U15564 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U15565 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13848) );
  NAND4_X1 U15566 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13852) );
  NOR2_X1 U15567 ( .A1(n13853), .A2(n13852), .ZN(n17118) );
  INV_X1 U15568 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13855) );
  INV_X1 U15569 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13854) );
  OAI22_X1 U15570 ( .A1(n13876), .A2(n13855), .B1(n13874), .B2(n13854), .ZN(
        n13856) );
  AOI21_X1 U15571 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n13856), .ZN(n13864) );
  INV_X1 U15572 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U15573 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13858) );
  NAND2_X1 U15574 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13857) );
  OAI211_X1 U15575 ( .C1(n13882), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        n13860) );
  INV_X1 U15576 ( .A(n13860), .ZN(n13863) );
  AOI22_X1 U15577 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U15578 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13861) );
  NAND4_X1 U15579 ( .A1(n13864), .A2(n13863), .A3(n13862), .A4(n13861), .ZN(
        n13871) );
  AOI22_X1 U15580 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U15581 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U15582 ( .A1(n13865), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13867) );
  NAND2_X1 U15583 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13866) );
  NAND4_X1 U15584 ( .A1(n13869), .A2(n13868), .A3(n13867), .A4(n13866), .ZN(
        n13870) );
  NOR2_X1 U15585 ( .A1(n13871), .A2(n13870), .ZN(n17135) );
  OR2_X1 U15586 ( .A1(n17118), .A2(n17135), .ZN(n17113) );
  OR2_X1 U15587 ( .A1(n17115), .A2(n17113), .ZN(n17104) );
  OR2_X1 U15588 ( .A1(n17107), .A2(n17104), .ZN(n15911) );
  NOR2_X1 U15589 ( .A1(n13872), .A2(n15911), .ZN(n15809) );
  AND2_X1 U15590 ( .A1(n15812), .A2(n15809), .ZN(n13899) );
  INV_X1 U15591 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13875) );
  INV_X1 U15592 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13873) );
  OAI22_X1 U15593 ( .A1(n13876), .A2(n13875), .B1(n13874), .B2(n13873), .ZN(
        n13877) );
  AOI21_X1 U15594 ( .B1(n13878), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n13877), .ZN(n13889) );
  NAND2_X1 U15595 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13881) );
  NAND2_X1 U15596 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13880) );
  OAI211_X1 U15597 ( .C1(n13882), .C2(n12717), .A(n13881), .B(n13880), .ZN(
        n13883) );
  INV_X1 U15598 ( .A(n13883), .ZN(n13888) );
  AOI22_X1 U15599 ( .A1(n12701), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U15600 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13886) );
  NAND4_X1 U15601 ( .A1(n13889), .A2(n13888), .A3(n13887), .A4(n13886), .ZN(
        n13898) );
  AOI22_X1 U15602 ( .A1(n11219), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12712), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U15603 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U15604 ( .A1(n13891), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13890), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13894) );
  NAND2_X1 U15605 ( .A1(n13892), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13893) );
  NAND4_X1 U15606 ( .A1(n13896), .A2(n13895), .A3(n13894), .A4(n13893), .ZN(
        n13897) );
  OR2_X1 U15607 ( .A1(n13898), .A2(n13897), .ZN(n15807) );
  AND2_X1 U15608 ( .A1(n13899), .A2(n15807), .ZN(n13900) );
  AND2_X1 U15609 ( .A1(n13900), .A2(n15703), .ZN(n13901) );
  XNOR2_X1 U15610 ( .A(n13903), .B(n13902), .ZN(n17100) );
  NAND2_X1 U15611 ( .A1(n13918), .A2(n13904), .ZN(n13908) );
  AOI22_X1 U15612 ( .A1(n13908), .A2(n13907), .B1(n13909), .B2(n19096), .ZN(
        n17096) );
  OAI211_X1 U15613 ( .C1(n13909), .C2(n13911), .A(n13914), .B(n13918), .ZN(
        n13913) );
  INV_X1 U15614 ( .A(n13913), .ZN(n13910) );
  INV_X1 U15615 ( .A(n13911), .ZN(n13912) );
  NOR2_X1 U15616 ( .A1(n19096), .A2(n13912), .ZN(n17086) );
  NAND2_X1 U15617 ( .A1(n17087), .A2(n17086), .ZN(n17085) );
  XNOR2_X1 U15618 ( .A(n13914), .B(n13916), .ZN(n13915) );
  NAND2_X1 U15619 ( .A1(n20227), .A2(n13916), .ZN(n17081) );
  NOR2_X2 U15620 ( .A1(n17082), .A2(n17081), .ZN(n17080) );
  NOR2_X2 U15621 ( .A1(n17080), .A2(n11276), .ZN(n13923) );
  OAI211_X1 U15622 ( .C1(n13919), .C2(n13920), .A(n17070), .B(n13918), .ZN(
        n13922) );
  INV_X1 U15623 ( .A(n13920), .ZN(n13921) );
  NOR2_X1 U15624 ( .A1(n19096), .A2(n13921), .ZN(n17077) );
  NAND2_X1 U15625 ( .A1(n13923), .A2(n13922), .ZN(n17075) );
  AOI22_X1 U15626 ( .A1(n13940), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13626), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U15627 ( .A1(n13941), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13925) );
  NAND2_X1 U15628 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13924) );
  NAND4_X1 U15629 ( .A1(n13926), .A2(n13925), .A3(n13924), .A4(n13950), .ZN(
        n13937) );
  AOI22_X1 U15630 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U15631 ( .A1(n19079), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U15632 ( .A1(n13928), .A2(n13927), .ZN(n13936) );
  INV_X1 U15633 ( .A(n19079), .ZN(n19084) );
  NOR2_X1 U15634 ( .A1(n19084), .A2(n13929), .ZN(n13930) );
  AOI211_X1 U15635 ( .C1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .C2(n13951), .A(
        n13950), .B(n13930), .ZN(n13934) );
  AOI22_X1 U15636 ( .A1(n13955), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U15637 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U15638 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13626), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13931) );
  NAND4_X1 U15639 ( .A1(n13934), .A2(n13933), .A3(n13932), .A4(n13931), .ZN(
        n13935) );
  OAI21_X1 U15640 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n13938) );
  NAND2_X1 U15641 ( .A1(n13939), .A2(n13938), .ZN(n16432) );
  NOR2_X1 U15642 ( .A1(n13939), .A2(n13938), .ZN(n16434) );
  AOI22_X1 U15643 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13626), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U15644 ( .A1(n19079), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13943) );
  NAND2_X1 U15645 ( .A1(n13941), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13942) );
  NAND4_X1 U15646 ( .A1(n13944), .A2(n13950), .A3(n13943), .A4(n13942), .ZN(
        n13962) );
  AOI22_X1 U15647 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13647), .B1(
        n13955), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U15648 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13954), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13946) );
  NAND2_X1 U15649 ( .A1(n13947), .A2(n13946), .ZN(n13961) );
  INV_X1 U15650 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13948) );
  NOR2_X1 U15651 ( .A1(n19084), .A2(n13948), .ZN(n13949) );
  AOI211_X1 U15652 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n13951), .A(
        n13950), .B(n13949), .ZN(n13959) );
  AOI22_X1 U15653 ( .A1(n12521), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13952), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U15654 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13954), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U15655 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13626), .B1(
        n13955), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13956) );
  NAND4_X1 U15656 ( .A1(n13959), .A2(n13958), .A3(n13957), .A4(n13956), .ZN(
        n13960) );
  OAI21_X1 U15657 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n13963) );
  XNOR2_X1 U15658 ( .A(n13964), .B(n13963), .ZN(n16446) );
  INV_X1 U15659 ( .A(n19192), .ZN(n13965) );
  NAND2_X1 U15660 ( .A1(n14274), .A2(n22264), .ZN(n19199) );
  NOR2_X1 U15661 ( .A1(n19202), .A2(n19199), .ZN(n13966) );
  AOI21_X1 U15662 ( .B1(n19197), .B2(n19185), .A(n13966), .ZN(n17611) );
  NAND2_X1 U15663 ( .A1(n17611), .A2(n13967), .ZN(n13968) );
  INV_X1 U15664 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17931) );
  AOI22_X1 U15665 ( .A1(n16414), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U15666 ( .B1(n13980), .B2(n17931), .A(n13969), .ZN(n17178) );
  NAND2_X1 U15667 ( .A1(n13970), .A2(n17178), .ZN(n17171) );
  NAND2_X1 U15668 ( .A1(n16415), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U15669 ( .A1(n16414), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13971) );
  AND2_X1 U15670 ( .A1(n13972), .A2(n13971), .ZN(n17172) );
  NOR2_X2 U15671 ( .A1(n17171), .A2(n17172), .ZN(n16937) );
  INV_X1 U15672 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19043) );
  AOI22_X1 U15673 ( .A1(n16414), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13973) );
  OAI21_X1 U15674 ( .B1(n13980), .B2(n19043), .A(n13973), .ZN(n17152) );
  INV_X1 U15675 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U15676 ( .A1(n16414), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13974) );
  OAI21_X1 U15677 ( .B1(n13980), .B2(n14238), .A(n13974), .ZN(n16919) );
  AND2_X1 U15678 ( .A1(n17152), .A2(n16919), .ZN(n13976) );
  INV_X1 U15679 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17933) );
  AOI22_X1 U15680 ( .A1(n16414), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13343), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13975) );
  OAI21_X1 U15681 ( .B1(n13980), .B2(n17933), .A(n13975), .ZN(n16938) );
  AND2_X1 U15682 ( .A1(n13976), .A2(n16938), .ZN(n13977) );
  AND2_X2 U15683 ( .A1(n16937), .A2(n13977), .ZN(n17155) );
  INV_X1 U15684 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U15685 ( .A1(n16414), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13345), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13978) );
  OAI21_X1 U15686 ( .B1(n13980), .B2(n17246), .A(n13978), .ZN(n16903) );
  NAND2_X1 U15687 ( .A1(n17155), .A2(n16903), .ZN(n16882) );
  INV_X1 U15688 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17935) );
  AOI22_X1 U15689 ( .A1(n16414), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13345), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13979) );
  OAI21_X1 U15690 ( .B1(n13980), .B2(n17935), .A(n13979), .ZN(n13981) );
  INV_X1 U15691 ( .A(n13981), .ZN(n16883) );
  AOI222_X1 U15692 ( .A1(n16415), .A2(P2_REIP_REG_28__SCAN_IN), .B1(n16414), 
        .B2(P2_EAX_REG_28__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C2(n13343), .ZN(n14263) );
  INV_X1 U15693 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19060) );
  AOI22_X1 U15694 ( .A1(n16414), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13345), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13982) );
  OAI21_X1 U15695 ( .B1(n13980), .B2(n19060), .A(n13982), .ZN(n16232) );
  AOI222_X1 U15696 ( .A1(n16415), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n16414), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), 
        .C2(n13345), .ZN(n16413) );
  INV_X1 U15697 ( .A(n16413), .ZN(n13984) );
  AND2_X1 U15698 ( .A1(n20026), .A2(n14347), .ZN(n13985) );
  NOR4_X1 U15699 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13989) );
  NOR4_X1 U15700 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13988) );
  NOR4_X1 U15701 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13987) );
  NOR4_X1 U15702 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13986) );
  NAND4_X1 U15703 ( .A1(n13989), .A2(n13988), .A3(n13987), .A4(n13986), .ZN(
        n13994) );
  NOR4_X1 U15704 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13992) );
  NOR4_X1 U15705 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13991) );
  NOR4_X1 U15706 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13990) );
  INV_X1 U15707 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17919) );
  NAND4_X1 U15708 ( .A1(n13992), .A2(n13991), .A3(n13990), .A4(n17919), .ZN(
        n13993) );
  OAI21_X1 U15709 ( .B1(n13994), .B2(n13993), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14531) );
  AOI22_X1 U15710 ( .A1(n19737), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19738), .ZN(n19713) );
  INV_X1 U15711 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n17915) );
  OAI22_X1 U15712 ( .A1(n20067), .A2(n19713), .B1(n20066), .B2(n17915), .ZN(
        n13995) );
  AOI21_X1 U15713 ( .B1(n20277), .B2(n11201), .A(n13995), .ZN(n13999) );
  INV_X1 U15714 ( .A(n13996), .ZN(n13997) );
  NAND2_X1 U15715 ( .A1(n20066), .A2(n13997), .ZN(n14489) );
  NOR2_X2 U15716 ( .A1(n14489), .A2(n19738), .ZN(n20169) );
  NOR2_X2 U15717 ( .A1(n14489), .A2(n19737), .ZN(n20170) );
  AOI22_X1 U15718 ( .A1(n20169), .A2(BUF1_REG_30__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U15719 ( .B1(n16446), .B2(n20222), .A(n14000), .ZN(P2_U2889) );
  AND2_X1 U15720 ( .A1(n20593), .A2(n16125), .ZN(n14001) );
  NOR2_X2 U15721 ( .A1(n14002), .A2(n14001), .ZN(n14014) );
  XNOR2_X1 U15722 ( .A(n16794), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14006) );
  INV_X1 U15723 ( .A(n14006), .ZN(n14004) );
  INV_X1 U15724 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14005) );
  AOI21_X1 U15725 ( .B1(n14005), .B2(n16125), .A(n20593), .ZN(n14010) );
  INV_X1 U15726 ( .A(n14010), .ZN(n14003) );
  NAND2_X1 U15727 ( .A1(n14004), .A2(n14003), .ZN(n14013) );
  NAND2_X1 U15728 ( .A1(n11597), .A2(n14005), .ZN(n14008) );
  NAND2_X1 U15729 ( .A1(n14014), .A2(n14007), .ZN(n14012) );
  INV_X1 U15730 ( .A(n14008), .ZN(n14009) );
  INV_X1 U15731 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16263) );
  OAI21_X1 U15732 ( .B1(n14010), .B2(n14009), .A(n16263), .ZN(n14011) );
  OAI211_X1 U15733 ( .C1(n14014), .C2(n14013), .A(n14012), .B(n14011), .ZN(
        n16266) );
  XNOR2_X1 U15734 ( .A(n14016), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14900) );
  INV_X1 U15735 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n16284) );
  NOR2_X1 U15736 ( .A1(n22016), .A2(n16284), .ZN(n16262) );
  AOI21_X1 U15737 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16262), .ZN(n14017) );
  OAI21_X1 U15738 ( .B1(n20633), .B2(n14900), .A(n14017), .ZN(n14018) );
  OAI21_X1 U15739 ( .B1(n16266), .B2(n22203), .A(n14019), .ZN(P1_U2968) );
  INV_X1 U15740 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20708) );
  INV_X1 U15741 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n15391) );
  NOR4_X1 U15742 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20708), .A4(n15391), .ZN(n14021) );
  NOR4_X1 U15743 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14020) );
  NAND3_X1 U15744 ( .A1(n15902), .A2(n14021), .A3(n14020), .ZN(U214) );
  NOR2_X1 U15745 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14023) );
  NOR4_X1 U15746 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14022) );
  NAND4_X1 U15747 ( .A1(n14023), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14022), .ZN(n14024) );
  OR2_X1 U15748 ( .A1(n19738), .A2(n14024), .ZN(n20640) );
  INV_X2 U15749 ( .A(U214), .ZN(n20693) );
  NOR2_X1 U15750 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14024), .ZN(n19275)
         );
  NAND2_X1 U15751 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18596) );
  INV_X1 U15752 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20871) );
  NOR2_X1 U15753 ( .A1(n18654), .A2(n20871), .ZN(n18649) );
  NAND4_X1 U15754 ( .A1(n18649), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20922) );
  NAND2_X1 U15755 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18697) );
  NAND3_X1 U15756 ( .A1(n20975), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18376), .ZN(n18353) );
  NAND2_X1 U15757 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18366) );
  NOR2_X2 U15758 ( .A1(n18353), .A2(n18366), .ZN(n21000) );
  CLKBUF_X1 U15759 ( .A(n14025), .Z(n18401) );
  INV_X1 U15760 ( .A(n18401), .ZN(n14026) );
  INV_X1 U15761 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14145) );
  INV_X1 U15762 ( .A(n14168), .ZN(n14167) );
  AOI21_X1 U15763 ( .B1(n14026), .B2(n14145), .A(n14167), .ZN(n18430) );
  AOI21_X1 U15764 ( .B1(n18327), .B2(n18400), .A(n18401), .ZN(n21028) );
  NAND2_X1 U15765 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18440) );
  NOR2_X4 U15766 ( .A1(n14168), .A2(n18440), .ZN(n18441) );
  INV_X1 U15767 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21073) );
  NAND2_X1 U15768 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18485) );
  NOR2_X4 U15769 ( .A1(n14163), .A2(n18485), .ZN(n14158) );
  NAND2_X2 U15770 ( .A1(n14158), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14159) );
  INV_X1 U15771 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21125) );
  INV_X1 U15772 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21150) );
  INV_X1 U15773 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21171) );
  XNOR2_X2 U15774 ( .A(n18552), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n18532) );
  INV_X1 U15775 ( .A(n21000), .ZN(n18575) );
  NOR2_X1 U15776 ( .A1(n18575), .A2(n18577), .ZN(n21014) );
  NAND2_X1 U15777 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n21014), .ZN(
        n18399) );
  INV_X1 U15778 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20892) );
  NAND2_X1 U15779 ( .A1(n20892), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20803) );
  NOR2_X1 U15780 ( .A1(n21027), .A2(n21151), .ZN(n14027) );
  NOR2_X1 U15781 ( .A1(n18430), .A2(n14027), .ZN(n14169) );
  INV_X1 U15782 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20711) );
  INV_X1 U15783 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22233) );
  NAND4_X1 U15784 ( .A1(n20715), .A2(n20711), .A3(n22233), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21882) );
  AOI211_X1 U15785 ( .C1(n18430), .C2(n14027), .A(n14169), .B(n21882), .ZN(
        n14153) );
  NOR3_X1 U15786 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20814) );
  INV_X1 U15787 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20813) );
  NAND2_X1 U15788 ( .A1(n20814), .A2(n20813), .ZN(n20818) );
  NOR2_X1 U15789 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20818), .ZN(n20840) );
  INV_X1 U15790 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U15791 ( .A1(n20840), .A2(n20847), .ZN(n20848) );
  INV_X1 U15792 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20867) );
  NAND2_X1 U15793 ( .A1(n20868), .A2(n20867), .ZN(n20878) );
  INV_X1 U15794 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20895) );
  NAND2_X1 U15795 ( .A1(n20893), .A2(n20895), .ZN(n20905) );
  INV_X1 U15796 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20933) );
  NAND2_X1 U15797 ( .A1(n20926), .A2(n20933), .ZN(n20934) );
  INV_X1 U15798 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20948) );
  NAND2_X1 U15799 ( .A1(n20946), .A2(n20948), .ZN(n20963) );
  INV_X1 U15800 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20971) );
  NAND2_X1 U15801 ( .A1(n20969), .A2(n20971), .ZN(n20984) );
  INV_X1 U15802 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21006) );
  NAND2_X1 U15803 ( .A1(n21004), .A2(n21006), .ZN(n21019) );
  INV_X1 U15804 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21032) );
  NAND2_X1 U15805 ( .A1(n21030), .A2(n21032), .ZN(n21029) );
  NAND2_X1 U15806 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21875) );
  INV_X2 U15807 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21403) );
  INV_X2 U15808 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21392) );
  AOI22_X1 U15809 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14042) );
  AOI22_X1 U15810 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14041) );
  INV_X1 U15811 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18159) );
  OR2_X2 U15812 ( .A1(n14031), .A2(n21404), .ZN(n18160) );
  INV_X2 U15813 ( .A(n18160), .ZN(n18234) );
  AOI22_X1 U15814 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18245), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14029) );
  OAI21_X1 U15815 ( .B1(n16062), .B2(n18159), .A(n14029), .ZN(n14039) );
  AOI22_X1 U15816 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14037) );
  INV_X2 U15817 ( .A(n15590), .ZN(n18006) );
  AOI22_X1 U15818 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14036) );
  INV_X2 U15819 ( .A(n18268), .ZN(n15556) );
  INV_X2 U15820 ( .A(n20790), .ZN(n21396) );
  NOR2_X4 U15821 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21396), .ZN(
        n18199) );
  AOI22_X1 U15822 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14035) );
  NOR2_X2 U15823 ( .A1(n21412), .A2(n14033), .ZN(n18279) );
  NOR2_X2 U15824 ( .A1(n21848), .A2(n21396), .ZN(n14066) );
  BUF_X2 U15825 ( .A(n14066), .Z(n18247) );
  AOI22_X1 U15826 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14034) );
  NAND4_X1 U15827 ( .A1(n14037), .A2(n14036), .A3(n14035), .A4(n14034), .ZN(
        n14038) );
  AOI211_X1 U15828 ( .C1(n18051), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n14039), .B(n14038), .ZN(n14040) );
  NAND3_X1 U15829 ( .A1(n14042), .A2(n14041), .A3(n14040), .ZN(n16010) );
  AOI22_X1 U15830 ( .A1(n18245), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U15831 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U15832 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U15833 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n21408), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14044) );
  NAND4_X1 U15834 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        n14053) );
  AOI22_X1 U15835 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U15836 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U15837 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U15838 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U15839 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14052) );
  AOI22_X1 U15840 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U15841 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14056) );
  AOI22_X1 U15842 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18279), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U15843 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14054) );
  NAND4_X1 U15844 ( .A1(n14057), .A2(n14056), .A3(n14055), .A4(n14054), .ZN(
        n14063) );
  AOI22_X1 U15845 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14061) );
  INV_X2 U15846 ( .A(n16022), .ZN(n18003) );
  AOI22_X1 U15847 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U15848 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U15849 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U15850 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14062) );
  AOI22_X1 U15851 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U15852 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U15853 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14065) );
  OAI21_X1 U15854 ( .B1(n16062), .B2(n18233), .A(n14065), .ZN(n14072) );
  AOI22_X1 U15855 ( .A1(n14043), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U15856 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U15857 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U15858 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14067) );
  NAND4_X1 U15859 ( .A1(n14070), .A2(n14069), .A3(n14068), .A4(n14067), .ZN(
        n14071) );
  AOI22_X1 U15860 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U15861 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U15862 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n21408), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U15863 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14076) );
  NAND4_X1 U15864 ( .A1(n14079), .A2(n14078), .A3(n14077), .A4(n14076), .ZN(
        n14085) );
  AOI22_X1 U15865 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U15866 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14082) );
  INV_X2 U15867 ( .A(n18160), .ZN(n18076) );
  AOI22_X1 U15868 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U15869 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U15870 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14084) );
  AOI22_X1 U15871 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U15872 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U15873 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14086) );
  OAI21_X1 U15874 ( .B1(n16062), .B2(n18267), .A(n14086), .ZN(n14094) );
  AOI22_X1 U15875 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U15876 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U15877 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U15878 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14089) );
  NAND4_X1 U15879 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14093) );
  AOI22_X1 U15880 ( .A1(n18245), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14101) );
  AOI22_X1 U15881 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U15882 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U15883 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18279), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14098) );
  NAND4_X1 U15884 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        n14107) );
  AOI22_X1 U15885 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U15886 ( .A1(n14108), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18262), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U15887 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U15888 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14102) );
  NAND4_X1 U15889 ( .A1(n14105), .A2(n14104), .A3(n14103), .A4(n14102), .ZN(
        n14106) );
  NAND2_X1 U15890 ( .A1(n18802), .A2(n19560), .ZN(n15543) );
  NOR2_X1 U15891 ( .A1(n21252), .A2(n19358), .ZN(n21378) );
  NOR2_X1 U15892 ( .A1(n21366), .A2(n21378), .ZN(n21195) );
  AOI22_X1 U15893 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U15894 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14117) );
  INV_X1 U15895 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18062) );
  AOI22_X1 U15896 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14109) );
  OAI21_X1 U15897 ( .B1(n16062), .B2(n18062), .A(n14109), .ZN(n14115) );
  AOI22_X1 U15898 ( .A1(n14043), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U15899 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U15900 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15901 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14110) );
  NAND4_X1 U15902 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        n14114) );
  AOI211_X1 U15903 ( .C1(n18272), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n14115), .B(n14114), .ZN(n14116) );
  NAND3_X1 U15904 ( .A1(n14118), .A2(n14117), .A3(n14116), .ZN(n14128) );
  NOR2_X1 U15905 ( .A1(n21252), .A2(n14128), .ZN(n15544) );
  NAND2_X1 U15906 ( .A1(n19519), .A2(n14120), .ZN(n15530) );
  AOI221_X1 U15907 ( .B1(n15544), .B2(n14126), .C1(n14129), .C2(n14126), .A(
        n14119), .ZN(n14125) );
  NAND2_X1 U15908 ( .A1(n21252), .A2(n19358), .ZN(n15525) );
  AOI21_X1 U15909 ( .B1(n19610), .B2(n19519), .A(n21378), .ZN(n15531) );
  NOR2_X1 U15910 ( .A1(n14120), .A2(n19358), .ZN(n21390) );
  NOR3_X1 U15911 ( .A1(n14127), .A2(n15531), .A3(n21390), .ZN(n14124) );
  NOR2_X1 U15912 ( .A1(n21366), .A2(n15536), .ZN(n14122) );
  NAND2_X1 U15913 ( .A1(n19610), .A2(n20710), .ZN(n15542) );
  NAND2_X1 U15914 ( .A1(n19519), .A2(n15542), .ZN(n15527) );
  INV_X1 U15915 ( .A(n15527), .ZN(n14121) );
  OAI22_X1 U15916 ( .A1(n14120), .A2(n14122), .B1(n15536), .B2(n14121), .ZN(
        n14123) );
  NOR4_X4 U15917 ( .A1(n15524), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n21410) );
  NAND2_X1 U15918 ( .A1(n19560), .A2(n19610), .ZN(n21192) );
  NOR2_X1 U15919 ( .A1(n21192), .A2(n21366), .ZN(n14130) );
  NAND2_X1 U15920 ( .A1(n15541), .A2(n14128), .ZN(n18224) );
  NAND2_X1 U15921 ( .A1(n21410), .A2(n15608), .ZN(n15540) );
  INV_X1 U15922 ( .A(n15540), .ZN(n21388) );
  NOR2_X1 U15923 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20715), .ZN(n21878) );
  NAND2_X1 U15924 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21878), .ZN(n21897) );
  NAND2_X1 U15925 ( .A1(n21852), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15518) );
  OAI22_X1 U15926 ( .A1(n21851), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21861), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14137) );
  OAI22_X1 U15927 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21865), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14134), .ZN(n14140) );
  NOR2_X1 U15928 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21865), .ZN(
        n14135) );
  NAND2_X1 U15929 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14134), .ZN(
        n14139) );
  AOI22_X1 U15930 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14140), .B1(
        n14135), .B2(n14139), .ZN(n15522) );
  OAI21_X1 U15931 ( .B1(n14138), .B2(n14137), .A(n15522), .ZN(n14136) );
  XOR2_X1 U15932 ( .A(n15518), .B(n15519), .Z(n14142) );
  OAI22_X1 U15933 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21846), .B1(
        n14141), .B2(n14140), .ZN(n15520) );
  NAND2_X1 U15934 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20710), .ZN(n14143) );
  AOI211_X4 U15935 ( .C1(n21875), .C2(n22233), .A(n14146), .B(n14143), .ZN(
        n21185) );
  AOI211_X1 U15936 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21029), .A(n21044), .B(
        n21160), .ZN(n14152) );
  INV_X1 U15937 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18746) );
  NAND2_X1 U15938 ( .A1(n18746), .A2(n20711), .ZN(n20714) );
  INV_X1 U15939 ( .A(n20714), .ZN(n21888) );
  NAND2_X1 U15940 ( .A1(n21888), .A2(n21885), .ZN(n18227) );
  OR2_X2 U15941 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18227), .ZN(n21808) );
  NAND2_X1 U15942 ( .A1(n20711), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21876) );
  INV_X1 U15943 ( .A(n21876), .ZN(n19347) );
  NAND2_X1 U15944 ( .A1(n21878), .A2(n19347), .ZN(n21894) );
  INV_X1 U15945 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n21169) );
  INV_X2 U15946 ( .A(n18842), .ZN(n22240) );
  INV_X1 U15947 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22287) );
  OAI211_X1 U15948 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n18839), .B(n22287), .ZN(n16116) );
  INV_X1 U15949 ( .A(n16116), .ZN(n20709) );
  OAI211_X1 U15950 ( .C1(n20709), .C2(n20710), .A(n21875), .B(n22233), .ZN(
        n21873) );
  OAI211_X2 U15951 ( .C1(n21169), .C2(n19560), .A(n21873), .B(n14144), .ZN(
        n21168) );
  INV_X1 U15952 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n18171) );
  OAI22_X1 U15953 ( .A1(n14145), .A2(n21170), .B1(n21168), .B2(n18171), .ZN(
        n14151) );
  NAND2_X1 U15954 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n21035) );
  INV_X1 U15955 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20993) );
  INV_X1 U15956 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21010) );
  INV_X1 U15957 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20986) );
  INV_X1 U15958 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20962) );
  INV_X1 U15959 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21535) );
  INV_X1 U15960 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21830) );
  INV_X1 U15961 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20877) );
  INV_X1 U15962 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20834) );
  INV_X1 U15963 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20801) );
  INV_X1 U15964 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20788) );
  INV_X1 U15965 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20787) );
  NOR2_X1 U15966 ( .A1(n20788), .A2(n20787), .ZN(n20786) );
  INV_X1 U15967 ( .A(n20786), .ZN(n20802) );
  NOR2_X1 U15968 ( .A1(n20801), .A2(n20802), .ZN(n20820) );
  NAND2_X1 U15969 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20820), .ZN(n20835) );
  NOR2_X1 U15970 ( .A1(n20834), .A2(n20835), .ZN(n20850) );
  NAND2_X1 U15971 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20850), .ZN(n20865) );
  NOR2_X1 U15972 ( .A1(n20877), .A2(n20865), .ZN(n20880) );
  NAND2_X1 U15973 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20880), .ZN(n20890) );
  NOR2_X1 U15974 ( .A1(n21830), .A2(n20890), .ZN(n20904) );
  NAND2_X1 U15975 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20904), .ZN(n20920) );
  NAND3_X1 U15976 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .A3(n21067), .ZN(n20961) );
  NOR4_X1 U15977 ( .A1(n20993), .A2(n21010), .A3(n20986), .A4(n21052), .ZN(
        n21036) );
  INV_X1 U15978 ( .A(n21036), .ZN(n21026) );
  NOR2_X1 U15979 ( .A1(n21035), .A2(n21026), .ZN(n14149) );
  INV_X1 U15980 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18833) );
  NAND3_X1 U15981 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n20999) );
  NOR3_X1 U15982 ( .A1(n18833), .A2(n20999), .A3(n21035), .ZN(n21050) );
  INV_X1 U15983 ( .A(n21050), .ZN(n14147) );
  INV_X1 U15984 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20954) );
  INV_X1 U15985 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20953) );
  NOR3_X1 U15986 ( .A1(n20962), .A2(n20954), .A3(n20953), .ZN(n14154) );
  NOR2_X1 U15987 ( .A1(n21535), .A2(n20920), .ZN(n20919) );
  NAND3_X1 U15988 ( .A1(n14154), .A2(n20919), .A3(n21184), .ZN(n20998) );
  NAND2_X1 U15989 ( .A1(n21081), .A2(n21184), .ZN(n21183) );
  OAI21_X1 U15990 ( .B1(n14147), .B2(n20998), .A(n21183), .ZN(n21064) );
  INV_X1 U15991 ( .A(n21064), .ZN(n14148) );
  MUX2_X1 U15992 ( .A(n14149), .B(n14148), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n14150) );
  INV_X1 U15993 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21046) );
  NAND2_X1 U15994 ( .A1(n21044), .A2(n21046), .ZN(n21057) );
  INV_X1 U15995 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21076) );
  NAND2_X1 U15996 ( .A1(n21077), .A2(n21076), .ZN(n21083) );
  NOR2_X1 U15997 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21083), .ZN(n21100) );
  INV_X1 U15998 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21099) );
  NAND2_X1 U15999 ( .A1(n21100), .A2(n21099), .ZN(n21110) );
  NOR2_X1 U16000 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21110), .ZN(n21130) );
  INV_X1 U16001 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21129) );
  NAND2_X1 U16002 ( .A1(n21130), .A2(n21129), .ZN(n21128) );
  NOR2_X1 U16003 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21128), .ZN(n21141) );
  AOI211_X1 U16004 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21128), .A(n21141), .B(
        n21160), .ZN(n14175) );
  INV_X1 U16005 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21136) );
  INV_X1 U16006 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18838) );
  INV_X1 U16007 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21066) );
  NAND2_X1 U16008 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n21050), .ZN(n21053) );
  INV_X1 U16009 ( .A(n14154), .ZN(n14155) );
  NOR3_X1 U16010 ( .A1(n21066), .A2(n21053), .A3(n14155), .ZN(n21068) );
  NAND3_X1 U16011 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20919), .A3(n21068), 
        .ZN(n21069) );
  NOR2_X1 U16012 ( .A1(n18838), .A2(n21069), .ZN(n21102) );
  AND2_X1 U16013 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21102), .ZN(n21109) );
  NAND2_X1 U16014 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21109), .ZN(n21124) );
  INV_X1 U16015 ( .A(n21124), .ZN(n14156) );
  NOR2_X1 U16016 ( .A1(n14156), .A2(n21081), .ZN(n21108) );
  NOR2_X1 U16017 ( .A1(n20879), .A2(n21108), .ZN(n21134) );
  INV_X1 U16018 ( .A(n21134), .ZN(n21116) );
  NOR2_X1 U16019 ( .A1(n21136), .A2(n21116), .ZN(n21137) );
  INV_X1 U16020 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21133) );
  NAND2_X1 U16021 ( .A1(n21103), .A2(n21133), .ZN(n21123) );
  NAND3_X1 U16022 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21103), .A3(n14156), 
        .ZN(n21135) );
  AOI22_X1 U16023 ( .A1(n21137), .A2(n21123), .B1(n21136), .B2(n21135), .ZN(
        n14174) );
  OAI21_X1 U16024 ( .B1(n14157), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n18568), .ZN(n18491) );
  INV_X1 U16025 ( .A(n18491), .ZN(n14171) );
  AOI21_X1 U16026 ( .B1(n14159), .B2(n21125), .A(n14157), .ZN(n21122) );
  OAI21_X1 U16027 ( .B1(n14158), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14159), .ZN(n14160) );
  INV_X1 U16028 ( .A(n14160), .ZN(n21113) );
  INV_X1 U16029 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U16030 ( .A1(n18458), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14161) );
  AOI21_X1 U16031 ( .B1(n14162), .B2(n14161), .A(n14158), .ZN(n21095) );
  INV_X1 U16032 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21091) );
  OAI22_X1 U16033 ( .A1(n14163), .A2(n21091), .B1(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18458), .ZN(n18475) );
  INV_X1 U16034 ( .A(n18475), .ZN(n21086) );
  INV_X1 U16035 ( .A(n18441), .ZN(n14164) );
  AOI21_X1 U16036 ( .B1(n14164), .B2(n21073), .A(n18458), .ZN(n21072) );
  INV_X1 U16037 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14166) );
  NAND2_X1 U16038 ( .A1(n14167), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14165) );
  AOI21_X1 U16039 ( .B1(n14166), .B2(n14165), .A(n18441), .ZN(n21056) );
  INV_X1 U16040 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18416) );
  OAI22_X1 U16041 ( .A1(n14168), .A2(n18416), .B1(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n14167), .ZN(n18413) );
  INV_X1 U16042 ( .A(n18413), .ZN(n21043) );
  NOR2_X1 U16043 ( .A1(n14169), .A2(n21151), .ZN(n21042) );
  NOR2_X1 U16044 ( .A1(n21043), .A2(n21042), .ZN(n21041) );
  NOR2_X1 U16045 ( .A1(n21041), .A2(n21151), .ZN(n21055) );
  NOR2_X1 U16046 ( .A1(n21056), .A2(n21055), .ZN(n21054) );
  NOR2_X1 U16047 ( .A1(n21054), .A2(n21151), .ZN(n21071) );
  NOR2_X1 U16048 ( .A1(n21072), .A2(n21071), .ZN(n21070) );
  NOR2_X1 U16049 ( .A1(n21070), .A2(n21151), .ZN(n21085) );
  NOR2_X1 U16050 ( .A1(n21086), .A2(n21085), .ZN(n21084) );
  NOR2_X1 U16051 ( .A1(n21084), .A2(n21151), .ZN(n21094) );
  NOR2_X1 U16052 ( .A1(n21095), .A2(n21094), .ZN(n21093) );
  NOR2_X1 U16053 ( .A1(n21093), .A2(n21151), .ZN(n21112) );
  NOR2_X1 U16054 ( .A1(n21113), .A2(n21112), .ZN(n21111) );
  NOR2_X1 U16055 ( .A1(n21111), .A2(n21151), .ZN(n21121) );
  NOR2_X1 U16056 ( .A1(n21122), .A2(n21121), .ZN(n21120) );
  NOR2_X1 U16057 ( .A1(n21120), .A2(n21151), .ZN(n14170) );
  NOR2_X1 U16058 ( .A1(n14171), .A2(n14170), .ZN(n21143) );
  AOI211_X1 U16059 ( .C1(n14171), .C2(n14170), .A(n21143), .B(n21882), .ZN(
        n14173) );
  INV_X1 U16060 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18489) );
  INV_X1 U16061 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18119) );
  OAI22_X1 U16062 ( .A1(n18489), .A2(n21170), .B1(n21168), .B2(n18119), .ZN(
        n14172) );
  OR4_X1 U16063 ( .A1(n14175), .A2(n14174), .A3(n14173), .A4(n14172), .ZN(
        P3_U2643) );
  INV_X1 U16064 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17271) );
  INV_X1 U16065 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19005) );
  INV_X1 U16066 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19044) );
  INV_X1 U16067 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16886) );
  INV_X1 U16068 ( .A(n14217), .ZN(n14177) );
  INV_X1 U16069 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14176) );
  OAI21_X1 U16070 ( .B1(n14177), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16852), .ZN(n17222) );
  INV_X1 U16071 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16423) );
  INV_X1 U16072 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n19062) );
  OAI21_X1 U16073 ( .B1(n14212), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14215), .ZN(n16897) );
  INV_X1 U16074 ( .A(n16897), .ZN(n17253) );
  OAI21_X1 U16075 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14209), .A(
        n14213), .ZN(n17826) );
  INV_X1 U16076 ( .A(n17826), .ZN(n14211) );
  OAI21_X1 U16077 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14206), .A(
        n14210), .ZN(n19026) );
  INV_X1 U16078 ( .A(n19026), .ZN(n14208) );
  INV_X1 U16079 ( .A(n14179), .ZN(n16951) );
  OAI21_X1 U16080 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14201), .A(
        n14205), .ZN(n17805) );
  INV_X1 U16081 ( .A(n17805), .ZN(n18980) );
  OAI21_X1 U16082 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14198), .A(
        n14202), .ZN(n17787) );
  INV_X1 U16083 ( .A(n17787), .ZN(n14200) );
  OAI21_X1 U16084 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14196), .A(
        n14199), .ZN(n17775) );
  INV_X1 U16085 ( .A(n17775), .ZN(n18944) );
  INV_X1 U16086 ( .A(n16973), .ZN(n14195) );
  OAI21_X1 U16087 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14180), .A(
        n14193), .ZN(n18900) );
  INV_X1 U16088 ( .A(n18900), .ZN(n14191) );
  AOI21_X1 U16089 ( .B1(n17751), .B2(n14187), .A(n14190), .ZN(n17740) );
  AOI21_X1 U16090 ( .B1(n15765), .B2(n14185), .A(n14188), .ZN(n18880) );
  AOI21_X1 U16091 ( .B1(n17027), .B2(n14183), .A(n14186), .ZN(n17025) );
  AOI21_X1 U16092 ( .B1(n17059), .B2(n14373), .A(n14184), .ZN(n17047) );
  AOI22_X1 U16093 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19237), .ZN(n14181) );
  INV_X1 U16094 ( .A(n14181), .ZN(n18870) );
  INV_X1 U16095 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14182) );
  OAI22_X1 U16096 ( .A1(n19237), .A2(n14182), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n17058) );
  OR2_X1 U16097 ( .A1(n18870), .A2(n17058), .ZN(n17046) );
  NOR2_X1 U16098 ( .A1(n17047), .A2(n17046), .ZN(n17035) );
  OAI21_X1 U16099 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14184), .A(
        n14183), .ZN(n17036) );
  NAND2_X1 U16100 ( .A1(n17035), .A2(n17036), .ZN(n17022) );
  NOR2_X1 U16101 ( .A1(n17025), .A2(n17022), .ZN(n17013) );
  OAI21_X1 U16102 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14186), .A(
        n14185), .ZN(n17739) );
  NAND2_X1 U16103 ( .A1(n17013), .A2(n17739), .ZN(n18878) );
  NOR2_X1 U16104 ( .A1(n18880), .A2(n18878), .ZN(n18886) );
  OAI21_X1 U16105 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14188), .A(
        n14187), .ZN(n18888) );
  NAND2_X1 U16106 ( .A1(n18886), .A2(n18888), .ZN(n16996) );
  NOR2_X1 U16107 ( .A1(n17740), .A2(n16996), .ZN(n16985) );
  OAI21_X1 U16108 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n14190), .A(
        n14189), .ZN(n17334) );
  NAND2_X1 U16109 ( .A1(n16985), .A2(n17334), .ZN(n18899) );
  NOR2_X1 U16110 ( .A1(n14191), .A2(n18899), .ZN(n18922) );
  AOI21_X1 U16111 ( .B1(n18913), .B2(n14193), .A(n14192), .ZN(n14194) );
  INV_X1 U16112 ( .A(n14194), .ZN(n18925) );
  NAND2_X1 U16113 ( .A1(n18922), .A2(n18925), .ZN(n18921) );
  NOR2_X1 U16114 ( .A1(n14195), .A2(n18921), .ZN(n18939) );
  AOI21_X1 U16115 ( .B1(n18930), .B2(n14197), .A(n14196), .ZN(n18933) );
  INV_X1 U16116 ( .A(n18933), .ZN(n18938) );
  NAND2_X1 U16117 ( .A1(n18939), .A2(n18938), .ZN(n18942) );
  NOR2_X1 U16118 ( .A1(n18944), .A2(n18942), .ZN(n18953) );
  AOI21_X1 U16119 ( .B1(n17784), .B2(n14199), .A(n14198), .ZN(n17776) );
  INV_X1 U16120 ( .A(n17776), .ZN(n18954) );
  NAND2_X1 U16121 ( .A1(n18953), .A2(n18954), .ZN(n16959) );
  NOR2_X1 U16122 ( .A1(n14200), .A2(n16959), .ZN(n18966) );
  AOI21_X1 U16123 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n17311) );
  INV_X1 U16124 ( .A(n17311), .ZN(n18968) );
  NAND2_X1 U16125 ( .A1(n18966), .A2(n18968), .ZN(n18978) );
  NOR2_X1 U16126 ( .A1(n18980), .A2(n18978), .ZN(n18992) );
  AOI21_X1 U16127 ( .B1(n17297), .B2(n14205), .A(n14204), .ZN(n17300) );
  INV_X1 U16128 ( .A(n17300), .ZN(n18994) );
  NAND2_X1 U16129 ( .A1(n18992), .A2(n18994), .ZN(n16949) );
  NOR2_X1 U16130 ( .A1(n16951), .A2(n16949), .ZN(n19015) );
  AOI21_X1 U16131 ( .B1(n14207), .B2(n19005), .A(n14206), .ZN(n19019) );
  INV_X1 U16132 ( .A(n19019), .ZN(n19017) );
  NAND2_X1 U16133 ( .A1(n19015), .A2(n19017), .ZN(n19023) );
  NOR2_X1 U16134 ( .A1(n14208), .A2(n19023), .ZN(n16929) );
  AOI21_X1 U16135 ( .B1(n17271), .B2(n14210), .A(n14209), .ZN(n16932) );
  INV_X1 U16136 ( .A(n16932), .ZN(n17274) );
  NAND2_X1 U16137 ( .A1(n16929), .A2(n17274), .ZN(n16912) );
  NOR2_X1 U16138 ( .A1(n14211), .A2(n16912), .ZN(n19039) );
  AOI21_X1 U16139 ( .B1(n19044), .B2(n14213), .A(n14212), .ZN(n19042) );
  INV_X1 U16140 ( .A(n19042), .ZN(n14214) );
  NAND2_X1 U16141 ( .A1(n19039), .A2(n14214), .ZN(n16894) );
  NOR2_X1 U16142 ( .A1(n17253), .A2(n16894), .ZN(n16875) );
  NAND2_X1 U16143 ( .A1(n14215), .A2(n16886), .ZN(n14216) );
  AND2_X1 U16144 ( .A1(n14217), .A2(n14216), .ZN(n17233) );
  INV_X1 U16145 ( .A(n17233), .ZN(n14218) );
  NAND2_X1 U16146 ( .A1(n16875), .A2(n14218), .ZN(n16849) );
  NAND2_X1 U16147 ( .A1(n11223), .A2(n16849), .ZN(n14220) );
  NAND4_X1 U16148 ( .A1(n19237), .A2(n19835), .A3(n22228), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19230) );
  OAI21_X1 U16149 ( .B1(n17222), .B2(n14220), .A(n19055), .ZN(n14219) );
  AOI21_X1 U16150 ( .B1(n17222), .B2(n14220), .A(n14219), .ZN(n14272) );
  INV_X1 U16151 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n19006) );
  NOR2_X1 U16152 ( .A1(n16391), .A2(n19006), .ZN(n16156) );
  NAND2_X1 U16153 ( .A1(n20026), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16181) );
  INV_X1 U16154 ( .A(n16181), .ZN(n14221) );
  NAND2_X1 U16155 ( .A1(n20026), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U16156 ( .A1(n20026), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U16157 ( .A1(n20026), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16195) );
  INV_X1 U16158 ( .A(n16192), .ZN(n14224) );
  INV_X1 U16159 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16904) );
  NOR2_X1 U16160 ( .A1(n16391), .A2(n16904), .ZN(n16191) );
  INV_X1 U16161 ( .A(n16191), .ZN(n14223) );
  NAND2_X1 U16162 ( .A1(n20026), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16199) );
  INV_X1 U16163 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14225) );
  NOR2_X1 U16164 ( .A1(n16391), .A2(n14225), .ZN(n14226) );
  NAND2_X1 U16165 ( .A1(n16203), .A2(n14226), .ZN(n14227) );
  NAND2_X1 U16166 ( .A1(n16353), .A2(n14227), .ZN(n16205) );
  NAND2_X1 U16167 ( .A1(n14228), .A2(n18852), .ZN(n14229) );
  INV_X1 U16168 ( .A(n14230), .ZN(n19098) );
  NAND2_X1 U16169 ( .A1(n19098), .A2(n18852), .ZN(n17665) );
  NAND2_X1 U16170 ( .A1(n14502), .A2(n17067), .ZN(n17731) );
  NOR2_X1 U16171 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n22275), .ZN(n14264) );
  INV_X1 U16172 ( .A(n14264), .ZN(n14231) );
  AND3_X1 U16173 ( .A1(n14261), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n14231), .ZN(
        n14232) );
  NAND2_X1 U16174 ( .A1(n17731), .A2(n14232), .ZN(n18996) );
  NOR2_X1 U16175 ( .A1(n16205), .A2(n18996), .ZN(n14271) );
  NOR4_X1 U16176 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n19237), .A4(n19834), .ZN(n19240) );
  INV_X1 U16177 ( .A(n19240), .ZN(n14233) );
  NAND3_X1 U16178 ( .A1(n19230), .A2(n17323), .A3(n14233), .ZN(n14234) );
  NAND2_X1 U16179 ( .A1(n19059), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19061) );
  AOI22_X1 U16180 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19009), .ZN(n14235) );
  INV_X1 U16181 ( .A(n14235), .ZN(n14270) );
  NAND2_X1 U16182 ( .A1(n12975), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14241) );
  NAND2_X1 U16183 ( .A1(n11221), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14237) );
  NAND2_X1 U16184 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14236) );
  OAI211_X1 U16185 ( .C1(n16236), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14239) );
  INV_X1 U16186 ( .A(n14239), .ZN(n14240) );
  NAND2_X1 U16187 ( .A1(n14241), .A2(n14240), .ZN(n16916) );
  NAND2_X1 U16188 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14243) );
  AOI22_X1 U16189 ( .A1(n16401), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n14242) );
  OAI211_X1 U16190 ( .C1(n16236), .C2(n17931), .A(n14243), .B(n14242), .ZN(
        n15917) );
  AND2_X2 U16191 ( .A1(n14244), .A2(n15917), .ZN(n15915) );
  INV_X1 U16192 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U16193 ( .A1(n12975), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14246) );
  AOI22_X1 U16194 ( .A1(n16401), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n14245) );
  OAI211_X1 U16195 ( .C1(n16236), .C2(n19031), .A(n14246), .B(n14245), .ZN(
        n15813) );
  NAND2_X1 U16196 ( .A1(n11221), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U16197 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14247) );
  OAI211_X1 U16198 ( .C1(n16236), .C2(n17933), .A(n14248), .B(n14247), .ZN(
        n14249) );
  AOI21_X1 U16199 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14249), .ZN(n16936) );
  NAND2_X1 U16200 ( .A1(n11194), .A2(n11196), .ZN(n17088) );
  NAND2_X1 U16201 ( .A1(n16401), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U16202 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14250) );
  OAI211_X1 U16203 ( .C1(n16236), .C2(n19043), .A(n14251), .B(n14250), .ZN(
        n14252) );
  AOI21_X1 U16204 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14252), .ZN(n17089) );
  OR2_X2 U16205 ( .A1(n17088), .A2(n17089), .ZN(n17090) );
  NAND2_X1 U16206 ( .A1(n11221), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U16207 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14253) );
  OAI211_X1 U16208 ( .C1(n16236), .C2(n17246), .A(n14254), .B(n14253), .ZN(
        n14255) );
  AOI21_X1 U16209 ( .B1(n12975), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14255), .ZN(n16900) );
  NAND2_X1 U16210 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14257) );
  AOI22_X1 U16211 ( .A1(n11221), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n14256) );
  OAI211_X1 U16212 ( .C1(n16236), .C2(n17935), .A(n14257), .B(n14256), .ZN(
        n16879) );
  INV_X1 U16213 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17219) );
  NAND2_X1 U16214 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14259) );
  AOI22_X1 U16215 ( .A1(n11221), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n14258) );
  OAI211_X1 U16216 ( .C1(n16236), .C2(n17219), .A(n14259), .B(n14258), .ZN(
        n16237) );
  NOR2_X1 U16217 ( .A1(n16881), .A2(n16237), .ZN(n14260) );
  AND3_X1 U16218 ( .A1(n14261), .A2(n22264), .A3(n22228), .ZN(n14262) );
  AOI21_X1 U16219 ( .B1(n14263), .B2(n16885), .A(n16233), .ZN(n17355) );
  NOR2_X1 U16220 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14266), .ZN(n19218) );
  OAI21_X1 U16221 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(n14264), .A(n19096), .ZN(
        n14265) );
  OAI21_X1 U16222 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n14266), .A(n14265), 
        .ZN(n14267) );
  AOI22_X1 U16223 ( .A1(n17355), .A2(n18916), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n11144), .ZN(n14268) );
  OAI21_X1 U16224 ( .B1(n17358), .B2(n19011), .A(n14268), .ZN(n14269) );
  INV_X1 U16225 ( .A(n17067), .ZN(n18869) );
  INV_X1 U16226 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14273) );
  OAI211_X1 U16227 ( .C1(n18869), .C2(n14273), .A(n17732), .B(n14502), .ZN(
        P2_U2814) );
  INV_X1 U16228 ( .A(n14274), .ZN(n14277) );
  INV_X1 U16229 ( .A(n17731), .ZN(n18850) );
  OAI21_X1 U16230 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n14275), .A(n18850), 
        .ZN(n14276) );
  OAI21_X1 U16231 ( .B1(n14277), .B2(n18850), .A(n14276), .ZN(P2_U3612) );
  NAND2_X1 U16232 ( .A1(n16447), .A2(n14278), .ZN(n14280) );
  INV_X1 U16233 ( .A(n21903), .ZN(n14283) );
  OR2_X1 U16234 ( .A1(n22465), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16450) );
  INV_X1 U16235 ( .A(n16450), .ZN(n14281) );
  OAI21_X1 U16236 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n14281), .A(n14283), 
        .ZN(n14282) );
  OAI21_X1 U16237 ( .B1(n14284), .B2(n14283), .A(n14282), .ZN(P1_U3487) );
  INV_X1 U16238 ( .A(n17718), .ZN(n14285) );
  INV_X1 U16239 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20474) );
  INV_X1 U16240 ( .A(n14909), .ZN(n21907) );
  INV_X1 U16241 ( .A(DATAI_15_), .ZN(n15172) );
  NOR2_X1 U16242 ( .A1(n15902), .A2(n15172), .ZN(n14288) );
  AOI21_X1 U16243 ( .B1(n15902), .B2(BUF1_REG_15__SCAN_IN), .A(n14288), .ZN(
        n15818) );
  INV_X1 U16244 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14289) );
  OAI222_X1 U16245 ( .A1(n22387), .A2(n20474), .B1(n22381), .B2(n15818), .C1(
        n22299), .C2(n14289), .ZN(P1_U2967) );
  INV_X1 U16246 ( .A(n11159), .ZN(n14292) );
  AOI21_X1 U16247 ( .B1(n14292), .B2(n14388), .A(n14291), .ZN(n14459) );
  INV_X1 U16248 ( .A(n14459), .ZN(n14298) );
  OR2_X1 U16249 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14293) );
  NAND2_X1 U16250 ( .A1(n14294), .A2(n14293), .ZN(n14600) );
  INV_X1 U16251 ( .A(n14600), .ZN(n15079) );
  INV_X1 U16252 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20526) );
  NOR2_X1 U16253 ( .A1(n22016), .A2(n20526), .ZN(n14458) );
  AOI21_X1 U16254 ( .B1(n14329), .B2(n15845), .A(n14388), .ZN(n14295) );
  AOI211_X1 U16255 ( .C1(n22037), .C2(n15079), .A(n14458), .B(n14295), .ZN(
        n14297) );
  OR2_X1 U16256 ( .A1(n14296), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14330) );
  OAI211_X1 U16257 ( .C1(n14298), .C2(n22033), .A(n14297), .B(n14330), .ZN(
        P1_U3031) );
  NAND3_X1 U16258 ( .A1(n11192), .A2(n14300), .A3(n14299), .ZN(n14301) );
  NOR2_X1 U16259 ( .A1(n14302), .A2(n14301), .ZN(n16826) );
  NOR2_X1 U16260 ( .A1(n14315), .A2(n14909), .ZN(n16465) );
  AND2_X1 U16261 ( .A1(n14303), .A2(n16465), .ZN(n16832) );
  XNOR2_X1 U16262 ( .A(n14304), .B(n17687), .ZN(n14311) );
  INV_X1 U16263 ( .A(n16826), .ZN(n16841) );
  NOR3_X1 U16264 ( .A1(n16841), .A2(n14305), .A3(n14311), .ZN(n14306) );
  AOI21_X1 U16265 ( .B1(n16832), .B2(n14311), .A(n14306), .ZN(n14310) );
  NAND2_X1 U16266 ( .A1(n16834), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14308) );
  NAND2_X1 U16267 ( .A1(n16834), .A2(n14307), .ZN(n16836) );
  MUX2_X1 U16268 ( .A(n14308), .B(n16836), .S(n17687), .Z(n14309) );
  OAI211_X1 U16269 ( .C1(n14822), .C2(n16826), .A(n14310), .B(n14309), .ZN(
        n17686) );
  NOR2_X1 U16270 ( .A1(n17727), .A2(n14388), .ZN(n16819) );
  OAI22_X1 U16271 ( .A1(n14444), .A2(n16263), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16820) );
  INV_X1 U16272 ( .A(n16820), .ZN(n14313) );
  INV_X1 U16273 ( .A(n16845), .ZN(n22215) );
  INV_X1 U16274 ( .A(n14311), .ZN(n14312) );
  AOI222_X1 U16275 ( .A1(n17686), .A2(n17648), .B1(n16819), .B2(n14313), .C1(
        n22215), .C2(n14312), .ZN(n14324) );
  INV_X1 U16276 ( .A(n14314), .ZN(n14321) );
  AOI22_X1 U16277 ( .A1(n16459), .A2(n16454), .B1(n11411), .B2(n14315), .ZN(
        n14320) );
  NOR2_X1 U16278 ( .A1(n22242), .A2(n22254), .ZN(n14316) );
  OAI211_X1 U16279 ( .C1(n16834), .C2(n14317), .A(n16461), .B(n14316), .ZN(
        n14318) );
  NAND4_X1 U16280 ( .A1(n14321), .A2(n14320), .A3(n14319), .A4(n14318), .ZN(
        n17697) );
  INV_X1 U16281 ( .A(n17697), .ZN(n17702) );
  NAND2_X1 U16282 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22209) );
  NOR2_X1 U16283 ( .A1(n22210), .A2(n22209), .ZN(n14477) );
  INV_X1 U16284 ( .A(n14477), .ZN(n14322) );
  INV_X1 U16285 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22204) );
  OAI22_X1 U16286 ( .A1(n17702), .A2(n22220), .B1(n14322), .B2(n22204), .ZN(
        n17647) );
  AOI21_X1 U16287 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22210), .A(n17647), 
        .ZN(n14390) );
  NAND2_X1 U16288 ( .A1(n17687), .A2(n14390), .ZN(n14323) );
  OAI21_X1 U16289 ( .B1(n14324), .B2(n14390), .A(n14323), .ZN(P1_U3472) );
  XNOR2_X1 U16290 ( .A(n16299), .B(n11229), .ZN(n16295) );
  INV_X1 U16291 ( .A(n16295), .ZN(n14337) );
  OR2_X1 U16292 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16292) );
  CLKBUF_X1 U16293 ( .A(n14327), .Z(n14328) );
  NAND3_X1 U16294 ( .A1(n16292), .A2(n14328), .A3(n22038), .ZN(n14336) );
  AOI21_X1 U16295 ( .B1(n14330), .B2(n14329), .A(n14444), .ZN(n14334) );
  INV_X1 U16296 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20527) );
  NOR2_X1 U16297 ( .A1(n22016), .A2(n20527), .ZN(n16289) );
  INV_X1 U16298 ( .A(n22015), .ZN(n14332) );
  AND3_X1 U16299 ( .A1(n14444), .A2(n14332), .A3(n14331), .ZN(n14333) );
  NOR3_X1 U16300 ( .A1(n14334), .A2(n16289), .A3(n14333), .ZN(n14335) );
  OAI211_X1 U16301 ( .C1(n22017), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        P1_U3030) );
  XNOR2_X1 U16302 ( .A(n18864), .B(n14339), .ZN(n14402) );
  NOR2_X1 U16303 ( .A1(n17323), .A2(n18862), .ZN(n14401) );
  AOI21_X1 U16304 ( .B1(n14339), .B2(n14338), .A(n11280), .ZN(n14403) );
  AND2_X1 U16305 ( .A1(n17820), .A2(n14403), .ZN(n14340) );
  AOI211_X1 U16306 ( .C1(n17818), .C2(n14402), .A(n14401), .B(n14340), .ZN(
        n14343) );
  OAI21_X1 U16307 ( .B1(n17814), .B2(n14341), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14342) );
  OAI211_X1 U16308 ( .C1(n13199), .C2(n14399), .A(n14343), .B(n14342), .ZN(
        P2_U3014) );
  INV_X1 U16309 ( .A(n19197), .ZN(n14345) );
  NAND2_X1 U16310 ( .A1(n14345), .A2(n19194), .ZN(n17610) );
  NAND2_X1 U16311 ( .A1(n17610), .A2(n13277), .ZN(n14346) );
  NAND2_X1 U16312 ( .A1(n17125), .A2(n14347), .ZN(n17128) );
  NAND2_X1 U16313 ( .A1(n19096), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14348) );
  NAND4_X1 U16314 ( .A1(n13736), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14348), 
        .A4(n19834), .ZN(n14349) );
  MUX2_X1 U16315 ( .A(n14399), .B(n14351), .S(n11163), .Z(n14352) );
  OAI21_X1 U16316 ( .B1(n17128), .B2(n19775), .A(n14352), .ZN(P2_U2887) );
  INV_X1 U16317 ( .A(n14356), .ZN(n14353) );
  AOI222_X1 U16318 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14356), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14355), .C1(n14354), .C2(
        n14353), .ZN(n17594) );
  OAI21_X1 U16319 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14358), .A(
        n14357), .ZN(n17590) );
  INV_X1 U16320 ( .A(n17590), .ZN(n14359) );
  NOR2_X1 U16321 ( .A1(n17323), .A2(n17918), .ZN(n17592) );
  AOI21_X1 U16322 ( .B1(n17820), .B2(n14359), .A(n17592), .ZN(n14361) );
  NAND2_X1 U16323 ( .A1(n17777), .A2(n17059), .ZN(n14360) );
  OAI211_X1 U16324 ( .C1(n17059), .C2(n17789), .A(n14361), .B(n14360), .ZN(
        n14362) );
  AOI21_X1 U16325 ( .B1(n17595), .B2(n17807), .A(n14362), .ZN(n14363) );
  OAI21_X1 U16326 ( .B1(n17594), .B2(n13196), .A(n14363), .ZN(P2_U3013) );
  XNOR2_X1 U16327 ( .A(n14365), .B(n14364), .ZN(n14420) );
  AOI22_X1 U16328 ( .A1(n17807), .A2(n17054), .B1(n17777), .B2(n17047), .ZN(
        n14372) );
  OAI21_X1 U16329 ( .B1(n14368), .B2(n14367), .A(n14366), .ZN(n14414) );
  INV_X1 U16330 ( .A(n14414), .ZN(n14370) );
  NOR2_X1 U16331 ( .A1(n17323), .A2(n14369), .ZN(n14416) );
  AOI21_X1 U16332 ( .B1(n17820), .B2(n14370), .A(n14416), .ZN(n14371) );
  OAI211_X1 U16333 ( .C1(n14373), .C2(n17789), .A(n14372), .B(n14371), .ZN(
        n14374) );
  INV_X1 U16334 ( .A(n14374), .ZN(n14375) );
  OAI21_X1 U16335 ( .B1(n13196), .B2(n14420), .A(n14375), .ZN(P2_U3012) );
  NOR2_X1 U16336 ( .A1(n11163), .A2(n17621), .ZN(n14380) );
  AOI21_X1 U16337 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n11163), .A(n14380), .ZN(
        n14381) );
  OAI21_X1 U16338 ( .B1(n19814), .B2(n17128), .A(n14381), .ZN(P2_U2886) );
  MUX2_X1 U16339 ( .A(n14411), .B(n13044), .S(n11164), .Z(n14386) );
  OAI21_X1 U16340 ( .B1(n20015), .B2(n17128), .A(n14386), .ZN(P2_U2885) );
  NOR2_X1 U16341 ( .A1(n11422), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14387) );
  AOI21_X1 U16342 ( .B1(n16804), .B2(n16841), .A(n14387), .ZN(n17700) );
  INV_X1 U16343 ( .A(n17648), .ZN(n16846) );
  AOI22_X1 U16344 ( .A1(n14391), .A2(n22215), .B1(n14388), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14389) );
  OAI21_X1 U16345 ( .B1(n17700), .B2(n16846), .A(n14389), .ZN(n14393) );
  INV_X1 U16346 ( .A(n14390), .ZN(n17650) );
  NAND2_X1 U16347 ( .A1(n16834), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17698) );
  OAI22_X1 U16348 ( .A1(n17698), .A2(n16846), .B1(n14391), .B2(n17650), .ZN(
        n14392) );
  AOI21_X1 U16349 ( .B1(n14393), .B2(n17650), .A(n14392), .ZN(n14394) );
  INV_X1 U16350 ( .A(n14394), .ZN(P1_U3474) );
  INV_X1 U16351 ( .A(n17598), .ZN(n17497) );
  INV_X1 U16352 ( .A(n14409), .ZN(n17593) );
  NOR2_X1 U16353 ( .A1(n14395), .A2(n14396), .ZN(n14397) );
  OR2_X1 U16354 ( .A1(n14398), .A2(n14397), .ZN(n20275) );
  OAI22_X1 U16355 ( .A1(n19130), .A2(n14399), .B1(n19134), .B2(n20275), .ZN(
        n14400) );
  AOI211_X1 U16356 ( .C1(n17593), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14401), .B(n14400), .ZN(n14405) );
  AOI22_X1 U16357 ( .A1(n19157), .A2(n14403), .B1(n19160), .B2(n14402), .ZN(
        n14404) );
  OAI211_X1 U16358 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17497), .A(
        n14405), .B(n14404), .ZN(P2_U3046) );
  XNOR2_X1 U16359 ( .A(n14407), .B(n14406), .ZN(n20012) );
  NOR2_X1 U16360 ( .A1(n14409), .A2(n14408), .ZN(n14413) );
  NOR2_X1 U16361 ( .A1(n14878), .A2(n14410), .ZN(n14417) );
  OAI22_X1 U16362 ( .A1(n14417), .A2(n17448), .B1(n19130), .B2(n14411), .ZN(
        n14412) );
  AOI211_X1 U16363 ( .C1(n19154), .C2(n20012), .A(n14413), .B(n14412), .ZN(
        n14419) );
  NOR2_X1 U16364 ( .A1(n19153), .A2(n14414), .ZN(n14415) );
  AOI211_X1 U16365 ( .C1(n14417), .C2(n17451), .A(n14416), .B(n14415), .ZN(
        n14418) );
  OAI211_X1 U16366 ( .C1(n19123), .C2(n14420), .A(n14419), .B(n14418), .ZN(
        P2_U3044) );
  XOR2_X1 U16367 ( .A(n14497), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14425)
         );
  AND2_X1 U16368 ( .A1(n14432), .A2(n14422), .ZN(n14423) );
  OR2_X1 U16369 ( .A1(n14423), .A2(n14494), .ZN(n15676) );
  MUX2_X1 U16370 ( .A(n15676), .B(n13073), .S(n11163), .Z(n14424) );
  OAI21_X1 U16371 ( .B1(n14425), .B2(n17128), .A(n14424), .ZN(P2_U2882) );
  OR2_X1 U16372 ( .A1(n14427), .A2(n14426), .ZN(n14428) );
  NAND2_X1 U16373 ( .A1(n14428), .A2(n14497), .ZN(n20076) );
  NAND2_X1 U16374 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  AND2_X1 U16375 ( .A1(n14432), .A2(n14431), .ZN(n17032) );
  INV_X1 U16376 ( .A(n17032), .ZN(n15073) );
  NOR2_X1 U16377 ( .A1(n15073), .A2(n11163), .ZN(n14433) );
  AOI21_X1 U16378 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n11163), .A(n14433), .ZN(
        n14434) );
  OAI21_X1 U16379 ( .B1(n20076), .B2(n17128), .A(n14434), .ZN(P2_U2883) );
  NAND2_X1 U16380 ( .A1(n14437), .A2(n14436), .ZN(n14438) );
  XOR2_X1 U16381 ( .A(n14439), .B(n14438), .Z(n16311) );
  NAND2_X1 U16382 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  AND2_X1 U16383 ( .A1(n14440), .A2(n14443), .ZN(n16321) );
  NOR2_X1 U16384 ( .A1(n14444), .A2(n15838), .ZN(n21926) );
  INV_X1 U16385 ( .A(n21926), .ZN(n14445) );
  INV_X1 U16386 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20476) );
  OR2_X1 U16387 ( .A1(n22016), .A2(n20476), .ZN(n16306) );
  OAI21_X1 U16388 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14445), .A(
        n16306), .ZN(n14446) );
  NOR2_X1 U16389 ( .A1(n15936), .A2(n21925), .ZN(n21923) );
  AOI211_X1 U16390 ( .C1(n22037), .C2(n16321), .A(n14446), .B(n21923), .ZN(
        n14450) );
  NAND2_X1 U16391 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14447) );
  OAI22_X1 U16392 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21944), .B1(
        n14447), .B2(n15936), .ZN(n14448) );
  OAI21_X1 U16393 ( .B1(n14448), .B2(n21979), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14449) );
  OAI211_X1 U16394 ( .C1(n16311), .C2(n22033), .A(n14450), .B(n14449), .ZN(
        P1_U3029) );
  INV_X1 U16395 ( .A(n14451), .ZN(n14454) );
  OAI21_X1 U16396 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n15085) );
  INV_X1 U16397 ( .A(n20627), .ZN(n15997) );
  INV_X1 U16398 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14455) );
  AOI21_X1 U16399 ( .B1(n15997), .B2(n14456), .A(n14455), .ZN(n14457) );
  AOI211_X1 U16400 ( .C1(n14459), .C2(n20629), .A(n14458), .B(n14457), .ZN(
        n14460) );
  OAI21_X1 U16401 ( .B1(n20599), .B2(n15085), .A(n14460), .ZN(P1_U2999) );
  INV_X1 U16402 ( .A(n19909), .ZN(n20018) );
  INV_X1 U16403 ( .A(n12643), .ZN(n19075) );
  MUX2_X1 U16404 ( .A(n19075), .B(n13048), .S(n11164), .Z(n14464) );
  OAI21_X1 U16405 ( .B1(n20018), .B2(n17128), .A(n14464), .ZN(P2_U2884) );
  XOR2_X1 U16406 ( .A(n14465), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14472)
         );
  NAND2_X1 U16407 ( .A1(n14466), .A2(n14495), .ZN(n14470) );
  CLKBUF_X1 U16408 ( .A(n14467), .Z(n14468) );
  INV_X1 U16409 ( .A(n14468), .ZN(n14469) );
  NAND2_X1 U16410 ( .A1(n14470), .A2(n14469), .ZN(n18891) );
  MUX2_X1 U16411 ( .A(n18891), .B(n13094), .S(n11163), .Z(n14471) );
  OAI21_X1 U16412 ( .B1(n14472), .B2(n17128), .A(n14471), .ZN(P2_U2880) );
  NAND2_X1 U16413 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22476), .ZN(n17722) );
  INV_X1 U16414 ( .A(n14473), .ZN(n14475) );
  AOI21_X1 U16415 ( .B1(n14475), .B2(n14474), .A(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14476) );
  NOR2_X1 U16416 ( .A1(n14476), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n16803) );
  OAI21_X1 U16417 ( .B1(n16803), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14477), .ZN(
        n14478) );
  NAND2_X1 U16418 ( .A1(n14966), .A2(n14478), .ZN(n17728) );
  INV_X1 U16419 ( .A(n14760), .ZN(n14821) );
  NAND2_X1 U16420 ( .A1(n16807), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22418) );
  INV_X1 U16421 ( .A(n22465), .ZN(n22417) );
  OAI21_X1 U16422 ( .B1(n14821), .B2(n22418), .A(n22417), .ZN(n16814) );
  INV_X1 U16423 ( .A(n22418), .ZN(n14681) );
  NOR2_X1 U16424 ( .A1(n14760), .A2(n14681), .ZN(n14480) );
  NAND2_X1 U16425 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22211), .ZN(n16811) );
  INV_X1 U16426 ( .A(n16811), .ZN(n16809) );
  OAI22_X1 U16427 ( .A1(n16814), .A2(n14480), .B1(n14822), .B2(n16809), .ZN(
        n14481) );
  NAND2_X1 U16428 ( .A1(n14481), .A2(n17728), .ZN(n14482) );
  OAI21_X1 U16429 ( .B1(n17707), .B2(n17728), .A(n14482), .ZN(P1_U3476) );
  INV_X1 U16430 ( .A(n14483), .ZN(n14486) );
  INV_X1 U16431 ( .A(n14484), .ZN(n14485) );
  NAND2_X1 U16432 ( .A1(n14486), .A2(n14485), .ZN(n14487) );
  NAND2_X1 U16433 ( .A1(n14488), .A2(n14487), .ZN(n20219) );
  INV_X1 U16434 ( .A(n20219), .ZN(n17589) );
  XNOR2_X1 U16435 ( .A(n19749), .B(n20219), .ZN(n20221) );
  NOR2_X1 U16436 ( .A1(n19775), .A2(n20275), .ZN(n20278) );
  NOR2_X1 U16437 ( .A1(n20221), .A2(n20278), .ZN(n20220) );
  AOI21_X1 U16438 ( .B1(n17589), .B2(n19814), .A(n20220), .ZN(n20013) );
  XNOR2_X1 U16439 ( .A(n20013), .B(n20012), .ZN(n20016) );
  XNOR2_X1 U16440 ( .A(n20016), .B(n20015), .ZN(n14492) );
  AOI22_X1 U16441 ( .A1(n20277), .A2(n20012), .B1(n20276), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U16442 ( .A1(n20067), .A2(n14489), .ZN(n20011) );
  OAI22_X1 U16443 ( .A1(n19738), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19737), .ZN(n20178) );
  INV_X1 U16444 ( .A(n20178), .ZN(n20167) );
  NAND2_X1 U16445 ( .A1(n20011), .A2(n20167), .ZN(n14490) );
  OAI211_X1 U16446 ( .C1(n14492), .C2(n20222), .A(n14491), .B(n14490), .ZN(
        P2_U2917) );
  OR2_X1 U16447 ( .A1(n14494), .A2(n14493), .ZN(n14496) );
  NAND2_X1 U16448 ( .A1(n14496), .A2(n14495), .ZN(n18881) );
  NOR2_X1 U16449 ( .A1(n14497), .A2(n13790), .ZN(n14498) );
  OAI211_X1 U16450 ( .C1(n14498), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17136), .B(n14465), .ZN(n14500) );
  NAND2_X1 U16451 ( .A1(n11163), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14499) );
  OAI211_X1 U16452 ( .C1(n18881), .C2(n11163), .A(n14500), .B(n14499), .ZN(
        P2_U2881) );
  INV_X1 U16453 ( .A(n14502), .ZN(n14501) );
  AOI22_X1 U16454 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n14503) );
  NOR3_X4 U16455 ( .A1(n14502), .A2(n20227), .A3(n22275), .ZN(n14576) );
  AOI22_X1 U16456 ( .A1(n19737), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19738), .ZN(n20226) );
  INV_X1 U16457 ( .A(n20226), .ZN(n17200) );
  NAND2_X1 U16458 ( .A1(n14576), .A2(n17200), .ZN(n14537) );
  NAND2_X1 U16459 ( .A1(n14503), .A2(n14537), .ZN(P2_U2968) );
  AOI22_X1 U16460 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n11245), .B1(n14550), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U16461 ( .A1(n14576), .A2(n20167), .ZN(n14529) );
  NAND2_X1 U16462 ( .A1(n14504), .A2(n14529), .ZN(P2_U2969) );
  AOI22_X1 U16463 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n14506) );
  INV_X1 U16464 ( .A(n19713), .ZN(n14505) );
  NAND2_X1 U16465 ( .A1(n14576), .A2(n14505), .ZN(n14533) );
  NAND2_X1 U16466 ( .A1(n14506), .A2(n14533), .ZN(P2_U2966) );
  AOI22_X1 U16467 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n11245), .B1(n14550), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n14508) );
  OAI22_X1 U16468 ( .A1(n19738), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19737), .ZN(n20080) );
  INV_X1 U16469 ( .A(n20080), .ZN(n14507) );
  NAND2_X1 U16470 ( .A1(n14576), .A2(n14507), .ZN(n14548) );
  NAND2_X1 U16471 ( .A1(n14508), .A2(n14548), .ZN(P2_U2971) );
  AOI22_X1 U16472 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U16473 ( .A1(n19737), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19738), .ZN(n19719) );
  INV_X1 U16474 ( .A(n19719), .ZN(n14509) );
  NAND2_X1 U16475 ( .A1(n14576), .A2(n14509), .ZN(n14520) );
  NAND2_X1 U16476 ( .A1(n14510), .A2(n14520), .ZN(P2_U2964) );
  AOI22_X1 U16477 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n11245), .B1(n14550), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U16478 ( .A1(n19737), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14531), .ZN(n19732) );
  INV_X1 U16479 ( .A(n19732), .ZN(n17162) );
  NAND2_X1 U16480 ( .A1(n14576), .A2(n17162), .ZN(n14551) );
  NAND2_X1 U16481 ( .A1(n14511), .A2(n14551), .ZN(P2_U2975) );
  AOI22_X1 U16482 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n14545), .B1(n14574), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n14512) );
  AOI22_X1 U16483 ( .A1(n19737), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n14531), .ZN(n19728) );
  INV_X1 U16484 ( .A(n19728), .ZN(n17157) );
  NAND2_X1 U16485 ( .A1(n14576), .A2(n17157), .ZN(n14517) );
  NAND2_X1 U16486 ( .A1(n14512), .A2(n14517), .ZN(P2_U2976) );
  AOI22_X1 U16487 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n14513) );
  AOI22_X1 U16488 ( .A1(n19737), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19738), .ZN(n20287) );
  INV_X1 U16489 ( .A(n20287), .ZN(n15735) );
  NAND2_X1 U16490 ( .A1(n14576), .A2(n15735), .ZN(n14546) );
  NAND2_X1 U16491 ( .A1(n14513), .A2(n14546), .ZN(P2_U2967) );
  AOI22_X1 U16492 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U16493 ( .A1(n19737), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19738), .ZN(n19722) );
  INV_X1 U16494 ( .A(n19722), .ZN(n14514) );
  NAND2_X1 U16495 ( .A1(n14576), .A2(n14514), .ZN(n14539) );
  NAND2_X1 U16496 ( .A1(n14515), .A2(n14539), .ZN(P2_U2963) );
  AOI22_X1 U16497 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n11245), .B1(n14550), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n14516) );
  INV_X1 U16498 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20652) );
  INV_X1 U16499 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21231) );
  OAI22_X1 U16500 ( .A1(n19738), .A2(n20652), .B1(n21231), .B2(n19737), .ZN(
        n20024) );
  NAND2_X1 U16501 ( .A1(n14576), .A2(n20024), .ZN(n14535) );
  NAND2_X1 U16502 ( .A1(n14516), .A2(n14535), .ZN(P2_U2972) );
  AOI22_X1 U16503 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n14518) );
  NAND2_X1 U16504 ( .A1(n14518), .A2(n14517), .ZN(P2_U2961) );
  AOI22_X1 U16505 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n11245), .B1(n14550), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U16506 ( .A1(n19737), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19738), .ZN(n20127) );
  INV_X1 U16507 ( .A(n20127), .ZN(n17191) );
  NAND2_X1 U16508 ( .A1(n14576), .A2(n17191), .ZN(n14527) );
  NAND2_X1 U16509 ( .A1(n14519), .A2(n14527), .ZN(P2_U2970) );
  AOI22_X1 U16510 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U16511 ( .A1(n14521), .A2(n14520), .ZN(P2_U2979) );
  AOI22_X1 U16512 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n14522) );
  AOI22_X1 U16513 ( .A1(n19737), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19738), .ZN(n19970) );
  INV_X1 U16514 ( .A(n19970), .ZN(n17174) );
  NAND2_X1 U16515 ( .A1(n14576), .A2(n17174), .ZN(n14541) );
  NAND2_X1 U16516 ( .A1(n14522), .A2(n14541), .ZN(P2_U2973) );
  AOI22_X1 U16517 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U16518 ( .A1(n19737), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19738), .ZN(n19741) );
  INV_X1 U16519 ( .A(n19741), .ZN(n14523) );
  NAND2_X1 U16520 ( .A1(n14576), .A2(n14523), .ZN(n14525) );
  NAND2_X1 U16521 ( .A1(n14524), .A2(n14525), .ZN(P2_U2959) );
  AOI22_X1 U16522 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U16523 ( .A1(n14526), .A2(n14525), .ZN(P2_U2974) );
  AOI22_X1 U16524 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n14528) );
  NAND2_X1 U16525 ( .A1(n14528), .A2(n14527), .ZN(P2_U2955) );
  AOI22_X1 U16526 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U16527 ( .A1(n14530), .A2(n14529), .ZN(P2_U2954) );
  AOI22_X1 U16528 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U16529 ( .A1(n19737), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n14531), .ZN(n19716) );
  INV_X1 U16530 ( .A(n19716), .ZN(n16440) );
  NAND2_X1 U16531 ( .A1(n14576), .A2(n16440), .ZN(n14543) );
  NAND2_X1 U16532 ( .A1(n14532), .A2(n14543), .ZN(P2_U2980) );
  AOI22_X1 U16533 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U16534 ( .A1(n14534), .A2(n14533), .ZN(P2_U2981) );
  AOI22_X1 U16535 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n14536) );
  NAND2_X1 U16536 ( .A1(n14536), .A2(n14535), .ZN(P2_U2957) );
  AOI22_X1 U16537 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U16538 ( .A1(n14538), .A2(n14537), .ZN(P2_U2953) );
  AOI22_X1 U16539 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n14545), .B1(n14574), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U16540 ( .A1(n14540), .A2(n14539), .ZN(P2_U2978) );
  AOI22_X1 U16541 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U16542 ( .A1(n14542), .A2(n14541), .ZN(P2_U2958) );
  AOI22_X1 U16543 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U16544 ( .A1(n14544), .A2(n14543), .ZN(P2_U2965) );
  AOI22_X1 U16545 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n11245), .B1(n14574), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U16546 ( .A1(n14547), .A2(n14546), .ZN(P2_U2952) );
  AOI22_X1 U16547 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U16548 ( .A1(n14549), .A2(n14548), .ZN(P2_U2956) );
  AOI22_X1 U16549 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n14545), .B1(n14550), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U16550 ( .A1(n14552), .A2(n14551), .ZN(P2_U2960) );
  INV_X1 U16551 ( .A(DATAI_29_), .ZN(n16575) );
  INV_X1 U16552 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20701) );
  OR2_X1 U16553 ( .A1(n14665), .A2(n20701), .ZN(n14553) );
  OAI21_X1 U16554 ( .B1(n14668), .B2(n16575), .A(n14553), .ZN(n22620) );
  INV_X1 U16555 ( .A(n22620), .ZN(n14983) );
  NAND2_X1 U16556 ( .A1(n14760), .A2(n14554), .ZN(n14706) );
  INV_X1 U16557 ( .A(n22403), .ZN(n14555) );
  NOR2_X2 U16558 ( .A1(n14706), .A2(n15006), .ZN(n22721) );
  INV_X1 U16559 ( .A(DATAI_21_), .ZN(n16004) );
  INV_X1 U16560 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20684) );
  OR2_X1 U16561 ( .A1(n14665), .A2(n20684), .ZN(n14556) );
  NOR2_X2 U16562 ( .A1(n14670), .A2(n14559), .ZN(n22619) );
  INV_X1 U16563 ( .A(n22619), .ZN(n14703) );
  INV_X1 U16564 ( .A(n14966), .ZN(n14660) );
  NOR2_X1 U16565 ( .A1(n15902), .A2(DATAI_5_), .ZN(n14560) );
  AOI21_X1 U16566 ( .B1(n15902), .B2(n20652), .A(n14560), .ZN(n16006) );
  NAND2_X1 U16567 ( .A1(n14660), .A2(n16006), .ZN(n22623) );
  INV_X1 U16568 ( .A(n14631), .ZN(n17644) );
  OR2_X1 U16569 ( .A1(n14822), .A2(n17644), .ZN(n22469) );
  AND2_X1 U16570 ( .A1(n14561), .A2(n16804), .ZN(n22420) );
  INV_X1 U16571 ( .A(n14615), .ZN(n22718) );
  AOI21_X1 U16572 ( .B1(n14934), .B2(n22420), .A(n22718), .ZN(n14564) );
  NOR2_X1 U16573 ( .A1(n17709), .A2(n22437), .ZN(n14566) );
  INV_X1 U16574 ( .A(n14566), .ZN(n14562) );
  OAI22_X1 U16575 ( .A1(n14564), .A2(n22465), .B1(n14562), .B2(n22476), .ZN(
        n22716) );
  INV_X1 U16576 ( .A(n22716), .ZN(n14614) );
  OAI22_X1 U16577 ( .A1(n14703), .A2(n14615), .B1(n22623), .B2(n14614), .ZN(
        n14563) );
  AOI21_X1 U16578 ( .B1(n22721), .B2(n14557), .A(n14563), .ZN(n14568) );
  OAI211_X1 U16579 ( .C1(n14706), .C2(n22418), .A(n22417), .B(n14564), .ZN(
        n14565) );
  OAI211_X1 U16580 ( .C1(n22417), .C2(n14566), .A(n14565), .B(n14824), .ZN(
        n22722) );
  NAND2_X1 U16581 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14567) );
  OAI211_X1 U16582 ( .C1(n14983), .C2(n22725), .A(n14568), .B(n14567), .ZN(
        P1_U3158) );
  INV_X1 U16583 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17874) );
  NAND2_X1 U16584 ( .A1(n19738), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14570) );
  INV_X1 U16585 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20662) );
  OR2_X1 U16586 ( .A1(n19738), .A2(n20662), .ZN(n14569) );
  NAND2_X1 U16587 ( .A1(n14570), .A2(n14569), .ZN(n19725) );
  NAND2_X1 U16588 ( .A1(n14576), .A2(n19725), .ZN(n14573) );
  NAND2_X1 U16589 ( .A1(n14545), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14571) );
  OAI211_X1 U16590 ( .C1(n17874), .C2(n17664), .A(n14573), .B(n14571), .ZN(
        P2_U2977) );
  INV_X1 U16591 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n17905) );
  NAND2_X1 U16592 ( .A1(n14545), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14572) );
  OAI211_X1 U16593 ( .C1(n17905), .C2(n17664), .A(n14573), .B(n14572), .ZN(
        P2_U2962) );
  AOI22_X1 U16594 ( .A1(n19737), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19738), .ZN(n19710) );
  INV_X1 U16595 ( .A(n19710), .ZN(n14575) );
  AOI222_X1 U16596 ( .A1(n14545), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n14576), 
        .B2(n14575), .C1(P2_EAX_REG_15__SCAN_IN), .C2(n14574), .ZN(n14577) );
  INV_X1 U16597 ( .A(n14577), .ZN(P2_U2982) );
  INV_X1 U16598 ( .A(DATAI_27_), .ZN(n16583) );
  INV_X1 U16599 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20697) );
  OR2_X1 U16600 ( .A1(n14665), .A2(n20697), .ZN(n14578) );
  OAI21_X1 U16601 ( .B1(n14668), .B2(n16583), .A(n14578), .ZN(n22576) );
  INV_X1 U16602 ( .A(n22576), .ZN(n14803) );
  INV_X1 U16603 ( .A(DATAI_19_), .ZN(n14579) );
  INV_X1 U16604 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20680) );
  NOR2_X2 U16605 ( .A1(n14670), .A2(n14580), .ZN(n22575) );
  INV_X1 U16606 ( .A(n22575), .ZN(n22564) );
  NAND2_X1 U16607 ( .A1(n14671), .A2(DATAI_3_), .ZN(n14582) );
  NAND2_X1 U16608 ( .A1(n15902), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14581) );
  AND2_X1 U16609 ( .A1(n14582), .A2(n14581), .ZN(n22314) );
  NOR2_X1 U16610 ( .A1(n14966), .A2(n22314), .ZN(n22573) );
  INV_X1 U16611 ( .A(n22573), .ZN(n22571) );
  OAI22_X1 U16612 ( .A1(n22564), .A2(n14615), .B1(n14614), .B2(n22571), .ZN(
        n14583) );
  AOI21_X1 U16613 ( .B1(n22568), .B2(n22721), .A(n14583), .ZN(n14585) );
  NAND2_X1 U16614 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14584) );
  OAI211_X1 U16615 ( .C1(n14803), .C2(n22725), .A(n14585), .B(n14584), .ZN(
        P1_U3156) );
  INV_X1 U16616 ( .A(DATAI_25_), .ZN(n16594) );
  INV_X1 U16617 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20692) );
  OR2_X1 U16618 ( .A1(n14665), .A2(n20692), .ZN(n14586) );
  OAI21_X1 U16619 ( .B1(n14668), .B2(n16594), .A(n14586), .ZN(n22516) );
  INV_X1 U16620 ( .A(n22516), .ZN(n14808) );
  INV_X1 U16621 ( .A(DATAI_17_), .ZN(n15744) );
  INV_X1 U16622 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20676) );
  OAI22_X1 U16623 ( .A1(n15744), .A2(n14668), .B1(n20676), .B2(n14665), .ZN(
        n22510) );
  NOR2_X2 U16624 ( .A1(n14670), .A2(n14587), .ZN(n22515) );
  INV_X1 U16625 ( .A(n22515), .ZN(n22506) );
  NAND2_X1 U16626 ( .A1(n14671), .A2(DATAI_1_), .ZN(n14589) );
  NAND2_X1 U16627 ( .A1(n15902), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14588) );
  AND2_X1 U16628 ( .A1(n14589), .A2(n14588), .ZN(n22305) );
  NOR2_X1 U16629 ( .A1(n14966), .A2(n22305), .ZN(n22514) );
  INV_X1 U16630 ( .A(n22514), .ZN(n22513) );
  OAI22_X1 U16631 ( .A1(n22506), .A2(n14615), .B1(n14614), .B2(n22513), .ZN(
        n14590) );
  AOI21_X1 U16632 ( .B1(n11247), .B2(n22721), .A(n14590), .ZN(n14592) );
  NAND2_X1 U16633 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14591) );
  OAI211_X1 U16634 ( .C1(n14808), .C2(n22725), .A(n14592), .B(n14591), .ZN(
        P1_U3154) );
  INV_X1 U16635 ( .A(DATAI_26_), .ZN(n16589) );
  INV_X1 U16636 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20695) );
  OR2_X1 U16637 ( .A1(n14665), .A2(n20695), .ZN(n14593) );
  OAI21_X1 U16638 ( .B1(n14668), .B2(n16589), .A(n14593), .ZN(n22541) );
  INV_X1 U16639 ( .A(n22541), .ZN(n14813) );
  INV_X1 U16640 ( .A(DATAI_18_), .ZN(n14594) );
  INV_X1 U16641 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20678) );
  OAI22_X1 U16642 ( .A1(n14594), .A2(n14668), .B1(n20678), .B2(n14665), .ZN(
        n22535) );
  NOR2_X2 U16643 ( .A1(n14670), .A2(n11411), .ZN(n22540) );
  INV_X1 U16644 ( .A(n22540), .ZN(n22531) );
  NAND2_X1 U16645 ( .A1(n14671), .A2(DATAI_2_), .ZN(n14596) );
  NAND2_X1 U16646 ( .A1(n15902), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14595) );
  AND2_X1 U16647 ( .A1(n14596), .A2(n14595), .ZN(n22309) );
  NOR2_X1 U16648 ( .A1(n14966), .A2(n22309), .ZN(n22539) );
  INV_X1 U16649 ( .A(n22539), .ZN(n22538) );
  OAI22_X1 U16650 ( .A1(n22531), .A2(n14615), .B1(n14614), .B2(n22538), .ZN(
        n14597) );
  AOI21_X1 U16651 ( .B1(n11249), .B2(n22721), .A(n14597), .ZN(n14599) );
  NAND2_X1 U16652 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14598) );
  OAI211_X1 U16653 ( .C1(n14813), .C2(n22725), .A(n14599), .B(n14598), .ZN(
        P1_U3155) );
  INV_X1 U16654 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n15318) );
  OAI222_X1 U16655 ( .A1(n14600), .A2(n20551), .B1(n15318), .B2(n20556), .C1(
        n16572), .C2(n15085), .ZN(P1_U2872) );
  OR2_X1 U16656 ( .A1(n14601), .A2(n14468), .ZN(n14602) );
  AND2_X1 U16657 ( .A1(n14602), .A2(n14750), .ZN(n19158) );
  INV_X1 U16658 ( .A(n19158), .ZN(n14608) );
  CLKBUF_X1 U16659 ( .A(n14603), .Z(n14747) );
  OAI211_X1 U16660 ( .C1(n14605), .C2(n14604), .A(n14747), .B(n17136), .ZN(
        n14607) );
  NAND2_X1 U16661 ( .A1(n11164), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14606) );
  OAI211_X1 U16662 ( .C1(n14608), .C2(n11164), .A(n14607), .B(n14606), .ZN(
        P2_U2879) );
  INV_X1 U16663 ( .A(DATAI_24_), .ZN(n16599) );
  INV_X1 U16664 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20690) );
  OR2_X1 U16665 ( .A1(n14665), .A2(n20690), .ZN(n14609) );
  INV_X1 U16666 ( .A(n22490), .ZN(n14771) );
  INV_X1 U16667 ( .A(DATAI_16_), .ZN(n14610) );
  INV_X1 U16668 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20674) );
  OAI22_X1 U16669 ( .A1(n14610), .A2(n14668), .B1(n20674), .B2(n14665), .ZN(
        n22475) );
  NOR2_X2 U16670 ( .A1(n14670), .A2(n14611), .ZN(n22489) );
  INV_X1 U16671 ( .A(n22489), .ZN(n22455) );
  NAND2_X1 U16672 ( .A1(n14671), .A2(DATAI_0_), .ZN(n14613) );
  NAND2_X1 U16673 ( .A1(n15902), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14612) );
  AND2_X1 U16674 ( .A1(n14613), .A2(n14612), .ZN(n22300) );
  NOR2_X1 U16675 ( .A1(n14966), .A2(n22300), .ZN(n22488) );
  OAI22_X1 U16676 ( .A1(n22455), .A2(n14615), .B1(n14614), .B2(n22487), .ZN(
        n14616) );
  AOI21_X1 U16677 ( .B1(n22475), .B2(n22721), .A(n14616), .ZN(n14618) );
  NAND2_X1 U16678 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14617) );
  OAI211_X1 U16679 ( .C1(n14771), .C2(n22725), .A(n14618), .B(n14617), .ZN(
        P1_U3153) );
  OAI21_X1 U16680 ( .B1(n14619), .B2(n14620), .A(n14627), .ZN(n16305) );
  NAND2_X1 U16681 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  NAND2_X2 U16682 ( .A1(n16612), .A2(n14623), .ZN(n16621) );
  OAI222_X1 U16683 ( .A1(n16305), .A2(n16621), .B1(n15819), .B2(n22305), .C1(
        n15817), .C2(n12070), .ZN(P1_U2903) );
  INV_X1 U16684 ( .A(n14624), .ZN(n14628) );
  INV_X1 U16685 ( .A(n14625), .ZN(n14626) );
  AOI21_X1 U16686 ( .B1(n14628), .B2(n14627), .A(n14626), .ZN(n16312) );
  INV_X1 U16687 ( .A(n16312), .ZN(n16330) );
  OAI222_X1 U16688 ( .A1(n16330), .A2(n16621), .B1(n15819), .B2(n22309), .C1(
        n15817), .C2(n12060), .ZN(P1_U2902) );
  INV_X1 U16689 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n22304) );
  OAI222_X1 U16690 ( .A1(n15085), .A2(n16621), .B1(n15819), .B2(n22300), .C1(
        n15817), .C2(n22304), .ZN(P1_U2904) );
  NAND2_X1 U16691 ( .A1(n14683), .A2(n14827), .ZN(n22431) );
  NOR3_X1 U16692 ( .A1(n17707), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14637) );
  INV_X1 U16693 ( .A(n14637), .ZN(n15009) );
  OR2_X1 U16694 ( .A1(n22454), .A2(n15009), .ZN(n14675) );
  OR2_X1 U16695 ( .A1(n14822), .A2(n14631), .ZN(n22433) );
  OAI21_X1 U16696 ( .B1(n22433), .B2(n14701), .A(n14675), .ZN(n14633) );
  AOI22_X1 U16697 ( .A1(n14633), .A2(n22417), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14637), .ZN(n14674) );
  OAI22_X1 U16698 ( .A1(n22455), .A2(n14675), .B1(n14674), .B2(n22487), .ZN(
        n14632) );
  AOI21_X1 U16699 ( .B1(n22475), .B2(n22673), .A(n14632), .ZN(n14639) );
  NAND2_X1 U16700 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n14683), .ZN(n14635) );
  INV_X1 U16701 ( .A(n14633), .ZN(n14634) );
  NAND3_X1 U16702 ( .A1(n14635), .A2(n22417), .A3(n14634), .ZN(n14636) );
  OAI211_X1 U16703 ( .C1(n22417), .C2(n14637), .A(n14636), .B(n14824), .ZN(
        n14678) );
  NAND2_X1 U16704 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14638) );
  OAI211_X1 U16705 ( .C1(n14771), .C2(n15049), .A(n14639), .B(n14638), .ZN(
        P1_U3073) );
  OAI22_X1 U16706 ( .A1(n22564), .A2(n14675), .B1(n14674), .B2(n22571), .ZN(
        n14640) );
  AOI21_X1 U16707 ( .B1(n22568), .B2(n22673), .A(n14640), .ZN(n14642) );
  NAND2_X1 U16708 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14641) );
  OAI211_X1 U16709 ( .C1(n14803), .C2(n15049), .A(n14642), .B(n14641), .ZN(
        P1_U3076) );
  INV_X1 U16710 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20705) );
  OAI22_X1 U16711 ( .A1(n15149), .A2(n14668), .B1(n20705), .B2(n14665), .ZN(
        n22702) );
  INV_X1 U16712 ( .A(n22702), .ZN(n22726) );
  INV_X1 U16713 ( .A(n14668), .ZN(n14643) );
  NAND2_X1 U16714 ( .A1(n14643), .A2(DATAI_23_), .ZN(n14645) );
  INV_X1 U16715 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20688) );
  OR2_X1 U16716 ( .A1(n14665), .A2(n20688), .ZN(n14644) );
  AND2_X1 U16717 ( .A1(n14645), .A2(n14644), .ZN(n22687) );
  INV_X1 U16718 ( .A(n22687), .ZN(n22720) );
  NOR2_X2 U16719 ( .A1(n14670), .A2(n15727), .ZN(n22719) );
  INV_X1 U16720 ( .A(n22719), .ZN(n22685) );
  MUX2_X1 U16721 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n15902), .Z(
        n16609) );
  NAND2_X1 U16722 ( .A1(n14660), .A2(n16609), .ZN(n22707) );
  OAI22_X1 U16723 ( .A1(n22685), .A2(n14675), .B1(n22707), .B2(n14674), .ZN(
        n14646) );
  AOI21_X1 U16724 ( .B1(n22673), .B2(n22720), .A(n14646), .ZN(n14648) );
  NAND2_X1 U16725 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14647) );
  OAI211_X1 U16726 ( .C1(n15049), .C2(n22726), .A(n14648), .B(n14647), .ZN(
        P1_U3080) );
  OAI22_X1 U16727 ( .A1(n22506), .A2(n14675), .B1(n14674), .B2(n22513), .ZN(
        n14649) );
  AOI21_X1 U16728 ( .B1(n11247), .B2(n22673), .A(n14649), .ZN(n14651) );
  NAND2_X1 U16729 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14650) );
  OAI211_X1 U16730 ( .C1(n14808), .C2(n15049), .A(n14651), .B(n14650), .ZN(
        P1_U3074) );
  OAI22_X1 U16731 ( .A1(n22531), .A2(n14675), .B1(n14674), .B2(n22538), .ZN(
        n14652) );
  AOI21_X1 U16732 ( .B1(n11249), .B2(n22673), .A(n14652), .ZN(n14654) );
  NAND2_X1 U16733 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14653) );
  OAI211_X1 U16734 ( .C1(n14813), .C2(n15049), .A(n14654), .B(n14653), .ZN(
        P1_U3075) );
  OAI22_X1 U16735 ( .A1(n14703), .A2(n14675), .B1(n22623), .B2(n14674), .ZN(
        n14655) );
  AOI21_X1 U16736 ( .B1(n22673), .B2(n14557), .A(n14655), .ZN(n14657) );
  NAND2_X1 U16737 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14656) );
  OAI211_X1 U16738 ( .C1(n14983), .C2(n15049), .A(n14657), .B(n14656), .ZN(
        P1_U3078) );
  INV_X1 U16739 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20703) );
  INV_X1 U16740 ( .A(DATAI_30_), .ZN(n14658) );
  OAI22_X1 U16741 ( .A1(n20703), .A2(n14665), .B1(n14658), .B2(n14668), .ZN(
        n22641) );
  INV_X1 U16742 ( .A(n22641), .ZN(n22652) );
  INV_X1 U16743 ( .A(DATAI_22_), .ZN(n16613) );
  INV_X1 U16744 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20686) );
  OR2_X1 U16745 ( .A1(n14665), .A2(n20686), .ZN(n14659) );
  OAI21_X2 U16746 ( .B1(n14668), .B2(n16613), .A(n14659), .ZN(n22649) );
  NOR2_X2 U16747 ( .A1(n14670), .A2(n12076), .ZN(n22648) );
  INV_X1 U16748 ( .A(n22648), .ZN(n22634) );
  MUX2_X1 U16749 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n15902), .Z(
        n16617) );
  NAND2_X1 U16750 ( .A1(n14660), .A2(n16617), .ZN(n22644) );
  OAI22_X1 U16751 ( .A1(n22634), .A2(n14675), .B1(n22644), .B2(n14674), .ZN(
        n14661) );
  AOI21_X1 U16752 ( .B1(n22673), .B2(n22649), .A(n14661), .ZN(n14663) );
  NAND2_X1 U16753 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14662) );
  OAI211_X1 U16754 ( .C1(n15049), .C2(n22652), .A(n14663), .B(n14662), .ZN(
        P1_U3079) );
  INV_X1 U16755 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20699) );
  INV_X1 U16756 ( .A(DATAI_28_), .ZN(n14664) );
  OAI22_X1 U16757 ( .A1(n20699), .A2(n14665), .B1(n14664), .B2(n14668), .ZN(
        n22595) );
  INV_X1 U16758 ( .A(n22595), .ZN(n22606) );
  INV_X1 U16759 ( .A(DATAI_20_), .ZN(n14667) );
  INV_X1 U16760 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20682) );
  OR2_X1 U16761 ( .A1(n14665), .A2(n20682), .ZN(n14666) );
  NOR2_X2 U16762 ( .A1(n14670), .A2(n11408), .ZN(n22603) );
  INV_X1 U16763 ( .A(n22603), .ZN(n14676) );
  NAND2_X1 U16764 ( .A1(n14671), .A2(DATAI_4_), .ZN(n14673) );
  NAND2_X1 U16765 ( .A1(n15902), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14672) );
  AND2_X1 U16766 ( .A1(n14673), .A2(n14672), .ZN(n22319) );
  INV_X1 U16767 ( .A(n22602), .ZN(n22598) );
  OAI22_X1 U16768 ( .A1(n14676), .A2(n14675), .B1(n14674), .B2(n22598), .ZN(
        n14677) );
  AOI21_X1 U16769 ( .B1(n22673), .B2(n14669), .A(n14677), .ZN(n14680) );
  NAND2_X1 U16770 ( .A1(n14678), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14679) );
  OAI211_X1 U16771 ( .C1(n15049), .C2(n22606), .A(n14680), .B(n14679), .ZN(
        P1_U3077) );
  NAND3_X1 U16772 ( .A1(n14683), .A2(n22417), .A3(n14681), .ZN(n16813) );
  OR2_X1 U16773 ( .A1(n22437), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14686) );
  INV_X1 U16774 ( .A(n14824), .ZN(n22424) );
  INV_X1 U16775 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14691) );
  INV_X1 U16776 ( .A(n15006), .ZN(n14682) );
  INV_X1 U16777 ( .A(n22674), .ZN(n14697) );
  NOR2_X1 U16778 ( .A1(n14684), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14741) );
  INV_X1 U16779 ( .A(n22433), .ZN(n14685) );
  AOI21_X1 U16780 ( .B1(n14685), .B2(n22420), .A(n14741), .ZN(n14687) );
  OAI22_X1 U16781 ( .A1(n14687), .A2(n22465), .B1(n14686), .B2(n22476), .ZN(
        n14740) );
  AOI22_X1 U16782 ( .A1(n22575), .A2(n14741), .B1(n22573), .B2(n14740), .ZN(
        n14688) );
  OAI21_X1 U16783 ( .B1(n14697), .B2(n14803), .A(n14688), .ZN(n14689) );
  AOI21_X1 U16784 ( .B1(n22568), .B2(n22560), .A(n14689), .ZN(n14690) );
  OAI21_X1 U16785 ( .B1(n14746), .B2(n14691), .A(n14690), .ZN(P1_U3092) );
  INV_X1 U16786 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U16787 ( .A1(n22540), .A2(n14741), .B1(n22539), .B2(n14740), .ZN(
        n14692) );
  OAI21_X1 U16788 ( .B1(n14697), .B2(n14813), .A(n14692), .ZN(n14693) );
  AOI21_X1 U16789 ( .B1(n11249), .B2(n22560), .A(n14693), .ZN(n14694) );
  OAI21_X1 U16790 ( .B1(n14746), .B2(n14695), .A(n14694), .ZN(P1_U3091) );
  INV_X1 U16791 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14700) );
  AOI22_X1 U16792 ( .A1(n22515), .A2(n14741), .B1(n22514), .B2(n14740), .ZN(
        n14696) );
  OAI21_X1 U16793 ( .B1(n14697), .B2(n14808), .A(n14696), .ZN(n14698) );
  AOI21_X1 U16794 ( .B1(n11247), .B2(n22560), .A(n14698), .ZN(n14699) );
  OAI21_X1 U16795 ( .B1(n14746), .B2(n14700), .A(n14699), .ZN(P1_U3090) );
  NOR3_X1 U16796 ( .A1(n17707), .A2(n17709), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14708) );
  INV_X1 U16797 ( .A(n14708), .ZN(n22474) );
  NOR2_X1 U16798 ( .A1(n22454), .A2(n22474), .ZN(n22709) );
  INV_X1 U16799 ( .A(n22709), .ZN(n14720) );
  INV_X1 U16800 ( .A(n14701), .ZN(n14823) );
  AOI21_X1 U16801 ( .B1(n14934), .B2(n14823), .A(n22709), .ZN(n14705) );
  INV_X1 U16802 ( .A(n14705), .ZN(n14702) );
  AOI22_X1 U16803 ( .A1(n14702), .A2(n22417), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14708), .ZN(n22599) );
  OAI22_X1 U16804 ( .A1(n14703), .A2(n14720), .B1(n22623), .B2(n22599), .ZN(
        n14704) );
  AOI21_X1 U16805 ( .B1(n22711), .B2(n14557), .A(n14704), .ZN(n14710) );
  OAI211_X1 U16806 ( .C1(n14706), .C2(n22223), .A(n22417), .B(n14705), .ZN(
        n14707) );
  OAI211_X1 U16807 ( .C1(n22417), .C2(n14708), .A(n14707), .B(n14824), .ZN(
        n22712) );
  NAND2_X1 U16808 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14709) );
  OAI211_X1 U16809 ( .C1(n14983), .C2(n22715), .A(n14710), .B(n14709), .ZN(
        P1_U3142) );
  OAI22_X1 U16810 ( .A1(n22564), .A2(n14720), .B1(n22599), .B2(n22571), .ZN(
        n14711) );
  AOI21_X1 U16811 ( .B1(n22711), .B2(n22568), .A(n14711), .ZN(n14713) );
  NAND2_X1 U16812 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14712) );
  OAI211_X1 U16813 ( .C1(n14803), .C2(n22715), .A(n14713), .B(n14712), .ZN(
        P1_U3140) );
  OAI22_X1 U16814 ( .A1(n22506), .A2(n14720), .B1(n22599), .B2(n22513), .ZN(
        n14714) );
  AOI21_X1 U16815 ( .B1(n22711), .B2(n11247), .A(n14714), .ZN(n14716) );
  NAND2_X1 U16816 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14715) );
  OAI211_X1 U16817 ( .C1(n14808), .C2(n22715), .A(n14716), .B(n14715), .ZN(
        P1_U3138) );
  OAI22_X1 U16818 ( .A1(n22531), .A2(n14720), .B1(n22599), .B2(n22538), .ZN(
        n14717) );
  AOI21_X1 U16819 ( .B1(n22711), .B2(n11249), .A(n14717), .ZN(n14719) );
  NAND2_X1 U16820 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14718) );
  OAI211_X1 U16821 ( .C1(n14813), .C2(n22715), .A(n14719), .B(n14718), .ZN(
        P1_U3139) );
  OAI22_X1 U16822 ( .A1(n22455), .A2(n14720), .B1(n22599), .B2(n22487), .ZN(
        n14721) );
  AOI21_X1 U16823 ( .B1(n22711), .B2(n22475), .A(n14721), .ZN(n14723) );
  NAND2_X1 U16824 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14722) );
  OAI211_X1 U16825 ( .C1(n14771), .C2(n22715), .A(n14723), .B(n14722), .ZN(
        P1_U3137) );
  INV_X1 U16826 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14727) );
  INV_X1 U16827 ( .A(n14669), .ZN(n15036) );
  AOI22_X1 U16828 ( .A1(n22603), .A2(n14741), .B1(n22602), .B2(n14740), .ZN(
        n14724) );
  OAI21_X1 U16829 ( .B1(n14984), .B2(n15036), .A(n14724), .ZN(n14725) );
  AOI21_X1 U16830 ( .B1(n22595), .B2(n22674), .A(n14725), .ZN(n14726) );
  OAI21_X1 U16831 ( .B1(n14746), .B2(n14727), .A(n14726), .ZN(P1_U3093) );
  INV_X1 U16832 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14731) );
  INV_X1 U16833 ( .A(n22649), .ZN(n22635) );
  AOI22_X1 U16834 ( .A1(n22648), .A2(n14741), .B1(n22647), .B2(n14740), .ZN(
        n14728) );
  OAI21_X1 U16835 ( .B1(n14984), .B2(n22635), .A(n14728), .ZN(n14729) );
  AOI21_X1 U16836 ( .B1(n22641), .B2(n22674), .A(n14729), .ZN(n14730) );
  OAI21_X1 U16837 ( .B1(n14746), .B2(n14731), .A(n14730), .ZN(P1_U3095) );
  INV_X1 U16838 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U16839 ( .A1(n22719), .A2(n14741), .B1(n22717), .B2(n14740), .ZN(
        n14732) );
  OAI21_X1 U16840 ( .B1(n14984), .B2(n22687), .A(n14732), .ZN(n14733) );
  AOI21_X1 U16841 ( .B1(n22702), .B2(n22674), .A(n14733), .ZN(n14734) );
  OAI21_X1 U16842 ( .B1(n14746), .B2(n14735), .A(n14734), .ZN(P1_U3096) );
  INV_X1 U16843 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14739) );
  INV_X1 U16844 ( .A(n14557), .ZN(n15042) );
  INV_X1 U16845 ( .A(n22623), .ZN(n15040) );
  AOI22_X1 U16846 ( .A1(n22619), .A2(n14741), .B1(n15040), .B2(n14740), .ZN(
        n14736) );
  OAI21_X1 U16847 ( .B1(n14984), .B2(n15042), .A(n14736), .ZN(n14737) );
  AOI21_X1 U16848 ( .B1(n22674), .B2(n22620), .A(n14737), .ZN(n14738) );
  OAI21_X1 U16849 ( .B1(n14746), .B2(n14739), .A(n14738), .ZN(P1_U3094) );
  INV_X1 U16850 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14745) );
  INV_X1 U16851 ( .A(n22475), .ZN(n22493) );
  AOI22_X1 U16852 ( .A1(n22489), .A2(n14741), .B1(n22488), .B2(n14740), .ZN(
        n14742) );
  OAI21_X1 U16853 ( .B1(n14984), .B2(n22493), .A(n14742), .ZN(n14743) );
  AOI21_X1 U16854 ( .B1(n22674), .B2(n22490), .A(n14743), .ZN(n14744) );
  OAI21_X1 U16855 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(P1_U3089) );
  OAI211_X1 U16856 ( .C1(n13765), .C2(n14748), .A(n17136), .B(n14858), .ZN(
        n14753) );
  INV_X1 U16857 ( .A(n14856), .ZN(n14749) );
  AOI21_X1 U16858 ( .B1(n14751), .B2(n14750), .A(n14749), .ZN(n17569) );
  NAND2_X1 U16859 ( .A1(n17125), .A2(n17569), .ZN(n14752) );
  OAI211_X1 U16860 ( .C1(n17125), .C2(n13105), .A(n14753), .B(n14752), .ZN(
        P2_U2878) );
  CLKBUF_X1 U16861 ( .A(n14754), .Z(n14755) );
  AND2_X1 U16862 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  OR2_X1 U16863 ( .A1(n14755), .A2(n14758), .ZN(n20561) );
  INV_X1 U16864 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n22324) );
  OAI222_X1 U16865 ( .A1(n20561), .A2(n16621), .B1(n15819), .B2(n22319), .C1(
        n22324), .C2(n16612), .ZN(P1_U2900) );
  NOR3_X1 U16866 ( .A1(n17709), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14762) );
  AND2_X1 U16867 ( .A1(n16842), .A2(n14822), .ZN(n22448) );
  INV_X1 U16868 ( .A(n14762), .ZN(n14964) );
  NOR2_X1 U16869 ( .A1(n22454), .A2(n14964), .ZN(n22680) );
  AOI21_X1 U16870 ( .B1(n22448), .B2(n14823), .A(n22680), .ZN(n14765) );
  OAI211_X1 U16871 ( .C1(n14789), .C2(n22223), .A(n22417), .B(n14765), .ZN(
        n14761) );
  OAI211_X1 U16872 ( .C1(n22417), .C2(n14762), .A(n14761), .B(n14824), .ZN(
        n22681) );
  INV_X1 U16873 ( .A(n22681), .ZN(n14787) );
  INV_X1 U16874 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14769) );
  OAI22_X1 U16875 ( .A1(n14765), .A2(n22465), .B1(n14964), .B2(n22476), .ZN(
        n22679) );
  AOI22_X1 U16876 ( .A1(n22619), .A2(n22680), .B1(n15040), .B2(n22679), .ZN(
        n14766) );
  OAI21_X1 U16877 ( .B1(n22684), .B2(n14983), .A(n14766), .ZN(n14767) );
  AOI21_X1 U16878 ( .B1(n22689), .B2(n14557), .A(n14767), .ZN(n14768) );
  OAI21_X1 U16879 ( .B1(n14787), .B2(n14769), .A(n14768), .ZN(P1_U3110) );
  INV_X1 U16880 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U16881 ( .A1(n22489), .A2(n22680), .B1(n22488), .B2(n22679), .ZN(
        n14770) );
  OAI21_X1 U16882 ( .B1(n22684), .B2(n14771), .A(n14770), .ZN(n14772) );
  AOI21_X1 U16883 ( .B1(n22475), .B2(n22689), .A(n14772), .ZN(n14773) );
  OAI21_X1 U16884 ( .B1(n14787), .B2(n14774), .A(n14773), .ZN(P1_U3105) );
  INV_X1 U16885 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U16886 ( .A1(n22575), .A2(n22680), .B1(n22573), .B2(n22679), .ZN(
        n14775) );
  OAI21_X1 U16887 ( .B1(n22684), .B2(n14803), .A(n14775), .ZN(n14776) );
  AOI21_X1 U16888 ( .B1(n22568), .B2(n22689), .A(n14776), .ZN(n14777) );
  OAI21_X1 U16889 ( .B1(n14787), .B2(n14778), .A(n14777), .ZN(P1_U3108) );
  INV_X1 U16890 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14782) );
  AOI22_X1 U16891 ( .A1(n22515), .A2(n22680), .B1(n22514), .B2(n22679), .ZN(
        n14779) );
  OAI21_X1 U16892 ( .B1(n22684), .B2(n14808), .A(n14779), .ZN(n14780) );
  AOI21_X1 U16893 ( .B1(n11247), .B2(n22689), .A(n14780), .ZN(n14781) );
  OAI21_X1 U16894 ( .B1(n14787), .B2(n14782), .A(n14781), .ZN(P1_U3106) );
  INV_X1 U16895 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16896 ( .A1(n22540), .A2(n22680), .B1(n22539), .B2(n22679), .ZN(
        n14783) );
  OAI21_X1 U16897 ( .B1(n22684), .B2(n14813), .A(n14783), .ZN(n14784) );
  AOI21_X1 U16898 ( .B1(n11249), .B2(n22689), .A(n14784), .ZN(n14785) );
  OAI21_X1 U16899 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(P1_U3107) );
  NOR3_X1 U16900 ( .A1(n17709), .A2(n22408), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22453) );
  INV_X1 U16901 ( .A(n22453), .ZN(n14791) );
  NOR2_X1 U16902 ( .A1(n22454), .A2(n14791), .ZN(n22695) );
  AOI21_X1 U16903 ( .B1(n22448), .B2(n22420), .A(n22695), .ZN(n14792) );
  OAI211_X1 U16904 ( .C1(n14789), .C2(n22418), .A(n22417), .B(n14792), .ZN(
        n14788) );
  OAI211_X1 U16905 ( .C1(n22417), .C2(n22453), .A(n14788), .B(n14824), .ZN(
        n22696) );
  INV_X1 U16906 ( .A(n22696), .ZN(n14853) );
  INV_X1 U16907 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14796) );
  OAI22_X1 U16908 ( .A1(n14792), .A2(n22465), .B1(n14791), .B2(n22476), .ZN(
        n22694) );
  AOI22_X1 U16909 ( .A1(n22619), .A2(n22695), .B1(n15040), .B2(n22694), .ZN(
        n14793) );
  OAI21_X1 U16910 ( .B1(n22699), .B2(n14983), .A(n14793), .ZN(n14794) );
  AOI21_X1 U16911 ( .B1(n22703), .B2(n14557), .A(n14794), .ZN(n14795) );
  OAI21_X1 U16912 ( .B1(n14853), .B2(n14796), .A(n14795), .ZN(P1_U3126) );
  XOR2_X1 U16913 ( .A(n14798), .B(n14797), .Z(n15004) );
  INV_X1 U16914 ( .A(n15004), .ZN(n14919) );
  INV_X1 U16915 ( .A(n14799), .ZN(n14800) );
  XNOR2_X1 U16916 ( .A(n14440), .B(n14800), .ZN(n21937) );
  INV_X1 U16917 ( .A(n20556), .ZN(n16562) );
  AOI22_X1 U16918 ( .A1(n21937), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14801) );
  OAI21_X1 U16919 ( .B1(n14919), .B2(n16572), .A(n14801), .ZN(P1_U2869) );
  INV_X1 U16920 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U16921 ( .A1(n22575), .A2(n22695), .B1(n22573), .B2(n22694), .ZN(
        n14802) );
  OAI21_X1 U16922 ( .B1(n22699), .B2(n14803), .A(n14802), .ZN(n14804) );
  AOI21_X1 U16923 ( .B1(n22568), .B2(n22703), .A(n14804), .ZN(n14805) );
  OAI21_X1 U16924 ( .B1(n14853), .B2(n14806), .A(n14805), .ZN(P1_U3124) );
  INV_X1 U16925 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16926 ( .A1(n22515), .A2(n22695), .B1(n22514), .B2(n22694), .ZN(
        n14807) );
  OAI21_X1 U16927 ( .B1(n22699), .B2(n14808), .A(n14807), .ZN(n14809) );
  AOI21_X1 U16928 ( .B1(n11247), .B2(n22703), .A(n14809), .ZN(n14810) );
  OAI21_X1 U16929 ( .B1(n14853), .B2(n14811), .A(n14810), .ZN(P1_U3122) );
  INV_X1 U16930 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14816) );
  AOI22_X1 U16931 ( .A1(n22540), .A2(n22695), .B1(n22539), .B2(n22694), .ZN(
        n14812) );
  OAI21_X1 U16932 ( .B1(n22699), .B2(n14813), .A(n14812), .ZN(n14814) );
  AOI21_X1 U16933 ( .B1(n11249), .B2(n22703), .A(n14814), .ZN(n14815) );
  OAI21_X1 U16934 ( .B1(n14853), .B2(n14816), .A(n14815), .ZN(P1_U3123) );
  OR2_X1 U16935 ( .A1(n14819), .A2(n14818), .ZN(n14820) );
  NAND2_X1 U16936 ( .A1(n14817), .A2(n14820), .ZN(n22062) );
  INV_X1 U16937 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n22056) );
  OAI222_X1 U16938 ( .A1(n22062), .A2(n20551), .B1(n22056), .B2(n20556), .C1(
        n20561), .C2(n16572), .ZN(P1_U2868) );
  NOR3_X1 U16939 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14826) );
  INV_X1 U16940 ( .A(n14822), .ZN(n16327) );
  OR2_X1 U16941 ( .A1(n16842), .A2(n16327), .ZN(n22406) );
  INV_X1 U16942 ( .A(n22406), .ZN(n22421) );
  INV_X1 U16943 ( .A(n14826), .ZN(n22392) );
  NOR2_X1 U16944 ( .A1(n22454), .A2(n22392), .ZN(n22547) );
  AOI21_X1 U16945 ( .B1(n22421), .B2(n14823), .A(n22547), .ZN(n14829) );
  OAI211_X1 U16946 ( .C1(n22419), .C2(n22223), .A(n22417), .B(n14829), .ZN(
        n14825) );
  OAI211_X1 U16947 ( .C1(n22417), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n22548) );
  INV_X1 U16948 ( .A(n22548), .ZN(n14847) );
  INV_X1 U16949 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14833) );
  INV_X1 U16950 ( .A(n22654), .ZN(n14843) );
  OAI22_X1 U16951 ( .A1(n14829), .A2(n22465), .B1(n22392), .B2(n22476), .ZN(
        n22546) );
  AOI22_X1 U16952 ( .A1(n22719), .A2(n22547), .B1(n22546), .B2(n22717), .ZN(
        n14830) );
  OAI21_X1 U16953 ( .B1(n14843), .B2(n22726), .A(n14830), .ZN(n14831) );
  AOI21_X1 U16954 ( .B1(n22660), .B2(n22720), .A(n14831), .ZN(n14832) );
  OAI21_X1 U16955 ( .B1(n14847), .B2(n14833), .A(n14832), .ZN(P1_U3048) );
  INV_X1 U16956 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16957 ( .A1(n22619), .A2(n22547), .B1(n22546), .B2(n15040), .ZN(
        n14834) );
  OAI21_X1 U16958 ( .B1(n14843), .B2(n14983), .A(n14834), .ZN(n14835) );
  AOI21_X1 U16959 ( .B1(n22660), .B2(n14557), .A(n14835), .ZN(n14836) );
  OAI21_X1 U16960 ( .B1(n14847), .B2(n14837), .A(n14836), .ZN(P1_U3046) );
  INV_X1 U16961 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16962 ( .A1(n22603), .A2(n22547), .B1(n22546), .B2(n22602), .ZN(
        n14838) );
  OAI21_X1 U16963 ( .B1(n14843), .B2(n22606), .A(n14838), .ZN(n14839) );
  AOI21_X1 U16964 ( .B1(n22660), .B2(n14669), .A(n14839), .ZN(n14840) );
  OAI21_X1 U16965 ( .B1(n14847), .B2(n14841), .A(n14840), .ZN(P1_U3045) );
  INV_X1 U16966 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U16967 ( .A1(n22648), .A2(n22547), .B1(n22546), .B2(n22647), .ZN(
        n14842) );
  OAI21_X1 U16968 ( .B1(n14843), .B2(n22652), .A(n14842), .ZN(n14844) );
  AOI21_X1 U16969 ( .B1(n22660), .B2(n22649), .A(n14844), .ZN(n14845) );
  OAI21_X1 U16970 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(P1_U3047) );
  INV_X1 U16971 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14852) );
  INV_X1 U16972 ( .A(n22703), .ZN(n14849) );
  AOI22_X1 U16973 ( .A1(n22489), .A2(n22695), .B1(n22488), .B2(n22694), .ZN(
        n14848) );
  OAI21_X1 U16974 ( .B1(n14849), .B2(n22493), .A(n14848), .ZN(n14850) );
  AOI21_X1 U16975 ( .B1(n22616), .B2(n22490), .A(n14850), .ZN(n14851) );
  OAI21_X1 U16976 ( .B1(n14853), .B2(n14852), .A(n14851), .ZN(P1_U3121) );
  AND2_X1 U16977 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  NOR2_X1 U16978 ( .A1(n14854), .A2(n14857), .ZN(n18902) );
  INV_X1 U16979 ( .A(n18902), .ZN(n14865) );
  INV_X1 U16980 ( .A(n14858), .ZN(n14862) );
  INV_X1 U16981 ( .A(n14859), .ZN(n14860) );
  OAI211_X1 U16982 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n17136), .ZN(
        n14864) );
  NAND2_X1 U16983 ( .A1(n11163), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14863) );
  OAI211_X1 U16984 ( .C1(n14865), .C2(n11163), .A(n14864), .B(n14863), .ZN(
        P2_U2877) );
  NOR2_X1 U16985 ( .A1(n14755), .A2(n14867), .ZN(n14868) );
  OR2_X1 U16986 ( .A1(n14866), .A2(n14868), .ZN(n20552) );
  INV_X1 U16987 ( .A(n16006), .ZN(n22325) );
  OAI222_X1 U16988 ( .A1(n20552), .A2(n16621), .B1(n15817), .B2(n14869), .C1(
        n15819), .C2(n22325), .ZN(P1_U2899) );
  OAI222_X1 U16989 ( .A1(n14919), .A2(n16621), .B1(n15819), .B2(n22314), .C1(
        n16612), .C2(n12090), .ZN(P1_U2901) );
  XNOR2_X1 U16990 ( .A(n14871), .B(n14870), .ZN(n14893) );
  XOR2_X1 U16991 ( .A(n14872), .B(n14873), .Z(n14890) );
  OR2_X1 U16992 ( .A1(n14875), .A2(n14874), .ZN(n14877) );
  NAND2_X1 U16993 ( .A1(n14877), .A2(n14876), .ZN(n20017) );
  INV_X1 U16994 ( .A(n14878), .ZN(n14881) );
  NOR2_X1 U16995 ( .A1(n17448), .A2(n14879), .ZN(n14880) );
  AOI211_X1 U16996 ( .C1(n17451), .C2(n14881), .A(n17593), .B(n14880), .ZN(
        n15772) );
  MUX2_X1 U16997 ( .A(n15771), .B(n15772), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n14883) );
  AOI22_X1 U16998 ( .A1(n12643), .A2(n19159), .B1(n19142), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n14882) );
  OAI211_X1 U16999 ( .C1(n19134), .C2(n20017), .A(n14883), .B(n14882), .ZN(
        n14884) );
  AOI21_X1 U17000 ( .B1(n14890), .B2(n19157), .A(n14884), .ZN(n14885) );
  OAI21_X1 U17001 ( .B1(n14893), .B2(n19123), .A(n14885), .ZN(P2_U3043) );
  INV_X1 U17002 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14887) );
  OAI22_X1 U17003 ( .A1(n17789), .A2(n14887), .B1(n14886), .B2(n17323), .ZN(
        n14889) );
  NOR2_X1 U17004 ( .A1(n17827), .A2(n17036), .ZN(n14888) );
  AOI211_X1 U17005 ( .C1(n17807), .C2(n12643), .A(n14889), .B(n14888), .ZN(
        n14892) );
  NAND2_X1 U17006 ( .A1(n14890), .A2(n17321), .ZN(n14891) );
  OAI211_X1 U17007 ( .C1(n14893), .C2(n13196), .A(n14892), .B(n14891), .ZN(
        P2_U3011) );
  OAI211_X1 U17008 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n17722), .A(n22210), 
        .B(n16450), .ZN(n14895) );
  NOR2_X1 U17009 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22214) );
  AOI21_X1 U17010 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22214), .A(n22210), 
        .ZN(n17721) );
  INV_X1 U17011 ( .A(n17721), .ZN(n14894) );
  AND2_X1 U17012 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  NOR2_X1 U17013 ( .A1(n14900), .A2(n17727), .ZN(n14897) );
  OAI21_X1 U17014 ( .B1(n14916), .B2(n14898), .A(n22181), .ZN(n22064) );
  INV_X1 U17015 ( .A(n22064), .ZN(n16329) );
  NAND2_X1 U17016 ( .A1(n22243), .A2(n22223), .ZN(n14906) );
  NAND3_X1 U17017 ( .A1(n11174), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n14906), 
        .ZN(n14899) );
  AND2_X1 U17018 ( .A1(n14900), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14901) );
  INV_X1 U17019 ( .A(n14916), .ZN(n14905) );
  INV_X1 U17020 ( .A(n14906), .ZN(n14902) );
  AND3_X1 U17021 ( .A1(n14903), .A2(n14902), .A3(n16332), .ZN(n14904) );
  INV_X1 U17022 ( .A(n22138), .ZN(n22153) );
  INV_X1 U17023 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U17024 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n16316) );
  XOR2_X1 U17025 ( .A(n15000), .B(n16316), .Z(n14911) );
  OR2_X1 U17026 ( .A1(n22254), .A2(n14906), .ZN(n17717) );
  INV_X1 U17027 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16268) );
  AND3_X1 U17028 ( .A1(n14907), .A2(n16268), .A3(n14906), .ZN(n14908) );
  AOI21_X1 U17029 ( .B1(n14909), .B2(n17717), .A(n14908), .ZN(n14910) );
  AOI22_X1 U17030 ( .A1(n22153), .A2(n14911), .B1(n11143), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14913) );
  NAND2_X1 U17031 ( .A1(n22095), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22188) );
  INV_X1 U17032 ( .A(n22095), .ZN(n16297) );
  AOI22_X1 U17033 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16297), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14912) );
  OAI211_X1 U17034 ( .C1(n15002), .C2(n22186), .A(n14913), .B(n14912), .ZN(
        n14914) );
  AOI21_X1 U17035 ( .B1(n16557), .B2(n21937), .A(n14914), .ZN(n14918) );
  NOR2_X1 U17036 ( .A1(n14916), .A2(n14915), .ZN(n22050) );
  NAND2_X1 U17037 ( .A1(n16842), .A2(n22050), .ZN(n14917) );
  OAI211_X1 U17038 ( .C1(n14919), .C2(n16329), .A(n14918), .B(n14917), .ZN(
        P1_U2837) );
  XNOR2_X1 U17039 ( .A(n11153), .B(n14921), .ZN(n14924) );
  NOR2_X1 U17040 ( .A1(n17125), .A2(n13114), .ZN(n14922) );
  AOI21_X1 U17041 ( .B1(n17520), .B2(n17125), .A(n14922), .ZN(n14923) );
  OAI21_X1 U17042 ( .B1(n14924), .B2(n17128), .A(n14923), .ZN(P2_U2875) );
  OAI21_X1 U17043 ( .B1(n14854), .B2(n14925), .A(n15127), .ZN(n18918) );
  INV_X1 U17044 ( .A(n11153), .ZN(n14926) );
  OAI211_X1 U17045 ( .C1(n14859), .C2(n14927), .A(n14926), .B(n17136), .ZN(
        n14929) );
  NAND2_X1 U17046 ( .A1(n11164), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14928) );
  OAI211_X1 U17047 ( .C1(n18918), .C2(n11164), .A(n14929), .B(n14928), .ZN(
        P2_U2876) );
  OAI21_X1 U17048 ( .B1(n14866), .B2(n14931), .A(n14930), .ZN(n20578) );
  INV_X1 U17049 ( .A(n16617), .ZN(n22330) );
  OAI222_X1 U17050 ( .A1(n20578), .A2(n16621), .B1(n15819), .B2(n22330), .C1(
        n15817), .C2(n12122), .ZN(P1_U2898) );
  OAI21_X1 U17051 ( .B1(n14956), .B2(n22711), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14935) );
  INV_X1 U17052 ( .A(n14933), .ZN(n22468) );
  NAND2_X1 U17053 ( .A1(n14934), .A2(n22468), .ZN(n14940) );
  AOI21_X1 U17054 ( .B1(n14935), .B2(n14940), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14937) );
  NOR3_X2 U17055 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17709), .A3(
        n22437), .ZN(n22574) );
  NOR2_X1 U17056 ( .A1(n14938), .A2(n22476), .ZN(n22450) );
  NOR2_X1 U17057 ( .A1(n22450), .A2(n14966), .ZN(n15010) );
  INV_X1 U17058 ( .A(n22477), .ZN(n14936) );
  NAND2_X1 U17059 ( .A1(n14936), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22449) );
  NAND2_X1 U17060 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22449), .ZN(n22457) );
  OAI211_X1 U17061 ( .C1(n14937), .C2(n22574), .A(n15010), .B(n22457), .ZN(
        n22577) );
  INV_X1 U17062 ( .A(n22577), .ZN(n14959) );
  INV_X1 U17063 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14944) );
  INV_X1 U17064 ( .A(n14938), .ZN(n14939) );
  NOR2_X1 U17065 ( .A1(n14939), .A2(n22476), .ZN(n22435) );
  INV_X1 U17066 ( .A(n22435), .ZN(n22471) );
  OAI22_X1 U17067 ( .A1(n14940), .A2(n22465), .B1(n22471), .B2(n22449), .ZN(
        n22572) );
  AOI22_X1 U17068 ( .A1(n22619), .A2(n22574), .B1(n22572), .B2(n15040), .ZN(
        n14941) );
  OAI21_X1 U17069 ( .B1(n14983), .B2(n14954), .A(n14941), .ZN(n14942) );
  AOI21_X1 U17070 ( .B1(n14956), .B2(n14557), .A(n14942), .ZN(n14943) );
  OAI21_X1 U17071 ( .B1(n14959), .B2(n14944), .A(n14943), .ZN(P1_U3150) );
  INV_X1 U17072 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U17073 ( .A1(n22648), .A2(n22574), .B1(n22572), .B2(n22647), .ZN(
        n14945) );
  OAI21_X1 U17074 ( .B1(n14954), .B2(n22652), .A(n14945), .ZN(n14946) );
  AOI21_X1 U17075 ( .B1(n14956), .B2(n22649), .A(n14946), .ZN(n14947) );
  OAI21_X1 U17076 ( .B1(n14959), .B2(n14948), .A(n14947), .ZN(P1_U3151) );
  INV_X1 U17077 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U17078 ( .A1(n22603), .A2(n22574), .B1(n22602), .B2(n22572), .ZN(
        n14949) );
  OAI21_X1 U17079 ( .B1(n14954), .B2(n22606), .A(n14949), .ZN(n14950) );
  AOI21_X1 U17080 ( .B1(n14956), .B2(n14669), .A(n14950), .ZN(n14951) );
  OAI21_X1 U17081 ( .B1(n14959), .B2(n14952), .A(n14951), .ZN(P1_U3149) );
  INV_X1 U17082 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U17083 ( .A1(n22719), .A2(n22574), .B1(n22572), .B2(n22717), .ZN(
        n14953) );
  OAI21_X1 U17084 ( .B1(n14954), .B2(n22726), .A(n14953), .ZN(n14955) );
  AOI21_X1 U17085 ( .B1(n14956), .B2(n22720), .A(n14955), .ZN(n14957) );
  OAI21_X1 U17086 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(P1_U3152) );
  NAND2_X1 U17087 ( .A1(n14960), .A2(n14961), .ZN(n14962) );
  NAND2_X1 U17088 ( .A1(n15120), .A2(n14962), .ZN(n21945) );
  OAI222_X1 U17089 ( .A1(n21945), .A2(n20551), .B1(n14963), .B2(n20556), .C1(
        n20578), .C2(n16572), .ZN(P1_U2866) );
  NOR2_X1 U17090 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14964), .ZN(
        n22559) );
  OAI21_X1 U17091 ( .B1(n14986), .B2(n22560), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14965) );
  AOI21_X1 U17092 ( .B1(n22448), .B2(n14933), .A(n22559), .ZN(n14969) );
  NAND2_X1 U17093 ( .A1(n14965), .A2(n14969), .ZN(n14967) );
  NOR2_X1 U17094 ( .A1(n22435), .A2(n14966), .ZN(n22411) );
  OAI211_X1 U17095 ( .C1(n22559), .C2(n22211), .A(n14967), .B(n22411), .ZN(
        n22561) );
  INV_X1 U17096 ( .A(n22561), .ZN(n14989) );
  INV_X1 U17097 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14973) );
  NAND3_X1 U17098 ( .A1(n22450), .A2(n22478), .A3(n22477), .ZN(n14968) );
  OAI21_X1 U17099 ( .B1(n14969), .B2(n22465), .A(n14968), .ZN(n22558) );
  AOI22_X1 U17100 ( .A1(n22719), .A2(n22559), .B1(n22717), .B2(n22558), .ZN(
        n14970) );
  OAI21_X1 U17101 ( .B1(n14984), .B2(n22726), .A(n14970), .ZN(n14971) );
  AOI21_X1 U17102 ( .B1(n14986), .B2(n22720), .A(n14971), .ZN(n14972) );
  OAI21_X1 U17103 ( .B1(n14989), .B2(n14973), .A(n14972), .ZN(P1_U3104) );
  INV_X1 U17104 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U17105 ( .A1(n22603), .A2(n22559), .B1(n22602), .B2(n22558), .ZN(
        n14974) );
  OAI21_X1 U17106 ( .B1(n14984), .B2(n22606), .A(n14974), .ZN(n14975) );
  AOI21_X1 U17107 ( .B1(n14986), .B2(n14669), .A(n14975), .ZN(n14976) );
  OAI21_X1 U17108 ( .B1(n14989), .B2(n14977), .A(n14976), .ZN(P1_U3101) );
  INV_X1 U17109 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14981) );
  AOI22_X1 U17110 ( .A1(n22648), .A2(n22559), .B1(n22647), .B2(n22558), .ZN(
        n14978) );
  OAI21_X1 U17111 ( .B1(n14984), .B2(n22652), .A(n14978), .ZN(n14979) );
  AOI21_X1 U17112 ( .B1(n14986), .B2(n22649), .A(n14979), .ZN(n14980) );
  OAI21_X1 U17113 ( .B1(n14989), .B2(n14981), .A(n14980), .ZN(P1_U3103) );
  INV_X1 U17114 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U17115 ( .A1(n22619), .A2(n22559), .B1(n15040), .B2(n22558), .ZN(
        n14982) );
  OAI21_X1 U17116 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14985) );
  AOI21_X1 U17117 ( .B1(n14986), .B2(n14557), .A(n14985), .ZN(n14987) );
  OAI21_X1 U17118 ( .B1(n14989), .B2(n14988), .A(n14987), .ZN(P1_U3102) );
  NAND2_X1 U17119 ( .A1(n14817), .A2(n14990), .ZN(n14991) );
  NAND2_X1 U17120 ( .A1(n14960), .A2(n14991), .ZN(n21955) );
  INV_X1 U17121 ( .A(n20552), .ZN(n20570) );
  NAND2_X1 U17122 ( .A1(n20570), .A2(n22064), .ZN(n14996) );
  NOR2_X1 U17123 ( .A1(n15000), .A2(n16316), .ZN(n22052) );
  NAND2_X1 U17124 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22052), .ZN(n15104) );
  NOR2_X1 U17125 ( .A1(n22138), .A2(n15104), .ZN(n15135) );
  NAND2_X1 U17126 ( .A1(n22138), .A2(n22095), .ZN(n22119) );
  INV_X1 U17127 ( .A(n22119), .ZN(n22155) );
  NOR2_X1 U17128 ( .A1(n15135), .A2(n22155), .ZN(n22059) );
  INV_X1 U17129 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21958) );
  AOI22_X1 U17130 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n22151), .B1(
        n15135), .B2(n21958), .ZN(n14992) );
  OAI211_X1 U17131 ( .C1(n22186), .C2(n20573), .A(n14992), .B(n22122), .ZN(
        n14994) );
  INV_X1 U17132 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20555) );
  NOR2_X1 U17133 ( .A1(n22191), .A2(n20555), .ZN(n14993) );
  AOI211_X1 U17134 ( .C1(n22059), .C2(P1_REIP_REG_5__SCAN_IN), .A(n14994), .B(
        n14993), .ZN(n14995) );
  OAI211_X1 U17135 ( .C1(n21955), .C2(n22202), .A(n14996), .B(n14995), .ZN(
        P1_U2835) );
  OAI21_X1 U17136 ( .B1(n14999), .B2(n14998), .A(n11209), .ZN(n21934) );
  NOR2_X1 U17137 ( .A1(n22016), .A2(n15000), .ZN(n21936) );
  AOI21_X1 U17138 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n21936), .ZN(n15001) );
  OAI21_X1 U17139 ( .B1(n20633), .B2(n15002), .A(n15001), .ZN(n15003) );
  AOI21_X1 U17140 ( .B1(n15004), .B2(n20628), .A(n15003), .ZN(n15005) );
  OAI21_X1 U17141 ( .B1(n22203), .B2(n21934), .A(n15005), .ZN(P1_U2996) );
  INV_X1 U17142 ( .A(n22667), .ZN(n15007) );
  AOI21_X1 U17143 ( .B1(n15007), .B2(n15049), .A(n22223), .ZN(n15008) );
  NOR2_X1 U17144 ( .A1(n22433), .A2(n22468), .ZN(n15013) );
  OAI21_X1 U17145 ( .B1(n15008), .B2(n15013), .A(n22211), .ZN(n15012) );
  NOR2_X1 U17146 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15009), .ZN(
        n15047) );
  INV_X1 U17147 ( .A(n15047), .ZN(n15011) );
  INV_X1 U17148 ( .A(n15010), .ZN(n22480) );
  INV_X1 U17149 ( .A(n22568), .ZN(n22580) );
  INV_X1 U17150 ( .A(n15013), .ZN(n15014) );
  INV_X1 U17151 ( .A(n22478), .ZN(n22470) );
  NAND2_X1 U17152 ( .A1(n22470), .A2(n22477), .ZN(n22394) );
  OAI22_X1 U17153 ( .A1(n15014), .A2(n22465), .B1(n22471), .B2(n22394), .ZN(
        n15046) );
  AOI22_X1 U17154 ( .A1(n22575), .A2(n15047), .B1(n22573), .B2(n15046), .ZN(
        n15015) );
  OAI21_X1 U17155 ( .B1(n15049), .B2(n22580), .A(n15015), .ZN(n15016) );
  AOI21_X1 U17156 ( .B1(n22667), .B2(n22576), .A(n15016), .ZN(n15017) );
  OAI21_X1 U17157 ( .B1(n15053), .B2(n15018), .A(n15017), .ZN(P1_U3068) );
  INV_X1 U17158 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U17159 ( .A1(n22489), .A2(n15047), .B1(n22488), .B2(n15046), .ZN(
        n15019) );
  OAI21_X1 U17160 ( .B1(n15049), .B2(n22493), .A(n15019), .ZN(n15020) );
  AOI21_X1 U17161 ( .B1(n22667), .B2(n22490), .A(n15020), .ZN(n15021) );
  OAI21_X1 U17162 ( .B1(n15053), .B2(n15022), .A(n15021), .ZN(P1_U3065) );
  INV_X1 U17163 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U17164 ( .A1(n22648), .A2(n15047), .B1(n22647), .B2(n15046), .ZN(
        n15023) );
  OAI21_X1 U17165 ( .B1(n22635), .B2(n15049), .A(n15023), .ZN(n15024) );
  AOI21_X1 U17166 ( .B1(n22667), .B2(n22641), .A(n15024), .ZN(n15025) );
  OAI21_X1 U17167 ( .B1(n15053), .B2(n15026), .A(n15025), .ZN(P1_U3071) );
  INV_X1 U17168 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15030) );
  AOI22_X1 U17169 ( .A1(n22540), .A2(n15047), .B1(n22539), .B2(n15046), .ZN(
        n15027) );
  OAI21_X1 U17170 ( .B1(n15049), .B2(n11248), .A(n15027), .ZN(n15028) );
  AOI21_X1 U17171 ( .B1(n22667), .B2(n22541), .A(n15028), .ZN(n15029) );
  OAI21_X1 U17172 ( .B1(n15053), .B2(n15030), .A(n15029), .ZN(P1_U3067) );
  INV_X1 U17173 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15034) );
  AOI22_X1 U17174 ( .A1(n22719), .A2(n15047), .B1(n22717), .B2(n15046), .ZN(
        n15031) );
  OAI21_X1 U17175 ( .B1(n22687), .B2(n15049), .A(n15031), .ZN(n15032) );
  AOI21_X1 U17176 ( .B1(n22667), .B2(n22702), .A(n15032), .ZN(n15033) );
  OAI21_X1 U17177 ( .B1(n15053), .B2(n15034), .A(n15033), .ZN(P1_U3072) );
  INV_X1 U17178 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U17179 ( .A1(n22603), .A2(n15047), .B1(n22602), .B2(n15046), .ZN(
        n15035) );
  OAI21_X1 U17180 ( .B1(n15036), .B2(n15049), .A(n15035), .ZN(n15037) );
  AOI21_X1 U17181 ( .B1(n22667), .B2(n22595), .A(n15037), .ZN(n15038) );
  OAI21_X1 U17182 ( .B1(n15053), .B2(n15039), .A(n15038), .ZN(P1_U3069) );
  INV_X1 U17183 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15045) );
  AOI22_X1 U17184 ( .A1(n22619), .A2(n15047), .B1(n15040), .B2(n15046), .ZN(
        n15041) );
  OAI21_X1 U17185 ( .B1(n15042), .B2(n15049), .A(n15041), .ZN(n15043) );
  AOI21_X1 U17186 ( .B1(n22667), .B2(n22620), .A(n15043), .ZN(n15044) );
  OAI21_X1 U17187 ( .B1(n15053), .B2(n15045), .A(n15044), .ZN(P1_U3070) );
  INV_X1 U17188 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U17189 ( .A1(n22515), .A2(n15047), .B1(n22514), .B2(n15046), .ZN(
        n15048) );
  OAI21_X1 U17190 ( .B1(n15049), .B2(n11246), .A(n15048), .ZN(n15050) );
  AOI21_X1 U17191 ( .B1(n22667), .B2(n22516), .A(n15050), .ZN(n15051) );
  OAI21_X1 U17192 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(P1_U3066) );
  XNOR2_X1 U17193 ( .A(n15054), .B(n15055), .ZN(n15077) );
  OAI21_X1 U17194 ( .B1(n15056), .B2(n15672), .A(n15057), .ZN(n15075) );
  OR2_X1 U17195 ( .A1(n15058), .A2(n15771), .ZN(n15671) );
  OAI21_X1 U17196 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17497), .A(
        n15772), .ZN(n15675) );
  INV_X1 U17197 ( .A(n15675), .ZN(n15060) );
  NAND2_X1 U17198 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19142), .ZN(n15059) );
  OAI221_X1 U17199 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15671), .C1(
        n15672), .C2(n15060), .A(n15059), .ZN(n15069) );
  INV_X1 U17200 ( .A(n14876), .ZN(n15061) );
  OR2_X1 U17201 ( .A1(n15062), .A2(n15061), .ZN(n15066) );
  CLKBUF_X1 U17202 ( .A(n15063), .Z(n15064) );
  INV_X1 U17203 ( .A(n15064), .ZN(n15065) );
  AND2_X1 U17204 ( .A1(n15066), .A2(n15065), .ZN(n20074) );
  INV_X1 U17205 ( .A(n20074), .ZN(n15067) );
  OAI22_X1 U17206 ( .A1(n15073), .A2(n19130), .B1(n19134), .B2(n15067), .ZN(
        n15068) );
  AOI211_X1 U17207 ( .C1(n15075), .C2(n19157), .A(n15069), .B(n15068), .ZN(
        n15070) );
  OAI21_X1 U17208 ( .B1(n15077), .B2(n19123), .A(n15070), .ZN(P2_U3042) );
  OAI22_X1 U17209 ( .A1(n17027), .A2(n17789), .B1(n13333), .B2(n18958), .ZN(
        n15071) );
  AOI21_X1 U17210 ( .B1(n17777), .B2(n17025), .A(n15071), .ZN(n15072) );
  OAI21_X1 U17211 ( .B1(n13199), .B2(n15073), .A(n15072), .ZN(n15074) );
  AOI21_X1 U17212 ( .B1(n15075), .B2(n17820), .A(n15074), .ZN(n15076) );
  OAI21_X1 U17213 ( .B1(n15077), .B2(n13196), .A(n15076), .ZN(P2_U3010) );
  NAND2_X1 U17214 ( .A1(n22188), .A2(n22186), .ZN(n15078) );
  AOI22_X1 U17215 ( .A1(n11143), .A2(P1_EBX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n15078), .ZN(n15082) );
  NAND2_X1 U17216 ( .A1(n22119), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15081) );
  NAND2_X1 U17217 ( .A1(n16557), .A2(n15079), .ZN(n15080) );
  NAND3_X1 U17218 ( .A1(n15082), .A2(n15081), .A3(n15080), .ZN(n15083) );
  AOI21_X1 U17219 ( .B1(n16804), .B2(n22050), .A(n15083), .ZN(n15084) );
  OAI21_X1 U17220 ( .B1(n15085), .B2(n16329), .A(n15084), .ZN(P1_U2840) );
  OAI21_X1 U17221 ( .B1(n15088), .B2(n15087), .A(n15086), .ZN(n15651) );
  INV_X1 U17222 ( .A(n15838), .ZN(n21953) );
  AOI22_X1 U17223 ( .A1(n21985), .A2(n15089), .B1(n15090), .B2(n21953), .ZN(
        n21951) );
  NOR4_X1 U17224 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21951), .A3(
        n21970), .A4(n21950), .ZN(n15097) );
  INV_X1 U17225 ( .A(n21951), .ZN(n15871) );
  NAND3_X1 U17226 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21970), .A3(
        n15871), .ZN(n21967) );
  INV_X1 U17227 ( .A(n15089), .ZN(n21954) );
  AOI21_X1 U17228 ( .B1(n21985), .B2(n21954), .A(n21979), .ZN(n21942) );
  OAI211_X1 U17229 ( .C1(n21944), .C2(n15090), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n21942), .ZN(n15091) );
  NAND2_X1 U17230 ( .A1(n16776), .A2(n15091), .ZN(n21969) );
  AOI21_X1 U17231 ( .B1(n21967), .B2(n21969), .A(n15092), .ZN(n15096) );
  OAI21_X1 U17232 ( .B1(n11186), .B2(n15094), .A(n15093), .ZN(n15684) );
  NAND2_X1 U17233 ( .A1(n22040), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15645) );
  OAI21_X1 U17234 ( .B1(n15684), .B2(n22017), .A(n15645), .ZN(n15095) );
  NOR3_X1 U17235 ( .A1(n15097), .A2(n15096), .A3(n15095), .ZN(n15098) );
  OAI21_X1 U17236 ( .B1(n15651), .B2(n22033), .A(n15098), .ZN(P1_U3023) );
  OAI21_X1 U17237 ( .B1(n11202), .B2(n15103), .A(n15102), .ZN(n15882) );
  INV_X1 U17238 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22074) );
  INV_X1 U17239 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n15137) );
  NOR4_X1 U17240 ( .A1(n22074), .A2(n15137), .A3(n21958), .A4(n15104), .ZN(
        n15635) );
  NAND2_X1 U17241 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15635), .ZN(n15106) );
  NOR2_X1 U17242 ( .A1(n22138), .A2(n15106), .ZN(n22080) );
  INV_X1 U17243 ( .A(n22080), .ZN(n15105) );
  INV_X1 U17244 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15690) );
  NOR2_X1 U17245 ( .A1(n15105), .A2(n15690), .ZN(n22089) );
  INV_X1 U17246 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15870) );
  NOR3_X1 U17247 ( .A1(n15870), .A2(n15690), .A3(n15106), .ZN(n15748) );
  INV_X1 U17248 ( .A(n15748), .ZN(n15952) );
  AOI21_X1 U17249 ( .B1(n22153), .B2(n15952), .A(n16297), .ZN(n15956) );
  INV_X1 U17250 ( .A(n15885), .ZN(n15113) );
  INV_X1 U17251 ( .A(n15699), .ZN(n15110) );
  NAND2_X1 U17252 ( .A1(n15108), .A2(n15107), .ZN(n15109) );
  NAND2_X1 U17253 ( .A1(n15110), .A2(n15109), .ZN(n15869) );
  AOI22_X1 U17254 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n22151), .B1(
        n11143), .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n15111) );
  OAI211_X1 U17255 ( .C1(n15869), .C2(n22202), .A(n15111), .B(n22122), .ZN(
        n15112) );
  AOI21_X1 U17256 ( .B1(n22195), .B2(n15113), .A(n15112), .ZN(n15114) );
  OAI21_X1 U17257 ( .B1(n15956), .B2(n15870), .A(n15114), .ZN(n15115) );
  AOI21_X1 U17258 ( .B1(n22089), .B2(n15952), .A(n15115), .ZN(n15116) );
  OAI21_X1 U17259 ( .B1(n15882), .B2(n22181), .A(n15116), .ZN(P1_U2830) );
  OR2_X1 U17260 ( .A1(n14930), .A2(n15117), .ZN(n15632) );
  INV_X1 U17261 ( .A(n15632), .ZN(n15118) );
  AOI21_X1 U17262 ( .B1(n15117), .B2(n14930), .A(n15118), .ZN(n22077) );
  INV_X1 U17263 ( .A(n22077), .ZN(n15133) );
  AND2_X1 U17264 ( .A1(n15120), .A2(n15119), .ZN(n15121) );
  NOR2_X1 U17265 ( .A1(n11186), .A2(n15121), .ZN(n22068) );
  AOI22_X1 U17266 ( .A1(n22068), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n15123) );
  OAI21_X1 U17267 ( .B1(n15133), .B2(n16572), .A(n15123), .ZN(P1_U2865) );
  AND2_X1 U17268 ( .A1(n15125), .A2(n15124), .ZN(n15128) );
  NOR2_X1 U17269 ( .A1(n15127), .A2(n15126), .ZN(n15655) );
  OAI211_X1 U17270 ( .C1(n11243), .C2(n15130), .A(n17136), .B(n15129), .ZN(
        n15132) );
  NAND2_X1 U17271 ( .A1(n11163), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n15131) );
  OAI211_X1 U17272 ( .C1(n19122), .C2(n11163), .A(n15132), .B(n15131), .ZN(
        P2_U2874) );
  INV_X1 U17273 ( .A(n16609), .ZN(n22335) );
  OAI222_X1 U17274 ( .A1(n15133), .A2(n16621), .B1(n15819), .B2(n22335), .C1(
        n16612), .C2(n12052), .ZN(P1_U2897) );
  MUX2_X1 U17275 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15902), .Z(
        n16591) );
  INV_X1 U17276 ( .A(n16591), .ZN(n22354) );
  OAI222_X1 U17277 ( .A1(n15882), .A2(n16621), .B1(n15819), .B2(n22354), .C1(
        n15134), .C2(n16612), .ZN(P1_U2894) );
  OAI222_X1 U17278 ( .A1(n15869), .A2(n20551), .B1(n15484), .B2(n20556), .C1(
        n15882), .C2(n16572), .ZN(P1_U2862) );
  AND2_X1 U17279 ( .A1(n15135), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15136) );
  NAND2_X1 U17280 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n15136), .ZN(n22075) );
  NAND2_X1 U17281 ( .A1(n22119), .A2(n22075), .ZN(n22073) );
  INV_X1 U17282 ( .A(n15136), .ZN(n15144) );
  NAND2_X1 U17283 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15140) );
  OAI22_X1 U17284 ( .A1(n15137), .A2(n22073), .B1(n22202), .B2(n21945), .ZN(
        n15138) );
  NOR2_X1 U17285 ( .A1(n22139), .A2(n15138), .ZN(n15139) );
  OAI211_X1 U17286 ( .C1(n22186), .C2(n20582), .A(n15140), .B(n15139), .ZN(
        n15142) );
  NOR2_X1 U17287 ( .A1(n20578), .A2(n22181), .ZN(n15141) );
  AOI211_X1 U17288 ( .C1(n11143), .C2(P1_EBX_REG_6__SCAN_IN), .A(n15142), .B(
        n15141), .ZN(n15143) );
  OAI21_X1 U17289 ( .B1(n22073), .B2(n15144), .A(n15143), .ZN(P1_U2834) );
  XOR2_X1 U17290 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .Z(n15148) );
  XNOR2_X1 U17291 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n15147)
         );
  XNOR2_X1 U17292 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .ZN(n15146)
         );
  XNOR2_X1 U17293 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .ZN(n15145)
         );
  NOR4_X1 U17294 ( .A1(n15148), .A2(n15147), .A3(n15146), .A4(n15145), .ZN(
        n15517) );
  XNOR2_X1 U17295 ( .A(n14664), .B(keyinput_4), .ZN(n15157) );
  XOR2_X1 U17296 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .Z(n15153)
         );
  XOR2_X1 U17297 ( .A(DATAI_30_), .B(keyinput_2), .Z(n15152) );
  XNOR2_X1 U17298 ( .A(n15149), .B(keyinput_1), .ZN(n15151) );
  XNOR2_X1 U17299 ( .A(DATAI_29_), .B(keyinput_3), .ZN(n15150) );
  NAND4_X1 U17300 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        n15156) );
  XNOR2_X1 U17301 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n15155) );
  XOR2_X1 U17302 ( .A(DATAI_27_), .B(keyinput_5), .Z(n15154) );
  AOI211_X1 U17303 ( .C1(n15157), .C2(n15156), .A(n15155), .B(n15154), .ZN(
        n15160) );
  XOR2_X1 U17304 ( .A(DATAI_25_), .B(keyinput_7), .Z(n15159) );
  XNOR2_X1 U17305 ( .A(DATAI_24_), .B(keyinput_8), .ZN(n15158) );
  OAI21_X1 U17306 ( .B1(n15160), .B2(n15159), .A(n15158), .ZN(n15164) );
  XNOR2_X1 U17307 ( .A(DATAI_23_), .B(keyinput_9), .ZN(n15163) );
  XNOR2_X1 U17308 ( .A(DATAI_21_), .B(keyinput_11), .ZN(n15162) );
  XNOR2_X1 U17309 ( .A(DATAI_22_), .B(keyinput_10), .ZN(n15161) );
  AOI211_X1 U17310 ( .C1(n15164), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15171) );
  XNOR2_X1 U17311 ( .A(DATAI_20_), .B(keyinput_12), .ZN(n15170) );
  XOR2_X1 U17312 ( .A(DATAI_17_), .B(keyinput_15), .Z(n15168) );
  XNOR2_X1 U17313 ( .A(DATAI_18_), .B(keyinput_14), .ZN(n15167) );
  XNOR2_X1 U17314 ( .A(DATAI_19_), .B(keyinput_13), .ZN(n15166) );
  XNOR2_X1 U17315 ( .A(DATAI_16_), .B(keyinput_16), .ZN(n15165) );
  NOR4_X1 U17316 ( .A1(n15168), .A2(n15167), .A3(n15166), .A4(n15165), .ZN(
        n15169) );
  OAI21_X1 U17317 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15176) );
  XNOR2_X1 U17318 ( .A(n15172), .B(keyinput_17), .ZN(n15175) );
  XOR2_X1 U17319 ( .A(DATAI_13_), .B(keyinput_19), .Z(n15174) );
  XOR2_X1 U17320 ( .A(DATAI_14_), .B(keyinput_18), .Z(n15173) );
  AOI211_X1 U17321 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15179) );
  XOR2_X1 U17322 ( .A(DATAI_12_), .B(keyinput_20), .Z(n15178) );
  XNOR2_X1 U17323 ( .A(DATAI_11_), .B(keyinput_21), .ZN(n15177) );
  NOR3_X1 U17324 ( .A1(n15179), .A2(n15178), .A3(n15177), .ZN(n15182) );
  XOR2_X1 U17325 ( .A(DATAI_10_), .B(keyinput_22), .Z(n15181) );
  XOR2_X1 U17326 ( .A(DATAI_9_), .B(keyinput_23), .Z(n15180) );
  OAI21_X1 U17327 ( .B1(n15182), .B2(n15181), .A(n15180), .ZN(n15186) );
  XOR2_X1 U17328 ( .A(DATAI_7_), .B(keyinput_25), .Z(n15185) );
  XOR2_X1 U17329 ( .A(DATAI_8_), .B(keyinput_24), .Z(n15184) );
  XNOR2_X1 U17330 ( .A(DATAI_6_), .B(keyinput_26), .ZN(n15183) );
  NAND4_X1 U17331 ( .A1(n15186), .A2(n15185), .A3(n15184), .A4(n15183), .ZN(
        n15190) );
  XNOR2_X1 U17332 ( .A(DATAI_5_), .B(keyinput_27), .ZN(n15189) );
  XNOR2_X1 U17333 ( .A(DATAI_3_), .B(keyinput_29), .ZN(n15188) );
  XNOR2_X1 U17334 ( .A(DATAI_4_), .B(keyinput_28), .ZN(n15187) );
  AOI211_X1 U17335 ( .C1(n15190), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15196) );
  XOR2_X1 U17336 ( .A(DATAI_2_), .B(keyinput_30), .Z(n15195) );
  XOR2_X1 U17337 ( .A(HOLD), .B(keyinput_33), .Z(n15193) );
  XNOR2_X1 U17338 ( .A(DATAI_1_), .B(keyinput_31), .ZN(n15192) );
  XNOR2_X1 U17339 ( .A(DATAI_0_), .B(keyinput_32), .ZN(n15191) );
  NOR3_X1 U17340 ( .A1(n15193), .A2(n15192), .A3(n15191), .ZN(n15194) );
  OAI21_X1 U17341 ( .B1(n15196), .B2(n15195), .A(n15194), .ZN(n15203) );
  XNOR2_X1 U17342 ( .A(NA), .B(keyinput_34), .ZN(n15202) );
  XNOR2_X1 U17343 ( .A(READY1), .B(keyinput_36), .ZN(n15200) );
  XNOR2_X1 U17344 ( .A(BS16), .B(keyinput_35), .ZN(n15199) );
  XNOR2_X1 U17345 ( .A(READY2), .B(keyinput_37), .ZN(n15198) );
  XNOR2_X1 U17346 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_38), .ZN(
        n15197) );
  NAND4_X1 U17347 ( .A1(n15200), .A2(n15199), .A3(n15198), .A4(n15197), .ZN(
        n15201) );
  AOI21_X1 U17348 ( .B1(n15203), .B2(n15202), .A(n15201), .ZN(n15206) );
  INV_X1 U17349 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17730) );
  XNOR2_X1 U17350 ( .A(n17730), .B(keyinput_39), .ZN(n15205) );
  XNOR2_X1 U17351 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_40), .ZN(n15204)
         );
  OAI21_X1 U17352 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15210) );
  XNOR2_X1 U17353 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n15209) );
  INV_X1 U17354 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20638) );
  XNOR2_X1 U17355 ( .A(n20638), .B(keyinput_42), .ZN(n15208) );
  XOR2_X1 U17356 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .Z(
        n15207) );
  AOI211_X1 U17357 ( .C1(n15210), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        n15217) );
  XNOR2_X1 U17358 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(keyinput_44), .ZN(n15216)
         );
  XOR2_X1 U17359 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .Z(n15214) );
  XOR2_X1 U17360 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .Z(n15213) );
  XNOR2_X1 U17361 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_45), .ZN(n15212) );
  XNOR2_X1 U17362 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .ZN(
        n15211) );
  NOR4_X1 U17363 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        n15215) );
  OAI21_X1 U17364 ( .B1(n15217), .B2(n15216), .A(n15215), .ZN(n15223) );
  INV_X1 U17365 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20535) );
  XNOR2_X1 U17366 ( .A(n20535), .B(keyinput_49), .ZN(n15222) );
  XOR2_X1 U17367 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .Z(
        n15220) );
  XNOR2_X1 U17368 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_50), .ZN(
        n15219) );
  XNOR2_X1 U17369 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .ZN(n15218)
         );
  NAND3_X1 U17370 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15221) );
  AOI21_X1 U17371 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15226) );
  XOR2_X1 U17372 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .Z(n15225) );
  XNOR2_X1 U17373 ( .A(n16480), .B(keyinput_54), .ZN(n15224) );
  NOR3_X1 U17374 ( .A1(n15226), .A2(n15225), .A3(n15224), .ZN(n15243) );
  INV_X1 U17375 ( .A(keyinput_55), .ZN(n15227) );
  XNOR2_X1 U17376 ( .A(n15227), .B(P1_REIP_REG_28__SCAN_IN), .ZN(n15231) );
  XNOR2_X1 U17377 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n15230)
         );
  XNOR2_X1 U17378 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .ZN(n15229)
         );
  XNOR2_X1 U17379 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_58), .ZN(n15228)
         );
  NAND4_X1 U17380 ( .A1(n15231), .A2(n15230), .A3(n15229), .A4(n15228), .ZN(
        n15242) );
  INV_X1 U17381 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n16672) );
  INV_X1 U17382 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n16679) );
  INV_X1 U17383 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n22131) );
  AOI22_X1 U17384 ( .A1(n16679), .A2(keyinput_60), .B1(keyinput_65), .B2(
        n22131), .ZN(n15234) );
  AOI22_X1 U17385 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_64), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .ZN(n15233) );
  INV_X1 U17386 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n16276) );
  AOI22_X1 U17387 ( .A1(n16672), .A2(keyinput_59), .B1(keyinput_61), .B2(
        n16276), .ZN(n15232) );
  AND3_X1 U17388 ( .A1(n15234), .A2(n15233), .A3(n15232), .ZN(n15235) );
  OAI21_X1 U17389 ( .B1(n16672), .B2(keyinput_59), .A(n15235), .ZN(n15239) );
  OAI22_X1 U17390 ( .A1(n16679), .A2(keyinput_60), .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .ZN(n15238) );
  OAI22_X1 U17391 ( .A1(n16276), .A2(keyinput_61), .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_64), .ZN(n15237) );
  NOR2_X1 U17392 ( .A1(n22131), .A2(keyinput_65), .ZN(n15236) );
  NOR4_X1 U17393 ( .A1(n15239), .A2(n15238), .A3(n15237), .A4(n15236), .ZN(
        n15241) );
  XNOR2_X1 U17394 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .ZN(n15240)
         );
  OAI211_X1 U17395 ( .C1(n15243), .C2(n15242), .A(n15241), .B(n15240), .ZN(
        n15247) );
  XOR2_X1 U17396 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_66), .Z(n15246) );
  XNOR2_X1 U17397 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_68), .ZN(n15245)
         );
  XNOR2_X1 U17398 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .ZN(n15244)
         );
  NAND4_X1 U17399 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15249) );
  XOR2_X1 U17400 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .Z(n15248) );
  NAND2_X1 U17401 ( .A1(n15249), .A2(n15248), .ZN(n15253) );
  INV_X1 U17402 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20589) );
  XNOR2_X1 U17403 ( .A(n20589), .B(keyinput_72), .ZN(n15252) );
  INV_X1 U17404 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15977) );
  XNOR2_X1 U17405 ( .A(n15977), .B(keyinput_70), .ZN(n15251) );
  XNOR2_X1 U17406 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_71), .ZN(n15250)
         );
  NAND4_X1 U17407 ( .A1(n15253), .A2(n15252), .A3(n15251), .A4(n15250), .ZN(
        n15256) );
  XOR2_X1 U17408 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .Z(n15255) );
  XNOR2_X1 U17409 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .ZN(n15254)
         );
  AOI21_X1 U17410 ( .B1(n15256), .B2(n15255), .A(n15254), .ZN(n15259) );
  XNOR2_X1 U17411 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .ZN(n15258)
         );
  XNOR2_X1 U17412 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .ZN(n15257)
         );
  NOR3_X1 U17413 ( .A1(n15259), .A2(n15258), .A3(n15257), .ZN(n15262) );
  XOR2_X1 U17414 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_77), .Z(n15261) );
  XNOR2_X1 U17415 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .ZN(n15260)
         );
  OAI21_X1 U17416 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15269) );
  XNOR2_X1 U17417 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .ZN(n15268)
         );
  XOR2_X1 U17418 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .Z(n15266) );
  XOR2_X1 U17419 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .Z(n15265) );
  XNOR2_X1 U17420 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .ZN(n15264)
         );
  XNOR2_X1 U17421 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .ZN(n15263)
         );
  NAND4_X1 U17422 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15267) );
  AOI21_X1 U17423 ( .B1(n15269), .B2(n15268), .A(n15267), .ZN(n15272) );
  XNOR2_X1 U17424 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .ZN(n15271)
         );
  XOR2_X1 U17425 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .Z(n15270) );
  OAI21_X1 U17426 ( .B1(n15272), .B2(n15271), .A(n15270), .ZN(n15275) );
  XOR2_X1 U17427 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .Z(n15274) );
  XNOR2_X1 U17428 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_87), .ZN(n15273)
         );
  NAND3_X1 U17429 ( .A1(n15275), .A2(n15274), .A3(n15273), .ZN(n15278) );
  XOR2_X1 U17430 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_88), .Z(n15277) );
  XOR2_X1 U17431 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .Z(n15276) );
  AOI21_X1 U17432 ( .B1(n15278), .B2(n15277), .A(n15276), .ZN(n15282) );
  XNOR2_X1 U17433 ( .A(n22190), .B(keyinput_91), .ZN(n15281) );
  XOR2_X1 U17434 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n15280) );
  XNOR2_X1 U17435 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .ZN(n15279)
         );
  NOR4_X1 U17436 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        n15286) );
  XNOR2_X1 U17437 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_93), .ZN(n15285)
         );
  XOR2_X1 U17438 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .Z(n15284) );
  XOR2_X1 U17439 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .Z(n15283) );
  OAI211_X1 U17440 ( .C1(n15286), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15289) );
  XOR2_X1 U17441 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_96), .Z(n15288) );
  XNOR2_X1 U17442 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_97), .ZN(n15287)
         );
  NAND3_X1 U17443 ( .A1(n15289), .A2(n15288), .A3(n15287), .ZN(n15292) );
  XOR2_X1 U17444 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .Z(n15291) );
  XNOR2_X1 U17445 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .ZN(n15290)
         );
  NAND3_X1 U17446 ( .A1(n15292), .A2(n15291), .A3(n15290), .ZN(n15295) );
  XNOR2_X1 U17447 ( .A(n22104), .B(keyinput_101), .ZN(n15294) );
  INV_X1 U17448 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15801) );
  XNOR2_X1 U17449 ( .A(n15801), .B(keyinput_100), .ZN(n15293) );
  NAND3_X1 U17450 ( .A1(n15295), .A2(n15294), .A3(n15293), .ZN(n15298) );
  XOR2_X1 U17451 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .Z(n15297) );
  XOR2_X1 U17452 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .Z(n15296) );
  NAND3_X1 U17453 ( .A1(n15298), .A2(n15297), .A3(n15296), .ZN(n15301) );
  XNOR2_X1 U17454 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .ZN(n15300)
         );
  XNOR2_X1 U17455 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_105), .ZN(n15299)
         );
  NAND3_X1 U17456 ( .A1(n15301), .A2(n15300), .A3(n15299), .ZN(n15304) );
  XOR2_X1 U17457 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_106), .Z(n15303) );
  XNOR2_X1 U17458 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n15302)
         );
  AOI21_X1 U17459 ( .B1(n15304), .B2(n15303), .A(n15302), .ZN(n15311) );
  XNOR2_X1 U17460 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .ZN(n15310)
         );
  XNOR2_X1 U17461 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_110), .ZN(n15309)
         );
  XOR2_X1 U17462 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .Z(n15307) );
  XNOR2_X1 U17463 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15306)
         );
  XNOR2_X1 U17464 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .ZN(n15305)
         );
  NAND3_X1 U17465 ( .A1(n15307), .A2(n15306), .A3(n15305), .ZN(n15308) );
  NOR4_X1 U17466 ( .A1(n15311), .A2(n15310), .A3(n15309), .A4(n15308), .ZN(
        n15313) );
  XNOR2_X1 U17467 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_113), .ZN(n15312)
         );
  NOR2_X1 U17468 ( .A1(n15313), .A2(n15312), .ZN(n15322) );
  INV_X1 U17469 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n15316) );
  AOI22_X1 U17470 ( .A1(n15316), .A2(keyinput_116), .B1(keyinput_114), .B2(
        n15315), .ZN(n15314) );
  OAI221_X1 U17471 ( .B1(n15316), .B2(keyinput_116), .C1(n15315), .C2(
        keyinput_114), .A(n15314), .ZN(n15321) );
  INV_X1 U17472 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n22375) );
  AOI22_X1 U17473 ( .A1(n15318), .A2(keyinput_115), .B1(n22375), .B2(
        keyinput_118), .ZN(n15317) );
  OAI221_X1 U17474 ( .B1(n15318), .B2(keyinput_115), .C1(n22375), .C2(
        keyinput_118), .A(n15317), .ZN(n15320) );
  XNOR2_X1 U17475 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n15319)
         );
  NOR4_X1 U17476 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        n15325) );
  XOR2_X1 U17477 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .Z(n15324) );
  XOR2_X1 U17478 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_120), .Z(n15323) );
  OAI21_X1 U17479 ( .B1(n15325), .B2(n15324), .A(n15323), .ZN(n15329) );
  XOR2_X1 U17480 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_123), .Z(n15328) );
  XNOR2_X1 U17481 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_121), .ZN(n15327)
         );
  XNOR2_X1 U17482 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_122), .ZN(n15326)
         );
  NAND4_X1 U17483 ( .A1(n15329), .A2(n15328), .A3(n15327), .A4(n15326), .ZN(
        n15516) );
  INV_X1 U17484 ( .A(keyinput_252), .ZN(n15330) );
  XNOR2_X1 U17485 ( .A(n15330), .B(P1_EAX_REG_23__SCAN_IN), .ZN(n15334) );
  XNOR2_X1 U17486 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .ZN(n15333)
         );
  XNOR2_X1 U17487 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .ZN(n15332)
         );
  XNOR2_X1 U17488 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n15331)
         );
  NAND4_X1 U17489 ( .A1(n15334), .A2(n15333), .A3(n15332), .A4(n15331), .ZN(
        n15515) );
  XOR2_X1 U17490 ( .A(DATAI_29_), .B(keyinput_131), .Z(n15338) );
  XNOR2_X1 U17491 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .ZN(
        n15337) );
  XNOR2_X1 U17492 ( .A(DATAI_31_), .B(keyinput_129), .ZN(n15336) );
  XNOR2_X1 U17493 ( .A(DATAI_30_), .B(keyinput_130), .ZN(n15335) );
  NOR4_X1 U17494 ( .A1(n15338), .A2(n15337), .A3(n15336), .A4(n15335), .ZN(
        n15342) );
  XNOR2_X1 U17495 ( .A(DATAI_28_), .B(keyinput_132), .ZN(n15341) );
  XOR2_X1 U17496 ( .A(DATAI_27_), .B(keyinput_133), .Z(n15340) );
  XNOR2_X1 U17497 ( .A(DATAI_26_), .B(keyinput_134), .ZN(n15339) );
  OAI211_X1 U17498 ( .C1(n15342), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        n15345) );
  XNOR2_X1 U17499 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n15344) );
  XOR2_X1 U17500 ( .A(DATAI_24_), .B(keyinput_136), .Z(n15343) );
  AOI21_X1 U17501 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15349) );
  XNOR2_X1 U17502 ( .A(DATAI_23_), .B(keyinput_137), .ZN(n15348) );
  XNOR2_X1 U17503 ( .A(DATAI_22_), .B(keyinput_138), .ZN(n15347) );
  XNOR2_X1 U17504 ( .A(DATAI_21_), .B(keyinput_139), .ZN(n15346) );
  OAI211_X1 U17505 ( .C1(n15349), .C2(n15348), .A(n15347), .B(n15346), .ZN(
        n15356) );
  XNOR2_X1 U17506 ( .A(DATAI_20_), .B(keyinput_140), .ZN(n15355) );
  XOR2_X1 U17507 ( .A(DATAI_17_), .B(keyinput_143), .Z(n15353) );
  XOR2_X1 U17508 ( .A(DATAI_18_), .B(keyinput_142), .Z(n15352) );
  XOR2_X1 U17509 ( .A(DATAI_16_), .B(keyinput_144), .Z(n15351) );
  XNOR2_X1 U17510 ( .A(n14579), .B(keyinput_141), .ZN(n15350) );
  NAND4_X1 U17511 ( .A1(n15353), .A2(n15352), .A3(n15351), .A4(n15350), .ZN(
        n15354) );
  AOI21_X1 U17512 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15360) );
  XNOR2_X1 U17513 ( .A(DATAI_15_), .B(keyinput_145), .ZN(n15359) );
  XOR2_X1 U17514 ( .A(DATAI_14_), .B(keyinput_146), .Z(n15358) );
  XOR2_X1 U17515 ( .A(DATAI_13_), .B(keyinput_147), .Z(n15357) );
  OAI211_X1 U17516 ( .C1(n15360), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15363) );
  XOR2_X1 U17517 ( .A(DATAI_12_), .B(keyinput_148), .Z(n15362) );
  XNOR2_X1 U17518 ( .A(DATAI_11_), .B(keyinput_149), .ZN(n15361) );
  NAND3_X1 U17519 ( .A1(n15363), .A2(n15362), .A3(n15361), .ZN(n15366) );
  XNOR2_X1 U17520 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n15365) );
  XNOR2_X1 U17521 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n15364) );
  AOI21_X1 U17522 ( .B1(n15366), .B2(n15365), .A(n15364), .ZN(n15370) );
  XOR2_X1 U17523 ( .A(DATAI_6_), .B(keyinput_154), .Z(n15369) );
  XNOR2_X1 U17524 ( .A(DATAI_7_), .B(keyinput_153), .ZN(n15368) );
  XNOR2_X1 U17525 ( .A(DATAI_8_), .B(keyinput_152), .ZN(n15367) );
  NOR4_X1 U17526 ( .A1(n15370), .A2(n15369), .A3(n15368), .A4(n15367), .ZN(
        n15374) );
  XOR2_X1 U17527 ( .A(DATAI_5_), .B(keyinput_155), .Z(n15373) );
  XOR2_X1 U17528 ( .A(DATAI_3_), .B(keyinput_157), .Z(n15372) );
  XNOR2_X1 U17529 ( .A(DATAI_4_), .B(keyinput_156), .ZN(n15371) );
  OAI211_X1 U17530 ( .C1(n15374), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15380) );
  XNOR2_X1 U17531 ( .A(DATAI_2_), .B(keyinput_158), .ZN(n15379) );
  XOR2_X1 U17532 ( .A(HOLD), .B(keyinput_161), .Z(n15377) );
  XOR2_X1 U17533 ( .A(DATAI_1_), .B(keyinput_159), .Z(n15376) );
  XNOR2_X1 U17534 ( .A(DATAI_0_), .B(keyinput_160), .ZN(n15375) );
  NAND3_X1 U17535 ( .A1(n15377), .A2(n15376), .A3(n15375), .ZN(n15378) );
  AOI21_X1 U17536 ( .B1(n15380), .B2(n15379), .A(n15378), .ZN(n15387) );
  XOR2_X1 U17537 ( .A(NA), .B(keyinput_162), .Z(n15386) );
  XOR2_X1 U17538 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_166), .Z(n15384) );
  XOR2_X1 U17539 ( .A(BS16), .B(keyinput_163), .Z(n15383) );
  XOR2_X1 U17540 ( .A(READY2), .B(keyinput_165), .Z(n15382) );
  XNOR2_X1 U17541 ( .A(READY1), .B(keyinput_164), .ZN(n15381) );
  NOR4_X1 U17542 ( .A1(n15384), .A2(n15383), .A3(n15382), .A4(n15381), .ZN(
        n15385) );
  OAI21_X1 U17543 ( .B1(n15387), .B2(n15386), .A(n15385), .ZN(n15390) );
  XNOR2_X1 U17544 ( .A(n17730), .B(keyinput_167), .ZN(n15389) );
  XNOR2_X1 U17545 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_168), .ZN(n15388) );
  AOI21_X1 U17546 ( .B1(n15390), .B2(n15389), .A(n15388), .ZN(n15395) );
  XNOR2_X1 U17547 ( .A(n15391), .B(keyinput_169), .ZN(n15394) );
  XNOR2_X1 U17548 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_171), .ZN(
        n15393) );
  XNOR2_X1 U17549 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_170), .ZN(n15392) );
  OAI211_X1 U17550 ( .C1(n15395), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15403) );
  XNOR2_X1 U17551 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(keyinput_172), .ZN(n15402) );
  INV_X1 U17552 ( .A(keyinput_176), .ZN(n15396) );
  XNOR2_X1 U17553 ( .A(n15396), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n15400)
         );
  XNOR2_X1 U17554 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_173), .ZN(n15399) );
  XNOR2_X1 U17555 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_175), .ZN(n15398) );
  XNOR2_X1 U17556 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_174), .ZN(n15397) );
  NAND4_X1 U17557 ( .A1(n15400), .A2(n15399), .A3(n15398), .A4(n15397), .ZN(
        n15401) );
  AOI21_X1 U17558 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(n15405) );
  XNOR2_X1 U17559 ( .A(n20535), .B(keyinput_177), .ZN(n15404) );
  NOR2_X1 U17560 ( .A1(n15405), .A2(n15404), .ZN(n15409) );
  XNOR2_X1 U17561 ( .A(n16284), .B(keyinput_180), .ZN(n15408) );
  XNOR2_X1 U17562 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_179), .ZN(
        n15407) );
  XNOR2_X1 U17563 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_178), .ZN(
        n15406) );
  NOR4_X1 U17564 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15412) );
  XNOR2_X1 U17565 ( .A(n16480), .B(keyinput_182), .ZN(n15411) );
  XOR2_X1 U17566 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .Z(n15410)
         );
  NOR3_X1 U17567 ( .A1(n15412), .A2(n15411), .A3(n15410), .ZN(n15418) );
  XNOR2_X1 U17568 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .ZN(n15414)
         );
  XNOR2_X1 U17569 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .ZN(n15413)
         );
  NAND2_X1 U17570 ( .A1(n15414), .A2(n15413), .ZN(n15417) );
  XNOR2_X1 U17571 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .ZN(n15416)
         );
  XNOR2_X1 U17572 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .ZN(n15415)
         );
  NOR4_X1 U17573 ( .A1(n15418), .A2(n15417), .A3(n15416), .A4(n15415), .ZN(
        n15428) );
  XNOR2_X1 U17574 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .ZN(n15427)
         );
  XNOR2_X1 U17575 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n15420)
         );
  XNOR2_X1 U17576 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .ZN(n15419)
         );
  NAND2_X1 U17577 ( .A1(n15420), .A2(n15419), .ZN(n15426) );
  XOR2_X1 U17578 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_193), .Z(n15424)
         );
  INV_X1 U17579 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n16702) );
  XNOR2_X1 U17580 ( .A(n16702), .B(keyinput_191), .ZN(n15423) );
  XNOR2_X1 U17581 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .ZN(n15422)
         );
  XNOR2_X1 U17582 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .ZN(n15421)
         );
  NAND4_X1 U17583 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15425) );
  NOR4_X1 U17584 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15432) );
  INV_X1 U17585 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15941) );
  XNOR2_X1 U17586 ( .A(n15941), .B(keyinput_195), .ZN(n15431) );
  XNOR2_X1 U17587 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_196), .ZN(n15430)
         );
  XNOR2_X1 U17588 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n15429)
         );
  NOR4_X1 U17589 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15438) );
  XOR2_X1 U17590 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .Z(n15437)
         );
  XOR2_X1 U17591 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_199), .Z(n15435)
         );
  XNOR2_X1 U17592 ( .A(n20589), .B(keyinput_200), .ZN(n15434) );
  XNOR2_X1 U17593 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_198), .ZN(n15433)
         );
  NOR3_X1 U17594 ( .A1(n15435), .A2(n15434), .A3(n15433), .ZN(n15436) );
  OAI21_X1 U17595 ( .B1(n15438), .B2(n15437), .A(n15436), .ZN(n15441) );
  XNOR2_X1 U17596 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .ZN(n15440)
         );
  XOR2_X1 U17597 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .Z(n15439) );
  AOI21_X1 U17598 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(n15444) );
  XOR2_X1 U17599 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_204), .Z(n15443) );
  XNOR2_X1 U17600 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .ZN(n15442)
         );
  NOR3_X1 U17601 ( .A1(n15444), .A2(n15443), .A3(n15442), .ZN(n15447) );
  XNOR2_X1 U17602 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .ZN(n15446)
         );
  XNOR2_X1 U17603 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_206), .ZN(n15445)
         );
  OAI21_X1 U17604 ( .B1(n15447), .B2(n15446), .A(n15445), .ZN(n15454) );
  XNOR2_X1 U17605 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .ZN(n15453)
         );
  XOR2_X1 U17606 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .Z(n15451) );
  XNOR2_X1 U17607 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .ZN(n15450)
         );
  XNOR2_X1 U17608 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .ZN(n15449)
         );
  XNOR2_X1 U17609 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .ZN(n15448)
         );
  NAND4_X1 U17610 ( .A1(n15451), .A2(n15450), .A3(n15449), .A4(n15448), .ZN(
        n15452) );
  AOI21_X1 U17611 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15457) );
  XNOR2_X1 U17612 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .ZN(n15456)
         );
  XOR2_X1 U17613 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .Z(n15455) );
  OAI21_X1 U17614 ( .B1(n15457), .B2(n15456), .A(n15455), .ZN(n15460) );
  XOR2_X1 U17615 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_214), .Z(n15459) );
  XNOR2_X1 U17616 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_215), .ZN(n15458)
         );
  NAND3_X1 U17617 ( .A1(n15460), .A2(n15459), .A3(n15458), .ZN(n15463) );
  XOR2_X1 U17618 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .Z(n15462) );
  XOR2_X1 U17619 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_217), .Z(n15461) );
  AOI21_X1 U17620 ( .B1(n15463), .B2(n15462), .A(n15461), .ZN(n15467) );
  XOR2_X1 U17621 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .Z(n15466) );
  XNOR2_X1 U17622 ( .A(n22190), .B(keyinput_219), .ZN(n15465) );
  XNOR2_X1 U17623 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_220), .ZN(n15464)
         );
  NOR4_X1 U17624 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15471) );
  XOR2_X1 U17625 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_221), .Z(n15470) );
  XOR2_X1 U17626 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_223), .Z(n15469) );
  XOR2_X1 U17627 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_222), .Z(n15468) );
  OAI211_X1 U17628 ( .C1(n15471), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15474) );
  XNOR2_X1 U17629 ( .A(n22127), .B(keyinput_225), .ZN(n15473) );
  XNOR2_X1 U17630 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .ZN(n15472)
         );
  NAND3_X1 U17631 ( .A1(n15474), .A2(n15473), .A3(n15472), .ZN(n15477) );
  XOR2_X1 U17632 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .Z(n15476) );
  XOR2_X1 U17633 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_227), .Z(n15475) );
  NAND3_X1 U17634 ( .A1(n15477), .A2(n15476), .A3(n15475), .ZN(n15480) );
  XNOR2_X1 U17635 ( .A(n15801), .B(keyinput_228), .ZN(n15479) );
  XNOR2_X1 U17636 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n15478)
         );
  NAND3_X1 U17637 ( .A1(n15480), .A2(n15479), .A3(n15478), .ZN(n15483) );
  XNOR2_X1 U17638 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .ZN(n15482)
         );
  XNOR2_X1 U17639 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n15481)
         );
  NAND3_X1 U17640 ( .A1(n15483), .A2(n15482), .A3(n15481), .ZN(n15487) );
  XOR2_X1 U17641 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .Z(n15486) );
  XNOR2_X1 U17642 ( .A(n15484), .B(keyinput_233), .ZN(n15485) );
  NAND3_X1 U17643 ( .A1(n15487), .A2(n15486), .A3(n15485), .ZN(n15490) );
  XOR2_X1 U17644 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .Z(n15489) );
  XNOR2_X1 U17645 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .ZN(n15488)
         );
  AOI21_X1 U17646 ( .B1(n15490), .B2(n15489), .A(n15488), .ZN(n15497) );
  XOR2_X1 U17647 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .Z(n15496) );
  XOR2_X1 U17648 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .Z(n15495) );
  XNOR2_X1 U17649 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n15493)
         );
  XNOR2_X1 U17650 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n15492)
         );
  XNOR2_X1 U17651 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_237), .ZN(n15491)
         );
  NAND3_X1 U17652 ( .A1(n15493), .A2(n15492), .A3(n15491), .ZN(n15494) );
  NOR4_X1 U17653 ( .A1(n15497), .A2(n15496), .A3(n15495), .A4(n15494), .ZN(
        n15506) );
  XNOR2_X1 U17654 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_241), .ZN(n15505)
         );
  XOR2_X1 U17655 ( .A(keyinput_242), .B(P1_EBX_REG_1__SCAN_IN), .Z(n15500) );
  XNOR2_X1 U17656 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .ZN(n15499)
         );
  XNOR2_X1 U17657 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n15498)
         );
  NAND3_X1 U17658 ( .A1(n15500), .A2(n15499), .A3(n15498), .ZN(n15503) );
  XNOR2_X1 U17659 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n15502)
         );
  XNOR2_X1 U17660 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .ZN(n15501)
         );
  NOR3_X1 U17661 ( .A1(n15503), .A2(n15502), .A3(n15501), .ZN(n15504) );
  OAI21_X1 U17662 ( .B1(n15506), .B2(n15505), .A(n15504), .ZN(n15509) );
  XNOR2_X1 U17663 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n15508)
         );
  XNOR2_X1 U17664 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .ZN(n15507)
         );
  AOI21_X1 U17665 ( .B1(n15509), .B2(n15508), .A(n15507), .ZN(n15513) );
  XOR2_X1 U17666 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .Z(n15512) );
  XNOR2_X1 U17667 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n15511)
         );
  XNOR2_X1 U17668 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .ZN(n15510)
         );
  NOR4_X1 U17669 ( .A1(n15513), .A2(n15512), .A3(n15511), .A4(n15510), .ZN(
        n15514) );
  AOI211_X1 U17670 ( .C1(n15517), .C2(n15516), .A(n15515), .B(n15514), .ZN(
        n15630) );
  OAI21_X1 U17671 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21852), .A(
        n15518), .ZN(n15533) );
  NOR2_X1 U17672 ( .A1(n15519), .A2(n15533), .ZN(n15521) );
  INV_X1 U17673 ( .A(n21839), .ZN(n18222) );
  XNOR2_X1 U17674 ( .A(n20710), .B(n19519), .ZN(n15523) );
  OAI21_X1 U17675 ( .B1(n15523), .B2(n20709), .A(n21875), .ZN(n21842) );
  NOR3_X1 U17676 ( .A1(n15544), .A2(n18222), .A3(n21842), .ZN(n15532) );
  INV_X1 U17677 ( .A(n15524), .ZN(n15529) );
  OAI211_X1 U17678 ( .C1(n21378), .C2(n14120), .A(n15545), .B(n15525), .ZN(
        n15526) );
  OAI21_X1 U17679 ( .B1(n15527), .B2(n15526), .A(n18224), .ZN(n15528) );
  OAI211_X1 U17680 ( .C1(n15531), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        n16118) );
  AOI211_X1 U17681 ( .C1(n21836), .C2(n16010), .A(n15532), .B(n16118), .ZN(
        n15539) );
  INV_X1 U17682 ( .A(n15533), .ZN(n15534) );
  AOI21_X1 U17683 ( .B1(n15535), .B2(n15534), .A(n18222), .ZN(n21840) );
  INV_X1 U17684 ( .A(n21840), .ZN(n18306) );
  NOR2_X1 U17685 ( .A1(n19560), .A2(n18306), .ZN(n15537) );
  OAI211_X1 U17686 ( .C1(n15537), .C2(n21836), .A(n15536), .B(n19519), .ZN(
        n15538) );
  INV_X1 U17687 ( .A(n21808), .ZN(n21801) );
  INV_X1 U17688 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20819) );
  NOR2_X1 U17689 ( .A1(n21808), .A2(n20819), .ZN(n18699) );
  NOR2_X1 U17690 ( .A1(n15541), .A2(n15540), .ZN(n21414) );
  NOR2_X1 U17691 ( .A1(n19560), .A2(n15545), .ZN(n21387) );
  NAND2_X1 U17692 ( .A1(n15543), .A2(n15542), .ZN(n20713) );
  NAND3_X1 U17693 ( .A1(n15545), .A2(n15544), .A3(n21390), .ZN(n16011) );
  INV_X1 U17694 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21471) );
  AOI22_X1 U17695 ( .A1(n14043), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U17696 ( .A1(n15574), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15548) );
  AOI22_X1 U17697 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18279), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15547) );
  AOI22_X1 U17698 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15546) );
  NAND4_X1 U17699 ( .A1(n15549), .A2(n15548), .A3(n15547), .A4(n15546), .ZN(
        n15555) );
  INV_X2 U17700 ( .A(n18063), .ZN(n18264) );
  AOI22_X1 U17701 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15590), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15553) );
  AOI22_X1 U17702 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15552) );
  AOI22_X1 U17703 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15563), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U17704 ( .A1(n14108), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15561), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15550) );
  NAND4_X1 U17705 ( .A1(n15553), .A2(n15552), .A3(n15551), .A4(n15550), .ZN(
        n15554) );
  AOI22_X1 U17706 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18254), .ZN(n15560) );
  AOI22_X1 U17707 ( .A1(n14108), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18076), .ZN(n15559) );
  AOI22_X1 U17708 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18199), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n18247), .ZN(n15558) );
  AOI22_X1 U17709 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18279), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15556), .ZN(n15557) );
  NAND4_X1 U17710 ( .A1(n15560), .A2(n15559), .A3(n15558), .A4(n15557), .ZN(
        n15569) );
  AOI22_X1 U17711 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U17712 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n14043), .B1(
        n15590), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U17713 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n15562), .B1(
        n15561), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15565) );
  AOI22_X1 U17714 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n15574), .B1(
        n15563), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15564) );
  NAND4_X1 U17715 ( .A1(n15567), .A2(n15566), .A3(n15565), .A4(n15564), .ZN(
        n15568) );
  OR2_X2 U17716 ( .A1(n15569), .A2(n15568), .ZN(n15581) );
  OR2_X1 U17717 ( .A1(n21471), .A2(n15583), .ZN(n15584) );
  AOI22_X1 U17718 ( .A1(n14108), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U17719 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U17720 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U17721 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15570) );
  NAND4_X1 U17722 ( .A1(n15573), .A2(n15572), .A3(n15571), .A4(n15570), .ZN(
        n15580) );
  AOI22_X1 U17723 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15574), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U17724 ( .A1(n14043), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U17725 ( .A1(n18245), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U17726 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15590), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15575) );
  NAND4_X1 U17727 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        n15579) );
  NOR2_X1 U17728 ( .A1(n15580), .A2(n15579), .ZN(n15620) );
  INV_X1 U17729 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21522) );
  NOR2_X1 U17730 ( .A1(n15620), .A2(n21522), .ZN(n18740) );
  INV_X1 U17731 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21462) );
  INV_X2 U17732 ( .A(n15581), .ZN(n15622) );
  XNOR2_X2 U17733 ( .A(n21462), .B(n15622), .ZN(n18733) );
  NAND2_X1 U17734 ( .A1(n18740), .A2(n18733), .ZN(n18730) );
  NAND2_X1 U17735 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15622), .ZN(
        n15582) );
  NAND2_X1 U17736 ( .A1(n18730), .A2(n15582), .ZN(n18721) );
  NAND2_X1 U17737 ( .A1(n18721), .A2(n18722), .ZN(n18720) );
  NAND2_X1 U17738 ( .A1(n15584), .A2(n18720), .ZN(n15585) );
  NAND2_X1 U17739 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15585), .ZN(
        n15597) );
  INV_X1 U17740 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21481) );
  XNOR2_X1 U17741 ( .A(n21481), .B(n15585), .ZN(n18715) );
  AOI22_X1 U17742 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U17743 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U17744 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U17745 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15586) );
  NAND4_X1 U17746 ( .A1(n15589), .A2(n15588), .A3(n15587), .A4(n15586), .ZN(
        n15596) );
  AOI22_X1 U17747 ( .A1(n14043), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U17748 ( .A1(n14108), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15593) );
  AOI22_X1 U17749 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U17750 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15590), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15591) );
  NAND4_X1 U17751 ( .A1(n15594), .A2(n15593), .A3(n15592), .A4(n15591), .ZN(
        n15595) );
  XOR2_X1 U17752 ( .A(n21237), .B(n15618), .Z(n18714) );
  NAND2_X1 U17753 ( .A1(n18715), .A2(n18714), .ZN(n18713) );
  NAND2_X1 U17754 ( .A1(n15597), .A2(n18713), .ZN(n18311) );
  AOI22_X1 U17755 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U17756 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U17757 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U17758 ( .A1(n15556), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15598) );
  NAND4_X1 U17759 ( .A1(n15601), .A2(n15600), .A3(n15599), .A4(n15598), .ZN(
        n15607) );
  AOI22_X1 U17760 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U17761 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U17762 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U17763 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15602) );
  NAND4_X1 U17764 ( .A1(n15605), .A2(n15604), .A3(n15603), .A4(n15602), .ZN(
        n15606) );
  XOR2_X1 U17765 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18309), .Z(
        n18310) );
  XOR2_X1 U17766 ( .A(n18311), .B(n18310), .Z(n18705) );
  INV_X1 U17767 ( .A(n21727), .ZN(n21783) );
  NOR2_X1 U17768 ( .A1(n21471), .A2(n21462), .ZN(n21427) );
  INV_X1 U17769 ( .A(n21427), .ZN(n15611) );
  INV_X1 U17770 ( .A(n15608), .ZN(n15612) );
  OAI21_X1 U17771 ( .B1(n15612), .B2(n15609), .A(n21410), .ZN(n21818) );
  NAND2_X1 U17772 ( .A1(n21818), .A2(n21522), .ZN(n21600) );
  INV_X1 U17773 ( .A(n21600), .ZN(n21763) );
  OAI21_X1 U17774 ( .B1(n21522), .B2(n21462), .A(n21471), .ZN(n21430) );
  OR2_X1 U17775 ( .A1(n21756), .A2(n21430), .ZN(n21460) );
  NAND2_X1 U17776 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21460), .ZN(
        n15610) );
  AOI211_X1 U17777 ( .C1(n21816), .C2(n15611), .A(n21763), .B(n15610), .ZN(
        n21474) );
  INV_X1 U17778 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21480) );
  NOR3_X1 U17779 ( .A1(n21783), .A2(n21474), .A3(n21480), .ZN(n15614) );
  NOR2_X1 U17780 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21805), .ZN(
        n21450) );
  NOR2_X1 U17781 ( .A1(n21764), .A2(n21450), .ZN(n21654) );
  AOI22_X1 U17782 ( .A1(n21835), .A2(n21430), .B1(n21427), .B2(n21654), .ZN(
        n21496) );
  NOR3_X1 U17783 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21496), .A3(
        n21481), .ZN(n15613) );
  AOI211_X1 U17784 ( .C1(n21483), .C2(n18705), .A(n15614), .B(n15613), .ZN(
        n15627) );
  NOR2_X1 U17785 ( .A1(n15622), .A2(n15620), .ZN(n15621) );
  NOR2_X1 U17786 ( .A1(n15615), .A2(n15621), .ZN(n15625) );
  INV_X1 U17787 ( .A(n15625), .ZN(n15617) );
  XNOR2_X1 U17788 ( .A(n21237), .B(n15617), .ZN(n15616) );
  NAND2_X1 U17789 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15616), .ZN(
        n15624) );
  XOR2_X1 U17790 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15616), .Z(
        n18710) );
  OAI21_X1 U17791 ( .B1(n15620), .B2(n15618), .A(n15617), .ZN(n15619) );
  NAND2_X1 U17792 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15619), .ZN(
        n15623) );
  XNOR2_X1 U17793 ( .A(n21471), .B(n15619), .ZN(n18725) );
  INV_X1 U17794 ( .A(n15620), .ZN(n21371) );
  NOR2_X1 U17795 ( .A1(n21371), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18741) );
  INV_X1 U17796 ( .A(n18741), .ZN(n18732) );
  NOR2_X1 U17797 ( .A1(n18733), .A2(n18732), .ZN(n18731) );
  AOI211_X1 U17798 ( .C1(n15622), .C2(n21462), .A(n18731), .B(n15621), .ZN(
        n18724) );
  NAND2_X1 U17799 ( .A1(n18725), .A2(n18724), .ZN(n18723) );
  NAND2_X1 U17800 ( .A1(n15623), .A2(n18723), .ZN(n18709) );
  NAND2_X1 U17801 ( .A1(n18710), .A2(n18709), .ZN(n18708) );
  NAND2_X1 U17802 ( .A1(n15624), .A2(n18708), .ZN(n18287) );
  XNOR2_X1 U17803 ( .A(n21480), .B(n18287), .ZN(n18286) );
  NOR2_X1 U17804 ( .A1(n21237), .A2(n15625), .ZN(n18290) );
  XOR2_X1 U17805 ( .A(n18290), .B(n18314), .Z(n18285) );
  XOR2_X1 U17806 ( .A(n18286), .B(n18285), .Z(n18701) );
  NAND2_X1 U17807 ( .A1(n21834), .A2(n18701), .ZN(n15626) );
  AOI21_X1 U17808 ( .B1(n15627), .B2(n15626), .A(n21685), .ZN(n15628) );
  AOI211_X1 U17809 ( .C1(n21803), .C2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18699), .B(n15628), .ZN(n15629) );
  XNOR2_X1 U17810 ( .A(n15630), .B(n15629), .ZN(P3_U2858) );
  INV_X1 U17811 ( .A(n15685), .ZN(n15631) );
  AOI21_X1 U17812 ( .B1(n15633), .B2(n15632), .A(n15631), .ZN(n15649) );
  INV_X1 U17813 ( .A(n15649), .ZN(n15682) );
  MUX2_X1 U17814 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n15902), .Z(
        n22340) );
  AOI22_X1 U17815 ( .A1(n15903), .A2(n22340), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15728), .ZN(n15634) );
  OAI21_X1 U17816 ( .B1(n15682), .B2(n16621), .A(n15634), .ZN(P1_U2896) );
  NAND2_X1 U17817 ( .A1(n15649), .A2(n22197), .ZN(n15643) );
  INV_X1 U17818 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15639) );
  NAND3_X1 U17819 ( .A1(n22153), .A2(n15639), .A3(n15635), .ZN(n15636) );
  OAI211_X1 U17820 ( .C1(n22188), .C2(n15647), .A(n22122), .B(n15636), .ZN(
        n15637) );
  AOI21_X1 U17821 ( .B1(n22195), .B2(n15644), .A(n15637), .ZN(n15638) );
  INV_X1 U17822 ( .A(n15638), .ZN(n15641) );
  NOR3_X1 U17823 ( .A1(n22080), .A2(n22155), .A3(n15639), .ZN(n15640) );
  AOI211_X1 U17824 ( .C1(n11143), .C2(P1_EBX_REG_8__SCAN_IN), .A(n15641), .B(
        n15640), .ZN(n15642) );
  OAI211_X1 U17825 ( .C1(n15684), .C2(n22202), .A(n15643), .B(n15642), .ZN(
        P1_U2832) );
  NAND2_X1 U17826 ( .A1(n20623), .A2(n15644), .ZN(n15646) );
  OAI211_X1 U17827 ( .C1(n15997), .C2(n15647), .A(n15646), .B(n15645), .ZN(
        n15648) );
  AOI21_X1 U17828 ( .B1(n15649), .B2(n20628), .A(n15648), .ZN(n15650) );
  OAI21_X1 U17829 ( .B1(n15651), .B2(n22203), .A(n15650), .ZN(P1_U2991) );
  AND2_X1 U17830 ( .A1(n15653), .A2(n15652), .ZN(n15705) );
  NOR2_X1 U17831 ( .A1(n15655), .A2(n15654), .ZN(n15656) );
  INV_X1 U17832 ( .A(n15129), .ZN(n15661) );
  INV_X1 U17833 ( .A(n15658), .ZN(n15659) );
  OAI211_X1 U17834 ( .C1(n15661), .C2(n15660), .A(n15659), .B(n17136), .ZN(
        n15663) );
  NAND2_X1 U17835 ( .A1(n11163), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15662) );
  OAI211_X1 U17836 ( .C1(n18948), .C2(n11164), .A(n15663), .B(n15662), .ZN(
        P2_U2873) );
  XNOR2_X1 U17837 ( .A(n15665), .B(n15664), .ZN(n17734) );
  XNOR2_X1 U17838 ( .A(n15666), .B(n15668), .ZN(n17733) );
  INV_X1 U17839 ( .A(n17733), .ZN(n15680) );
  OAI21_X1 U17840 ( .B1(n15064), .B2(n15670), .A(n11146), .ZN(n20022) );
  AOI221_X1 U17841 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n15664), .C2(n15672), .A(
        n15671), .ZN(n15674) );
  NOR2_X1 U17842 ( .A1(n12980), .A2(n18958), .ZN(n15673) );
  AOI211_X1 U17843 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15675), .A(
        n15674), .B(n15673), .ZN(n15678) );
  INV_X1 U17844 ( .A(n15676), .ZN(n17736) );
  NAND2_X1 U17845 ( .A1(n17736), .A2(n19159), .ZN(n15677) );
  OAI211_X1 U17846 ( .C1(n20022), .C2(n19134), .A(n15678), .B(n15677), .ZN(
        n15679) );
  AOI21_X1 U17847 ( .B1(n15680), .B2(n19160), .A(n15679), .ZN(n15681) );
  OAI21_X1 U17848 ( .B1(n19153), .B2(n17734), .A(n15681), .ZN(P2_U3041) );
  INV_X1 U17849 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15683) );
  OAI222_X1 U17850 ( .A1(n15684), .A2(n20551), .B1(n15683), .B2(n20556), .C1(
        n15682), .C2(n16572), .ZN(P1_U2864) );
  XOR2_X1 U17851 ( .A(n15686), .B(n15685), .Z(n22085) );
  INV_X1 U17852 ( .A(n22085), .ZN(n15715) );
  MUX2_X1 U17853 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n15902), .Z(
        n22347) );
  AOI22_X1 U17854 ( .A1(n15903), .A2(n22347), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15728), .ZN(n15687) );
  OAI21_X1 U17855 ( .B1(n15715), .B2(n16621), .A(n15687), .ZN(P1_U2895) );
  OAI21_X1 U17856 ( .B1(n15689), .B2(n15688), .A(n11158), .ZN(n21971) );
  NOR2_X1 U17857 ( .A1(n22016), .A2(n15690), .ZN(n21973) );
  AND2_X1 U17858 ( .A1(n20627), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15691) );
  AOI211_X1 U17859 ( .C1(n20623), .C2(n22084), .A(n21973), .B(n15691), .ZN(
        n15693) );
  NAND2_X1 U17860 ( .A1(n22085), .A2(n20628), .ZN(n15692) );
  OAI211_X1 U17861 ( .C1(n21971), .C2(n22203), .A(n15693), .B(n15692), .ZN(
        P1_U2990) );
  OAI21_X1 U17862 ( .B1(n15101), .B2(n15695), .A(n15694), .ZN(n15857) );
  XNOR2_X1 U17863 ( .A(n15857), .B(n15856), .ZN(n20598) );
  MUX2_X1 U17864 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n15902), .Z(
        n16585) );
  INV_X1 U17865 ( .A(n16585), .ZN(n22359) );
  OAI222_X1 U17866 ( .A1(n20598), .A2(n16621), .B1(n15819), .B2(n22359), .C1(
        n15696), .C2(n16612), .ZN(P1_U2893) );
  NOR2_X1 U17867 ( .A1(n15699), .A2(n15698), .ZN(n15700) );
  OR2_X1 U17868 ( .A1(n15697), .A2(n15700), .ZN(n21997) );
  INV_X1 U17869 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15701) );
  OAI222_X1 U17870 ( .A1(n20598), .A2(n16572), .B1(n20551), .B2(n21997), .C1(
        n15701), .C2(n20556), .ZN(P1_U2861) );
  INV_X1 U17871 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n15712) );
  INV_X1 U17872 ( .A(n15808), .ZN(n15702) );
  OAI211_X1 U17873 ( .C1(n15658), .C2(n15703), .A(n15702), .B(n17136), .ZN(
        n15711) );
  INV_X1 U17874 ( .A(n15705), .ZN(n15708) );
  INV_X1 U17875 ( .A(n15706), .ZN(n15707) );
  NAND2_X1 U17876 ( .A1(n15708), .A2(n15707), .ZN(n15709) );
  AND2_X1 U17877 ( .A1(n15704), .A2(n15709), .ZN(n18956) );
  NAND2_X1 U17878 ( .A1(n18956), .A2(n17125), .ZN(n15710) );
  OAI211_X1 U17879 ( .C1(n17125), .C2(n15712), .A(n15711), .B(n15710), .ZN(
        P2_U2872) );
  INV_X1 U17880 ( .A(n15713), .ZN(n15714) );
  XNOR2_X1 U17881 ( .A(n15093), .B(n15714), .ZN(n21974) );
  INV_X1 U17882 ( .A(n21974), .ZN(n22082) );
  INV_X1 U17883 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n22081) );
  OAI222_X1 U17884 ( .A1(n22082), .A2(n20551), .B1(n20556), .B2(n22081), .C1(
        n16572), .C2(n15715), .ZN(P1_U2863) );
  OAI21_X1 U17885 ( .B1(n15808), .B2(n15807), .A(n17134), .ZN(n15738) );
  NAND2_X1 U17886 ( .A1(n15704), .A2(n15717), .ZN(n15718) );
  NAND2_X1 U17887 ( .A1(n15716), .A2(n15718), .ZN(n19131) );
  NOR2_X1 U17888 ( .A1(n19131), .A2(n11164), .ZN(n15719) );
  AOI21_X1 U17889 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n11164), .A(n15719), .ZN(
        n15720) );
  OAI21_X1 U17890 ( .B1(n15738), .B2(n17128), .A(n15720), .ZN(P2_U2871) );
  NAND2_X1 U17891 ( .A1(n15790), .A2(n15722), .ZN(n15741) );
  AND2_X1 U17892 ( .A1(n15790), .A2(n15723), .ZN(n15794) );
  OR2_X1 U17893 ( .A1(n15794), .A2(n15724), .ZN(n15725) );
  NAND2_X1 U17894 ( .A1(n15741), .A2(n15725), .ZN(n22115) );
  INV_X1 U17895 ( .A(n16614), .ZN(n16381) );
  AOI22_X1 U17896 ( .A1(n16381), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15728), .ZN(n15731) );
  NOR3_X2 U17897 ( .A1(n15728), .A2(n15727), .A3(n15726), .ZN(n16618) );
  INV_X1 U17898 ( .A(n22300), .ZN(n15729) );
  AOI22_X1 U17899 ( .A1(n16618), .A2(n15729), .B1(n16616), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15730) );
  OAI211_X1 U17900 ( .C1(n22115), .C2(n16621), .A(n15731), .B(n15730), .ZN(
        P1_U2888) );
  XNOR2_X1 U17901 ( .A(n15733), .B(n15732), .ZN(n19133) );
  INV_X1 U17902 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n17885) );
  OAI22_X1 U17903 ( .A1(n20172), .A2(n19133), .B1(n20066), .B2(n17885), .ZN(
        n15734) );
  AOI21_X1 U17904 ( .B1(n20168), .B2(n15735), .A(n15734), .ZN(n15737) );
  AOI22_X1 U17905 ( .A1(n20169), .A2(BUF1_REG_16__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n15736) );
  OAI211_X1 U17906 ( .C1(n15738), .C2(n20222), .A(n15737), .B(n15736), .ZN(
        P2_U2903) );
  NAND2_X1 U17907 ( .A1(n15741), .A2(n15740), .ZN(n15742) );
  AND2_X1 U17908 ( .A1(n15739), .A2(n15742), .ZN(n20624) );
  INV_X1 U17909 ( .A(n20624), .ZN(n15760) );
  INV_X1 U17910 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15743) );
  OAI22_X1 U17911 ( .A1(n16614), .A2(n15744), .B1(n15743), .B2(n16612), .ZN(
        n15746) );
  INV_X1 U17912 ( .A(n16618), .ZN(n15966) );
  NOR2_X1 U17913 ( .A1(n15966), .A2(n22305), .ZN(n15745) );
  AOI211_X1 U17914 ( .C1(n16616), .C2(BUF1_REG_17__SCAN_IN), .A(n15746), .B(
        n15745), .ZN(n15747) );
  OAI21_X1 U17915 ( .B1(n15760), .B2(n16621), .A(n15747), .ZN(P1_U2887) );
  INV_X1 U17916 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20493) );
  INV_X1 U17917 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20491) );
  INV_X1 U17918 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22094) );
  NAND2_X1 U17919 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15748), .ZN(n22091) );
  NOR2_X1 U17920 ( .A1(n22094), .A2(n22091), .ZN(n22090) );
  NAND2_X1 U17921 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n22090), .ZN(n16270) );
  NOR2_X1 U17922 ( .A1(n22138), .A2(n16270), .ZN(n22103) );
  NAND2_X1 U17923 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n22103), .ZN(n15803) );
  NOR2_X1 U17924 ( .A1(n20491), .A2(n15803), .ZN(n22120) );
  NAND2_X1 U17925 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22120), .ZN(n22118) );
  NOR2_X1 U17926 ( .A1(n20493), .A2(n22118), .ZN(n22125) );
  OR2_X1 U17927 ( .A1(n22125), .A2(n22155), .ZN(n22130) );
  INV_X1 U17928 ( .A(n22130), .ZN(n22147) );
  NAND2_X1 U17929 ( .A1(n20493), .A2(n22118), .ZN(n15758) );
  INV_X1 U17930 ( .A(n15749), .ZN(n15864) );
  NAND2_X1 U17931 ( .A1(n15750), .A2(n15751), .ZN(n15752) );
  NAND2_X1 U17932 ( .A1(n15864), .A2(n15752), .ZN(n22027) );
  OAI21_X1 U17933 ( .B1(n22188), .B2(n15753), .A(n22122), .ZN(n15755) );
  INV_X1 U17934 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20543) );
  NOR2_X1 U17935 ( .A1(n22191), .A2(n20543), .ZN(n15754) );
  AOI211_X1 U17936 ( .C1(n20622), .C2(n22195), .A(n15755), .B(n15754), .ZN(
        n15756) );
  OAI21_X1 U17937 ( .B1(n22027), .B2(n22202), .A(n15756), .ZN(n15757) );
  AOI21_X1 U17938 ( .B1(n22147), .B2(n15758), .A(n15757), .ZN(n15759) );
  OAI21_X1 U17939 ( .B1(n15760), .B2(n22181), .A(n15759), .ZN(P1_U2823) );
  XNOR2_X1 U17940 ( .A(n15761), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15784) );
  XOR2_X1 U17941 ( .A(n15762), .B(n15764), .Z(n15782) );
  OAI22_X1 U17942 ( .A1(n15765), .A2(n17789), .B1(n12984), .B2(n18958), .ZN(
        n15766) );
  AOI21_X1 U17943 ( .B1(n17777), .B2(n18880), .A(n15766), .ZN(n15767) );
  OAI21_X1 U17944 ( .B1(n18881), .B2(n13199), .A(n15767), .ZN(n15768) );
  AOI21_X1 U17945 ( .B1(n15782), .B2(n17818), .A(n15768), .ZN(n15769) );
  OAI21_X1 U17946 ( .B1(n15784), .B2(n17779), .A(n15769), .ZN(P2_U3008) );
  NAND3_X1 U17947 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15770) );
  NOR2_X1 U17948 ( .A1(n15771), .A2(n15770), .ZN(n15775) );
  OAI21_X1 U17949 ( .B1(n17497), .B2(n15773), .A(n15772), .ZN(n19155) );
  NOR2_X1 U17950 ( .A1(n12984), .A2(n18958), .ZN(n15774) );
  AOI221_X1 U17951 ( .B1(n15775), .B2(n13089), .C1(n19155), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n15774), .ZN(n15776) );
  INV_X1 U17952 ( .A(n15776), .ZN(n15781) );
  NAND2_X1 U17953 ( .A1(n11146), .A2(n15777), .ZN(n15779) );
  XNOR2_X1 U17954 ( .A(n15779), .B(n15778), .ZN(n19969) );
  OAI22_X1 U17955 ( .A1(n19969), .A2(n19134), .B1(n19130), .B2(n18881), .ZN(
        n15780) );
  AOI211_X1 U17956 ( .C1(n15782), .C2(n19160), .A(n15781), .B(n15780), .ZN(
        n15783) );
  OAI21_X1 U17957 ( .B1(n15784), .B2(n19153), .A(n15783), .ZN(P2_U3040) );
  OR2_X1 U17958 ( .A1(n15798), .A2(n15785), .ZN(n15786) );
  AND2_X1 U17959 ( .A1(n15750), .A2(n15786), .ZN(n15942) );
  INV_X1 U17960 ( .A(n15942), .ZN(n22114) );
  INV_X1 U17961 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15787) );
  OAI222_X1 U17962 ( .A1(n22114), .A2(n20551), .B1(n15787), .B2(n20556), .C1(
        n22115), .C2(n16572), .ZN(P1_U2856) );
  NAND2_X1 U17963 ( .A1(n15790), .A2(n15788), .ZN(n15891) );
  NAND2_X1 U17964 ( .A1(n15790), .A2(n15789), .ZN(n15795) );
  INV_X1 U17965 ( .A(n15795), .ZN(n15791) );
  AOI21_X1 U17966 ( .B1(n15792), .B2(n15891), .A(n15791), .ZN(n22110) );
  INV_X1 U17967 ( .A(n22110), .ZN(n15890) );
  MUX2_X1 U17968 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n15902), .Z(
        n22379) );
  AOI22_X1 U17969 ( .A1(n15903), .A2(n22379), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15728), .ZN(n15793) );
  OAI21_X1 U17970 ( .B1(n15890), .B2(n16621), .A(n15793), .ZN(P1_U2890) );
  AOI21_X1 U17971 ( .B1(n15796), .B2(n15795), .A(n15794), .ZN(n20611) );
  INV_X1 U17972 ( .A(n20611), .ZN(n15820) );
  INV_X1 U17973 ( .A(n15797), .ZN(n15799) );
  AOI21_X1 U17974 ( .B1(n15799), .B2(n11875), .A(n15798), .ZN(n22008) );
  OAI22_X1 U17975 ( .A1(n22191), .A2(n15801), .B1(n22186), .B2(n15800), .ZN(
        n15805) );
  NAND2_X1 U17976 ( .A1(n22119), .A2(n15803), .ZN(n22105) );
  AOI21_X1 U17977 ( .B1(n22151), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n22139), .ZN(n15802) );
  OAI221_X1 U17978 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15803), .C1(n20491), 
        .C2(n22105), .A(n15802), .ZN(n15804) );
  AOI211_X1 U17979 ( .C1(n22008), .C2(n16557), .A(n15805), .B(n15804), .ZN(
        n15806) );
  OAI21_X1 U17980 ( .B1(n15820), .B2(n22181), .A(n15806), .ZN(P1_U2825) );
  AND2_X1 U17981 ( .A1(n15808), .A2(n15807), .ZN(n15810) );
  AND2_X1 U17982 ( .A1(n15810), .A2(n15809), .ZN(n15912) );
  OAI21_X1 U17983 ( .B1(n15912), .B2(n15812), .A(n15811), .ZN(n17177) );
  NAND2_X1 U17984 ( .A1(n11164), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15816) );
  OR2_X1 U17985 ( .A1(n15915), .A2(n15813), .ZN(n15814) );
  AND2_X1 U17986 ( .A1(n15814), .A2(n16935), .ZN(n19027) );
  NAND2_X1 U17987 ( .A1(n19027), .A2(n17125), .ZN(n15815) );
  OAI211_X1 U17988 ( .C1(n17177), .C2(n17128), .A(n15816), .B(n15815), .ZN(
        P2_U2865) );
  OAI222_X1 U17989 ( .A1(n15820), .A2(n16621), .B1(n15819), .B2(n15818), .C1(
        n15817), .C2(n20474), .ZN(P1_U2889) );
  AND2_X1 U17990 ( .A1(n15739), .A2(n15821), .ZN(n15823) );
  OR2_X1 U17991 ( .A1(n15823), .A2(n15822), .ZN(n22132) );
  AOI22_X1 U17992 ( .A1(n16381), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15728), .ZN(n15826) );
  INV_X1 U17993 ( .A(n22309), .ZN(n15824) );
  AOI22_X1 U17994 ( .A1(n16618), .A2(n15824), .B1(n16616), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15825) );
  OAI211_X1 U17995 ( .C1(n22132), .C2(n16621), .A(n15826), .B(n15825), .ZN(
        P1_U2886) );
  INV_X1 U17996 ( .A(n20590), .ZN(n15828) );
  OAI21_X1 U17997 ( .B1(n15829), .B2(n20593), .A(n15828), .ZN(n20618) );
  INV_X1 U17998 ( .A(n15830), .ZN(n15831) );
  AOI21_X1 U17999 ( .B1(n20618), .B2(n15832), .A(n15831), .ZN(n15834) );
  MUX2_X1 U18000 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n11870), .S(
        n20593), .Z(n15833) );
  XNOR2_X1 U18001 ( .A(n15834), .B(n15833), .ZN(n15855) );
  AOI22_X1 U18002 ( .A1(n20627), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n22040), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15835) );
  OAI21_X1 U18003 ( .B1(n20633), .B2(n22108), .A(n15835), .ZN(n15836) );
  AOI21_X1 U18004 ( .B1(n22110), .B2(n20628), .A(n15836), .ZN(n15837) );
  OAI21_X1 U18005 ( .B1(n15855), .B2(n22203), .A(n15837), .ZN(P1_U2985) );
  NOR2_X1 U18006 ( .A1(n21980), .A2(n15838), .ZN(n21986) );
  INV_X1 U18007 ( .A(n15839), .ZN(n15840) );
  NOR2_X1 U18008 ( .A1(n15936), .A2(n15840), .ZN(n15841) );
  NOR3_X1 U18009 ( .A1(n21987), .A2(n21993), .A3(n22003), .ZN(n22012) );
  NAND3_X1 U18010 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n22012), .A3(
        n11870), .ZN(n15854) );
  INV_X1 U18011 ( .A(n11185), .ZN(n15894) );
  AND2_X1 U18012 ( .A1(n15894), .A2(n15843), .ZN(n15844) );
  OR2_X1 U18013 ( .A1(n15844), .A2(n11184), .ZN(n22113) );
  INV_X1 U18014 ( .A(n22113), .ZN(n15852) );
  INV_X1 U18015 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n16271) );
  NOR2_X1 U18016 ( .A1(n22016), .A2(n16271), .ZN(n15851) );
  AOI21_X1 U18017 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21916), .A(
        n15845), .ZN(n21915) );
  OAI22_X1 U18018 ( .A1(n15937), .A2(n15936), .B1(n15846), .B2(n21916), .ZN(
        n15847) );
  NOR3_X1 U18019 ( .A1(n21915), .A2(n21979), .A3(n15847), .ZN(n21922) );
  AND3_X1 U18020 ( .A1(n15848), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n21916), .ZN(n15849) );
  OAI211_X1 U18021 ( .C1(n21985), .C2(n15849), .A(n15937), .B(n21921), .ZN(
        n21912) );
  AOI21_X1 U18022 ( .B1(n21922), .B2(n21912), .A(n11870), .ZN(n15850) );
  AOI211_X1 U18023 ( .C1(n22037), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        n15853) );
  OAI211_X1 U18024 ( .C1(n15855), .C2(n22033), .A(n15854), .B(n15853), .ZN(
        P1_U3017) );
  OAI21_X1 U18025 ( .B1(n15857), .B2(n15856), .A(n15694), .ZN(n15859) );
  INV_X1 U18026 ( .A(n15859), .ZN(n15861) );
  INV_X1 U18027 ( .A(n15858), .ZN(n15860) );
  AOI21_X1 U18028 ( .B1(n15861), .B2(n15860), .A(n15893), .ZN(n22098) );
  INV_X1 U18029 ( .A(n22098), .ZN(n15909) );
  MUX2_X1 U18030 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n15902), .Z(
        n22365) );
  AOI22_X1 U18031 ( .A1(n15903), .A2(n22365), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15728), .ZN(n15862) );
  OAI21_X1 U18032 ( .B1(n15909), .B2(n16621), .A(n15862), .ZN(P1_U2892) );
  NAND2_X1 U18033 ( .A1(n15864), .A2(n15863), .ZN(n15865) );
  NAND2_X1 U18034 ( .A1(n15984), .A2(n15865), .ZN(n22136) );
  OAI222_X1 U18035 ( .A1(n22136), .A2(n20551), .B1(n22127), .B2(n20556), .C1(
        n22132), .C2(n16572), .ZN(P1_U2854) );
  MUX2_X1 U18036 ( .A(n11158), .B(n20590), .S(n11595), .Z(n15867) );
  INV_X1 U18037 ( .A(n15867), .ZN(n15868) );
  OAI21_X1 U18038 ( .B1(n15868), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20591), .ZN(n15889) );
  INV_X1 U18039 ( .A(n15869), .ZN(n15880) );
  NOR2_X1 U18040 ( .A1(n22016), .A2(n15870), .ZN(n15883) );
  NAND2_X1 U18041 ( .A1(n15872), .A2(n15871), .ZN(n21978) );
  XOR2_X1 U18042 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21977), .Z(
        n15878) );
  OAI21_X1 U18043 ( .B1(n21944), .B2(n15874), .A(n15873), .ZN(n15875) );
  AOI21_X1 U18044 ( .B1(n21985), .B2(n15876), .A(n15875), .ZN(n21976) );
  OAI22_X1 U18045 ( .A1(n21978), .A2(n15878), .B1(n15877), .B2(n21976), .ZN(
        n15879) );
  AOI211_X1 U18046 ( .C1(n22037), .C2(n15880), .A(n15883), .B(n15879), .ZN(
        n15881) );
  OAI21_X1 U18047 ( .B1(n15889), .B2(n22033), .A(n15881), .ZN(P1_U3021) );
  INV_X1 U18048 ( .A(n15882), .ZN(n15887) );
  AOI21_X1 U18049 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15883), .ZN(n15884) );
  OAI21_X1 U18050 ( .B1(n20633), .B2(n15885), .A(n15884), .ZN(n15886) );
  AOI21_X1 U18051 ( .B1(n15887), .B2(n20628), .A(n15886), .ZN(n15888) );
  OAI21_X1 U18052 ( .B1(n15889), .B2(n22203), .A(n15888), .ZN(P1_U2989) );
  OAI222_X1 U18053 ( .A1(n22113), .A2(n20551), .B1(n22104), .B2(n20556), .C1(
        n15890), .C2(n16572), .ZN(P1_U2858) );
  AOI21_X1 U18054 ( .B1(n15895), .B2(n15908), .A(n11185), .ZN(n21917) );
  INV_X1 U18055 ( .A(n15979), .ZN(n15897) );
  AOI22_X1 U18056 ( .A1(n11143), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n22151), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15896) );
  OAI21_X1 U18057 ( .B1(n22186), .B2(n15897), .A(n15896), .ZN(n15900) );
  OAI211_X1 U18058 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n22090), .A(n22153), 
        .B(n16270), .ZN(n15898) );
  OAI211_X1 U18059 ( .C1(n22095), .C2(n15977), .A(n22122), .B(n15898), .ZN(
        n15899) );
  AOI211_X1 U18060 ( .C1(n21917), .C2(n16557), .A(n15900), .B(n15899), .ZN(
        n15901) );
  OAI21_X1 U18061 ( .B1(n15982), .B2(n22181), .A(n15901), .ZN(P1_U2827) );
  MUX2_X1 U18062 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n15902), .Z(
        n22372) );
  AOI22_X1 U18063 ( .A1(n15903), .A2(n22372), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15728), .ZN(n15904) );
  OAI21_X1 U18064 ( .B1(n15982), .B2(n16621), .A(n15904), .ZN(P1_U2891) );
  AOI22_X1 U18065 ( .A1(n21917), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15905) );
  OAI21_X1 U18066 ( .B1(n15982), .B2(n16572), .A(n15905), .ZN(P1_U2859) );
  OR2_X1 U18067 ( .A1(n15697), .A2(n15906), .ZN(n15907) );
  NAND2_X1 U18068 ( .A1(n15908), .A2(n15907), .ZN(n22102) );
  INV_X1 U18069 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15910) );
  OAI222_X1 U18070 ( .A1(n22102), .A2(n20551), .B1(n15910), .B2(n20556), .C1(
        n15909), .C2(n16572), .ZN(P1_U2860) );
  NOR2_X1 U18071 ( .A1(n17134), .A2(n15911), .ZN(n17105) );
  INV_X1 U18072 ( .A(n15912), .ZN(n15913) );
  OAI21_X1 U18073 ( .B1(n17105), .B2(n15914), .A(n15913), .ZN(n17184) );
  INV_X1 U18074 ( .A(n15915), .ZN(n15916) );
  OAI21_X1 U18075 ( .B1(n14244), .B2(n15917), .A(n15916), .ZN(n19012) );
  NOR2_X1 U18076 ( .A1(n19012), .A2(n11163), .ZN(n15918) );
  AOI21_X1 U18077 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n11164), .A(n15918), .ZN(
        n15919) );
  OAI21_X1 U18078 ( .B1(n17184), .B2(n17128), .A(n15919), .ZN(P2_U2866) );
  OAI21_X1 U18079 ( .B1(n15921), .B2(n15924), .A(n15923), .ZN(n22159) );
  NOR2_X1 U18080 ( .A1(n16612), .A2(n22321), .ZN(n15927) );
  INV_X1 U18081 ( .A(n16616), .ZN(n15925) );
  OAI22_X1 U18082 ( .A1(n15966), .A2(n22319), .B1(n15925), .B2(n20682), .ZN(
        n15926) );
  AOI211_X1 U18083 ( .C1(DATAI_20_), .C2(n16381), .A(n15927), .B(n15926), .ZN(
        n15928) );
  OAI21_X1 U18084 ( .B1(n22159), .B2(n16621), .A(n15928), .ZN(P1_U2884) );
  AOI21_X1 U18085 ( .B1(n20590), .B2(n15930), .A(n15929), .ZN(n20608) );
  AND2_X1 U18086 ( .A1(n15931), .A2(n15932), .ZN(n20607) );
  NAND2_X1 U18087 ( .A1(n20608), .A2(n20607), .ZN(n20606) );
  NAND2_X1 U18088 ( .A1(n20606), .A2(n15932), .ZN(n15934) );
  XNOR2_X1 U18089 ( .A(n15934), .B(n15933), .ZN(n15957) );
  INV_X1 U18090 ( .A(n15957), .ZN(n15947) );
  NAND2_X1 U18091 ( .A1(n15938), .A2(n22012), .ZN(n22025) );
  NOR2_X1 U18092 ( .A1(n15935), .A2(n22025), .ZN(n15945) );
  AOI21_X1 U18093 ( .B1(n21916), .B2(n15938), .A(n21944), .ZN(n15940) );
  AOI21_X1 U18094 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15939) );
  NOR3_X1 U18095 ( .A1(n15940), .A2(n15939), .A3(n21979), .ZN(n22013) );
  NOR2_X1 U18096 ( .A1(n22016), .A2(n15941), .ZN(n15960) );
  AOI21_X1 U18097 ( .B1(n15942), .B2(n22037), .A(n15960), .ZN(n15943) );
  OAI21_X1 U18098 ( .B1(n22013), .B2(n20614), .A(n15943), .ZN(n15944) );
  AOI21_X1 U18099 ( .B1(n15945), .B2(n22026), .A(n15944), .ZN(n15946) );
  OAI21_X1 U18100 ( .B1(n15947), .B2(n22033), .A(n15946), .ZN(P1_U3015) );
  INV_X1 U18101 ( .A(n21997), .ZN(n15948) );
  AOI22_X1 U18102 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n22151), .B1(
        n16557), .B2(n15948), .ZN(n15949) );
  INV_X1 U18103 ( .A(n15949), .ZN(n15951) );
  OAI22_X1 U18104 ( .A1(n20595), .A2(n22186), .B1(n22181), .B2(n20598), .ZN(
        n15950) );
  NOR3_X1 U18105 ( .A1(n22139), .A2(n15951), .A3(n15950), .ZN(n15955) );
  NOR2_X1 U18106 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15952), .ZN(n15953) );
  AOI22_X1 U18107 ( .A1(n22153), .A2(n15953), .B1(n11143), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15954) );
  OAI211_X1 U18108 ( .C1(n15956), .C2(n20589), .A(n15955), .B(n15954), .ZN(
        P1_U2829) );
  NAND2_X1 U18109 ( .A1(n15957), .A2(n20629), .ZN(n15962) );
  INV_X1 U18110 ( .A(n22117), .ZN(n15958) );
  NOR2_X1 U18111 ( .A1(n15958), .A2(n20633), .ZN(n15959) );
  AOI211_X1 U18112 ( .C1(n20627), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15960), .B(n15959), .ZN(n15961) );
  OAI211_X1 U18113 ( .C1(n20599), .C2(n22115), .A(n15962), .B(n15961), .ZN(
        P1_U2983) );
  INV_X1 U18114 ( .A(n15963), .ZN(n15965) );
  INV_X1 U18115 ( .A(n15822), .ZN(n15964) );
  AOI21_X1 U18116 ( .B1(n15965), .B2(n15964), .A(n15921), .ZN(n22145) );
  INV_X1 U18117 ( .A(n22145), .ZN(n15987) );
  OAI22_X1 U18118 ( .A1(n16614), .A2(n14579), .B1(n22316), .B2(n16612), .ZN(
        n15968) );
  NOR2_X1 U18119 ( .A1(n15966), .A2(n22314), .ZN(n15967) );
  AOI211_X1 U18120 ( .C1(n16616), .C2(BUF1_REG_19__SCAN_IN), .A(n15968), .B(
        n15967), .ZN(n15969) );
  OAI21_X1 U18121 ( .B1(n15987), .B2(n16621), .A(n15969), .ZN(P1_U2885) );
  INV_X1 U18122 ( .A(n15970), .ZN(n15971) );
  AOI22_X1 U18123 ( .A1(n20590), .A2(n15972), .B1(n11595), .B2(n15971), .ZN(
        n20602) );
  INV_X1 U18124 ( .A(n15974), .ZN(n15973) );
  AOI21_X1 U18125 ( .B1(n11595), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15973), .ZN(n20601) );
  NAND2_X1 U18126 ( .A1(n20602), .A2(n20601), .ZN(n20600) );
  NAND2_X1 U18127 ( .A1(n20600), .A2(n15974), .ZN(n15975) );
  XOR2_X1 U18128 ( .A(n15976), .B(n15975), .Z(n21918) );
  NAND2_X1 U18129 ( .A1(n21918), .A2(n20629), .ZN(n15981) );
  OAI22_X1 U18130 ( .A1(n15997), .A2(n12226), .B1(n22016), .B2(n15977), .ZN(
        n15978) );
  AOI21_X1 U18131 ( .B1(n20623), .B2(n15979), .A(n15978), .ZN(n15980) );
  OAI211_X1 U18132 ( .C1(n20599), .C2(n15982), .A(n15981), .B(n15980), .ZN(
        P1_U2986) );
  INV_X1 U18133 ( .A(n15991), .ZN(n15986) );
  NAND2_X1 U18134 ( .A1(n15984), .A2(n15983), .ZN(n15985) );
  NAND2_X1 U18135 ( .A1(n15986), .A2(n15985), .ZN(n22150) );
  INV_X1 U18136 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15988) );
  OAI222_X1 U18137 ( .A1(n22150), .A2(n20551), .B1(n15988), .B2(n20556), .C1(
        n15987), .C2(n16572), .ZN(P1_U2853) );
  INV_X1 U18138 ( .A(n22159), .ZN(n16706) );
  NOR2_X1 U18139 ( .A1(n15991), .A2(n15990), .ZN(n15992) );
  OR2_X1 U18140 ( .A1(n15989), .A2(n15992), .ZN(n22163) );
  OAI22_X1 U18141 ( .A1(n22163), .A2(n20551), .B1(n15993), .B2(n20556), .ZN(
        n15994) );
  AOI21_X1 U18142 ( .B1(n16706), .B2(n13591), .A(n15994), .ZN(n15995) );
  INV_X1 U18143 ( .A(n15995), .ZN(P1_U2852) );
  XNOR2_X1 U18144 ( .A(n20593), .B(n22011), .ZN(n16692) );
  XNOR2_X1 U18145 ( .A(n16693), .B(n16692), .ZN(n22018) );
  OAI22_X1 U18146 ( .A1(n15997), .A2(n15996), .B1(n22016), .B2(n22131), .ZN(
        n15999) );
  NOR2_X1 U18147 ( .A1(n22132), .A2(n20599), .ZN(n15998) );
  AOI211_X1 U18148 ( .C1(n20623), .C2(n22129), .A(n15999), .B(n15998), .ZN(
        n16000) );
  OAI21_X1 U18149 ( .B1(n22018), .B2(n22203), .A(n16000), .ZN(P1_U2981) );
  NAND2_X1 U18150 ( .A1(n15923), .A2(n16002), .ZN(n16003) );
  INV_X1 U18151 ( .A(n22171), .ZN(n16009) );
  OAI22_X1 U18152 ( .A1(n16614), .A2(n16004), .B1(n22327), .B2(n16612), .ZN(
        n16005) );
  INV_X1 U18153 ( .A(n16005), .ZN(n16008) );
  AOI22_X1 U18154 ( .A1(n16618), .A2(n16006), .B1(n16616), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16007) );
  OAI211_X1 U18155 ( .C1(n16009), .C2(n16621), .A(n16008), .B(n16007), .ZN(
        P1_U2883) );
  NOR2_X1 U18156 ( .A1(n21290), .A2(n16010), .ZN(n16012) );
  NAND4_X1 U18157 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17945) );
  NAND2_X1 U18158 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n18058) );
  NAND2_X1 U18159 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n17964) );
  NAND4_X1 U18160 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n16014) );
  NOR4_X1 U18161 ( .A1(n17945), .A2(n18058), .A3(n17964), .A4(n16014), .ZN(
        n18002) );
  NAND3_X1 U18162 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17998) );
  NOR2_X1 U18163 ( .A1(n20971), .A2(n17998), .ZN(n17976) );
  NAND3_X1 U18164 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18002), .A3(n17976), 
        .ZN(n18211) );
  NOR2_X1 U18165 ( .A1(n21006), .A2(n18211), .ZN(n18210) );
  NAND2_X1 U18166 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18210), .ZN(n18183) );
  NOR2_X1 U18167 ( .A1(n18218), .A2(n18183), .ZN(n18197) );
  NAND2_X1 U18168 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18197), .ZN(n18196) );
  NOR2_X1 U18169 ( .A1(n18171), .A2(n18196), .ZN(n18093) );
  INV_X1 U18170 ( .A(n18093), .ZN(n18094) );
  NAND4_X1 U18171 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .A4(P3_EBX_REG_25__SCAN_IN), .ZN(n16016)
         );
  NAND4_X1 U18172 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16015)
         );
  NOR3_X1 U18173 ( .A1(n18094), .A2(n16016), .A3(n16015), .ZN(n18112) );
  NAND3_X1 U18174 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(n18112), .ZN(n18092) );
  INV_X1 U18175 ( .A(n18092), .ZN(n18091) );
  AOI21_X1 U18176 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n18112), .A(
        P3_EBX_REG_30__SCAN_IN), .ZN(n16017) );
  NOR2_X1 U18177 ( .A1(n18091), .A2(n16017), .ZN(n16114) );
  AOI22_X1 U18178 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18051), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U18179 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16020) );
  AOI22_X1 U18180 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U18181 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16018) );
  NAND4_X1 U18182 ( .A1(n16021), .A2(n16020), .A3(n16019), .A4(n16018), .ZN(
        n16029) );
  INV_X2 U18183 ( .A(n16022), .ZN(n18263) );
  AOI22_X1 U18184 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U18185 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16026) );
  CLKBUF_X1 U18186 ( .A(n18248), .Z(n20808) );
  AOI22_X1 U18187 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16025) );
  AOI22_X1 U18188 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16024) );
  NAND4_X1 U18189 ( .A1(n16027), .A2(n16026), .A3(n16025), .A4(n16024), .ZN(
        n16028) );
  NOR2_X1 U18190 ( .A1(n16029), .A2(n16028), .ZN(n16112) );
  AOI22_X1 U18191 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16033) );
  AOI22_X1 U18192 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16032) );
  AOI22_X1 U18193 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U18194 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16030) );
  NAND4_X1 U18195 ( .A1(n16033), .A2(n16032), .A3(n16031), .A4(n16030), .ZN(
        n16039) );
  AOI22_X1 U18196 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U18197 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U18198 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16035) );
  AOI22_X1 U18199 ( .A1(n18245), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16034) );
  NAND4_X1 U18200 ( .A1(n16037), .A2(n16036), .A3(n16035), .A4(n16034), .ZN(
        n16038) );
  NOR2_X1 U18201 ( .A1(n16039), .A2(n16038), .ZN(n18117) );
  AOI22_X1 U18202 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16043) );
  AOI22_X1 U18203 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16042) );
  AOI22_X1 U18204 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16041) );
  AOI22_X1 U18205 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16040) );
  NAND4_X1 U18206 ( .A1(n16043), .A2(n16042), .A3(n16041), .A4(n16040), .ZN(
        n16049) );
  AOI22_X1 U18207 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16047) );
  AOI22_X1 U18208 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U18209 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16045) );
  AOI22_X1 U18210 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16044) );
  NAND4_X1 U18211 ( .A1(n16047), .A2(n16046), .A3(n16045), .A4(n16044), .ZN(
        n16048) );
  NOR2_X1 U18212 ( .A1(n16049), .A2(n16048), .ZN(n18124) );
  AOI22_X1 U18213 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16053) );
  AOI22_X1 U18214 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18234), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16052) );
  AOI22_X1 U18215 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n18265), .ZN(n16051) );
  AOI22_X1 U18216 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18247), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16050) );
  NAND4_X1 U18217 ( .A1(n16053), .A2(n16052), .A3(n16051), .A4(n16050), .ZN(
        n16059) );
  AOI22_X1 U18218 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11171), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18245), .ZN(n16057) );
  AOI22_X1 U18219 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18263), .ZN(n16056) );
  AOI22_X1 U18220 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18254), .ZN(n16055) );
  AOI22_X1 U18221 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16054) );
  NAND4_X1 U18222 ( .A1(n16057), .A2(n16056), .A3(n16055), .A4(n16054), .ZN(
        n16058) );
  NOR2_X1 U18223 ( .A1(n16059), .A2(n16058), .ZN(n18134) );
  AOI22_X1 U18224 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U18225 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16070) );
  INV_X1 U18226 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U18227 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16060) );
  OAI21_X1 U18228 ( .B1(n16062), .B2(n16061), .A(n16060), .ZN(n16068) );
  AOI22_X1 U18229 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U18230 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U18231 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16064) );
  AOI22_X1 U18232 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16063) );
  NAND4_X1 U18233 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n16063), .ZN(
        n16067) );
  AOI211_X1 U18234 ( .C1(n18246), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n16068), .B(n16067), .ZN(n16069) );
  NAND3_X1 U18235 ( .A1(n16071), .A2(n16070), .A3(n16069), .ZN(n18140) );
  AOI22_X1 U18236 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16081) );
  AOI22_X1 U18237 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16080) );
  AOI22_X1 U18238 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16072) );
  OAI21_X1 U18239 ( .B1(n18160), .B2(n18233), .A(n16072), .ZN(n16078) );
  AOI22_X1 U18240 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U18241 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16075) );
  AOI22_X1 U18242 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U18243 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16073) );
  NAND4_X1 U18244 ( .A1(n16076), .A2(n16075), .A3(n16074), .A4(n16073), .ZN(
        n16077) );
  AOI211_X1 U18245 ( .C1(n18051), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n16078), .B(n16077), .ZN(n16079) );
  NAND3_X1 U18246 ( .A1(n16081), .A2(n16080), .A3(n16079), .ZN(n18141) );
  NAND2_X1 U18247 ( .A1(n18140), .A2(n18141), .ZN(n18139) );
  NOR2_X1 U18248 ( .A1(n18134), .A2(n18139), .ZN(n18133) );
  AOI22_X1 U18249 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16091) );
  AOI22_X1 U18250 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U18251 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16082) );
  OAI21_X1 U18252 ( .B1(n18006), .B2(n18062), .A(n16082), .ZN(n16088) );
  AOI22_X1 U18253 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U18254 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16085) );
  AOI22_X1 U18255 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16084) );
  AOI22_X1 U18256 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16083) );
  NAND4_X1 U18257 ( .A1(n16086), .A2(n16085), .A3(n16084), .A4(n16083), .ZN(
        n16087) );
  AOI211_X1 U18258 ( .C1(n18262), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n16088), .B(n16087), .ZN(n16089) );
  NAND3_X1 U18259 ( .A1(n16091), .A2(n16090), .A3(n16089), .ZN(n18130) );
  NAND2_X1 U18260 ( .A1(n18133), .A2(n18130), .ZN(n18129) );
  NOR2_X1 U18261 ( .A1(n18124), .A2(n18129), .ZN(n18123) );
  AOI22_X1 U18262 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U18263 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16100) );
  AOI22_X1 U18264 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16092) );
  OAI21_X1 U18265 ( .B1(n18006), .B2(n18159), .A(n16092), .ZN(n16098) );
  AOI22_X1 U18266 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16096) );
  AOI22_X1 U18267 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16095) );
  AOI22_X1 U18268 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16094) );
  AOI22_X1 U18269 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16093) );
  NAND4_X1 U18270 ( .A1(n16096), .A2(n16095), .A3(n16094), .A4(n16093), .ZN(
        n16097) );
  AOI211_X1 U18271 ( .C1(n18272), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n16098), .B(n16097), .ZN(n16099) );
  NAND3_X1 U18272 ( .A1(n16101), .A2(n16100), .A3(n16099), .ZN(n18107) );
  NAND2_X1 U18273 ( .A1(n18123), .A2(n18107), .ZN(n18116) );
  NOR2_X1 U18274 ( .A1(n18117), .A2(n18116), .ZN(n18115) );
  AOI22_X1 U18275 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16111) );
  AOI22_X1 U18276 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16110) );
  AOI22_X1 U18277 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16102) );
  OAI21_X1 U18278 ( .B1(n18006), .B2(n18267), .A(n16102), .ZN(n16108) );
  AOI22_X1 U18279 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U18280 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16105) );
  AOI22_X1 U18281 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16104) );
  AOI22_X1 U18282 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16103) );
  NAND4_X1 U18283 ( .A1(n16106), .A2(n16105), .A3(n16104), .A4(n16103), .ZN(
        n16107) );
  AOI211_X1 U18284 ( .C1(n18272), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16108), .B(n16107), .ZN(n16109) );
  NAND3_X1 U18285 ( .A1(n16111), .A2(n16110), .A3(n16109), .ZN(n18110) );
  NAND2_X1 U18286 ( .A1(n18115), .A2(n18110), .ZN(n18109) );
  XNOR2_X1 U18287 ( .A(n16112), .B(n18109), .ZN(n21307) );
  INV_X1 U18288 ( .A(n21307), .ZN(n16113) );
  MUX2_X1 U18289 ( .A(n16114), .B(n16113), .S(n18219), .Z(P3_U2673) );
  OAI21_X1 U18290 ( .B1(n21412), .B2(n21848), .A(n21846), .ZN(n16115) );
  NAND2_X1 U18291 ( .A1(n16121), .A2(n16115), .ZN(n21845) );
  NAND2_X1 U18292 ( .A1(n18746), .A2(n21885), .ZN(n21423) );
  NOR2_X1 U18293 ( .A1(n21845), .A2(n21423), .ZN(n16124) );
  NAND2_X1 U18294 ( .A1(n20715), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19278) );
  INV_X1 U18295 ( .A(n21875), .ZN(n22292) );
  NOR2_X1 U18296 ( .A1(n22292), .A2(n18222), .ZN(n16120) );
  AOI211_X1 U18297 ( .C1(n16120), .C2(n17655), .A(n16119), .B(n16118), .ZN(
        n16122) );
  NAND2_X1 U18298 ( .A1(n16122), .A2(n21193), .ZN(n21849) );
  NAND2_X1 U18299 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18228) );
  NOR2_X1 U18300 ( .A1(n20715), .A2(n18228), .ZN(n17653) );
  AOI22_X1 U18301 ( .A1(n21849), .A2(n21872), .B1(P3_FLUSH_REG_SCAN_IN), .B2(
        n17653), .ZN(n16123) );
  NAND2_X1 U18302 ( .A1(n19278), .A2(n16123), .ZN(n21424) );
  MUX2_X1 U18303 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n16124), .S(
        n21424), .Z(P3_U3284) );
  INV_X1 U18304 ( .A(n16478), .ZN(n16139) );
  NOR2_X1 U18305 ( .A1(n22015), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16258) );
  OAI21_X1 U18306 ( .B1(n16132), .B2(n16258), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16137) );
  INV_X1 U18307 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n16133) );
  NOR2_X1 U18308 ( .A1(n22016), .A2(n16133), .ZN(n16142) );
  INV_X1 U18309 ( .A(n16142), .ZN(n16136) );
  NAND2_X1 U18310 ( .A1(n16134), .A2(n16776), .ZN(n16722) );
  NAND2_X1 U18311 ( .A1(n16722), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16259) );
  NAND3_X1 U18312 ( .A1(n16259), .A2(n16264), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16135) );
  NAND3_X1 U18313 ( .A1(n16137), .A2(n16136), .A3(n16135), .ZN(n16138) );
  AOI21_X1 U18314 ( .B1(n16139), .B2(n22037), .A(n16138), .ZN(n16140) );
  OAI21_X1 U18315 ( .B1(n16146), .B2(n22033), .A(n16140), .ZN(P1_U3001) );
  INV_X1 U18316 ( .A(n16141), .ZN(n16470) );
  AOI21_X1 U18317 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16142), .ZN(n16143) );
  OAI21_X1 U18318 ( .B1(n20633), .B2(n16470), .A(n16143), .ZN(n16144) );
  AOI21_X1 U18319 ( .B1(n16468), .B2(n20628), .A(n16144), .ZN(n16145) );
  OAI21_X1 U18320 ( .B1(n16146), .B2(n22203), .A(n16145), .ZN(P1_U2969) );
  NAND2_X1 U18321 ( .A1(n20026), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16351) );
  INV_X1 U18322 ( .A(n16353), .ZN(n16147) );
  XOR2_X1 U18323 ( .A(n16351), .B(n16147), .Z(n19069) );
  NAND2_X1 U18324 ( .A1(n19069), .A2(n16393), .ZN(n16148) );
  INV_X1 U18325 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16244) );
  NAND2_X1 U18326 ( .A1(n16148), .A2(n16244), .ZN(n16349) );
  INV_X1 U18327 ( .A(n16148), .ZN(n16149) );
  NAND2_X1 U18328 ( .A1(n16149), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16385) );
  NAND2_X1 U18329 ( .A1(n16349), .A2(n16385), .ZN(n16215) );
  INV_X1 U18330 ( .A(n16150), .ZN(n16152) );
  AND2_X1 U18331 ( .A1(n16153), .A2(n17463), .ZN(n16154) );
  NAND2_X1 U18332 ( .A1(n16157), .A2(n16156), .ZN(n16158) );
  NAND2_X1 U18333 ( .A1(n19014), .A2(n16393), .ZN(n16170) );
  INV_X1 U18334 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17269) );
  NAND2_X1 U18335 ( .A1(n16170), .A2(n17269), .ZN(n17280) );
  INV_X1 U18336 ( .A(n16159), .ZN(n17304) );
  INV_X1 U18337 ( .A(n16160), .ZN(n16161) );
  NAND3_X1 U18338 ( .A1(n17304), .A2(n16161), .A3(n17786), .ZN(n16162) );
  NOR2_X1 U18339 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  OAI211_X1 U18340 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n16177), .A(
        n17280), .B(n16164), .ZN(n16165) );
  INV_X1 U18341 ( .A(n16165), .ZN(n16167) );
  AND2_X1 U18342 ( .A1(n16167), .A2(n16166), .ZN(n16168) );
  NAND2_X1 U18343 ( .A1(n16169), .A2(n16168), .ZN(n16180) );
  INV_X1 U18344 ( .A(n16170), .ZN(n16171) );
  NAND2_X1 U18345 ( .A1(n16171), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17281) );
  INV_X1 U18346 ( .A(n16172), .ZN(n17800) );
  INV_X1 U18347 ( .A(n16173), .ZN(n16174) );
  NAND4_X1 U18348 ( .A1(n17800), .A2(n16175), .A3(n17290), .A4(n16174), .ZN(
        n16176) );
  AOI21_X1 U18349 ( .B1(n16177), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16176), .ZN(n16178) );
  AND2_X1 U18350 ( .A1(n17281), .A2(n16178), .ZN(n16179) );
  XNOR2_X1 U18351 ( .A(n11233), .B(n16181), .ZN(n19033) );
  NAND2_X1 U18352 ( .A1(n19033), .A2(n16393), .ZN(n17416) );
  INV_X1 U18353 ( .A(n16182), .ZN(n16185) );
  INV_X1 U18354 ( .A(n16183), .ZN(n16184) );
  NAND2_X1 U18355 ( .A1(n16185), .A2(n16184), .ZN(n16186) );
  NAND2_X1 U18356 ( .A1(n16190), .A2(n16186), .ZN(n16946) );
  OR2_X1 U18357 ( .A1(n16946), .A2(n13093), .ZN(n16187) );
  INV_X1 U18358 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17398) );
  NAND2_X1 U18359 ( .A1(n16187), .A2(n17398), .ZN(n17266) );
  NAND2_X1 U18360 ( .A1(n17267), .A2(n17266), .ZN(n16188) );
  XNOR2_X1 U18361 ( .A(n16190), .B(n16189), .ZN(n16911) );
  NAND2_X1 U18362 ( .A1(n16911), .A2(n16393), .ZN(n17816) );
  INV_X1 U18363 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19112) );
  XNOR2_X1 U18364 ( .A(n16192), .B(n16191), .ZN(n16910) );
  INV_X1 U18365 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17213) );
  OAI21_X1 U18366 ( .B1(n16910), .B2(n13093), .A(n17213), .ZN(n16193) );
  AND2_X1 U18367 ( .A1(n16193), .A2(n16213), .ZN(n17242) );
  INV_X1 U18368 ( .A(n16194), .ZN(n16196) );
  XNOR2_X1 U18369 ( .A(n16196), .B(n16195), .ZN(n19049) );
  NAND2_X1 U18370 ( .A1(n19049), .A2(n16393), .ZN(n16212) );
  INV_X1 U18371 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16211) );
  NAND2_X1 U18372 ( .A1(n16212), .A2(n16211), .ZN(n17258) );
  NAND2_X1 U18373 ( .A1(n16197), .A2(n11286), .ZN(n17212) );
  INV_X1 U18374 ( .A(n16198), .ZN(n16201) );
  INV_X1 U18375 ( .A(n16199), .ZN(n16200) );
  NAND2_X1 U18376 ( .A1(n16201), .A2(n16200), .ZN(n16202) );
  NAND2_X1 U18377 ( .A1(n16203), .A2(n16202), .ZN(n16893) );
  INV_X1 U18378 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17230) );
  NOR2_X1 U18379 ( .A1(n16204), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16208) );
  INV_X1 U18380 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17353) );
  OR2_X2 U18381 ( .A1(n16205), .A2(n13093), .ZN(n17216) );
  INV_X1 U18382 ( .A(n16206), .ZN(n16207) );
  NAND2_X1 U18383 ( .A1(n17216), .A2(n17353), .ZN(n16209) );
  NAND2_X1 U18384 ( .A1(n16210), .A2(n16209), .ZN(n16214) );
  XOR2_X1 U18385 ( .A(n16215), .B(n16350), .Z(n17211) );
  AND2_X1 U18386 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19114) );
  NAND2_X1 U18387 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19114), .ZN(
        n17255) );
  NAND2_X1 U18388 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16216) );
  OR2_X1 U18389 ( .A1(n17255), .A2(n16216), .ZN(n16217) );
  NOR2_X2 U18390 ( .A1(n16218), .A2(n16217), .ZN(n17249) );
  AND2_X1 U18391 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16219) );
  NAND2_X1 U18392 ( .A1(n17249), .A2(n16219), .ZN(n16221) );
  INV_X1 U18393 ( .A(n17232), .ZN(n16220) );
  NAND2_X1 U18394 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16418) );
  NOR2_X2 U18395 ( .A1(n16221), .A2(n16418), .ZN(n16397) );
  NOR2_X1 U18396 ( .A1(n16222), .A2(n16397), .ZN(n17209) );
  NAND2_X1 U18397 ( .A1(n17451), .A2(n16223), .ZN(n16224) );
  INV_X1 U18398 ( .A(n16226), .ZN(n16227) );
  NOR2_X1 U18399 ( .A1(n16228), .A2(n16227), .ZN(n16229) );
  NAND2_X1 U18400 ( .A1(n17571), .A2(n16229), .ZN(n17425) );
  NOR2_X1 U18401 ( .A1(n17425), .A2(n17269), .ZN(n17400) );
  AND2_X1 U18402 ( .A1(n19114), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16241) );
  NAND2_X1 U18403 ( .A1(n17400), .A2(n16241), .ZN(n16230) );
  OR2_X1 U18404 ( .A1(n17598), .A2(n17593), .ZN(n17424) );
  NAND2_X1 U18405 ( .A1(n16230), .A2(n17424), .ZN(n19104) );
  NAND2_X1 U18406 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16242) );
  AOI21_X1 U18407 ( .B1(n17598), .B2(n16242), .A(n17230), .ZN(n16231) );
  AND2_X1 U18408 ( .A1(n19104), .A2(n16231), .ZN(n17371) );
  INV_X1 U18409 ( .A(n17424), .ZN(n17527) );
  NOR3_X1 U18410 ( .A1(n17371), .A2(n17527), .A3(n16244), .ZN(n16248) );
  OAI21_X1 U18411 ( .B1(n16233), .B2(n16232), .A(n16412), .ZN(n19073) );
  NAND2_X1 U18412 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16235) );
  AOI22_X1 U18413 ( .A1(n16401), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n16234) );
  OAI211_X1 U18414 ( .C1(n16236), .C2(n19060), .A(n16235), .B(n16234), .ZN(
        n16239) );
  AND2_X1 U18415 ( .A1(n16239), .A2(n16237), .ZN(n16238) );
  INV_X1 U18416 ( .A(n16400), .ZN(n16364) );
  INV_X1 U18417 ( .A(n17207), .ZN(n19066) );
  NOR2_X1 U18418 ( .A1(n17323), .A2(n19060), .ZN(n17204) );
  INV_X1 U18419 ( .A(n16418), .ZN(n16243) );
  NAND3_X1 U18420 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n17438), .ZN(n17426) );
  NOR2_X1 U18421 ( .A1(n17269), .A2(n17426), .ZN(n19113) );
  NAND2_X1 U18422 ( .A1(n16241), .A2(n19113), .ZN(n17388) );
  NOR2_X1 U18423 ( .A1(n17388), .A2(n16242), .ZN(n17364) );
  NAND2_X1 U18424 ( .A1(n17364), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17351) );
  AOI211_X1 U18425 ( .C1(n17353), .C2(n16244), .A(n16243), .B(n17351), .ZN(
        n16245) );
  AOI211_X1 U18426 ( .C1(n19066), .C2(n19159), .A(n17204), .B(n16245), .ZN(
        n16246) );
  OAI21_X1 U18427 ( .B1(n19134), .B2(n19073), .A(n16246), .ZN(n16247) );
  AOI211_X1 U18428 ( .C1(n17209), .C2(n19157), .A(n16248), .B(n16247), .ZN(
        n16249) );
  OAI21_X1 U18429 ( .B1(n17211), .B2(n19123), .A(n16249), .ZN(P2_U3017) );
  NAND2_X1 U18430 ( .A1(n16251), .A2(n16250), .ZN(n16253) );
  NAND2_X1 U18431 ( .A1(n16253), .A2(n16252), .ZN(n16256) );
  OAI22_X1 U18432 ( .A1(n16254), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n11229), .ZN(n16255) );
  NOR3_X1 U18433 ( .A1(n16259), .A2(n16258), .A3(n16257), .ZN(n16261) );
  INV_X1 U18434 ( .A(n16262), .ZN(n16265) );
  OAI21_X1 U18435 ( .B1(n16266), .B2(n22033), .A(n11278), .ZN(P1_U3000) );
  OAI22_X1 U18436 ( .A1(n16267), .A2(n20551), .B1(n16268), .B2(n20556), .ZN(
        P1_U2841) );
  NAND2_X1 U18437 ( .A1(n11208), .A2(n22197), .ZN(n16288) );
  INV_X1 U18438 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16274) );
  INV_X1 U18439 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20498) );
  NOR3_X1 U18440 ( .A1(n22131), .A2(n16271), .A3(n16270), .ZN(n16272) );
  NAND4_X1 U18441 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_17__SCAN_IN), .A4(n16272), .ZN(n22137) );
  NOR2_X1 U18442 ( .A1(n20498), .A2(n22137), .ZN(n22152) );
  NAND2_X1 U18443 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n22152), .ZN(n16275) );
  NOR2_X1 U18444 ( .A1(n22138), .A2(n16275), .ZN(n22167) );
  NAND2_X1 U18445 ( .A1(n22167), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16554) );
  NOR2_X1 U18446 ( .A1(n16276), .A2(n16554), .ZN(n22179) );
  NAND3_X1 U18447 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(n22179), .ZN(n16533) );
  NAND2_X1 U18448 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n16278) );
  NOR2_X1 U18449 ( .A1(n16533), .A2(n16278), .ZN(n16506) );
  NAND3_X1 U18450 ( .A1(n16506), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n16471) );
  NAND3_X1 U18451 ( .A1(n16284), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .ZN(n16273) );
  OAI22_X1 U18452 ( .A1(n22188), .A2(n16274), .B1(n16471), .B2(n16273), .ZN(
        n16286) );
  NAND2_X1 U18453 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n16283) );
  NOR2_X1 U18454 ( .A1(n16297), .A2(n16275), .ZN(n22154) );
  NAND2_X1 U18455 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22154), .ZN(n16549) );
  NOR3_X1 U18456 ( .A1(n16549), .A2(n16679), .A3(n16276), .ZN(n16277) );
  OR2_X1 U18457 ( .A1(n16277), .A2(n22155), .ZN(n22175) );
  OAI21_X1 U18458 ( .B1(n16672), .B2(n16278), .A(n22119), .ZN(n16279) );
  NAND2_X1 U18459 ( .A1(n22175), .A2(n16279), .ZN(n16525) );
  INV_X1 U18460 ( .A(n16525), .ZN(n16282) );
  NAND2_X1 U18461 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n16280) );
  NAND2_X1 U18462 ( .A1(n22119), .A2(n16280), .ZN(n16281) );
  NAND2_X1 U18463 ( .A1(n16282), .A2(n16281), .ZN(n16501) );
  AOI21_X1 U18464 ( .B1(n16283), .B2(n22119), .A(n16501), .ZN(n16473) );
  NOR2_X1 U18465 ( .A1(n16473), .A2(n16284), .ZN(n16285) );
  AOI211_X1 U18466 ( .C1(P1_EBX_REG_31__SCAN_IN), .C2(n11143), .A(n16286), .B(
        n16285), .ZN(n16287) );
  OAI211_X1 U18467 ( .C1(n16267), .C2(n22202), .A(n16288), .B(n16287), .ZN(
        P1_U2809) );
  AOI21_X1 U18468 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16289), .ZN(n16290) );
  OAI21_X1 U18469 ( .B1(n20633), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16290), .ZN(n16291) );
  INV_X1 U18470 ( .A(n16291), .ZN(n16294) );
  NAND3_X1 U18471 ( .A1(n16292), .A2(n14328), .A3(n20629), .ZN(n16293) );
  OAI211_X1 U18472 ( .C1(n16305), .C2(n20599), .A(n16294), .B(n16293), .ZN(
        P1_U2998) );
  AOI22_X1 U18473 ( .A1(n16295), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n16296) );
  OAI21_X1 U18474 ( .B1(n16305), .B2(n16572), .A(n16296), .ZN(P1_U2871) );
  AOI22_X1 U18475 ( .A1(n16297), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n11143), 
        .B2(P1_EBX_REG_1__SCAN_IN), .ZN(n16298) );
  OAI21_X1 U18476 ( .B1(n16299), .B2(n22202), .A(n16298), .ZN(n16301) );
  NOR2_X1 U18477 ( .A1(n22186), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16300) );
  AOI211_X1 U18478 ( .C1(n22151), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16301), .B(n16300), .ZN(n16302) );
  OAI21_X1 U18479 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n22138), .A(n16302), .ZN(
        n16303) );
  AOI21_X1 U18480 ( .B1(n22468), .B2(n22050), .A(n16303), .ZN(n16304) );
  OAI21_X1 U18481 ( .B1(n16305), .B2(n16329), .A(n16304), .ZN(P1_U2839) );
  INV_X1 U18482 ( .A(n16306), .ZN(n16307) );
  AOI21_X1 U18483 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16307), .ZN(n16308) );
  OAI21_X1 U18484 ( .B1(n20633), .B2(n16318), .A(n16308), .ZN(n16309) );
  AOI21_X1 U18485 ( .B1(n16312), .B2(n20628), .A(n16309), .ZN(n16310) );
  OAI21_X1 U18486 ( .B1(n16311), .B2(n22203), .A(n16310), .ZN(P1_U2997) );
  NAND2_X1 U18487 ( .A1(n16312), .A2(n13591), .ZN(n16314) );
  NAND2_X1 U18488 ( .A1(n16321), .A2(n20544), .ZN(n16313) );
  OAI211_X1 U18489 ( .C1(n16315), .C2(n20556), .A(n16314), .B(n16313), .ZN(
        P1_U2870) );
  OAI211_X1 U18490 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), 
        .A(n22153), .B(n16316), .ZN(n16325) );
  INV_X1 U18491 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16317) );
  OAI22_X1 U18492 ( .A1(n22188), .A2(n16317), .B1(n22095), .B2(n20476), .ZN(
        n16320) );
  NOR2_X1 U18493 ( .A1(n22186), .A2(n16318), .ZN(n16319) );
  NOR2_X1 U18494 ( .A1(n16320), .A2(n16319), .ZN(n16324) );
  NAND2_X1 U18495 ( .A1(n16557), .A2(n16321), .ZN(n16323) );
  NAND2_X1 U18496 ( .A1(n11143), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n16322) );
  NAND4_X1 U18497 ( .A1(n16325), .A2(n16324), .A3(n16323), .A4(n16322), .ZN(
        n16326) );
  AOI21_X1 U18498 ( .B1(n16327), .B2(n22050), .A(n16326), .ZN(n16328) );
  OAI21_X1 U18499 ( .B1(n16330), .B2(n16329), .A(n16328), .ZN(P1_U2838) );
  NAND2_X1 U18500 ( .A1(n20453), .A2(n14907), .ZN(n16348) );
  NOR2_X1 U18501 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22209), .ZN(n20464) );
  AOI22_X1 U18502 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20471), .B1(n20464), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n16333) );
  OAI21_X1 U18503 ( .B1(n12191), .B2(n16348), .A(n16333), .ZN(P1_U2920) );
  AOI22_X1 U18504 ( .A1(n21905), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n16334) );
  OAI21_X1 U18505 ( .B1(n15743), .B2(n16348), .A(n16334), .ZN(P1_U2919) );
  INV_X1 U18506 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n22311) );
  AOI22_X1 U18507 ( .A1(n21905), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n16335) );
  OAI21_X1 U18508 ( .B1(n22311), .B2(n16348), .A(n16335), .ZN(P1_U2918) );
  AOI22_X1 U18509 ( .A1(n21905), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n16336) );
  OAI21_X1 U18510 ( .B1(n22316), .B2(n16348), .A(n16336), .ZN(P1_U2917) );
  AOI22_X1 U18511 ( .A1(n21905), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n16337) );
  OAI21_X1 U18512 ( .B1(n22321), .B2(n16348), .A(n16337), .ZN(P1_U2916) );
  AOI22_X1 U18513 ( .A1(n21905), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n16338) );
  OAI21_X1 U18514 ( .B1(n22327), .B2(n16348), .A(n16338), .ZN(P1_U2915) );
  INV_X1 U18515 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n22332) );
  AOI22_X1 U18516 ( .A1(n21905), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n16339) );
  OAI21_X1 U18517 ( .B1(n22332), .B2(n16348), .A(n16339), .ZN(P1_U2914) );
  AOI22_X1 U18518 ( .A1(n21905), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n16340) );
  OAI21_X1 U18519 ( .B1(n22337), .B2(n16348), .A(n16340), .ZN(P1_U2913) );
  AOI22_X1 U18520 ( .A1(n21905), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n16341) );
  OAI21_X1 U18521 ( .B1(n22343), .B2(n16348), .A(n16341), .ZN(P1_U2912) );
  INV_X1 U18522 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n22350) );
  AOI22_X1 U18523 ( .A1(n21905), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n16342) );
  OAI21_X1 U18524 ( .B1(n22350), .B2(n16348), .A(n16342), .ZN(P1_U2911) );
  AOI22_X1 U18525 ( .A1(n21905), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n16343) );
  OAI21_X1 U18526 ( .B1(n22356), .B2(n16348), .A(n16343), .ZN(P1_U2910) );
  INV_X1 U18527 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n22361) );
  AOI22_X1 U18528 ( .A1(n21905), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n16344) );
  OAI21_X1 U18529 ( .B1(n22361), .B2(n16348), .A(n16344), .ZN(P1_U2909) );
  AOI22_X1 U18530 ( .A1(n21905), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n16345) );
  OAI21_X1 U18531 ( .B1(n22368), .B2(n16348), .A(n16345), .ZN(P1_U2908) );
  AOI22_X1 U18532 ( .A1(n21905), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n16346) );
  OAI21_X1 U18533 ( .B1(n22375), .B2(n16348), .A(n16346), .ZN(P1_U2907) );
  INV_X1 U18534 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n22383) );
  AOI22_X1 U18535 ( .A1(n21905), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n16347) );
  OAI21_X1 U18536 ( .B1(n22383), .B2(n16348), .A(n16347), .ZN(P1_U2906) );
  NAND2_X1 U18537 ( .A1(n16389), .A2(n16385), .ZN(n16357) );
  INV_X1 U18538 ( .A(n16351), .ZN(n16352) );
  NAND2_X1 U18539 ( .A1(n20026), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16354) );
  XNOR2_X1 U18540 ( .A(n16390), .B(n16354), .ZN(n16862) );
  AOI21_X1 U18541 ( .B1(n16862), .B2(n16393), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16388) );
  AND2_X1 U18542 ( .A1(n16393), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16355) );
  NOR2_X1 U18543 ( .A1(n16388), .A2(n11288), .ZN(n16356) );
  XNOR2_X1 U18544 ( .A(n16357), .B(n16356), .ZN(n16380) );
  XNOR2_X1 U18545 ( .A(n16397), .B(n16358), .ZN(n16378) );
  NAND2_X1 U18546 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17371), .ZN(
        n16359) );
  OAI21_X1 U18547 ( .B1(n16359), .B2(n16418), .A(n17424), .ZN(n16424) );
  NOR2_X1 U18548 ( .A1(n16424), .A2(n16358), .ZN(n16369) );
  INV_X1 U18549 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17937) );
  NAND2_X1 U18550 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16362) );
  AOI22_X1 U18551 ( .A1(n11221), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n16361) );
  OAI211_X1 U18552 ( .C1(n16236), .C2(n17937), .A(n16362), .B(n16361), .ZN(
        n16399) );
  NOR3_X1 U18553 ( .A1(n17351), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16418), .ZN(n16365) );
  NOR2_X1 U18554 ( .A1(n18958), .A2(n17937), .ZN(n16372) );
  OAI21_X1 U18555 ( .B1(n16373), .B2(n19130), .A(n16367), .ZN(n16368) );
  OAI21_X1 U18556 ( .B1(n16380), .B2(n19123), .A(n16370), .ZN(P2_U3016) );
  INV_X1 U18557 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16371) );
  XNOR2_X1 U18558 ( .A(n16851), .B(n16371), .ZN(n16854) );
  INV_X1 U18559 ( .A(n16854), .ZN(n16866) );
  INV_X1 U18560 ( .A(n16372), .ZN(n16374) );
  INV_X1 U18561 ( .A(n16375), .ZN(n16376) );
  OAI21_X1 U18562 ( .B1(n16866), .B2(n17827), .A(n16376), .ZN(n16377) );
  OAI21_X1 U18563 ( .B1(n16380), .B2(n13196), .A(n16379), .ZN(P2_U2984) );
  AOI22_X1 U18564 ( .A1(n16381), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15728), .ZN(n16383) );
  AOI22_X1 U18565 ( .A1(n16618), .A2(n22379), .B1(n16616), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n16382) );
  OAI211_X1 U18566 ( .C1(n16384), .C2(n16621), .A(n16383), .B(n16382), .ZN(
        P1_U2874) );
  INV_X1 U18567 ( .A(n16385), .ZN(n16386) );
  NOR2_X1 U18568 ( .A1(n16390), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16392) );
  MUX2_X1 U18569 ( .A(n16392), .B(n13103), .S(n16391), .Z(n16848) );
  NAND2_X1 U18570 ( .A1(n16848), .A2(n16393), .ZN(n16394) );
  XNOR2_X1 U18571 ( .A(n16394), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16395) );
  XNOR2_X1 U18572 ( .A(n16396), .B(n16395), .ZN(n16431) );
  NAND2_X1 U18573 ( .A1(n16397), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16398) );
  INV_X1 U18574 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17938) );
  NOR2_X1 U18575 ( .A1(n18958), .A2(n17938), .ZN(n16419) );
  NAND2_X1 U18576 ( .A1(n16400), .A2(n16399), .ZN(n16406) );
  AOI22_X1 U18577 ( .A1(n16401), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n16402) );
  OAI21_X1 U18578 ( .B1(n16236), .B2(n17938), .A(n16402), .ZN(n16403) );
  AOI21_X1 U18579 ( .B1(n16404), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16403), .ZN(n16405) );
  NOR2_X1 U18580 ( .A1(n16422), .A2(n13199), .ZN(n16407) );
  OAI21_X1 U18581 ( .B1(n16409), .B2(n17827), .A(n16408), .ZN(n16410) );
  OAI21_X1 U18582 ( .B1(n16431), .B2(n13196), .A(n16411), .ZN(P2_U2983) );
  AOI222_X1 U18583 ( .A1(n16415), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n16414), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), 
        .C2(n13345), .ZN(n16416) );
  XNOR2_X1 U18584 ( .A(n16417), .B(n16416), .ZN(n19707) );
  NOR4_X1 U18585 ( .A1(n17351), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16358), .A4(n16418), .ZN(n16420) );
  OAI21_X1 U18586 ( .B1(n16431), .B2(n19123), .A(n16430), .ZN(P2_U3015) );
  INV_X1 U18587 ( .A(n16432), .ZN(n16433) );
  XNOR2_X1 U18588 ( .A(n16436), .B(n16435), .ZN(n16443) );
  NOR2_X1 U18589 ( .A1(n17207), .A2(n11164), .ZN(n16437) );
  AOI21_X1 U18590 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n11163), .A(n16437), .ZN(
        n16438) );
  OAI21_X1 U18591 ( .B1(n16443), .B2(n17128), .A(n16438), .ZN(P2_U2858) );
  INV_X1 U18592 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n17911) );
  OAI22_X1 U18593 ( .A1(n20172), .A2(n19073), .B1(n20066), .B2(n17911), .ZN(
        n16439) );
  AOI21_X1 U18594 ( .B1(n20168), .B2(n16440), .A(n16439), .ZN(n16442) );
  AOI22_X1 U18595 ( .A1(n20169), .A2(BUF1_REG_29__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n16441) );
  OAI211_X1 U18596 ( .C1(n16443), .C2(n20222), .A(n16442), .B(n16441), .ZN(
        P2_U2890) );
  NOR2_X1 U18597 ( .A1(n16373), .A2(n11163), .ZN(n16444) );
  AOI21_X1 U18598 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n11164), .A(n16444), .ZN(
        n16445) );
  OAI21_X1 U18599 ( .B1(n16446), .B2(n17128), .A(n16445), .ZN(P2_U2857) );
  INV_X1 U18600 ( .A(n16447), .ZN(n16453) );
  NOR2_X1 U18601 ( .A1(n16448), .A2(n16453), .ZN(n16464) );
  INV_X1 U18602 ( .A(n16464), .ZN(n16449) );
  OAI21_X1 U18603 ( .B1(n16449), .B2(n22220), .A(P1_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n16452) );
  NAND3_X1 U18604 ( .A1(n16452), .A2(n16451), .A3(n16450), .ZN(P1_U2801) );
  NAND2_X1 U18605 ( .A1(n16459), .A2(n16463), .ZN(n16457) );
  NAND2_X1 U18606 ( .A1(n11712), .A2(n16453), .ZN(n16456) );
  NAND2_X1 U18607 ( .A1(n16454), .A2(n16461), .ZN(n16455) );
  NAND3_X1 U18608 ( .A1(n16457), .A2(n16456), .A3(n16455), .ZN(n16458) );
  AOI21_X1 U18609 ( .B1(n16460), .B2(n16459), .A(n16458), .ZN(n17693) );
  INV_X1 U18610 ( .A(n17693), .ZN(n16467) );
  OAI22_X1 U18611 ( .A1(n16464), .A2(n16463), .B1(n16462), .B2(n16461), .ZN(
        n20634) );
  INV_X1 U18612 ( .A(n16465), .ZN(n16466) );
  AOI21_X1 U18613 ( .B1(n16466), .B2(n22254), .A(n22242), .ZN(n21906) );
  NOR2_X1 U18614 ( .A1(n20634), .A2(n21906), .ZN(n17689) );
  NOR2_X1 U18615 ( .A1(n17689), .A2(n22220), .ZN(n22205) );
  MUX2_X1 U18616 ( .A(P1_MORE_REG_SCAN_IN), .B(n16467), .S(n22205), .Z(
        P1_U3484) );
  NAND2_X1 U18617 ( .A1(n16468), .A2(n22197), .ZN(n16477) );
  OAI22_X1 U18618 ( .A1(n16470), .A2(n22186), .B1(n22188), .B2(n16469), .ZN(
        n16475) );
  INV_X1 U18619 ( .A(n16471), .ZN(n16481) );
  AOI21_X1 U18620 ( .B1(n16481), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n16472) );
  NOR2_X1 U18621 ( .A1(n16473), .A2(n16472), .ZN(n16474) );
  AOI211_X1 U18622 ( .C1(P1_EBX_REG_30__SCAN_IN), .C2(n11143), .A(n16475), .B(
        n16474), .ZN(n16476) );
  OAI211_X1 U18623 ( .C1(n16478), .C2(n22202), .A(n16477), .B(n16476), .ZN(
        P1_U2810) );
  INV_X1 U18624 ( .A(n16479), .ZN(n16579) );
  AOI22_X1 U18625 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n16481), .B2(n16480), .ZN(n16483) );
  NAND2_X1 U18626 ( .A1(n11143), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n16482) );
  OAI211_X1 U18627 ( .C1(n22186), .C2(n16484), .A(n16483), .B(n16482), .ZN(
        n16485) );
  AOI21_X1 U18628 ( .B1(n16501), .B2(P1_REIP_REG_29__SCAN_IN), .A(n16485), 
        .ZN(n16487) );
  NAND2_X1 U18629 ( .A1(n16559), .A2(n16557), .ZN(n16486) );
  OAI211_X1 U18630 ( .C1(n16579), .C2(n22181), .A(n16487), .B(n16486), .ZN(
        P1_U2811) );
  BUF_X1 U18631 ( .A(n16488), .Z(n16489) );
  INV_X1 U18632 ( .A(n16492), .ZN(n16634) );
  INV_X1 U18633 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16641) );
  NOR2_X1 U18634 ( .A1(n16641), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16493) );
  AOI22_X1 U18635 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n16506), .B2(n16493), .ZN(n16495) );
  NAND2_X1 U18636 ( .A1(n11143), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n16494) );
  OAI211_X1 U18637 ( .C1(n22186), .C2(n16634), .A(n16495), .B(n16494), .ZN(
        n16500) );
  OAI21_X1 U18638 ( .B1(n16496), .B2(n16498), .A(n16497), .ZN(n16712) );
  NOR2_X1 U18639 ( .A1(n16712), .A2(n22202), .ZN(n16499) );
  AOI211_X1 U18640 ( .C1(P1_REIP_REG_28__SCAN_IN), .C2(n16501), .A(n16500), 
        .B(n16499), .ZN(n16502) );
  OAI21_X1 U18641 ( .B1(n16631), .B2(n22181), .A(n16502), .ZN(P1_U2812) );
  BUF_X1 U18642 ( .A(n16503), .Z(n16504) );
  AOI21_X1 U18643 ( .B1(n16505), .B2(n16504), .A(n16489), .ZN(n16645) );
  INV_X1 U18644 ( .A(n16645), .ZN(n16588) );
  AOI22_X1 U18645 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n16506), .B2(n16641), .ZN(n16508) );
  NAND2_X1 U18646 ( .A1(n11143), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n16507) );
  OAI211_X1 U18647 ( .C1(n22186), .C2(n16643), .A(n16508), .B(n16507), .ZN(
        n16509) );
  AOI21_X1 U18648 ( .B1(n16525), .B2(P1_REIP_REG_27__SCAN_IN), .A(n16509), 
        .ZN(n16513) );
  AOI21_X1 U18649 ( .B1(n16511), .B2(n16521), .A(n16496), .ZN(n16724) );
  NAND2_X1 U18650 ( .A1(n16724), .A2(n16557), .ZN(n16512) );
  OAI211_X1 U18651 ( .C1(n16588), .C2(n22181), .A(n16513), .B(n16512), .ZN(
        P1_U2813) );
  OAI21_X1 U18652 ( .B1(n16515), .B2(n16516), .A(n16504), .ZN(n16647) );
  INV_X1 U18653 ( .A(n16653), .ZN(n16520) );
  NAND2_X1 U18654 ( .A1(n11143), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n16519) );
  INV_X1 U18655 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n16662) );
  NOR3_X1 U18656 ( .A1(n16533), .A2(n16662), .A3(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n16517) );
  AOI21_X1 U18657 ( .B1(n22151), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16517), .ZN(n16518) );
  OAI211_X1 U18658 ( .C1(n22186), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        n16524) );
  OAI21_X1 U18659 ( .B1(n16530), .B2(n16522), .A(n16521), .ZN(n16738) );
  NOR2_X1 U18660 ( .A1(n16738), .A2(n22202), .ZN(n16523) );
  AOI211_X1 U18661 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n16525), .A(n16524), 
        .B(n16523), .ZN(n16526) );
  OAI21_X1 U18662 ( .B1(n16647), .B2(n22181), .A(n16526), .ZN(P1_U2814) );
  NOR2_X1 U18663 ( .A1(n16527), .A2(n16528), .ZN(n16529) );
  OR2_X1 U18664 ( .A1(n16530), .A2(n16529), .ZN(n16743) );
  AOI21_X1 U18665 ( .B1(n16532), .B2(n16571), .A(n16515), .ZN(n16666) );
  NAND2_X1 U18666 ( .A1(n16666), .A2(n22197), .ZN(n16542) );
  INV_X1 U18667 ( .A(n16533), .ZN(n16534) );
  AOI22_X1 U18668 ( .A1(n22151), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n16534), .B2(n16662), .ZN(n16535) );
  OAI21_X1 U18669 ( .B1(n16664), .B2(n22186), .A(n16535), .ZN(n16540) );
  INV_X1 U18670 ( .A(n22179), .ZN(n16536) );
  NOR2_X1 U18671 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n16536), .ZN(n16537) );
  AND2_X1 U18672 ( .A1(n16537), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n22193) );
  INV_X1 U18673 ( .A(n22193), .ZN(n16538) );
  AOI21_X1 U18674 ( .B1(n22175), .B2(n16538), .A(n16662), .ZN(n16539) );
  AOI211_X1 U18675 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n11143), .A(n16540), .B(
        n16539), .ZN(n16541) );
  OAI211_X1 U18676 ( .C1(n22202), .C2(n16743), .A(n16542), .B(n16541), .ZN(
        P1_U2815) );
  AOI21_X1 U18677 ( .B1(n16544), .B2(n16001), .A(n16605), .ZN(n16690) );
  INV_X1 U18678 ( .A(n16690), .ZN(n16622) );
  OR2_X1 U18679 ( .A1(n16546), .A2(n16547), .ZN(n16548) );
  NAND2_X1 U18680 ( .A1(n11183), .A2(n16548), .ZN(n16574) );
  INV_X1 U18681 ( .A(n16574), .ZN(n22036) );
  AND3_X1 U18682 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n22119), .A3(n16549), 
        .ZN(n16556) );
  INV_X1 U18683 ( .A(n16550), .ZN(n16688) );
  OAI22_X1 U18684 ( .A1(n16551), .A2(n22188), .B1(n22186), .B2(n16688), .ZN(
        n16552) );
  AOI21_X1 U18685 ( .B1(n11143), .B2(P1_EBX_REG_22__SCAN_IN), .A(n16552), .ZN(
        n16553) );
  OAI21_X1 U18686 ( .B1(n16554), .B2(P1_REIP_REG_22__SCAN_IN), .A(n16553), 
        .ZN(n16555) );
  AOI211_X1 U18687 ( .C1(n22036), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        n16558) );
  OAI21_X1 U18688 ( .B1(n16622), .B2(n22181), .A(n16558), .ZN(P1_U2818) );
  AOI22_X1 U18689 ( .A1(n16559), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n16560) );
  OAI21_X1 U18690 ( .B1(n16579), .B2(n16572), .A(n16560), .ZN(P1_U2843) );
  INV_X1 U18691 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16561) );
  OAI222_X1 U18692 ( .A1(n16561), .A2(n20556), .B1(n20551), .B2(n16712), .C1(
        n16631), .C2(n16572), .ZN(P1_U2844) );
  AOI22_X1 U18693 ( .A1(n16724), .A2(n20544), .B1(n16562), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n16563) );
  OAI21_X1 U18694 ( .B1(n16588), .B2(n16572), .A(n16563), .ZN(P1_U2845) );
  INV_X1 U18695 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16564) );
  OAI222_X1 U18696 ( .A1(n16738), .A2(n20551), .B1(n16564), .B2(n20556), .C1(
        n16647), .C2(n16572), .ZN(P1_U2846) );
  INV_X1 U18697 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16565) );
  INV_X1 U18698 ( .A(n16666), .ZN(n16598) );
  OAI222_X1 U18699 ( .A1(n16565), .A2(n20556), .B1(n20551), .B2(n16743), .C1(
        n16598), .C2(n16572), .ZN(P1_U2847) );
  AND2_X1 U18700 ( .A1(n16760), .A2(n16566), .ZN(n16567) );
  OR2_X1 U18701 ( .A1(n16567), .A2(n16527), .ZN(n22201) );
  OR2_X1 U18702 ( .A1(n16568), .A2(n16569), .ZN(n16570) );
  AND2_X1 U18703 ( .A1(n16571), .A2(n16570), .ZN(n22198) );
  INV_X1 U18704 ( .A(n22198), .ZN(n16603) );
  OAI222_X1 U18705 ( .A1(n22201), .A2(n20551), .B1(n22190), .B2(n20556), .C1(
        n16603), .C2(n16572), .ZN(P1_U2848) );
  INV_X1 U18706 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16573) );
  OAI222_X1 U18707 ( .A1(n16574), .A2(n20551), .B1(n16573), .B2(n20556), .C1(
        n16622), .C2(n16572), .ZN(P1_U2850) );
  OAI22_X1 U18708 ( .A1(n16614), .A2(n16575), .B1(n22375), .B2(n16612), .ZN(
        n16576) );
  INV_X1 U18709 ( .A(n16576), .ZN(n16578) );
  AOI22_X1 U18710 ( .A1(n16618), .A2(n22372), .B1(n16616), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16577) );
  OAI211_X1 U18711 ( .C1(n16579), .C2(n16621), .A(n16578), .B(n16577), .ZN(
        P1_U2875) );
  OAI22_X1 U18712 ( .A1(n16614), .A2(n14664), .B1(n22368), .B2(n16612), .ZN(
        n16580) );
  INV_X1 U18713 ( .A(n16580), .ZN(n16582) );
  AOI22_X1 U18714 ( .A1(n16618), .A2(n22365), .B1(n16616), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16581) );
  OAI211_X1 U18715 ( .C1(n16631), .C2(n16621), .A(n16582), .B(n16581), .ZN(
        P1_U2876) );
  OAI22_X1 U18716 ( .A1(n16614), .A2(n16583), .B1(n22361), .B2(n16612), .ZN(
        n16584) );
  INV_X1 U18717 ( .A(n16584), .ZN(n16587) );
  AOI22_X1 U18718 ( .A1(n16618), .A2(n16585), .B1(n16616), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16586) );
  OAI211_X1 U18719 ( .C1(n16588), .C2(n16621), .A(n16587), .B(n16586), .ZN(
        P1_U2877) );
  OAI22_X1 U18720 ( .A1(n16614), .A2(n16589), .B1(n22356), .B2(n16612), .ZN(
        n16590) );
  INV_X1 U18721 ( .A(n16590), .ZN(n16593) );
  AOI22_X1 U18722 ( .A1(n16618), .A2(n16591), .B1(n16616), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16592) );
  OAI211_X1 U18723 ( .C1(n16647), .C2(n16621), .A(n16593), .B(n16592), .ZN(
        P1_U2878) );
  OAI22_X1 U18724 ( .A1(n16614), .A2(n16594), .B1(n22350), .B2(n16612), .ZN(
        n16595) );
  INV_X1 U18725 ( .A(n16595), .ZN(n16597) );
  AOI22_X1 U18726 ( .A1(n16618), .A2(n22347), .B1(n16616), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16596) );
  OAI211_X1 U18727 ( .C1(n16598), .C2(n16621), .A(n16597), .B(n16596), .ZN(
        P1_U2879) );
  OAI22_X1 U18728 ( .A1(n16614), .A2(n16599), .B1(n22343), .B2(n16612), .ZN(
        n16600) );
  INV_X1 U18729 ( .A(n16600), .ZN(n16602) );
  AOI22_X1 U18730 ( .A1(n16618), .A2(n22340), .B1(n16616), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16601) );
  OAI211_X1 U18731 ( .C1(n16603), .C2(n16621), .A(n16602), .B(n16601), .ZN(
        P1_U2880) );
  NOR2_X1 U18732 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  OR2_X1 U18733 ( .A1(n16568), .A2(n16606), .ZN(n22182) );
  INV_X1 U18734 ( .A(DATAI_23_), .ZN(n16607) );
  OAI22_X1 U18735 ( .A1(n16614), .A2(n16607), .B1(n22337), .B2(n16612), .ZN(
        n16608) );
  INV_X1 U18736 ( .A(n16608), .ZN(n16611) );
  AOI22_X1 U18737 ( .A1(n16618), .A2(n16609), .B1(n16616), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16610) );
  OAI211_X1 U18738 ( .C1(n22182), .C2(n16621), .A(n16611), .B(n16610), .ZN(
        P1_U2881) );
  OAI22_X1 U18739 ( .A1(n16614), .A2(n16613), .B1(n22332), .B2(n16612), .ZN(
        n16615) );
  INV_X1 U18740 ( .A(n16615), .ZN(n16620) );
  AOI22_X1 U18741 ( .A1(n16618), .A2(n16617), .B1(n16616), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16619) );
  OAI211_X1 U18742 ( .C1(n16622), .C2(n16621), .A(n16620), .B(n16619), .ZN(
        P1_U2882) );
  INV_X1 U18743 ( .A(n16678), .ZN(n16668) );
  NAND2_X1 U18744 ( .A1(n16668), .A2(n16624), .ZN(n16629) );
  INV_X1 U18745 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U18746 ( .A1(n16625), .A2(n16721), .ZN(n16626) );
  MUX2_X1 U18747 ( .A(n16626), .B(n16734), .S(n20593), .Z(n16628) );
  NOR2_X1 U18748 ( .A1(n16629), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16627) );
  AOI211_X1 U18749 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16629), .A(
        n16628), .B(n16627), .ZN(n16630) );
  XNOR2_X1 U18750 ( .A(n16630), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16716) );
  INV_X1 U18751 ( .A(n16631), .ZN(n16636) );
  INV_X1 U18752 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n16632) );
  NOR2_X1 U18753 ( .A1(n22016), .A2(n16632), .ZN(n16710) );
  AOI21_X1 U18754 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16710), .ZN(n16633) );
  OAI21_X1 U18755 ( .B1(n20633), .B2(n16634), .A(n16633), .ZN(n16635) );
  AOI21_X1 U18756 ( .B1(n16636), .B2(n20628), .A(n16635), .ZN(n16637) );
  OAI21_X1 U18757 ( .B1(n22203), .B2(n16716), .A(n16637), .ZN(P1_U2971) );
  XNOR2_X1 U18758 ( .A(n16794), .B(n16721), .ZN(n16640) );
  XNOR2_X1 U18759 ( .A(n16639), .B(n16640), .ZN(n16726) );
  NOR2_X1 U18760 ( .A1(n22016), .A2(n16641), .ZN(n16718) );
  AOI21_X1 U18761 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16718), .ZN(n16642) );
  OAI21_X1 U18762 ( .B1(n20633), .B2(n16643), .A(n16642), .ZN(n16644) );
  AOI21_X1 U18763 ( .B1(n16645), .B2(n20628), .A(n16644), .ZN(n16646) );
  OAI21_X1 U18764 ( .B1(n16726), .B2(n22203), .A(n16646), .ZN(P1_U2972) );
  INV_X1 U18765 ( .A(n16647), .ZN(n16648) );
  NAND2_X1 U18766 ( .A1(n16648), .A2(n20628), .ZN(n16657) );
  INV_X1 U18767 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16649) );
  NOR2_X1 U18768 ( .A1(n22016), .A2(n16649), .ZN(n16733) );
  AOI21_X1 U18769 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16733), .ZN(n16656) );
  NAND2_X1 U18771 ( .A1(n16652), .A2(n16734), .ZN(n16727) );
  NAND3_X1 U18772 ( .A1(n22731), .A2(n20629), .A3(n16727), .ZN(n16655) );
  NAND2_X1 U18773 ( .A1(n20623), .A2(n16653), .ZN(n16654) );
  NAND4_X1 U18774 ( .A1(n16657), .A2(n16656), .A3(n16655), .A4(n16654), .ZN(
        P1_U2973) );
  MUX2_X1 U18775 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n16658), .S(
        n20593), .Z(n16660) );
  NOR2_X1 U18776 ( .A1(n16678), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16659) );
  AOI211_X1 U18777 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16750), .A(
        n16660), .B(n16659), .ZN(n16661) );
  XNOR2_X1 U18778 ( .A(n16661), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16747) );
  NOR2_X1 U18779 ( .A1(n22016), .A2(n16662), .ZN(n16741) );
  AOI21_X1 U18780 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16741), .ZN(n16663) );
  OAI21_X1 U18781 ( .B1(n20633), .B2(n16664), .A(n16663), .ZN(n16665) );
  AOI21_X1 U18782 ( .B1(n16666), .B2(n20628), .A(n16665), .ZN(n16667) );
  OAI21_X1 U18783 ( .B1(n16747), .B2(n22203), .A(n16667), .ZN(P1_U2974) );
  NAND3_X1 U18784 ( .A1(n16668), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n11597), .ZN(n16670) );
  NAND3_X1 U18785 ( .A1(n16678), .A2(n11595), .A3(n16750), .ZN(n16669) );
  NAND2_X1 U18786 ( .A1(n16670), .A2(n16669), .ZN(n16671) );
  XNOR2_X1 U18787 ( .A(n16671), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16757) );
  INV_X1 U18788 ( .A(n22196), .ZN(n16674) );
  NOR2_X1 U18789 ( .A1(n22016), .A2(n16672), .ZN(n16752) );
  AOI21_X1 U18790 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16752), .ZN(n16673) );
  OAI21_X1 U18791 ( .B1(n20633), .B2(n16674), .A(n16673), .ZN(n16675) );
  AOI21_X1 U18792 ( .B1(n22198), .B2(n20628), .A(n16675), .ZN(n16676) );
  OAI21_X1 U18793 ( .B1(n16757), .B2(n22203), .A(n16676), .ZN(P1_U2975) );
  XNOR2_X1 U18794 ( .A(n16794), .B(n16750), .ZN(n16677) );
  XNOR2_X1 U18795 ( .A(n16678), .B(n16677), .ZN(n16768) );
  INV_X1 U18796 ( .A(n22182), .ZN(n16682) );
  NOR2_X1 U18797 ( .A1(n22016), .A2(n16679), .ZN(n16761) );
  AOI21_X1 U18798 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16761), .ZN(n16680) );
  OAI21_X1 U18799 ( .B1(n20633), .B2(n22187), .A(n16680), .ZN(n16681) );
  AOI21_X1 U18800 ( .B1(n16682), .B2(n20628), .A(n16681), .ZN(n16683) );
  OAI21_X1 U18801 ( .B1(n16768), .B2(n22203), .A(n16683), .ZN(P1_U2976) );
  NOR2_X1 U18802 ( .A1(n16685), .A2(n16684), .ZN(n16686) );
  XNOR2_X1 U18803 ( .A(n16686), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n22035) );
  AOI22_X1 U18804 ( .A1(n20627), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n22040), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16687) );
  OAI21_X1 U18805 ( .B1(n20633), .B2(n16688), .A(n16687), .ZN(n16689) );
  AOI21_X1 U18806 ( .B1(n16690), .B2(n20628), .A(n16689), .ZN(n16691) );
  OAI21_X1 U18807 ( .B1(n22203), .B2(n22035), .A(n16691), .ZN(P1_U2977) );
  NOR2_X1 U18808 ( .A1(n16693), .A2(n16692), .ZN(n16694) );
  AOI21_X1 U18809 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n11595), .A(
        n16694), .ZN(n16796) );
  OAI22_X1 U18810 ( .A1(n16796), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11595), .B2(n16694), .ZN(n16700) );
  MUX2_X1 U18811 ( .A(n11595), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n16785), .Z(n16695) );
  NOR2_X1 U18812 ( .A1(n16700), .A2(n16695), .ZN(n16696) );
  XNOR2_X1 U18813 ( .A(n16696), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16769) );
  INV_X1 U18814 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22166) );
  NOR2_X1 U18815 ( .A1(n22016), .A2(n22166), .ZN(n16779) );
  AOI21_X1 U18816 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16779), .ZN(n16697) );
  OAI21_X1 U18817 ( .B1(n20633), .B2(n22174), .A(n16697), .ZN(n16698) );
  AOI21_X1 U18818 ( .B1(n22171), .B2(n20628), .A(n16698), .ZN(n16699) );
  OAI21_X1 U18819 ( .B1(n16769), .B2(n22203), .A(n16699), .ZN(P1_U2978) );
  AOI21_X1 U18820 ( .B1(n11595), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16700), .ZN(n16701) );
  XNOR2_X1 U18821 ( .A(n16701), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16793) );
  INV_X1 U18822 ( .A(n22161), .ZN(n16704) );
  NOR2_X1 U18823 ( .A1(n22016), .A2(n16702), .ZN(n16788) );
  AOI21_X1 U18824 ( .B1(n20627), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16788), .ZN(n16703) );
  OAI21_X1 U18825 ( .B1(n20633), .B2(n16704), .A(n16703), .ZN(n16705) );
  AOI21_X1 U18826 ( .B1(n16706), .B2(n20628), .A(n16705), .ZN(n16707) );
  OAI21_X1 U18827 ( .B1(n16793), .B2(n22203), .A(n16707), .ZN(P1_U2979) );
  INV_X1 U18828 ( .A(n16722), .ZN(n16711) );
  NOR3_X1 U18829 ( .A1(n16717), .A2(n16708), .A3(n11700), .ZN(n16709) );
  AOI211_X1 U18830 ( .C1(n16711), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16710), .B(n16709), .ZN(n16715) );
  INV_X1 U18831 ( .A(n16712), .ZN(n16713) );
  NAND2_X1 U18832 ( .A1(n16713), .A2(n22037), .ZN(n16714) );
  OAI211_X1 U18833 ( .C1(n16716), .C2(n22033), .A(n16715), .B(n16714), .ZN(
        P1_U3003) );
  INV_X1 U18834 ( .A(n16717), .ZN(n16719) );
  AOI21_X1 U18835 ( .B1(n16719), .B2(n16721), .A(n16718), .ZN(n16720) );
  OAI21_X1 U18836 ( .B1(n16722), .B2(n16721), .A(n16720), .ZN(n16723) );
  AOI21_X1 U18837 ( .B1(n16724), .B2(n22037), .A(n16723), .ZN(n16725) );
  OAI21_X1 U18838 ( .B1(n16726), .B2(n22033), .A(n16725), .ZN(P1_U3004) );
  NAND3_X1 U18839 ( .A1(n22731), .A2(n22038), .A3(n16727), .ZN(n16737) );
  INV_X1 U18840 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16728) );
  NAND2_X1 U18841 ( .A1(n16729), .A2(n16728), .ZN(n16730) );
  NOR2_X1 U18842 ( .A1(n16764), .A2(n16730), .ZN(n16740) );
  INV_X1 U18843 ( .A(n16740), .ZN(n16731) );
  AOI21_X1 U18844 ( .B1(n16739), .B2(n16731), .A(n16734), .ZN(n16732) );
  AOI211_X1 U18845 ( .C1(n16735), .C2(n16734), .A(n16733), .B(n16732), .ZN(
        n16736) );
  OAI211_X1 U18846 ( .C1(n22017), .C2(n16738), .A(n16737), .B(n16736), .ZN(
        P1_U3005) );
  INV_X1 U18847 ( .A(n16739), .ZN(n16742) );
  AOI211_X1 U18848 ( .C1(n16742), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16741), .B(n16740), .ZN(n16746) );
  INV_X1 U18849 ( .A(n16743), .ZN(n16744) );
  NAND2_X1 U18850 ( .A1(n16744), .A2(n22037), .ZN(n16745) );
  OAI211_X1 U18851 ( .C1(n16747), .C2(n22033), .A(n16746), .B(n16745), .ZN(
        P1_U3006) );
  INV_X1 U18852 ( .A(n16762), .ZN(n16748) );
  OAI21_X1 U18853 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16749), .A(
        n16748), .ZN(n16753) );
  NOR3_X1 U18854 ( .A1(n16764), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16750), .ZN(n16751) );
  AOI211_X1 U18855 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16753), .A(
        n16752), .B(n16751), .ZN(n16756) );
  INV_X1 U18856 ( .A(n22201), .ZN(n16754) );
  NAND2_X1 U18857 ( .A1(n16754), .A2(n22037), .ZN(n16755) );
  OAI211_X1 U18858 ( .C1(n16757), .C2(n22033), .A(n16756), .B(n16755), .ZN(
        P1_U3007) );
  NAND2_X1 U18859 ( .A1(n11183), .A2(n16758), .ZN(n16759) );
  NAND2_X1 U18860 ( .A1(n16760), .A2(n16759), .ZN(n22180) );
  INV_X1 U18861 ( .A(n22180), .ZN(n16766) );
  AOI21_X1 U18862 ( .B1(n16762), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16761), .ZN(n16763) );
  OAI21_X1 U18863 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16764), .A(
        n16763), .ZN(n16765) );
  AOI21_X1 U18864 ( .B1(n16766), .B2(n22037), .A(n16765), .ZN(n16767) );
  OAI21_X1 U18865 ( .B1(n16768), .B2(n22033), .A(n16767), .ZN(P1_U3008) );
  NOR2_X1 U18866 ( .A1(n16769), .A2(n22033), .ZN(n16782) );
  INV_X1 U18867 ( .A(n16770), .ZN(n16771) );
  NOR2_X1 U18868 ( .A1(n16784), .A2(n16771), .ZN(n16775) );
  INV_X1 U18869 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16772) );
  AND3_X1 U18870 ( .A1(n21999), .A2(n16775), .A3(n16772), .ZN(n22041) );
  NOR2_X1 U18871 ( .A1(n15989), .A2(n16773), .ZN(n16774) );
  OR2_X1 U18872 ( .A1(n16546), .A2(n16774), .ZN(n22169) );
  INV_X1 U18873 ( .A(n16775), .ZN(n16777) );
  OAI21_X1 U18874 ( .B1(n16783), .B2(n16777), .A(n16776), .ZN(n16778) );
  INV_X1 U18875 ( .A(n16778), .ZN(n22042) );
  AOI21_X1 U18876 ( .B1(n22042), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16779), .ZN(n16780) );
  OAI21_X1 U18877 ( .B1(n22169), .B2(n22017), .A(n16780), .ZN(n16781) );
  OR3_X1 U18878 ( .A1(n16782), .A2(n22041), .A3(n16781), .ZN(P1_U3010) );
  NOR2_X1 U18879 ( .A1(n21987), .A2(n16784), .ZN(n22044) );
  INV_X1 U18880 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16799) );
  NOR2_X1 U18881 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16799), .ZN(
        n16787) );
  AOI21_X1 U18882 ( .B1(n21985), .B2(n16784), .A(n16783), .ZN(n16798) );
  NAND2_X1 U18883 ( .A1(n22044), .A2(n16799), .ZN(n16797) );
  AOI21_X1 U18884 ( .B1(n16798), .B2(n16797), .A(n16785), .ZN(n16786) );
  AOI21_X1 U18885 ( .B1(n22044), .B2(n16787), .A(n16786), .ZN(n16790) );
  INV_X1 U18886 ( .A(n16788), .ZN(n16789) );
  OAI211_X1 U18887 ( .C1(n22163), .C2(n22017), .A(n16790), .B(n16789), .ZN(
        n16791) );
  INV_X1 U18888 ( .A(n16791), .ZN(n16792) );
  OAI21_X1 U18889 ( .B1(n16793), .B2(n22033), .A(n16792), .ZN(P1_U3011) );
  XNOR2_X1 U18890 ( .A(n16794), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16795) );
  XNOR2_X1 U18891 ( .A(n16796), .B(n16795), .ZN(n20630) );
  NAND2_X1 U18892 ( .A1(n20630), .A2(n22038), .ZN(n16802) );
  OAI21_X1 U18893 ( .B1(n16799), .B2(n16798), .A(n16797), .ZN(n16800) );
  AOI21_X1 U18894 ( .B1(n22040), .B2(P1_REIP_REG_19__SCAN_IN), .A(n16800), 
        .ZN(n16801) );
  OAI211_X1 U18895 ( .C1(n22017), .C2(n22150), .A(n16802), .B(n16801), .ZN(
        P1_U3012) );
  NOR2_X1 U18896 ( .A1(n16803), .A2(n22209), .ZN(n22218) );
  AOI21_X1 U18897 ( .B1(n16804), .B2(n16811), .A(n22218), .ZN(n16805) );
  OAI21_X1 U18898 ( .B1(n12075), .B2(n22465), .A(n16805), .ZN(n16806) );
  MUX2_X1 U18899 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16806), .S(
        n17728), .Z(P1_U3478) );
  OAI211_X1 U18900 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n16807), .A(n22418), 
        .B(n22417), .ZN(n16808) );
  OAI21_X1 U18901 ( .B1(n16809), .B2(n14933), .A(n16808), .ZN(n16810) );
  MUX2_X1 U18902 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16810), .S(
        n17728), .Z(P1_U3477) );
  NAND2_X1 U18903 ( .A1(n16842), .A2(n16811), .ZN(n16812) );
  OAI211_X1 U18904 ( .C1(n16814), .C2(n14759), .A(n16813), .B(n16812), .ZN(
        n16815) );
  MUX2_X1 U18905 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16815), .S(
        n17728), .Z(P1_U3475) );
  INV_X1 U18906 ( .A(n16836), .ZN(n16817) );
  NOR3_X1 U18907 ( .A1(n11422), .A2(n14304), .A3(n14473), .ZN(n16816) );
  AOI211_X1 U18908 ( .C1(n22468), .C2(n16841), .A(n16817), .B(n16816), .ZN(
        n17701) );
  NOR3_X1 U18909 ( .A1(n14473), .A2(n14304), .A3(n16845), .ZN(n16818) );
  AOI21_X1 U18910 ( .B1(n16820), .B2(n16819), .A(n16818), .ZN(n16821) );
  OAI21_X1 U18911 ( .B1(n17701), .B2(n16846), .A(n16821), .ZN(n16822) );
  MUX2_X1 U18912 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16822), .S(
        n17650), .Z(P1_U3473) );
  AOI21_X1 U18913 ( .B1(n14304), .B2(n17687), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16823) );
  NOR2_X1 U18914 ( .A1(n16824), .A2(n16823), .ZN(n16843) );
  NAND3_X1 U18915 ( .A1(n16826), .A2(n16825), .A3(n16843), .ZN(n16839) );
  NOR3_X1 U18916 ( .A1(n16829), .A2(n14304), .A3(n17687), .ZN(n16827) );
  AOI21_X1 U18917 ( .B1(n16828), .B2(n16834), .A(n16827), .ZN(n16838) );
  AND2_X1 U18918 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n17687), .ZN(
        n16833) );
  INV_X1 U18919 ( .A(n14304), .ZN(n16830) );
  NAND2_X1 U18920 ( .A1(n16830), .A2(n16829), .ZN(n16831) );
  AOI22_X1 U18921 ( .A1(n16834), .A2(n16833), .B1(n16832), .B2(n16831), .ZN(
        n16835) );
  MUX2_X1 U18922 ( .A(n16836), .B(n16835), .S(n17685), .Z(n16837) );
  NAND3_X1 U18923 ( .A1(n16839), .A2(n16838), .A3(n16837), .ZN(n16840) );
  AOI21_X1 U18924 ( .B1(n16842), .B2(n16841), .A(n16840), .ZN(n17684) );
  INV_X1 U18925 ( .A(n16843), .ZN(n16844) );
  OAI22_X1 U18926 ( .A1(n17684), .A2(n16846), .B1(n16845), .B2(n16844), .ZN(
        n16847) );
  MUX2_X1 U18927 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16847), .S(
        n17650), .Z(P1_U3469) );
  INV_X1 U18928 ( .A(n16848), .ZN(n16861) );
  NOR2_X2 U18929 ( .A1(n19230), .A2(n19054), .ZN(n18937) );
  INV_X1 U18930 ( .A(n18937), .ZN(n16948) );
  INV_X1 U18931 ( .A(n17222), .ZN(n16850) );
  NOR2_X1 U18932 ( .A1(n16850), .A2(n16849), .ZN(n19053) );
  AOI21_X1 U18933 ( .B1(n19062), .B2(n16852), .A(n16851), .ZN(n19058) );
  INV_X1 U18934 ( .A(n19058), .ZN(n16853) );
  NAND2_X1 U18935 ( .A1(n19053), .A2(n16853), .ZN(n16863) );
  NOR3_X1 U18936 ( .A1(n16854), .A2(n16948), .A3(n16863), .ZN(n16857) );
  INV_X1 U18937 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16855) );
  OAI22_X1 U18938 ( .A1(n16855), .A2(n19007), .B1(n17938), .B2(n19059), .ZN(
        n16856) );
  AOI211_X1 U18939 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19028), .A(
        n16857), .B(n16856), .ZN(n16860) );
  INV_X1 U18940 ( .A(n16858), .ZN(n17068) );
  AOI22_X1 U18941 ( .A1(n17068), .A2(n19067), .B1(n18916), .B2(n19707), .ZN(
        n16859) );
  OAI211_X1 U18942 ( .C1(n16861), .C2(n18996), .A(n16860), .B(n16859), .ZN(
        P2_U2824) );
  INV_X1 U18943 ( .A(n16862), .ZN(n16874) );
  NAND2_X1 U18944 ( .A1(n11223), .A2(n16863), .ZN(n16865) );
  OAI21_X1 U18945 ( .B1(n16866), .B2(n16865), .A(n19055), .ZN(n16864) );
  AOI21_X1 U18946 ( .B1(n16866), .B2(n16865), .A(n16864), .ZN(n16869) );
  AOI22_X1 U18947 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n11144), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19009), .ZN(n16867) );
  INV_X1 U18948 ( .A(n16867), .ZN(n16868) );
  AOI211_X1 U18949 ( .C1(n19028), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16869), .B(n16868), .ZN(n16873) );
  INV_X1 U18950 ( .A(n16373), .ZN(n16871) );
  AOI22_X1 U18951 ( .A1(n16871), .A2(n19067), .B1(n18916), .B2(n11201), .ZN(
        n16872) );
  OAI211_X1 U18952 ( .C1(n16874), .C2(n18996), .A(n16873), .B(n16872), .ZN(
        P2_U2825) );
  NOR2_X1 U18953 ( .A1(n19054), .A2(n16875), .ZN(n16877) );
  OAI21_X1 U18954 ( .B1(n17233), .B2(n16877), .A(n19055), .ZN(n16876) );
  AOI21_X1 U18955 ( .B1(n17233), .B2(n16877), .A(n16876), .ZN(n16878) );
  INV_X1 U18956 ( .A(n16878), .ZN(n16892) );
  NOR2_X1 U18957 ( .A1(n16899), .A2(n16879), .ZN(n16880) );
  OR2_X1 U18958 ( .A1(n16881), .A2(n16880), .ZN(n17236) );
  INV_X1 U18959 ( .A(n17236), .ZN(n17367) );
  NAND2_X1 U18960 ( .A1(n16882), .A2(n16883), .ZN(n16884) );
  INV_X1 U18961 ( .A(n17366), .ZN(n16889) );
  OAI22_X1 U18962 ( .A1(n16886), .A2(n19061), .B1(n17935), .B2(n19059), .ZN(
        n16887) );
  AOI21_X1 U18963 ( .B1(n11144), .B2(P2_EBX_REG_27__SCAN_IN), .A(n16887), .ZN(
        n16888) );
  OAI21_X1 U18964 ( .B1(n19072), .B2(n16889), .A(n16888), .ZN(n16890) );
  AOI21_X1 U18965 ( .B1(n17367), .B2(n19067), .A(n16890), .ZN(n16891) );
  OAI211_X1 U18966 ( .C1(n18996), .C2(n16893), .A(n16892), .B(n16891), .ZN(
        P2_U2828) );
  NAND2_X1 U18967 ( .A1(n11223), .A2(n16894), .ZN(n16896) );
  OAI21_X1 U18968 ( .B1(n16897), .B2(n16896), .A(n19055), .ZN(n16895) );
  AOI21_X1 U18969 ( .B1(n16897), .B2(n16896), .A(n16895), .ZN(n16898) );
  INV_X1 U18970 ( .A(n16898), .ZN(n16909) );
  INV_X1 U18971 ( .A(n16899), .ZN(n16902) );
  NAND2_X1 U18972 ( .A1(n17090), .A2(n16900), .ZN(n16901) );
  NAND2_X1 U18973 ( .A1(n16902), .A2(n16901), .ZN(n17248) );
  INV_X1 U18974 ( .A(n17248), .ZN(n17379) );
  OAI21_X1 U18975 ( .B1(n17155), .B2(n16903), .A(n16882), .ZN(n17381) );
  OAI22_X1 U18976 ( .A1(n16904), .A2(n19007), .B1(n19072), .B2(n17381), .ZN(
        n16907) );
  AOI22_X1 U18977 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19009), .ZN(n16905) );
  INV_X1 U18978 ( .A(n16905), .ZN(n16906) );
  AOI211_X1 U18979 ( .C1(n19067), .C2(n17379), .A(n16907), .B(n16906), .ZN(
        n16908) );
  OAI211_X1 U18980 ( .C1(n16910), .C2(n18996), .A(n16909), .B(n16908), .ZN(
        P2_U2829) );
  INV_X1 U18981 ( .A(n16911), .ZN(n16928) );
  NAND2_X1 U18982 ( .A1(n11223), .A2(n16912), .ZN(n16914) );
  OAI21_X1 U18983 ( .B1(n17826), .B2(n16914), .A(n19055), .ZN(n16913) );
  AOI21_X1 U18984 ( .B1(n17826), .B2(n16914), .A(n16913), .ZN(n16915) );
  INV_X1 U18985 ( .A(n16915), .ZN(n16927) );
  OR2_X1 U18986 ( .A1(n16916), .A2(n16934), .ZN(n16917) );
  NAND2_X1 U18987 ( .A1(n17088), .A2(n16917), .ZN(n19110) );
  INV_X1 U18988 ( .A(n19110), .ZN(n16925) );
  INV_X1 U18989 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16921) );
  NAND2_X1 U18990 ( .A1(n16937), .A2(n16938), .ZN(n16939) );
  INV_X1 U18991 ( .A(n16939), .ZN(n16918) );
  NOR2_X1 U18992 ( .A1(n16919), .A2(n16918), .ZN(n16920) );
  OAI22_X1 U18993 ( .A1(n16921), .A2(n19007), .B1(n19072), .B2(n19103), .ZN(
        n16924) );
  AOI22_X1 U18994 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19009), .ZN(n16922) );
  INV_X1 U18995 ( .A(n16922), .ZN(n16923) );
  AOI211_X1 U18996 ( .C1(n19067), .C2(n16925), .A(n16924), .B(n16923), .ZN(
        n16926) );
  OAI211_X1 U18997 ( .C1(n16928), .C2(n18996), .A(n16927), .B(n16926), .ZN(
        P2_U2831) );
  NOR2_X1 U18998 ( .A1(n19054), .A2(n16929), .ZN(n16931) );
  OAI21_X1 U18999 ( .B1(n16932), .B2(n16931), .A(n19055), .ZN(n16930) );
  AOI21_X1 U19000 ( .B1(n16932), .B2(n16931), .A(n16930), .ZN(n16933) );
  INV_X1 U19001 ( .A(n16933), .ZN(n16945) );
  AOI21_X1 U19002 ( .B1(n16936), .B2(n16935), .A(n16934), .ZN(n17404) );
  INV_X1 U19003 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16941) );
  OR2_X1 U19004 ( .A1(n16938), .A2(n16937), .ZN(n16940) );
  NAND2_X1 U19005 ( .A1(n16940), .A2(n16939), .ZN(n17407) );
  OAI22_X1 U19006 ( .A1(n16941), .A2(n19007), .B1(n19072), .B2(n17407), .ZN(
        n16943) );
  OAI22_X1 U19007 ( .A1(n17271), .A2(n19061), .B1(n17933), .B2(n19059), .ZN(
        n16942) );
  AOI211_X1 U19008 ( .C1(n19067), .C2(n17404), .A(n16943), .B(n16942), .ZN(
        n16944) );
  OAI211_X1 U19009 ( .C1(n18996), .C2(n16946), .A(n16945), .B(n16944), .ZN(
        P2_U2832) );
  INV_X1 U19010 ( .A(n16947), .ZN(n16958) );
  NAND2_X1 U19011 ( .A1(n19055), .A2(n19054), .ZN(n18926) );
  AOI21_X1 U19012 ( .B1(n16951), .B2(n18932), .A(n16950), .ZN(n16957) );
  INV_X1 U19013 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16954) );
  NAND2_X1 U19014 ( .A1(n18916), .A2(n20069), .ZN(n16953) );
  AOI22_X1 U19015 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n11144), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19009), .ZN(n16952) );
  OAI211_X1 U19016 ( .C1(n19061), .C2(n16954), .A(n16953), .B(n16952), .ZN(
        n16955) );
  AOI21_X1 U19017 ( .B1(n17103), .B2(n19067), .A(n16955), .ZN(n16956) );
  OAI211_X1 U19018 ( .C1(n16958), .C2(n18996), .A(n16957), .B(n16956), .ZN(
        P2_U2835) );
  NAND2_X1 U19019 ( .A1(n11223), .A2(n16959), .ZN(n16960) );
  XOR2_X1 U19020 ( .A(n17787), .B(n16960), .Z(n16970) );
  INV_X1 U19021 ( .A(n19131), .ZN(n16966) );
  INV_X1 U19022 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17788) );
  OAI22_X1 U19023 ( .A1(n17788), .A2(n19061), .B1(n13018), .B2(n19059), .ZN(
        n16961) );
  INV_X1 U19024 ( .A(n16961), .ZN(n16962) );
  NAND2_X1 U19025 ( .A1(n17323), .A2(n16962), .ZN(n16963) );
  AOI21_X1 U19026 ( .B1(n11144), .B2(P2_EBX_REG_16__SCAN_IN), .A(n16963), .ZN(
        n16964) );
  OAI21_X1 U19027 ( .B1(n19072), .B2(n19133), .A(n16964), .ZN(n16965) );
  AOI21_X1 U19028 ( .B1(n16966), .B2(n19067), .A(n16965), .ZN(n16967) );
  OAI21_X1 U19029 ( .B1(n16968), .B2(n18996), .A(n16967), .ZN(n16969) );
  AOI21_X1 U19030 ( .B1(n16970), .B2(n19055), .A(n16969), .ZN(n16971) );
  INV_X1 U19031 ( .A(n16971), .ZN(P2_U2839) );
  NAND2_X1 U19032 ( .A1(n11222), .A2(n18921), .ZN(n16972) );
  XOR2_X1 U19033 ( .A(n16973), .B(n16972), .Z(n16974) );
  NAND2_X1 U19034 ( .A1(n16974), .A2(n19055), .ZN(n16983) );
  INV_X1 U19035 ( .A(n16975), .ZN(n16976) );
  XNOR2_X1 U19036 ( .A(n16977), .B(n16976), .ZN(n19721) );
  AOI22_X1 U19037 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19009), .ZN(n16978) );
  NAND2_X1 U19038 ( .A1(n18958), .A2(n16978), .ZN(n16979) );
  AOI21_X1 U19039 ( .B1(n11144), .B2(P2_EBX_REG_12__SCAN_IN), .A(n16979), .ZN(
        n16980) );
  OAI21_X1 U19040 ( .B1(n19072), .B2(n19721), .A(n16980), .ZN(n16981) );
  AOI21_X1 U19041 ( .B1(n17520), .B2(n19067), .A(n16981), .ZN(n16982) );
  OAI211_X1 U19042 ( .C1(n18996), .C2(n16984), .A(n16983), .B(n16982), .ZN(
        P2_U2843) );
  NOR2_X1 U19043 ( .A1(n19054), .A2(n16985), .ZN(n16986) );
  XNOR2_X1 U19044 ( .A(n16986), .B(n17334), .ZN(n16987) );
  NAND2_X1 U19045 ( .A1(n16987), .A2(n19055), .ZN(n16995) );
  AOI22_X1 U19046 ( .A1(n16988), .A2(n19068), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19028), .ZN(n16989) );
  OAI211_X1 U19047 ( .C1(n13105), .C2(n19007), .A(n16989), .B(n17323), .ZN(
        n16990) );
  AOI21_X1 U19048 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n19009), .A(n16990), .ZN(
        n16994) );
  XNOR2_X1 U19049 ( .A(n16991), .B(n11200), .ZN(n19730) );
  INV_X1 U19050 ( .A(n19730), .ZN(n16992) );
  AOI22_X1 U19051 ( .A1(n17569), .A2(n19067), .B1(n18916), .B2(n16992), .ZN(
        n16993) );
  NAND3_X1 U19052 ( .A1(n16995), .A2(n16994), .A3(n16993), .ZN(P2_U2846) );
  NAND2_X1 U19053 ( .A1(n11223), .A2(n16996), .ZN(n16997) );
  XNOR2_X1 U19054 ( .A(n17740), .B(n16997), .ZN(n16998) );
  NAND2_X1 U19055 ( .A1(n16998), .A2(n19055), .ZN(n17012) );
  INV_X1 U19056 ( .A(n16999), .ZN(n17000) );
  OR2_X1 U19057 ( .A1(n17001), .A2(n17000), .ZN(n17004) );
  INV_X1 U19058 ( .A(n11200), .ZN(n17003) );
  AND2_X1 U19059 ( .A1(n17004), .A2(n17003), .ZN(n19731) );
  NAND2_X1 U19060 ( .A1(n18916), .A2(n19731), .ZN(n17005) );
  OAI211_X1 U19061 ( .C1(n17006), .C2(n19007), .A(n17005), .B(n17323), .ZN(
        n17010) );
  AOI22_X1 U19062 ( .A1(n17007), .A2(n19068), .B1(n19009), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n17008) );
  OAI21_X1 U19063 ( .B1(n17751), .B2(n19061), .A(n17008), .ZN(n17009) );
  AOI211_X1 U19064 ( .C1(n19067), .C2(n19158), .A(n17010), .B(n17009), .ZN(
        n17011) );
  NAND2_X1 U19065 ( .A1(n17012), .A2(n17011), .ZN(P2_U2847) );
  NOR2_X1 U19066 ( .A1(n19054), .A2(n17013), .ZN(n17014) );
  XNOR2_X1 U19067 ( .A(n17739), .B(n17014), .ZN(n17015) );
  NAND2_X1 U19068 ( .A1(n17015), .A2(n19055), .ZN(n17021) );
  NOR2_X1 U19069 ( .A1(n18996), .A2(n17016), .ZN(n17019) );
  AOI22_X1 U19070 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19009), .ZN(n17017) );
  OAI211_X1 U19071 ( .C1(n19007), .C2(n13073), .A(n17017), .B(n17323), .ZN(
        n17018) );
  AOI211_X1 U19072 ( .C1(n17736), .C2(n19067), .A(n17019), .B(n17018), .ZN(
        n17020) );
  OAI211_X1 U19073 ( .C1(n20022), .C2(n19072), .A(n17021), .B(n17020), .ZN(
        P2_U2850) );
  AND2_X1 U19074 ( .A1(n11223), .A2(n17022), .ZN(n17024) );
  AOI21_X1 U19075 ( .B1(n17025), .B2(n17024), .A(n19230), .ZN(n17023) );
  OAI21_X1 U19076 ( .B1(n17025), .B2(n17024), .A(n17023), .ZN(n17034) );
  AOI22_X1 U19077 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n11144), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19009), .ZN(n17026) );
  OAI211_X1 U19078 ( .C1(n19061), .C2(n17027), .A(n17323), .B(n17026), .ZN(
        n17028) );
  AOI21_X1 U19079 ( .B1(n18916), .B2(n20074), .A(n17028), .ZN(n17029) );
  OAI21_X1 U19080 ( .B1(n17030), .B2(n18996), .A(n17029), .ZN(n17031) );
  AOI21_X1 U19081 ( .B1(n17032), .B2(n19067), .A(n17031), .ZN(n17033) );
  OAI211_X1 U19082 ( .C1(n17067), .C2(n20076), .A(n17034), .B(n17033), .ZN(
        P2_U2851) );
  NOR2_X1 U19083 ( .A1(n19054), .A2(n17035), .ZN(n17037) );
  XNOR2_X1 U19084 ( .A(n17037), .B(n17036), .ZN(n17038) );
  NAND2_X1 U19085 ( .A1(n17038), .A2(n19055), .ZN(n17045) );
  OAI22_X1 U19086 ( .A1(n13048), .A2(n19007), .B1(n14886), .B2(n19059), .ZN(
        n17039) );
  AOI21_X1 U19087 ( .B1(n19028), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n17039), .ZN(n17040) );
  OAI21_X1 U19088 ( .B1(n18996), .B2(n17041), .A(n17040), .ZN(n17043) );
  NOR2_X1 U19089 ( .A1(n20017), .A2(n19072), .ZN(n17042) );
  AOI211_X1 U19090 ( .C1(n19067), .C2(n12643), .A(n17043), .B(n17042), .ZN(
        n17044) );
  OAI211_X1 U19091 ( .C1(n20018), .C2(n17067), .A(n17045), .B(n17044), .ZN(
        P2_U2852) );
  NAND2_X1 U19092 ( .A1(n11222), .A2(n17046), .ZN(n17057) );
  XNOR2_X1 U19093 ( .A(n17047), .B(n17057), .ZN(n17048) );
  NAND2_X1 U19094 ( .A1(n17048), .A2(n19055), .ZN(n17056) );
  NAND2_X1 U19095 ( .A1(n20012), .A2(n18916), .ZN(n17051) );
  OAI22_X1 U19096 ( .A1(n13044), .A2(n19007), .B1(n14369), .B2(n19059), .ZN(
        n17049) );
  AOI21_X1 U19097 ( .B1(n19028), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17049), .ZN(n17050) );
  OAI211_X1 U19098 ( .C1(n18996), .C2(n17052), .A(n17051), .B(n17050), .ZN(
        n17053) );
  AOI21_X1 U19099 ( .B1(n17054), .B2(n19067), .A(n17053), .ZN(n17055) );
  OAI211_X1 U19100 ( .C1(n17067), .C2(n20015), .A(n17056), .B(n17055), .ZN(
        P2_U2853) );
  AOI21_X1 U19101 ( .B1(n18870), .B2(n17058), .A(n17057), .ZN(n17623) );
  AOI22_X1 U19102 ( .A1(n17623), .A2(n19055), .B1(n18932), .B2(n17059), .ZN(
        n17066) );
  AOI22_X1 U19103 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19009), .ZN(n17061) );
  NAND2_X1 U19104 ( .A1(n11144), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n17060) );
  OAI211_X1 U19105 ( .C1(n19072), .C2(n17589), .A(n17061), .B(n17060), .ZN(
        n17063) );
  NOR2_X1 U19106 ( .A1(n17621), .A2(n19011), .ZN(n17062) );
  AOI211_X1 U19107 ( .C1(n19068), .C2(n17064), .A(n17063), .B(n17062), .ZN(
        n17065) );
  OAI211_X1 U19108 ( .C1(n19814), .C2(n17067), .A(n17066), .B(n17065), .ZN(
        P2_U2854) );
  MUX2_X1 U19109 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n17068), .S(n17125), .Z(
        P2_U2856) );
  NAND2_X1 U19110 ( .A1(n11213), .A2(n17070), .ZN(n17072) );
  XNOR2_X1 U19111 ( .A(n17072), .B(n17071), .ZN(n17142) );
  NOR2_X1 U19112 ( .A1(n17358), .A2(n11164), .ZN(n17073) );
  AOI21_X1 U19113 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n11164), .A(n17073), .ZN(
        n17074) );
  OAI21_X1 U19114 ( .B1(n17142), .B2(n17128), .A(n17074), .ZN(P2_U2859) );
  NAND2_X1 U19115 ( .A1(n11213), .A2(n17075), .ZN(n17076) );
  XOR2_X1 U19116 ( .A(n17077), .B(n17076), .Z(n17146) );
  NOR2_X1 U19117 ( .A1(n17236), .A2(n11163), .ZN(n17078) );
  AOI21_X1 U19118 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n11164), .A(n17078), .ZN(
        n17079) );
  OAI21_X1 U19119 ( .B1(n17146), .B2(n17128), .A(n17079), .ZN(P2_U2860) );
  AOI21_X1 U19120 ( .B1(n17082), .B2(n17081), .A(n17080), .ZN(n17150) );
  NAND2_X1 U19121 ( .A1(n17150), .A2(n17136), .ZN(n17084) );
  NAND2_X1 U19122 ( .A1(n11163), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n17083) );
  OAI211_X1 U19123 ( .C1(n17248), .C2(n11163), .A(n17084), .B(n17083), .ZN(
        P2_U2861) );
  OAI21_X1 U19124 ( .B1(n17087), .B2(n17086), .A(n17085), .ZN(n17160) );
  INV_X1 U19125 ( .A(n17088), .ZN(n17092) );
  INV_X1 U19126 ( .A(n17089), .ZN(n17091) );
  OAI21_X1 U19127 ( .B1(n17092), .B2(n17091), .A(n17090), .ZN(n19047) );
  INV_X1 U19128 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n17093) );
  MUX2_X1 U19129 ( .A(n19047), .B(n17093), .S(n11164), .Z(n17094) );
  OAI21_X1 U19130 ( .B1(n17160), .B2(n17128), .A(n17094), .ZN(P2_U2862) );
  OAI21_X1 U19131 ( .B1(n17097), .B2(n17096), .A(n11214), .ZN(n17165) );
  NOR2_X1 U19132 ( .A1(n11164), .A2(n19110), .ZN(n17098) );
  AOI21_X1 U19133 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n11163), .A(n17098), .ZN(
        n17099) );
  OAI21_X1 U19134 ( .B1(n17165), .B2(n17128), .A(n17099), .ZN(P2_U2863) );
  XNOR2_X1 U19135 ( .A(n15811), .B(n17100), .ZN(n17170) );
  NAND2_X1 U19136 ( .A1(n11163), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n17102) );
  NAND2_X1 U19137 ( .A1(n17125), .A2(n17404), .ZN(n17101) );
  OAI211_X1 U19138 ( .C1(n17170), .C2(n17128), .A(n17102), .B(n17101), .ZN(
        P2_U2864) );
  INV_X1 U19139 ( .A(n17103), .ZN(n17110) );
  NOR2_X1 U19140 ( .A1(n17134), .A2(n17104), .ZN(n17114) );
  INV_X1 U19141 ( .A(n17114), .ZN(n17106) );
  AOI21_X1 U19142 ( .B1(n17107), .B2(n17106), .A(n17105), .ZN(n20070) );
  NAND2_X1 U19143 ( .A1(n20070), .A2(n17136), .ZN(n17109) );
  NAND2_X1 U19144 ( .A1(n11164), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n17108) );
  OAI211_X1 U19145 ( .C1(n17110), .C2(n11164), .A(n17109), .B(n17108), .ZN(
        P2_U2867) );
  NOR2_X1 U19146 ( .A1(n17111), .A2(n17122), .ZN(n17112) );
  OR2_X1 U19147 ( .A1(n13034), .A2(n17112), .ZN(n19000) );
  OR2_X1 U19148 ( .A1(n17134), .A2(n17113), .ZN(n17120) );
  AOI21_X1 U19149 ( .B1(n17115), .B2(n17120), .A(n17114), .ZN(n17185) );
  NAND2_X1 U19150 ( .A1(n17185), .A2(n17136), .ZN(n17117) );
  NAND2_X1 U19151 ( .A1(n11164), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n17116) );
  OAI211_X1 U19152 ( .C1(n19000), .C2(n11163), .A(n17117), .B(n17116), .ZN(
        P2_U2868) );
  NAND2_X1 U19153 ( .A1(n17132), .A2(n17118), .ZN(n17119) );
  NAND2_X1 U19154 ( .A1(n17120), .A2(n17119), .ZN(n20173) );
  OR2_X1 U19155 ( .A1(n17131), .A2(n17121), .ZN(n17124) );
  INV_X1 U19156 ( .A(n17122), .ZN(n17123) );
  AND2_X1 U19157 ( .A1(n17124), .A2(n17123), .ZN(n19148) );
  NAND2_X1 U19158 ( .A1(n19148), .A2(n17125), .ZN(n17127) );
  NAND2_X1 U19159 ( .A1(n11164), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U19160 ( .C1(n20173), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        P2_U2869) );
  AND2_X1 U19161 ( .A1(n15716), .A2(n17129), .ZN(n17130) );
  OR2_X1 U19162 ( .A1(n17131), .A2(n17130), .ZN(n18973) );
  INV_X1 U19163 ( .A(n17132), .ZN(n17133) );
  AOI21_X1 U19164 ( .B1(n17135), .B2(n17134), .A(n17133), .ZN(n17195) );
  NAND2_X1 U19165 ( .A1(n17195), .A2(n17136), .ZN(n17138) );
  NAND2_X1 U19166 ( .A1(n11163), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n17137) );
  OAI211_X1 U19167 ( .C1(n18973), .C2(n11164), .A(n17138), .B(n17137), .ZN(
        P2_U2870) );
  INV_X1 U19168 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n17909) );
  OAI22_X1 U19169 ( .A1(n20067), .A2(n19719), .B1(n20066), .B2(n17909), .ZN(
        n17139) );
  AOI21_X1 U19170 ( .B1(n17355), .B2(n20277), .A(n17139), .ZN(n17141) );
  AOI22_X1 U19171 ( .A1(n20169), .A2(BUF1_REG_28__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n17140) );
  OAI211_X1 U19172 ( .C1(n17142), .C2(n20222), .A(n17141), .B(n17140), .ZN(
        P2_U2891) );
  INV_X1 U19173 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n17907) );
  OAI22_X1 U19174 ( .A1(n20067), .A2(n19722), .B1(n20066), .B2(n17907), .ZN(
        n17143) );
  AOI21_X1 U19175 ( .B1(n20277), .B2(n17366), .A(n17143), .ZN(n17145) );
  AOI22_X1 U19176 ( .A1(n20169), .A2(BUF1_REG_27__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n17144) );
  OAI211_X1 U19177 ( .C1(n17146), .C2(n20222), .A(n17145), .B(n17144), .ZN(
        P2_U2892) );
  AOI22_X1 U19178 ( .A1(n20169), .A2(BUF1_REG_26__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U19179 ( .A1(n20168), .A2(n19725), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20276), .ZN(n17147) );
  OAI211_X1 U19180 ( .C1(n20172), .C2(n17381), .A(n17148), .B(n17147), .ZN(
        n17149) );
  AOI21_X1 U19181 ( .B1(n17150), .B2(n20279), .A(n17149), .ZN(n17151) );
  INV_X1 U19182 ( .A(n17151), .ZN(P2_U2893) );
  NOR2_X1 U19183 ( .A1(n17153), .A2(n17152), .ZN(n17154) );
  OR2_X1 U19184 ( .A1(n17155), .A2(n17154), .ZN(n19052) );
  INV_X1 U19185 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n17903) );
  OAI22_X1 U19186 ( .A1(n20172), .A2(n19052), .B1(n17903), .B2(n20066), .ZN(
        n17156) );
  AOI21_X1 U19187 ( .B1(n20168), .B2(n17157), .A(n17156), .ZN(n17159) );
  AOI22_X1 U19188 ( .A1(n20169), .A2(BUF1_REG_25__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n17158) );
  OAI211_X1 U19189 ( .C1(n17160), .C2(n20222), .A(n17159), .B(n17158), .ZN(
        P2_U2894) );
  INV_X1 U19190 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n17900) );
  OAI22_X1 U19191 ( .A1(n20172), .A2(n19103), .B1(n20066), .B2(n17900), .ZN(
        n17161) );
  AOI21_X1 U19192 ( .B1(n20168), .B2(n17162), .A(n17161), .ZN(n17164) );
  AOI22_X1 U19193 ( .A1(n20169), .A2(BUF1_REG_24__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n17163) );
  OAI211_X1 U19194 ( .C1(n17165), .C2(n20222), .A(n17164), .B(n17163), .ZN(
        P2_U2895) );
  INV_X1 U19195 ( .A(n17407), .ZN(n17167) );
  INV_X1 U19196 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17898) );
  OAI22_X1 U19197 ( .A1(n20067), .A2(n19741), .B1(n20066), .B2(n17898), .ZN(
        n17166) );
  AOI21_X1 U19198 ( .B1(n20277), .B2(n17167), .A(n17166), .ZN(n17169) );
  AOI22_X1 U19199 ( .A1(n20169), .A2(BUF1_REG_23__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n17168) );
  OAI211_X1 U19200 ( .C1(n17170), .C2(n20222), .A(n17169), .B(n17168), .ZN(
        P2_U2896) );
  XNOR2_X1 U19201 ( .A(n17172), .B(n17179), .ZN(n19038) );
  INV_X1 U19202 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n17896) );
  OAI22_X1 U19203 ( .A1(n20172), .A2(n19038), .B1(n20066), .B2(n17896), .ZN(
        n17173) );
  AOI21_X1 U19204 ( .B1(n20168), .B2(n17174), .A(n17173), .ZN(n17176) );
  AOI22_X1 U19205 ( .A1(n20169), .A2(BUF1_REG_22__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n17175) );
  OAI211_X1 U19206 ( .C1(n17177), .C2(n20222), .A(n17176), .B(n17175), .ZN(
        P2_U2897) );
  OR2_X1 U19207 ( .A1(n17178), .A2(n13970), .ZN(n17180) );
  NAND2_X1 U19208 ( .A1(n17180), .A2(n17179), .ZN(n19022) );
  INV_X1 U19209 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n17894) );
  OAI22_X1 U19210 ( .A1(n20172), .A2(n19022), .B1(n20066), .B2(n17894), .ZN(
        n17181) );
  AOI21_X1 U19211 ( .B1(n20168), .B2(n20024), .A(n17181), .ZN(n17183) );
  AOI22_X1 U19212 ( .A1(n20169), .A2(BUF1_REG_21__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n17182) );
  OAI211_X1 U19213 ( .C1(n17184), .C2(n20222), .A(n17183), .B(n17182), .ZN(
        P2_U2898) );
  INV_X1 U19214 ( .A(n17185), .ZN(n17194) );
  OR2_X1 U19215 ( .A1(n17187), .A2(n17186), .ZN(n17189) );
  NAND2_X1 U19216 ( .A1(n17189), .A2(n17188), .ZN(n18999) );
  INV_X1 U19217 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n17891) );
  OAI22_X1 U19218 ( .A1(n20172), .A2(n18999), .B1(n20066), .B2(n17891), .ZN(
        n17190) );
  AOI21_X1 U19219 ( .B1(n20168), .B2(n17191), .A(n17190), .ZN(n17193) );
  AOI22_X1 U19220 ( .A1(n20169), .A2(BUF1_REG_19__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n17192) );
  OAI211_X1 U19221 ( .C1(n17194), .C2(n20222), .A(n17193), .B(n17192), .ZN(
        P2_U2900) );
  INV_X1 U19222 ( .A(n17195), .ZN(n17203) );
  XNOR2_X1 U19223 ( .A(n17198), .B(n17197), .ZN(n18972) );
  INV_X1 U19224 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n17887) );
  OAI22_X1 U19225 ( .A1(n20172), .A2(n18972), .B1(n20066), .B2(n17887), .ZN(
        n17199) );
  AOI21_X1 U19226 ( .B1(n20168), .B2(n17200), .A(n17199), .ZN(n17202) );
  AOI22_X1 U19227 ( .A1(n20169), .A2(BUF1_REG_17__SCAN_IN), .B1(n20170), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n17201) );
  OAI211_X1 U19228 ( .C1(n17203), .C2(n20222), .A(n17202), .B(n17201), .ZN(
        P2_U2902) );
  NAND2_X1 U19229 ( .A1(n19058), .A2(n17777), .ZN(n17206) );
  AOI21_X1 U19230 ( .B1(n17814), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17204), .ZN(n17205) );
  OAI211_X1 U19231 ( .C1(n13199), .C2(n17207), .A(n17206), .B(n17205), .ZN(
        n17208) );
  AOI21_X1 U19232 ( .B1(n17209), .B2(n17321), .A(n17208), .ZN(n17210) );
  OAI21_X1 U19233 ( .B1(n17211), .B2(n13196), .A(n17210), .ZN(P2_U2985) );
  NAND3_X1 U19234 ( .A1(n17212), .A2(n17213), .A3(n17259), .ZN(n17214) );
  NAND2_X1 U19235 ( .A1(n17214), .A2(n16204), .ZN(n17226) );
  NAND2_X1 U19236 ( .A1(n17226), .A2(n17230), .ZN(n17225) );
  NAND2_X1 U19237 ( .A1(n17244), .A2(n17215), .ZN(n17227) );
  NAND2_X1 U19238 ( .A1(n17225), .A2(n17227), .ZN(n17218) );
  XNOR2_X1 U19239 ( .A(n17216), .B(n17353), .ZN(n17217) );
  XNOR2_X1 U19240 ( .A(n17218), .B(n17217), .ZN(n17363) );
  XNOR2_X1 U19241 ( .A(n17232), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17361) );
  NOR2_X1 U19242 ( .A1(n18958), .A2(n17219), .ZN(n17352) );
  NOR2_X1 U19243 ( .A1(n13199), .A2(n17358), .ZN(n17220) );
  OAI21_X1 U19244 ( .B1(n17222), .B2(n17827), .A(n17221), .ZN(n17223) );
  AOI21_X1 U19245 ( .B1(n17361), .B2(n17321), .A(n17223), .ZN(n17224) );
  OAI21_X1 U19246 ( .B1(n17363), .B2(n13196), .A(n17224), .ZN(P2_U2986) );
  INV_X1 U19247 ( .A(n17225), .ZN(n17229) );
  AOI21_X1 U19248 ( .B1(n17226), .B2(n17227), .A(n17230), .ZN(n17228) );
  OAI22_X1 U19249 ( .A1(n17229), .A2(n17228), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17227), .ZN(n17375) );
  NAND2_X1 U19250 ( .A1(n17249), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17250) );
  NAND2_X1 U19251 ( .A1(n17250), .A2(n17230), .ZN(n17231) );
  AND2_X1 U19252 ( .A1(n17232), .A2(n17231), .ZN(n17373) );
  NAND2_X1 U19253 ( .A1(n17233), .A2(n17777), .ZN(n17235) );
  NOR2_X1 U19254 ( .A1(n17323), .A2(n17935), .ZN(n17365) );
  AOI21_X1 U19255 ( .B1(n17814), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17365), .ZN(n17234) );
  OAI211_X1 U19256 ( .C1(n17236), .C2(n13199), .A(n17235), .B(n17234), .ZN(
        n17237) );
  AOI21_X1 U19257 ( .B1(n17373), .B2(n17321), .A(n17237), .ZN(n17238) );
  OAI21_X1 U19258 ( .B1(n17375), .B2(n13196), .A(n17238), .ZN(P2_U2987) );
  INV_X1 U19259 ( .A(n17258), .ZN(n17241) );
  AOI21_X1 U19260 ( .B1(n17240), .B2(n17259), .A(n17241), .ZN(n17243) );
  MUX2_X1 U19261 ( .A(n17243), .B(n17259), .S(n17242), .Z(n17245) );
  NAND2_X1 U19262 ( .A1(n17245), .A2(n17244), .ZN(n17386) );
  NOR2_X1 U19263 ( .A1(n17323), .A2(n17246), .ZN(n17378) );
  AOI21_X1 U19264 ( .B1(n17814), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17378), .ZN(n17247) );
  OAI21_X1 U19265 ( .B1(n13199), .B2(n17248), .A(n17247), .ZN(n17252) );
  NOR2_X1 U19266 ( .A1(n17382), .A2(n17779), .ZN(n17251) );
  OAI21_X1 U19267 ( .B1(n13196), .B2(n17386), .A(n17254), .ZN(P2_U2988) );
  NOR2_X2 U19268 ( .A1(n17285), .A2(n17255), .ZN(n17819) );
  AOI21_X1 U19269 ( .B1(n17819), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17256) );
  OR2_X1 U19270 ( .A1(n17257), .A2(n17256), .ZN(n17396) );
  NAND2_X1 U19271 ( .A1(n17259), .A2(n17258), .ZN(n17260) );
  XOR2_X1 U19272 ( .A(n17260), .B(n17240), .Z(n17387) );
  NAND2_X1 U19273 ( .A1(n17387), .A2(n17818), .ZN(n17264) );
  OAI22_X1 U19274 ( .A1(n19044), .A2(n17789), .B1(n19043), .B2(n18958), .ZN(
        n17262) );
  NOR2_X1 U19275 ( .A1(n13199), .A2(n19047), .ZN(n17261) );
  AOI211_X1 U19276 ( .C1(n17777), .C2(n19042), .A(n17262), .B(n17261), .ZN(
        n17263) );
  OAI211_X1 U19277 ( .C1(n17779), .C2(n17396), .A(n17264), .B(n17263), .ZN(
        P2_U2989) );
  NAND2_X1 U19278 ( .A1(n17266), .A2(n17265), .ZN(n17268) );
  XOR2_X1 U19279 ( .A(n17268), .B(n17267), .Z(n17410) );
  AOI21_X1 U19280 ( .B1(n17422), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17270) );
  NOR2_X1 U19281 ( .A1(n17270), .A2(n17819), .ZN(n17397) );
  OAI22_X1 U19282 ( .A1(n17271), .A2(n17789), .B1(n17933), .B2(n18958), .ZN(
        n17272) );
  AOI21_X1 U19283 ( .B1(n17807), .B2(n17404), .A(n17272), .ZN(n17273) );
  OAI21_X1 U19284 ( .B1(n17274), .B2(n17827), .A(n17273), .ZN(n17275) );
  AOI21_X1 U19285 ( .B1(n17397), .B2(n17321), .A(n17275), .ZN(n17276) );
  OAI21_X1 U19286 ( .B1(n17410), .B2(n13196), .A(n17276), .ZN(P2_U2991) );
  INV_X1 U19287 ( .A(n11188), .ZN(n17278) );
  NAND2_X1 U19288 ( .A1(n17281), .A2(n17280), .ZN(n17282) );
  XNOR2_X1 U19289 ( .A(n17283), .B(n17282), .ZN(n17435) );
  NOR2_X1 U19290 ( .A1(n17323), .A2(n17931), .ZN(n17428) );
  AOI21_X1 U19291 ( .B1(n17814), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17428), .ZN(n17284) );
  OAI21_X1 U19292 ( .B1(n13199), .B2(n19012), .A(n17284), .ZN(n17288) );
  INV_X1 U19293 ( .A(n17285), .ZN(n17286) );
  NOR2_X1 U19294 ( .A1(n17286), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17423) );
  NOR3_X1 U19295 ( .A1(n17423), .A2(n17422), .A3(n17779), .ZN(n17287) );
  AOI211_X1 U19296 ( .C1(n17777), .C2(n19019), .A(n17288), .B(n17287), .ZN(
        n17289) );
  OAI21_X1 U19297 ( .B1(n17435), .B2(n13196), .A(n17289), .ZN(P2_U2993) );
  NAND2_X1 U19298 ( .A1(n17291), .A2(n17290), .ZN(n17295) );
  INV_X1 U19299 ( .A(n17799), .ZN(n17292) );
  NOR2_X1 U19300 ( .A1(n17293), .A2(n17292), .ZN(n17294) );
  XOR2_X1 U19301 ( .A(n17295), .B(n17294), .Z(n17445) );
  AOI21_X1 U19302 ( .B1(n17437), .B2(n17796), .A(n17296), .ZN(n17436) );
  NAND2_X1 U19303 ( .A1(n17436), .A2(n17321), .ZN(n17302) );
  OAI22_X1 U19304 ( .A1(n17297), .A2(n17789), .B1(n17929), .B2(n18958), .ZN(
        n17299) );
  NOR2_X1 U19305 ( .A1(n13199), .A2(n19000), .ZN(n17298) );
  AOI211_X1 U19306 ( .C1(n17300), .C2(n17777), .A(n17299), .B(n17298), .ZN(
        n17301) );
  OAI211_X1 U19307 ( .C1(n13196), .C2(n17445), .A(n17302), .B(n17301), .ZN(
        P2_U2995) );
  NAND2_X1 U19308 ( .A1(n17304), .A2(n17303), .ZN(n17308) );
  NAND2_X1 U19309 ( .A1(n11189), .A2(n17305), .ZN(n17307) );
  XOR2_X1 U19310 ( .A(n17308), .B(n17307), .Z(n17462) );
  INV_X1 U19311 ( .A(n17792), .ZN(n17310) );
  INV_X1 U19312 ( .A(n17797), .ZN(n17309) );
  OAI211_X1 U19313 ( .C1(n17310), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17321), .B(n17309), .ZN(n17315) );
  INV_X1 U19314 ( .A(n18973), .ZN(n17459) );
  AOI22_X1 U19315 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17814), .B1(
        n17777), .B2(n17311), .ZN(n17312) );
  OAI21_X1 U19316 ( .B1(n17457), .B2(n17323), .A(n17312), .ZN(n17313) );
  AOI21_X1 U19317 ( .B1(n17459), .B2(n17807), .A(n17313), .ZN(n17314) );
  OAI211_X1 U19318 ( .C1(n17462), .C2(n13196), .A(n17315), .B(n17314), .ZN(
        P2_U2997) );
  NOR3_X1 U19319 ( .A1(n17316), .A2(n17331), .A3(n17556), .ZN(n17320) );
  NAND2_X1 U19320 ( .A1(n17318), .A2(n17317), .ZN(n17319) );
  XNOR2_X1 U19321 ( .A(n17320), .B(n17319), .ZN(n17540) );
  AOI21_X1 U19322 ( .B1(n17544), .B2(n17533), .A(n17510), .ZN(n17542) );
  NAND2_X1 U19323 ( .A1(n17542), .A2(n17321), .ZN(n17326) );
  INV_X1 U19324 ( .A(n18918), .ZN(n17537) );
  NOR2_X1 U19325 ( .A1(n17323), .A2(n17322), .ZN(n17531) );
  OAI22_X1 U19326 ( .A1(n18913), .A2(n17789), .B1(n17827), .B2(n18925), .ZN(
        n17324) );
  AOI211_X1 U19327 ( .C1(n17807), .C2(n17537), .A(n17531), .B(n17324), .ZN(
        n17325) );
  OAI211_X1 U19328 ( .C1(n17540), .C2(n13196), .A(n17326), .B(n17325), .ZN(
        P2_U3003) );
  NAND2_X1 U19329 ( .A1(n17329), .A2(n17328), .ZN(n17555) );
  INV_X1 U19330 ( .A(n17331), .ZN(n17554) );
  AND2_X1 U19331 ( .A1(n17554), .A2(n17328), .ZN(n17330) );
  OAI22_X1 U19332 ( .A1(n17555), .A2(n17331), .B1(n17330), .B2(n17329), .ZN(
        n17577) );
  INV_X1 U19333 ( .A(n17332), .ZN(n17565) );
  NAND2_X1 U19334 ( .A1(n17333), .A2(n17573), .ZN(n17564) );
  NAND3_X1 U19335 ( .A1(n17565), .A2(n17820), .A3(n17564), .ZN(n17339) );
  NAND2_X1 U19336 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19142), .ZN(n17567) );
  INV_X1 U19337 ( .A(n17567), .ZN(n17337) );
  INV_X1 U19338 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17335) );
  OAI22_X1 U19339 ( .A1(n17335), .A2(n17789), .B1(n17827), .B2(n17334), .ZN(
        n17336) );
  AOI211_X1 U19340 ( .C1(n17569), .C2(n17807), .A(n17337), .B(n17336), .ZN(
        n17338) );
  OAI211_X1 U19341 ( .C1(n17577), .C2(n13196), .A(n17339), .B(n17338), .ZN(
        P2_U3005) );
  XNOR2_X1 U19342 ( .A(n17341), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17342) );
  XNOR2_X1 U19343 ( .A(n17340), .B(n17342), .ZN(n17588) );
  XOR2_X1 U19344 ( .A(n17345), .B(n17344), .Z(n17586) );
  INV_X1 U19345 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17346) );
  OAI22_X1 U19346 ( .A1(n17346), .A2(n17789), .B1(n17827), .B2(n18888), .ZN(
        n17349) );
  OAI22_X1 U19347 ( .A1(n13199), .A2(n18891), .B1(n18958), .B2(n17347), .ZN(
        n17348) );
  AOI211_X1 U19348 ( .C1(n17586), .C2(n17818), .A(n17349), .B(n17348), .ZN(
        n17350) );
  OAI21_X1 U19349 ( .B1(n17588), .B2(n17779), .A(n17350), .ZN(P2_U3007) );
  NOR3_X1 U19350 ( .A1(n17371), .A2(n17527), .A3(n17353), .ZN(n17360) );
  INV_X1 U19351 ( .A(n17351), .ZN(n17354) );
  AOI21_X1 U19352 ( .B1(n17354), .B2(n17353), .A(n17352), .ZN(n17357) );
  NAND2_X1 U19353 ( .A1(n19154), .A2(n17355), .ZN(n17356) );
  OAI211_X1 U19354 ( .C1(n19130), .C2(n17358), .A(n17357), .B(n17356), .ZN(
        n17359) );
  AOI211_X1 U19355 ( .C1(n17361), .C2(n19157), .A(n17360), .B(n17359), .ZN(
        n17362) );
  OAI21_X1 U19356 ( .B1(n17363), .B2(n19123), .A(n17362), .ZN(P2_U3018) );
  NOR2_X1 U19357 ( .A1(n17364), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17370) );
  AOI21_X1 U19358 ( .B1(n19154), .B2(n17366), .A(n17365), .ZN(n17369) );
  NAND2_X1 U19359 ( .A1(n19159), .A2(n17367), .ZN(n17368) );
  OAI211_X1 U19360 ( .C1(n17371), .C2(n17370), .A(n17369), .B(n17368), .ZN(
        n17372) );
  AOI21_X1 U19361 ( .B1(n17373), .B2(n19157), .A(n17372), .ZN(n17374) );
  OAI21_X1 U19362 ( .B1(n17375), .B2(n19123), .A(n17374), .ZN(P2_U3019) );
  INV_X1 U19363 ( .A(n19104), .ZN(n17393) );
  XNOR2_X1 U19364 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17376) );
  NOR2_X1 U19365 ( .A1(n17388), .A2(n17376), .ZN(n17377) );
  AOI211_X1 U19366 ( .C1(n19159), .C2(n17379), .A(n17378), .B(n17377), .ZN(
        n17380) );
  OAI21_X1 U19367 ( .B1(n19134), .B2(n17381), .A(n17380), .ZN(n17384) );
  NOR2_X1 U19368 ( .A1(n17382), .A2(n19153), .ZN(n17383) );
  AOI211_X1 U19369 ( .C1(n17393), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17384), .B(n17383), .ZN(n17385) );
  OAI21_X1 U19370 ( .B1(n19123), .B2(n17386), .A(n17385), .ZN(P2_U3020) );
  NAND2_X1 U19371 ( .A1(n17387), .A2(n19160), .ZN(n17395) );
  INV_X1 U19372 ( .A(n19052), .ZN(n17390) );
  OAI22_X1 U19373 ( .A1(n17388), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n19043), .B2(n17323), .ZN(n17389) );
  AOI21_X1 U19374 ( .B1(n19154), .B2(n17390), .A(n17389), .ZN(n17391) );
  OAI21_X1 U19375 ( .B1(n19130), .B2(n19047), .A(n17391), .ZN(n17392) );
  AOI21_X1 U19376 ( .B1(n17393), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17392), .ZN(n17394) );
  OAI211_X1 U19377 ( .C1(n17396), .C2(n19153), .A(n17395), .B(n17394), .ZN(
        P2_U3021) );
  NAND2_X1 U19378 ( .A1(n17397), .A2(n19157), .ZN(n17406) );
  XNOR2_X1 U19379 ( .A(n17398), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17399) );
  NAND2_X1 U19380 ( .A1(n17399), .A2(n19113), .ZN(n17402) );
  NOR2_X1 U19381 ( .A1(n17527), .A2(n17400), .ZN(n17413) );
  NAND2_X1 U19382 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17413), .ZN(
        n17401) );
  OAI211_X1 U19383 ( .C1(n17933), .C2(n17323), .A(n17402), .B(n17401), .ZN(
        n17403) );
  AOI21_X1 U19384 ( .B1(n19159), .B2(n17404), .A(n17403), .ZN(n17405) );
  OAI211_X1 U19385 ( .C1(n19134), .C2(n17407), .A(n17406), .B(n17405), .ZN(
        n17408) );
  INV_X1 U19386 ( .A(n17408), .ZN(n17409) );
  OAI21_X1 U19387 ( .B1(n17410), .B2(n19123), .A(n17409), .ZN(P2_U3023) );
  NAND2_X1 U19388 ( .A1(n17811), .A2(n19157), .ZN(n17421) );
  NOR2_X1 U19389 ( .A1(n19031), .A2(n18958), .ZN(n17412) );
  AOI221_X1 U19390 ( .B1(n17413), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n19113), .C2(n17411), .A(n17412), .ZN(n17420) );
  INV_X1 U19391 ( .A(n19038), .ZN(n17414) );
  AOI22_X1 U19392 ( .A1(n19154), .A2(n17414), .B1(n19159), .B2(n19027), .ZN(
        n17419) );
  XNOR2_X1 U19393 ( .A(n17416), .B(n17411), .ZN(n17417) );
  XNOR2_X1 U19394 ( .A(n17415), .B(n17417), .ZN(n17806) );
  NAND2_X1 U19395 ( .A1(n17806), .A2(n19160), .ZN(n17418) );
  NAND4_X1 U19396 ( .A1(n17421), .A2(n17420), .A3(n17419), .A4(n17418), .ZN(
        P2_U3024) );
  NOR3_X1 U19397 ( .A1(n17423), .A2(n17422), .A3(n19153), .ZN(n17433) );
  NAND3_X1 U19398 ( .A1(n17425), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17424), .ZN(n17431) );
  INV_X1 U19399 ( .A(n19022), .ZN(n17429) );
  NOR2_X1 U19400 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17426), .ZN(
        n17427) );
  AOI211_X1 U19401 ( .C1(n19154), .C2(n17429), .A(n17428), .B(n17427), .ZN(
        n17430) );
  OAI211_X1 U19402 ( .C1(n19012), .C2(n19130), .A(n17431), .B(n17430), .ZN(
        n17432) );
  NOR2_X1 U19403 ( .A1(n17433), .A2(n17432), .ZN(n17434) );
  OAI21_X1 U19404 ( .B1(n17435), .B2(n19123), .A(n17434), .ZN(P2_U3025) );
  NAND2_X1 U19405 ( .A1(n17436), .A2(n19157), .ZN(n17444) );
  NOR2_X1 U19406 ( .A1(n19130), .A2(n19000), .ZN(n17441) );
  AOI22_X1 U19407 ( .A1(n19142), .A2(P2_REIP_REG_19__SCAN_IN), .B1(n17438), 
        .B2(n17437), .ZN(n17439) );
  OAI21_X1 U19408 ( .B1(n19134), .B2(n18999), .A(n17439), .ZN(n17440) );
  AOI211_X1 U19409 ( .C1(n17442), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n17441), .B(n17440), .ZN(n17443) );
  OAI211_X1 U19410 ( .C1(n17445), .C2(n19123), .A(n17444), .B(n17443), .ZN(
        P2_U3027) );
  AOI22_X1 U19411 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17480), .B1(
        n19157), .B2(n17793), .ZN(n19141) );
  INV_X1 U19412 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U19413 ( .B1(n19141), .B2(n19140), .A(n17446), .ZN(n17456) );
  NAND2_X1 U19414 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17449), .ZN(
        n17450) );
  NAND2_X1 U19415 ( .A1(n17451), .A2(n17450), .ZN(n17452) );
  NAND2_X1 U19416 ( .A1(n17453), .A2(n17452), .ZN(n17486) );
  OAI211_X1 U19417 ( .C1(n17497), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n19139), .ZN(n17455) );
  NAND2_X1 U19418 ( .A1(n17456), .A2(n17455), .ZN(n17461) );
  OAI22_X1 U19419 ( .A1(n19134), .A2(n18972), .B1(n18958), .B2(n17457), .ZN(
        n17458) );
  AOI21_X1 U19420 ( .B1(n17459), .B2(n19159), .A(n17458), .ZN(n17460) );
  OAI211_X1 U19421 ( .C1(n17462), .C2(n19123), .A(n17461), .B(n17460), .ZN(
        P2_U3029) );
  NAND2_X1 U19422 ( .A1(n17464), .A2(n17463), .ZN(n17466) );
  NAND2_X1 U19423 ( .A1(n17466), .A2(n17465), .ZN(n17761) );
  INV_X1 U19424 ( .A(n17759), .ZN(n17467) );
  AOI21_X1 U19425 ( .B1(n17761), .B2(n17758), .A(n17467), .ZN(n17491) );
  NOR3_X1 U19426 ( .A1(n17493), .A2(n17492), .A3(n17491), .ZN(n17494) );
  NOR2_X1 U19427 ( .A1(n17493), .A2(n17494), .ZN(n17471) );
  NOR2_X1 U19428 ( .A1(n17469), .A2(n17468), .ZN(n17470) );
  XNOR2_X1 U19429 ( .A(n17471), .B(n17470), .ZN(n17780) );
  NAND2_X1 U19430 ( .A1(n17769), .A2(n17473), .ZN(n17474) );
  NAND2_X1 U19431 ( .A1(n17475), .A2(n17474), .ZN(n17778) );
  CLKBUF_X1 U19432 ( .A(n17476), .Z(n17477) );
  OR2_X1 U19433 ( .A1(n17478), .A2(n17477), .ZN(n17479) );
  NAND2_X1 U19434 ( .A1(n17479), .A2(n15732), .ZN(n19712) );
  NOR2_X1 U19435 ( .A1(n13505), .A2(n18958), .ZN(n17483) );
  INV_X1 U19436 ( .A(n17480), .ZN(n17481) );
  NOR2_X1 U19437 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17481), .ZN(
        n17482) );
  NOR2_X1 U19438 ( .A1(n17483), .A2(n17482), .ZN(n17484) );
  OAI21_X1 U19439 ( .B1(n19134), .B2(n19712), .A(n17484), .ZN(n17485) );
  AOI21_X1 U19440 ( .B1(n18956), .B2(n19159), .A(n17485), .ZN(n17488) );
  NAND2_X1 U19441 ( .A1(n17486), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17487) );
  OAI211_X1 U19442 ( .C1(n17778), .C2(n19153), .A(n17488), .B(n17487), .ZN(
        n17489) );
  INV_X1 U19443 ( .A(n17489), .ZN(n17490) );
  OAI21_X1 U19444 ( .B1(n17780), .B2(n19123), .A(n17490), .ZN(P2_U3031) );
  OAI21_X1 U19445 ( .B1(n17493), .B2(n17492), .A(n17491), .ZN(n17496) );
  INV_X1 U19446 ( .A(n17494), .ZN(n17495) );
  NAND2_X1 U19447 ( .A1(n17496), .A2(n17495), .ZN(n17772) );
  INV_X1 U19448 ( .A(n17772), .ZN(n17514) );
  NOR3_X1 U19449 ( .A1(n17573), .A2(n17546), .A3(n17566), .ZN(n17532) );
  NAND2_X1 U19450 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17532), .ZN(
        n17500) );
  NOR2_X1 U19451 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17500), .ZN(
        n17518) );
  OAI21_X1 U19452 ( .B1(n17498), .B2(n17497), .A(n17571), .ZN(n17519) );
  NOR2_X1 U19453 ( .A1(n17518), .A2(n17519), .ZN(n19119) );
  OR2_X1 U19454 ( .A1(n17500), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19128) );
  NAND2_X1 U19455 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19142), .ZN(n17499) );
  OAI221_X1 U19456 ( .B1(n17511), .B2(n19119), .C1(n17511), .C2(n19128), .A(
        n17499), .ZN(n17509) );
  NAND2_X1 U19457 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17501) );
  NOR3_X1 U19458 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17501), .A3(
        n17500), .ZN(n17508) );
  INV_X1 U19459 ( .A(n17502), .ZN(n17503) );
  OR2_X1 U19460 ( .A1(n17504), .A2(n17503), .ZN(n17506) );
  INV_X1 U19461 ( .A(n17477), .ZN(n17505) );
  NAND2_X1 U19462 ( .A1(n17506), .A2(n17505), .ZN(n19715) );
  OAI22_X1 U19463 ( .A1(n18948), .A2(n19130), .B1(n19134), .B2(n19715), .ZN(
        n17507) );
  NOR3_X1 U19464 ( .A1(n17509), .A2(n17508), .A3(n17507), .ZN(n17513) );
  NAND3_X1 U19465 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n17510), .ZN(n17756) );
  NAND2_X1 U19466 ( .A1(n17511), .A2(n17756), .ZN(n17768) );
  NAND3_X1 U19467 ( .A1(n17769), .A2(n19157), .A3(n17768), .ZN(n17512) );
  OAI211_X1 U19468 ( .C1(n17514), .C2(n19123), .A(n17513), .B(n17512), .ZN(
        P2_U3032) );
  NAND2_X1 U19469 ( .A1(n17516), .A2(n19157), .ZN(n17526) );
  NOR2_X1 U19470 ( .A1(n13443), .A2(n18958), .ZN(n17517) );
  AOI211_X1 U19471 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17519), .A(
        n17518), .B(n17517), .ZN(n17525) );
  INV_X1 U19472 ( .A(n19721), .ZN(n17521) );
  AOI22_X1 U19473 ( .A1(n19154), .A2(n17521), .B1(n19159), .B2(n17520), .ZN(
        n17524) );
  NAND2_X1 U19474 ( .A1(n17522), .A2(n19160), .ZN(n17523) );
  NAND4_X1 U19475 ( .A1(n17526), .A2(n17525), .A3(n17524), .A4(n17523), .ZN(
        P2_U3034) );
  AOI21_X1 U19476 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17571), .A(
        n17527), .ZN(n17549) );
  NOR3_X1 U19477 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17573), .A3(
        n17566), .ZN(n17548) );
  OAI21_X1 U19478 ( .B1(n17549), .B2(n17548), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17539) );
  OR2_X1 U19479 ( .A1(n17529), .A2(n17528), .ZN(n17530) );
  NAND2_X1 U19480 ( .A1(n17530), .A2(n16975), .ZN(n19724) );
  INV_X1 U19481 ( .A(n17531), .ZN(n17535) );
  NAND2_X1 U19482 ( .A1(n17533), .A2(n17532), .ZN(n17534) );
  OAI211_X1 U19483 ( .C1(n19134), .C2(n19724), .A(n17535), .B(n17534), .ZN(
        n17536) );
  AOI21_X1 U19484 ( .B1(n19159), .B2(n17537), .A(n17536), .ZN(n17538) );
  OAI211_X1 U19485 ( .C1(n17540), .C2(n19123), .A(n17539), .B(n17538), .ZN(
        n17541) );
  AOI21_X1 U19486 ( .B1(n17542), .B2(n19157), .A(n17541), .ZN(n17543) );
  INV_X1 U19487 ( .A(n17543), .ZN(P2_U3035) );
  INV_X1 U19488 ( .A(n17544), .ZN(n17545) );
  AOI21_X1 U19489 ( .B1(n17546), .B2(n17565), .A(n17545), .ZN(n17752) );
  NAND2_X1 U19490 ( .A1(n17752), .A2(n19157), .ZN(n17563) );
  NOR2_X1 U19491 ( .A1(n13405), .A2(n18958), .ZN(n17547) );
  AOI211_X1 U19492 ( .C1(n17549), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17548), .B(n17547), .ZN(n17562) );
  INV_X1 U19493 ( .A(n17550), .ZN(n17551) );
  XNOR2_X1 U19494 ( .A(n17552), .B(n17551), .ZN(n19727) );
  INV_X1 U19495 ( .A(n19727), .ZN(n17553) );
  AOI22_X1 U19496 ( .A1(n19154), .A2(n17553), .B1(n19159), .B2(n18902), .ZN(
        n17561) );
  NAND2_X1 U19497 ( .A1(n17555), .A2(n17554), .ZN(n17559) );
  OR2_X1 U19498 ( .A1(n17557), .A2(n17556), .ZN(n17558) );
  XNOR2_X1 U19499 ( .A(n17559), .B(n17558), .ZN(n17753) );
  NAND2_X1 U19500 ( .A1(n17753), .A2(n19160), .ZN(n17560) );
  NAND4_X1 U19501 ( .A1(n17563), .A2(n17562), .A3(n17561), .A4(n17560), .ZN(
        P2_U3036) );
  NAND3_X1 U19502 ( .A1(n17565), .A2(n19157), .A3(n17564), .ZN(n17576) );
  INV_X1 U19503 ( .A(n17566), .ZN(n17574) );
  OAI21_X1 U19504 ( .B1(n19134), .B2(n19730), .A(n17567), .ZN(n17568) );
  AOI21_X1 U19505 ( .B1(n19159), .B2(n17569), .A(n17568), .ZN(n17570) );
  OAI21_X1 U19506 ( .B1(n17571), .B2(n17573), .A(n17570), .ZN(n17572) );
  AOI21_X1 U19507 ( .B1(n17574), .B2(n17573), .A(n17572), .ZN(n17575) );
  OAI211_X1 U19508 ( .C1(n19123), .C2(n17577), .A(n17576), .B(n17575), .ZN(
        P2_U3037) );
  OR2_X1 U19509 ( .A1(n17579), .A2(n17578), .ZN(n17580) );
  NAND2_X1 U19510 ( .A1(n17580), .A2(n16999), .ZN(n19736) );
  NAND2_X1 U19511 ( .A1(n19163), .A2(n17581), .ZN(n17584) );
  OAI22_X1 U19512 ( .A1(n19130), .A2(n18891), .B1(n17347), .B2(n17323), .ZN(
        n17582) );
  AOI21_X1 U19513 ( .B1(n19155), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17582), .ZN(n17583) );
  OAI211_X1 U19514 ( .C1(n19134), .C2(n19736), .A(n17584), .B(n17583), .ZN(
        n17585) );
  AOI21_X1 U19515 ( .B1(n17586), .B2(n19160), .A(n17585), .ZN(n17587) );
  OAI21_X1 U19516 ( .B1(n17588), .B2(n19153), .A(n17587), .ZN(P2_U3039) );
  OAI22_X1 U19517 ( .A1(n19153), .A2(n17590), .B1(n17589), .B2(n19134), .ZN(
        n17591) );
  AOI211_X1 U19518 ( .C1(n17593), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17592), .B(n17591), .ZN(n17601) );
  INV_X1 U19519 ( .A(n17594), .ZN(n17596) );
  AOI22_X1 U19520 ( .A1(n17596), .A2(n19160), .B1(n17595), .B2(n19159), .ZN(
        n17600) );
  OAI211_X1 U19521 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n17598), .B(n17597), .ZN(n17599) );
  NAND3_X1 U19522 ( .A1(n17601), .A2(n17600), .A3(n17599), .ZN(P2_U3045) );
  INV_X1 U19523 ( .A(n19074), .ZN(n17606) );
  INV_X1 U19524 ( .A(n17602), .ZN(n17603) );
  NAND2_X1 U19525 ( .A1(n17604), .A2(n17603), .ZN(n17617) );
  MUX2_X1 U19526 ( .A(n17617), .B(n19082), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n17605) );
  AOI21_X1 U19527 ( .B1(n18865), .B2(n17606), .A(n17605), .ZN(n19170) );
  AOI22_X1 U19528 ( .A1(n19054), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18870), .B2(n11223), .ZN(n17622) );
  INV_X1 U19529 ( .A(n17622), .ZN(n17607) );
  OAI222_X1 U19530 ( .A1(n19775), .A2(n19236), .B1(n19224), .B2(n19170), .C1(
        n17661), .C2(n17607), .ZN(n17616) );
  NOR2_X1 U19531 ( .A1(n19237), .A2(n17668), .ZN(n19243) );
  INV_X1 U19532 ( .A(n17608), .ZN(n17609) );
  AND3_X1 U19533 ( .A1(n17611), .A2(n17610), .A3(n17609), .ZN(n17614) );
  NAND3_X1 U19534 ( .A1(n17612), .A2(n19098), .A3(n19201), .ZN(n17613) );
  OAI22_X1 U19535 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19834), .B1(n19184), 
        .B2(n19247), .ZN(n17615) );
  AOI21_X1 U19536 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n19243), .A(n17615), .ZN(
        n19099) );
  MUX2_X1 U19537 ( .A(n17616), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n19099), .Z(P2_U3601) );
  OAI21_X1 U19538 ( .B1(n12663), .B2(n12664), .A(n17617), .ZN(n17619) );
  INV_X1 U19539 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17618) );
  NAND2_X1 U19540 ( .A1(n19082), .A2(n17618), .ZN(n19077) );
  AND2_X1 U19541 ( .A1(n17619), .A2(n19077), .ZN(n17620) );
  OAI21_X1 U19542 ( .B1(n17621), .B2(n19074), .A(n17620), .ZN(n19172) );
  NOR2_X1 U19543 ( .A1(n17622), .A2(n17661), .ZN(n17635) );
  AOI21_X1 U19544 ( .B1(n19054), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17623), .ZN(n17636) );
  INV_X1 U19545 ( .A(n19236), .ZN(n17624) );
  AOI222_X1 U19546 ( .A1(n19172), .A2(n17625), .B1(n17635), .B2(n17636), .C1(
        n19749), .C2(n17624), .ZN(n17627) );
  NAND2_X1 U19547 ( .A1(n19099), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17626) );
  OAI21_X1 U19548 ( .B1(n17627), .B2(n19099), .A(n17626), .ZN(P2_U3600) );
  INV_X1 U19549 ( .A(n13277), .ZN(n17628) );
  NOR2_X1 U19550 ( .A1(n17629), .A2(n17628), .ZN(n19080) );
  NOR2_X1 U19551 ( .A1(n19185), .A2(n19194), .ZN(n19086) );
  INV_X1 U19552 ( .A(n12660), .ZN(n19076) );
  NAND2_X1 U19553 ( .A1(n19076), .A2(n17630), .ZN(n19081) );
  NAND2_X1 U19554 ( .A1(n19084), .A2(n19081), .ZN(n17631) );
  MUX2_X1 U19555 ( .A(n19080), .B(n19086), .S(n17631), .Z(n17634) );
  NAND2_X1 U19556 ( .A1(n19082), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17632) );
  MUX2_X1 U19557 ( .A(n17632), .B(n19077), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17633) );
  OAI211_X1 U19558 ( .C1(n14411), .C2(n19074), .A(n17634), .B(n17633), .ZN(
        n19174) );
  INV_X1 U19559 ( .A(n19174), .ZN(n17638) );
  INV_X1 U19560 ( .A(n17635), .ZN(n17637) );
  OAI222_X1 U19561 ( .A1(n20015), .A2(n19236), .B1(n19224), .B2(n17638), .C1(
        n17637), .C2(n17636), .ZN(n17639) );
  MUX2_X1 U19562 ( .A(n17639), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19099), .Z(P2_U3599) );
  NAND2_X1 U19563 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19277) );
  NAND2_X1 U19564 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18702) );
  INV_X1 U19565 ( .A(n18702), .ZN(n18653) );
  NAND2_X1 U19566 ( .A1(n21885), .A2(n18228), .ZN(n20717) );
  NOR2_X1 U19567 ( .A1(n18653), .A2(n20717), .ZN(n17642) );
  NOR2_X1 U19568 ( .A1(n21885), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19280) );
  INV_X1 U19569 ( .A(n19280), .ZN(n17641) );
  OAI211_X1 U19570 ( .C1(n21848), .C2(n21412), .A(n18160), .B(n21846), .ZN(
        n18229) );
  NOR2_X1 U19571 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18229), .ZN(n17640) );
  INV_X1 U19572 ( .A(n17653), .ZN(n21883) );
  NAND2_X1 U19573 ( .A1(n21846), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21421) );
  AOI21_X1 U19574 ( .B1(n20714), .B2(n18228), .A(n21887), .ZN(n19279) );
  OAI21_X1 U19575 ( .B1(n17640), .B2(n21883), .A(n19518), .ZN(n18231) );
  NAND2_X1 U19576 ( .A1(n17641), .A2(n18231), .ZN(n18755) );
  AOI221_X1 U19577 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19277), .C1(n17642), 
        .C2(n19277), .A(n18755), .ZN(n18753) );
  NAND3_X1 U19578 ( .A1(n20711), .A2(n21885), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19333) );
  INV_X1 U19579 ( .A(n19333), .ZN(n18754) );
  NOR2_X1 U19580 ( .A1(n21885), .A2(n21852), .ZN(n19284) );
  OAI21_X1 U19581 ( .B1(n17642), .B2(n19284), .A(n18231), .ZN(n18757) );
  INV_X1 U19582 ( .A(n18757), .ZN(n18751) );
  OAI22_X1 U19583 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18754), .B1(
        n18751), .B2(n18750), .ZN(n17643) );
  AOI22_X1 U19584 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18753), .B1(
        n17643), .B2(n21861), .ZN(P3_U2865) );
  NOR2_X1 U19585 ( .A1(n17645), .A2(n17644), .ZN(n17646) );
  XNOR2_X1 U19586 ( .A(n17646), .B(n17696), .ZN(n22051) );
  NAND4_X1 U19587 ( .A1(n22051), .A2(n17648), .A3(n17688), .A4(n17647), .ZN(
        n17649) );
  OAI21_X1 U19588 ( .B1(n17650), .B2(n17696), .A(n17649), .ZN(P1_U3468) );
  INV_X1 U19589 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17651) );
  AOI221_X1 U19590 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n22288), .C1(
        P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n22240), 
        .ZN(n22236) );
  INV_X1 U19591 ( .A(BS16), .ZN(n17682) );
  INV_X1 U19592 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22285) );
  NAND2_X1 U19593 ( .A1(n22285), .A2(n22288), .ZN(n22238) );
  AOI21_X1 U19594 ( .B1(n17682), .B2(n22238), .A(n17652), .ZN(n22232) );
  AOI21_X1 U19595 ( .B1(n17651), .B2(n17652), .A(n22232), .ZN(P3_U3280) );
  AND2_X1 U19596 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17652), .ZN(P3_U3028) );
  AND2_X1 U19597 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17652), .ZN(P3_U3027) );
  AND2_X1 U19598 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17652), .ZN(P3_U3026) );
  AND2_X1 U19599 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17652), .ZN(P3_U3025) );
  AND2_X1 U19600 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17652), .ZN(P3_U3024) );
  AND2_X1 U19601 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17652), .ZN(P3_U3023) );
  AND2_X1 U19602 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17652), .ZN(P3_U3022) );
  AND2_X1 U19603 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17652), .ZN(P3_U3021) );
  AND2_X1 U19604 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17652), .ZN(
        P3_U3020) );
  AND2_X1 U19605 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17652), .ZN(
        P3_U3019) );
  AND2_X1 U19606 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17652), .ZN(
        P3_U3018) );
  AND2_X1 U19607 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17652), .ZN(
        P3_U3017) );
  AND2_X1 U19608 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17652), .ZN(
        P3_U3016) );
  AND2_X1 U19609 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17652), .ZN(
        P3_U3015) );
  AND2_X1 U19610 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17652), .ZN(
        P3_U3014) );
  AND2_X1 U19611 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17652), .ZN(
        P3_U3013) );
  AND2_X1 U19612 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17652), .ZN(
        P3_U3012) );
  AND2_X1 U19613 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17652), .ZN(
        P3_U3011) );
  AND2_X1 U19614 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17652), .ZN(
        P3_U3010) );
  AND2_X1 U19615 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17652), .ZN(
        P3_U3009) );
  AND2_X1 U19616 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17652), .ZN(
        P3_U3008) );
  AND2_X1 U19617 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17652), .ZN(
        P3_U3007) );
  AND2_X1 U19618 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17652), .ZN(
        P3_U3006) );
  AND2_X1 U19619 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17652), .ZN(
        P3_U3005) );
  AND2_X1 U19620 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17652), .ZN(
        P3_U3004) );
  AND2_X1 U19621 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17652), .ZN(
        P3_U3003) );
  AND2_X1 U19622 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17652), .ZN(
        P3_U3002) );
  AND2_X1 U19623 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17652), .ZN(
        P3_U3001) );
  AND2_X1 U19624 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17652), .ZN(
        P3_U3000) );
  AND2_X1 U19625 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17652), .ZN(
        P3_U2999) );
  AOI21_X1 U19626 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17654)
         );
  NOR4_X1 U19627 ( .A1(n18746), .A2(n20715), .A3(n21875), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21833) );
  AOI211_X1 U19628 ( .C1(n18702), .C2(n17654), .A(n17653), .B(n21833), .ZN(
        P3_U2998) );
  NOR2_X1 U19629 ( .A1(n21865), .A2(n18231), .ZN(P3_U2867) );
  NAND2_X1 U19630 ( .A1(n20715), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18744) );
  AND2_X1 U19631 ( .A1(n18812), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AND2_X1 U19632 ( .A1(n18227), .A2(n20720), .ZN(n17657) );
  INV_X1 U19633 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18782) );
  AOI22_X1 U19634 ( .A1(n17657), .A2(n18782), .B1(n17656), .B2(n20713), .ZN(
        P3_U3298) );
  INV_X1 U19635 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18781) );
  NAND2_X1 U19636 ( .A1(n19610), .A2(n17656), .ZN(n20809) );
  INV_X1 U19637 ( .A(n20809), .ZN(n21182) );
  AOI21_X1 U19638 ( .B1(n17657), .B2(n18781), .A(n21182), .ZN(P3_U3299) );
  NOR2_X1 U19639 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22263), .ZN(n22274) );
  INV_X1 U19640 ( .A(n22266), .ZN(n17658) );
  AOI21_X1 U19641 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22274), .A(n17658), 
        .ZN(n17659) );
  INV_X1 U19642 ( .A(n17659), .ZN(n22231) );
  INV_X1 U19643 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17679) );
  NAND2_X1 U19644 ( .A1(n22270), .A2(n22263), .ZN(n22261) );
  AOI21_X1 U19645 ( .B1(n17682), .B2(n22261), .A(n17660), .ZN(n22227) );
  AOI21_X1 U19646 ( .B1(n17660), .B2(n17679), .A(n22227), .ZN(P2_U3591) );
  AND2_X1 U19647 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17660), .ZN(P2_U3208) );
  AND2_X1 U19648 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17660), .ZN(P2_U3207) );
  AND2_X1 U19649 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17660), .ZN(P2_U3206) );
  AND2_X1 U19650 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17660), .ZN(P2_U3205) );
  AND2_X1 U19651 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17660), .ZN(P2_U3204) );
  AND2_X1 U19652 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17660), .ZN(P2_U3203) );
  AND2_X1 U19653 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17660), .ZN(P2_U3202) );
  AND2_X1 U19654 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17660), .ZN(P2_U3201) );
  AND2_X1 U19655 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17660), .ZN(
        P2_U3200) );
  AND2_X1 U19656 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17660), .ZN(
        P2_U3199) );
  AND2_X1 U19657 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17660), .ZN(
        P2_U3198) );
  AND2_X1 U19658 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17660), .ZN(
        P2_U3197) );
  AND2_X1 U19659 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17660), .ZN(
        P2_U3196) );
  AND2_X1 U19660 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17660), .ZN(
        P2_U3195) );
  AND2_X1 U19661 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17659), .ZN(
        P2_U3194) );
  AND2_X1 U19662 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17659), .ZN(
        P2_U3193) );
  AND2_X1 U19663 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17659), .ZN(
        P2_U3192) );
  AND2_X1 U19664 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17659), .ZN(
        P2_U3191) );
  AND2_X1 U19665 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17659), .ZN(
        P2_U3190) );
  AND2_X1 U19666 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17659), .ZN(
        P2_U3189) );
  AND2_X1 U19667 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17659), .ZN(
        P2_U3188) );
  AND2_X1 U19668 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17659), .ZN(
        P2_U3187) );
  AND2_X1 U19669 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17659), .ZN(
        P2_U3186) );
  AND2_X1 U19670 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17659), .ZN(
        P2_U3185) );
  AND2_X1 U19671 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17659), .ZN(
        P2_U3184) );
  AND2_X1 U19672 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17659), .ZN(
        P2_U3183) );
  AND2_X1 U19673 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17660), .ZN(
        P2_U3182) );
  AND2_X1 U19674 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17660), .ZN(
        P2_U3181) );
  AND2_X1 U19675 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17660), .ZN(
        P2_U3180) );
  AND2_X1 U19676 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17660), .ZN(
        P2_U3179) );
  NAND2_X1 U19677 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n22264), .ZN(n19223) );
  NOR2_X1 U19678 ( .A1(n17661), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18848) );
  AOI21_X1 U19679 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n18848), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17662) );
  AOI221_X1 U19680 ( .B1(n19223), .B2(n17662), .C1(n17661), .C2(n17662), .A(
        n19243), .ZN(P2_U3178) );
  INV_X1 U19681 ( .A(n19243), .ZN(n19232) );
  INV_X1 U19682 ( .A(n18848), .ZN(n17663) );
  NAND2_X1 U19683 ( .A1(n19215), .A2(n17663), .ZN(n19235) );
  NAND2_X1 U19684 ( .A1(n17668), .A2(n19235), .ZN(n19744) );
  OAI221_X1 U19685 ( .B1(n12926), .B2(n19232), .C1(n19242), .C2(n19232), .A(
        n20286), .ZN(n17844) );
  NOR2_X1 U19686 ( .A1(n19181), .A2(n17844), .ZN(P2_U3047) );
  OAI21_X1 U19687 ( .B1(n17666), .B2(n17665), .A(n17664), .ZN(n17667) );
  NOR2_X1 U19688 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17668), .ZN(n17876) );
  NOR2_X4 U19689 ( .A1(n17883), .A2(n17912), .ZN(n17901) );
  AND2_X1 U19690 ( .A1(n17901), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19691 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17672) );
  NOR4_X1 U19692 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17671) );
  NOR4_X1 U19693 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17670) );
  NOR4_X1 U19694 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17669) );
  NAND4_X1 U19695 ( .A1(n17672), .A2(n17671), .A3(n17670), .A4(n17669), .ZN(
        n17678) );
  NOR4_X1 U19696 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17676) );
  AOI211_X1 U19697 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17675) );
  NOR4_X1 U19698 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17674) );
  NOR4_X1 U19699 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17673) );
  NAND4_X1 U19700 ( .A1(n17676), .A2(n17675), .A3(n17674), .A4(n17673), .ZN(
        n17677) );
  NOR2_X1 U19701 ( .A1(n17678), .A2(n17677), .ZN(n17854) );
  INV_X1 U19702 ( .A(n17854), .ZN(n17852) );
  NOR2_X1 U19703 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17852), .ZN(n17847) );
  INV_X1 U19704 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22230) );
  NAND3_X1 U19705 ( .A1(n18862), .A2(n22230), .A3(n17679), .ZN(n17851) );
  INV_X1 U19706 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U19707 ( .A1(n17847), .A2(n17851), .B1(n17852), .B2(n17680), .ZN(
        P2_U2821) );
  INV_X1 U19708 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17681) );
  AOI22_X1 U19709 ( .A1(n17847), .A2(n18862), .B1(n17852), .B2(n17681), .ZN(
        P2_U2820) );
  INV_X1 U19710 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20530) );
  AOI21_X1 U19711 ( .B1(n22251), .B2(P1_STATE_REG_1__SCAN_IN), .A(n11714), 
        .ZN(n22241) );
  INV_X1 U19712 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22250) );
  NOR2_X2 U19713 ( .A1(n22250), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22727) );
  NOR2_X1 U19714 ( .A1(n22241), .A2(n22727), .ZN(n22226) );
  NAND2_X1 U19715 ( .A1(n22251), .A2(n11714), .ZN(n20639) );
  AOI21_X1 U19716 ( .B1(n17682), .B2(n20639), .A(n17683), .ZN(n22222) );
  AOI21_X1 U19717 ( .B1(n20530), .B2(n17683), .A(n22222), .ZN(P1_U3464) );
  AND2_X1 U19718 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17683), .ZN(P1_U3193) );
  AND2_X1 U19719 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17683), .ZN(P1_U3192) );
  AND2_X1 U19720 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17683), .ZN(P1_U3191) );
  AND2_X1 U19721 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17683), .ZN(P1_U3190) );
  AND2_X1 U19722 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17683), .ZN(P1_U3189) );
  AND2_X1 U19723 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17683), .ZN(P1_U3188) );
  AND2_X1 U19724 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17683), .ZN(P1_U3187) );
  AND2_X1 U19725 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17683), .ZN(P1_U3186) );
  AND2_X1 U19726 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17683), .ZN(
        P1_U3185) );
  AND2_X1 U19727 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17683), .ZN(
        P1_U3184) );
  AND2_X1 U19728 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17683), .ZN(
        P1_U3183) );
  AND2_X1 U19729 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17683), .ZN(
        P1_U3182) );
  AND2_X1 U19730 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17683), .ZN(
        P1_U3181) );
  AND2_X1 U19731 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17683), .ZN(
        P1_U3180) );
  AND2_X1 U19732 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17683), .ZN(
        P1_U3179) );
  AND2_X1 U19733 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17683), .ZN(
        P1_U3178) );
  AND2_X1 U19734 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17683), .ZN(
        P1_U3177) );
  AND2_X1 U19735 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17683), .ZN(
        P1_U3176) );
  AND2_X1 U19736 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17683), .ZN(
        P1_U3175) );
  AND2_X1 U19737 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17683), .ZN(
        P1_U3174) );
  AND2_X1 U19738 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17683), .ZN(
        P1_U3173) );
  AND2_X1 U19739 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17683), .ZN(
        P1_U3172) );
  AND2_X1 U19740 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17683), .ZN(
        P1_U3171) );
  AND2_X1 U19741 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17683), .ZN(
        P1_U3170) );
  AND2_X1 U19742 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17683), .ZN(
        P1_U3169) );
  AND2_X1 U19743 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17683), .ZN(
        P1_U3168) );
  AND2_X1 U19744 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17683), .ZN(
        P1_U3167) );
  AND2_X1 U19745 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17683), .ZN(
        P1_U3166) );
  AND2_X1 U19746 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17683), .ZN(
        P1_U3165) );
  AND2_X1 U19747 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17683), .ZN(
        P1_U3164) );
  MUX2_X1 U19748 ( .A(n17685), .B(n17684), .S(n17697), .Z(n17708) );
  INV_X1 U19749 ( .A(n17708), .ZN(n17716) );
  MUX2_X1 U19750 ( .A(n17687), .B(n17686), .S(n17697), .Z(n17715) );
  NAND2_X1 U19751 ( .A1(n17688), .A2(n22051), .ZN(n17695) );
  OAI21_X1 U19752 ( .B1(P1_MORE_REG_SCAN_IN), .B2(P1_FLUSH_REG_SCAN_IN), .A(
        n17689), .ZN(n17692) );
  INV_X1 U19753 ( .A(n17690), .ZN(n17691) );
  AND3_X1 U19754 ( .A1(n17693), .A2(n17692), .A3(n17691), .ZN(n17694) );
  OAI211_X1 U19755 ( .C1(n17697), .C2(n17696), .A(n17695), .B(n17694), .ZN(
        n17714) );
  AND2_X1 U19756 ( .A1(n17698), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17699) );
  AND2_X1 U19757 ( .A1(n17700), .A2(n17699), .ZN(n17705) );
  AOI211_X1 U19758 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n17705), .A(
        n17702), .B(n17701), .ZN(n17703) );
  INV_X1 U19759 ( .A(n17703), .ZN(n17704) );
  OAI21_X1 U19760 ( .B1(n17705), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17704), .ZN(n17706) );
  AOI222_X1 U19761 ( .A1(n17715), .A2(n17707), .B1(n17715), .B2(n17706), .C1(
        n17707), .C2(n17706), .ZN(n17712) );
  OR2_X1 U19762 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17708), .ZN(
        n17711) );
  NOR2_X1 U19763 ( .A1(n17716), .A2(n17709), .ZN(n17710) );
  AOI211_X1 U19764 ( .C1(n17712), .C2(n17711), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n17710), .ZN(n17713) );
  AOI211_X1 U19765 ( .C1(n17716), .C2(n17715), .A(n17714), .B(n17713), .ZN(
        n22221) );
  NOR2_X1 U19766 ( .A1(n17718), .A2(n17717), .ZN(n17719) );
  AOI221_X1 U19767 ( .B1(n17720), .B2(n22207), .C1(n22243), .C2(n22207), .A(
        n17719), .ZN(n17725) );
  OAI221_X1 U19768 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n22221), 
        .A(n17725), .ZN(n22206) );
  OAI211_X1 U19769 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22243), .A(n17721), 
        .B(n22206), .ZN(n22217) );
  OR3_X1 U19770 ( .A1(n22242), .A2(n22210), .A3(n17722), .ZN(n17724) );
  AND2_X1 U19771 ( .A1(n17724), .A2(n17723), .ZN(n22208) );
  AOI21_X1 U19772 ( .B1(n22208), .B2(n22209), .A(n17725), .ZN(n17726) );
  AOI21_X1 U19773 ( .B1(n17727), .B2(n22217), .A(n17726), .ZN(P1_U3162) );
  NOR2_X1 U19774 ( .A1(n17729), .A2(n17728), .ZN(P1_U3032) );
  AND2_X1 U19775 ( .A1(n20469), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI21_X1 U19776 ( .B1(n22241), .B2(n17730), .A(n22727), .ZN(P1_U2802) );
  INV_X1 U19777 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17916) );
  OAI22_X1 U19778 ( .A1(n19237), .A2(n17732), .B1(n17731), .B2(n17916), .ZN(
        P2_U2816) );
  AOI22_X1 U19779 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19142), .ZN(n17738) );
  OAI22_X1 U19780 ( .A1(n17734), .A2(n17779), .B1(n13196), .B2(n17733), .ZN(
        n17735) );
  AOI21_X1 U19781 ( .B1(n17807), .B2(n17736), .A(n17735), .ZN(n17737) );
  OAI211_X1 U19782 ( .C1(n17827), .C2(n17739), .A(n17738), .B(n17737), .ZN(
        P2_U3009) );
  AOI22_X1 U19783 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19142), .B1(n17777), 
        .B2(n17740), .ZN(n17750) );
  NAND2_X1 U19784 ( .A1(n17742), .A2(n17741), .ZN(n17743) );
  XNOR2_X1 U19785 ( .A(n17744), .B(n17743), .ZN(n19161) );
  OAI21_X1 U19786 ( .B1(n11181), .B2(n17746), .A(n17745), .ZN(n17748) );
  INV_X1 U19787 ( .A(n17748), .ZN(n19156) );
  AOI222_X1 U19788 ( .A1(n19161), .A2(n17818), .B1(n17807), .B2(n19158), .C1(
        n17820), .C2(n19156), .ZN(n17749) );
  OAI211_X1 U19789 ( .C1(n17751), .C2(n17789), .A(n17750), .B(n17749), .ZN(
        P2_U3006) );
  AOI22_X1 U19790 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19142), .ZN(n17755) );
  AOI222_X1 U19791 ( .A1(n17753), .A2(n17818), .B1(n17807), .B2(n18902), .C1(
        n17820), .C2(n17752), .ZN(n17754) );
  OAI211_X1 U19792 ( .C1(n17827), .C2(n18900), .A(n17755), .B(n17754), .ZN(
        P2_U3004) );
  AOI22_X1 U19793 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19142), .B1(n17777), 
        .B2(n18933), .ZN(n17767) );
  OAI21_X1 U19794 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17757), .A(
        n17756), .ZN(n19121) );
  NAND2_X1 U19795 ( .A1(n17759), .A2(n17758), .ZN(n17760) );
  XNOR2_X1 U19796 ( .A(n17761), .B(n17760), .ZN(n19124) );
  INV_X1 U19797 ( .A(n19122), .ZN(n17762) );
  NAND2_X1 U19798 ( .A1(n17762), .A2(n17807), .ZN(n17763) );
  OAI211_X1 U19799 ( .C1(n18930), .C2(n17789), .A(n17767), .B(n17766), .ZN(
        P2_U3001) );
  AOI22_X1 U19800 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19142), .ZN(n17774) );
  NAND3_X1 U19801 ( .A1(n17769), .A2(n17820), .A3(n17768), .ZN(n17770) );
  OAI21_X1 U19802 ( .B1(n13199), .B2(n18948), .A(n17770), .ZN(n17771) );
  AOI21_X1 U19803 ( .B1(n17772), .B2(n17818), .A(n17771), .ZN(n17773) );
  OAI211_X1 U19804 ( .C1(n17827), .C2(n17775), .A(n17774), .B(n17773), .ZN(
        P2_U3000) );
  AOI22_X1 U19805 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19142), .B1(n17777), 
        .B2(n17776), .ZN(n17783) );
  OAI22_X1 U19806 ( .A1(n17780), .A2(n13196), .B1(n17779), .B2(n17778), .ZN(
        n17781) );
  AOI21_X1 U19807 ( .B1(n17807), .B2(n18956), .A(n17781), .ZN(n17782) );
  OAI211_X1 U19808 ( .C1(n17784), .C2(n17789), .A(n17783), .B(n17782), .ZN(
        P2_U2999) );
  XOR2_X1 U19809 ( .A(n17785), .B(n17786), .Z(n19137) );
  NOR2_X1 U19810 ( .A1(n17827), .A2(n17787), .ZN(n17791) );
  OR2_X1 U19811 ( .A1(n18958), .A2(n13018), .ZN(n19132) );
  OAI21_X1 U19812 ( .B1(n17789), .B2(n17788), .A(n19132), .ZN(n17790) );
  AOI211_X1 U19813 ( .C1(n19137), .C2(n17818), .A(n17791), .B(n17790), .ZN(
        n17795) );
  OAI211_X1 U19814 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17793), .A(
        n17792), .B(n17820), .ZN(n17794) );
  OAI211_X1 U19815 ( .C1(n19131), .C2(n13199), .A(n17795), .B(n17794), .ZN(
        P2_U2998) );
  AOI22_X1 U19816 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19142), .ZN(n17804) );
  OAI21_X1 U19817 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17797), .A(
        n17796), .ZN(n19152) );
  INV_X1 U19818 ( .A(n19152), .ZN(n17802) );
  NAND2_X1 U19819 ( .A1(n17800), .A2(n17799), .ZN(n17801) );
  XNOR2_X1 U19820 ( .A(n11193), .B(n17801), .ZN(n19149) );
  AOI222_X1 U19821 ( .A1(n17802), .A2(n17820), .B1(n17807), .B2(n19148), .C1(
        n17818), .C2(n19149), .ZN(n17803) );
  OAI211_X1 U19822 ( .C1(n17827), .C2(n17805), .A(n17804), .B(n17803), .ZN(
        P2_U2996) );
  AOI22_X1 U19823 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19142), .ZN(n17813) );
  NAND2_X1 U19824 ( .A1(n19027), .A2(n17807), .ZN(n17808) );
  OAI211_X1 U19825 ( .C1(n17827), .C2(n19026), .A(n17813), .B(n17812), .ZN(
        P2_U2992) );
  AOI22_X1 U19826 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17814), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19142), .ZN(n17825) );
  XNOR2_X1 U19827 ( .A(n17816), .B(n19112), .ZN(n17817) );
  XNOR2_X1 U19828 ( .A(n17815), .B(n17817), .ZN(n19106) );
  NAND2_X1 U19829 ( .A1(n19106), .A2(n17818), .ZN(n17822) );
  XNOR2_X1 U19830 ( .A(n17819), .B(n19112), .ZN(n19107) );
  NAND2_X1 U19831 ( .A1(n19107), .A2(n17820), .ZN(n17821) );
  OAI211_X1 U19832 ( .C1(n13199), .C2(n19110), .A(n17822), .B(n17821), .ZN(
        n17823) );
  INV_X1 U19833 ( .A(n17823), .ZN(n17824) );
  OAI211_X1 U19834 ( .C1(n17827), .C2(n17826), .A(n17825), .B(n17824), .ZN(
        P2_U2990) );
  INV_X1 U19835 ( .A(n17844), .ZN(n17846) );
  INV_X1 U19836 ( .A(n17828), .ZN(n18851) );
  NAND3_X1 U19837 ( .A1(n17829), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U19838 ( .B1(n19775), .B2(n18851), .A(n17830), .ZN(n17831) );
  AOI21_X1 U19839 ( .B1(n19856), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17831), 
        .ZN(n17832) );
  OAI22_X1 U19840 ( .A1(n19856), .A2(n17844), .B1(n17846), .B2(n17832), .ZN(
        P2_U3605) );
  NAND2_X1 U19841 ( .A1(n19749), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19845) );
  INV_X1 U19842 ( .A(n19845), .ZN(n17833) );
  NAND2_X1 U19843 ( .A1(n20015), .A2(n17833), .ZN(n19908) );
  NAND2_X1 U19844 ( .A1(n19845), .A2(n19939), .ZN(n17834) );
  NAND2_X1 U19845 ( .A1(n17834), .A2(n19224), .ZN(n17843) );
  NAND2_X1 U19846 ( .A1(n19883), .A2(n17843), .ZN(n17836) );
  NAND2_X1 U19847 ( .A1(n20012), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17835) );
  OAI211_X1 U19848 ( .C1(n19908), .C2(n19953), .A(n17836), .B(n17835), .ZN(
        n17837) );
  INV_X1 U19849 ( .A(n17837), .ZN(n17838) );
  AOI22_X1 U19850 ( .A1(n17846), .A2(n19906), .B1(n17838), .B2(n17844), .ZN(
        P2_U3603) );
  NOR2_X1 U19851 ( .A1(n19953), .A2(n22228), .ZN(n17841) );
  OR2_X1 U19852 ( .A1(n19749), .A2(n17841), .ZN(n17839) );
  AOI22_X1 U19853 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20219), .B1(n17843), 
        .B2(n17839), .ZN(n17840) );
  AOI22_X1 U19854 ( .A1(n17846), .A2(n19910), .B1(n17840), .B2(n17844), .ZN(
        P2_U3604) );
  INV_X1 U19855 ( .A(n20017), .ZN(n20120) );
  OAI21_X1 U19856 ( .B1(n19872), .B2(n19814), .A(n19821), .ZN(n17842) );
  AOI222_X1 U19857 ( .A1(n17843), .A2(n19909), .B1(n20120), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n17842), .C2(n17841), .ZN(n17845) );
  AOI22_X1 U19858 ( .A1(n17846), .A2(n19905), .B1(n17845), .B2(n17844), .ZN(
        P2_U3602) );
  NAND2_X1 U19859 ( .A1(n17847), .A2(n22230), .ZN(n17850) );
  OAI21_X1 U19860 ( .B1(n17918), .B2(n18862), .A(n17854), .ZN(n17848) );
  OAI21_X1 U19861 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17854), .A(n17848), 
        .ZN(n17849) );
  OAI221_X1 U19862 ( .B1(n17850), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17850), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17849), .ZN(P2_U2822) );
  INV_X1 U19863 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17853) );
  OAI221_X1 U19864 ( .B1(n17854), .B2(n17853), .C1(n17852), .C2(n17851), .A(
        n17850), .ZN(P2_U2823) );
  INV_X1 U19865 ( .A(n17855), .ZN(n22262) );
  MUX2_X1 U19866 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n22262), .Z(P2_U3611) );
  INV_X2 U19867 ( .A(n22262), .ZN(n17942) );
  INV_X1 U19868 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17856) );
  AOI22_X1 U19869 ( .A1(n17942), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17856), 
        .B2(n22262), .ZN(P2_U3608) );
  AOI21_X1 U19870 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22231), .ZN(n17857) );
  INV_X1 U19871 ( .A(n17857), .ZN(P2_U2815) );
  AOI22_X1 U19872 ( .A1(n17912), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17858) );
  OAI21_X1 U19873 ( .B1(n13307), .B2(n17881), .A(n17858), .ZN(P2_U2951) );
  INV_X1 U19874 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U19875 ( .A1(n17876), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17859) );
  OAI21_X1 U19876 ( .B1(n17860), .B2(n17881), .A(n17859), .ZN(P2_U2950) );
  INV_X1 U19877 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17862) );
  AOI22_X1 U19878 ( .A1(n17912), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17861) );
  OAI21_X1 U19879 ( .B1(n17862), .B2(n17881), .A(n17861), .ZN(P2_U2949) );
  INV_X1 U19880 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17864) );
  AOI22_X1 U19881 ( .A1(n17876), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17863) );
  OAI21_X1 U19882 ( .B1(n17864), .B2(n17881), .A(n17863), .ZN(P2_U2948) );
  INV_X1 U19883 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17866) );
  AOI22_X1 U19884 ( .A1(n17876), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17865) );
  OAI21_X1 U19885 ( .B1(n17866), .B2(n17881), .A(n17865), .ZN(P2_U2947) );
  INV_X1 U19886 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U19887 ( .A1(n17876), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17867) );
  OAI21_X1 U19888 ( .B1(n17868), .B2(n17881), .A(n17867), .ZN(P2_U2946) );
  INV_X1 U19889 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U19890 ( .A1(n17876), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17869) );
  OAI21_X1 U19891 ( .B1(n19968), .B2(n17881), .A(n17869), .ZN(P2_U2945) );
  INV_X1 U19892 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U19893 ( .A1(n17876), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17870) );
  OAI21_X1 U19894 ( .B1(n19735), .B2(n17881), .A(n17870), .ZN(P2_U2944) );
  INV_X1 U19895 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19733) );
  AOI22_X1 U19896 ( .A1(n17876), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17871) );
  OAI21_X1 U19897 ( .B1(n19733), .B2(n17881), .A(n17871), .ZN(P2_U2943) );
  INV_X1 U19898 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19729) );
  AOI22_X1 U19899 ( .A1(n17876), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17872) );
  OAI21_X1 U19900 ( .B1(n19729), .B2(n17881), .A(n17872), .ZN(P2_U2942) );
  AOI22_X1 U19901 ( .A1(n17876), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17873) );
  OAI21_X1 U19902 ( .B1(n17874), .B2(n17881), .A(n17873), .ZN(P2_U2941) );
  INV_X1 U19903 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19723) );
  AOI22_X1 U19904 ( .A1(n17912), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17875) );
  OAI21_X1 U19905 ( .B1(n19723), .B2(n17881), .A(n17875), .ZN(P2_U2940) );
  INV_X1 U19906 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U19907 ( .A1(n17876), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17877) );
  OAI21_X1 U19908 ( .B1(n19720), .B2(n17881), .A(n17877), .ZN(P2_U2939) );
  INV_X1 U19909 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19717) );
  AOI22_X1 U19910 ( .A1(n17912), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17878) );
  OAI21_X1 U19911 ( .B1(n19717), .B2(n17881), .A(n17878), .ZN(P2_U2938) );
  INV_X1 U19912 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U19913 ( .A1(n17912), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17879) );
  OAI21_X1 U19914 ( .B1(n19714), .B2(n17881), .A(n17879), .ZN(P2_U2937) );
  INV_X1 U19915 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19711) );
  AOI22_X1 U19916 ( .A1(n17912), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17880) );
  OAI21_X1 U19917 ( .B1(n19711), .B2(n17881), .A(n17880), .ZN(P2_U2936) );
  NAND2_X1 U19918 ( .A1(n17883), .A2(n17882), .ZN(n17914) );
  AOI22_X1 U19919 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17901), .B1(n17912), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n17884) );
  OAI21_X1 U19920 ( .B1(n17885), .B2(n17914), .A(n17884), .ZN(P2_U2935) );
  AOI22_X1 U19921 ( .A1(n17912), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n17886) );
  OAI21_X1 U19922 ( .B1(n17887), .B2(n17914), .A(n17886), .ZN(P2_U2934) );
  INV_X1 U19923 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n17889) );
  AOI22_X1 U19924 ( .A1(n17912), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n17888) );
  OAI21_X1 U19925 ( .B1(n17889), .B2(n17914), .A(n17888), .ZN(P2_U2933) );
  AOI22_X1 U19926 ( .A1(n17912), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n17890) );
  OAI21_X1 U19927 ( .B1(n17891), .B2(n17914), .A(n17890), .ZN(P2_U2932) );
  INV_X1 U19928 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U19929 ( .A1(n17912), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n17892) );
  OAI21_X1 U19930 ( .B1(n20065), .B2(n17914), .A(n17892), .ZN(P2_U2931) );
  AOI22_X1 U19931 ( .A1(n17912), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n17893) );
  OAI21_X1 U19932 ( .B1(n17894), .B2(n17914), .A(n17893), .ZN(P2_U2930) );
  AOI22_X1 U19933 ( .A1(n17912), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n17895) );
  OAI21_X1 U19934 ( .B1(n17896), .B2(n17914), .A(n17895), .ZN(P2_U2929) );
  AOI22_X1 U19935 ( .A1(n17912), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n17897) );
  OAI21_X1 U19936 ( .B1(n17898), .B2(n17914), .A(n17897), .ZN(P2_U2928) );
  AOI22_X1 U19937 ( .A1(n17912), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n17899) );
  OAI21_X1 U19938 ( .B1(n17900), .B2(n17914), .A(n17899), .ZN(P2_U2927) );
  AOI22_X1 U19939 ( .A1(n17912), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n17902) );
  OAI21_X1 U19940 ( .B1(n17903), .B2(n17914), .A(n17902), .ZN(P2_U2926) );
  AOI22_X1 U19941 ( .A1(n17912), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n17904) );
  OAI21_X1 U19942 ( .B1(n17905), .B2(n17914), .A(n17904), .ZN(P2_U2925) );
  AOI22_X1 U19943 ( .A1(n17912), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n17906) );
  OAI21_X1 U19944 ( .B1(n17907), .B2(n17914), .A(n17906), .ZN(P2_U2924) );
  AOI22_X1 U19945 ( .A1(n17912), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n17908) );
  OAI21_X1 U19946 ( .B1(n17909), .B2(n17914), .A(n17908), .ZN(P2_U2923) );
  AOI22_X1 U19947 ( .A1(n17912), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n17910) );
  OAI21_X1 U19948 ( .B1(n17911), .B2(n17914), .A(n17910), .ZN(P2_U2922) );
  AOI22_X1 U19949 ( .A1(n17912), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17901), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n17913) );
  OAI21_X1 U19950 ( .B1(n17915), .B2(n17914), .A(n17913), .ZN(P2_U2921) );
  AOI22_X1 U19951 ( .A1(n17942), .A2(n17916), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n22262), .ZN(n17917) );
  OAI21_X1 U19952 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22261), .A(n17917), 
        .ZN(P2_U2817) );
  OAI222_X1 U19953 ( .A1(n17939), .A2(n14369), .B1(n17919), .B2(n17942), .C1(
        n17918), .C2(n17936), .ZN(P2_U3212) );
  INV_X1 U19954 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17920) );
  OAI222_X1 U19955 ( .A1(n17939), .A2(n14886), .B1(n17920), .B2(n17942), .C1(
        n14369), .C2(n17936), .ZN(P2_U3213) );
  INV_X1 U19956 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n17921) );
  OAI222_X1 U19957 ( .A1(n17939), .A2(n13333), .B1(n17921), .B2(n17942), .C1(
        n14886), .C2(n17936), .ZN(P2_U3214) );
  INV_X1 U19958 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n17922) );
  OAI222_X1 U19959 ( .A1(n17939), .A2(n12980), .B1(n17922), .B2(n17942), .C1(
        n13333), .C2(n17936), .ZN(P2_U3215) );
  INV_X1 U19960 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n17923) );
  OAI222_X1 U19961 ( .A1(n17939), .A2(n12984), .B1(n17923), .B2(n17942), .C1(
        n12980), .C2(n17936), .ZN(P2_U3216) );
  INV_X1 U19962 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n17924) );
  OAI222_X1 U19963 ( .A1(n17939), .A2(n17347), .B1(n17924), .B2(n17942), .C1(
        n12984), .C2(n17936), .ZN(P2_U3217) );
  INV_X1 U19964 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n17925) );
  OAI222_X1 U19965 ( .A1(n17939), .A2(n13363), .B1(n17925), .B2(n17942), .C1(
        n17347), .C2(n17936), .ZN(P2_U3218) );
  INV_X1 U19966 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n17926) );
  OAI222_X1 U19967 ( .A1(n17939), .A2(n13384), .B1(n17926), .B2(n17942), .C1(
        n13363), .C2(n17936), .ZN(P2_U3219) );
  INV_X1 U19968 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n17927) );
  OAI222_X1 U19969 ( .A1(n17936), .A2(n13384), .B1(n17927), .B2(n17942), .C1(
        n13405), .C2(n17939), .ZN(P2_U3220) );
  INV_X1 U19970 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n17928) );
  OAI222_X1 U19971 ( .A1(n17936), .A2(n13405), .B1(n17928), .B2(n17942), .C1(
        n17322), .C2(n17939), .ZN(P2_U3221) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20413) );
  OAI222_X1 U19973 ( .A1(n17936), .A2(n17322), .B1(n20413), .B2(n17942), .C1(
        n13443), .C2(n17939), .ZN(P2_U3222) );
  INV_X1 U19974 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20415) );
  OAI222_X1 U19975 ( .A1(n17936), .A2(n13443), .B1(n20415), .B2(n17942), .C1(
        n13461), .C2(n17939), .ZN(P2_U3223) );
  INV_X1 U19976 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20417) );
  OAI222_X1 U19977 ( .A1(n17936), .A2(n13461), .B1(n20417), .B2(n17942), .C1(
        n13484), .C2(n17939), .ZN(P2_U3224) );
  INV_X1 U19978 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20419) );
  OAI222_X1 U19979 ( .A1(n17936), .A2(n13484), .B1(n20419), .B2(n17942), .C1(
        n13505), .C2(n17939), .ZN(P2_U3225) );
  INV_X1 U19980 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20421) );
  OAI222_X1 U19981 ( .A1(n17936), .A2(n13505), .B1(n20421), .B2(n17942), .C1(
        n13018), .C2(n17939), .ZN(P2_U3226) );
  INV_X1 U19982 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20423) );
  OAI222_X1 U19983 ( .A1(n17936), .A2(n13018), .B1(n20423), .B2(n17942), .C1(
        n17457), .C2(n17939), .ZN(P2_U3227) );
  INV_X1 U19984 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20425) );
  OAI222_X1 U19985 ( .A1(n17936), .A2(n17457), .B1(n20425), .B2(n17942), .C1(
        n13027), .C2(n17939), .ZN(P2_U3228) );
  INV_X1 U19986 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20427) );
  OAI222_X1 U19987 ( .A1(n17939), .A2(n17929), .B1(n20427), .B2(n17942), .C1(
        n13027), .C2(n17936), .ZN(P2_U3229) );
  INV_X1 U19988 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20429) );
  INV_X1 U19989 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17930) );
  OAI222_X1 U19990 ( .A1(n17936), .A2(n17929), .B1(n20429), .B2(n17942), .C1(
        n17930), .C2(n17939), .ZN(P2_U3230) );
  INV_X1 U19991 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20431) );
  OAI222_X1 U19992 ( .A1(n17939), .A2(n17931), .B1(n20431), .B2(n17942), .C1(
        n17930), .C2(n17936), .ZN(P2_U3231) );
  INV_X1 U19993 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20433) );
  OAI222_X1 U19994 ( .A1(n17939), .A2(n19031), .B1(n20433), .B2(n17942), .C1(
        n17931), .C2(n17936), .ZN(P2_U3232) );
  INV_X1 U19995 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n17932) );
  OAI222_X1 U19996 ( .A1(n17939), .A2(n17933), .B1(n17932), .B2(n17942), .C1(
        n19031), .C2(n17936), .ZN(P2_U3233) );
  INV_X1 U19997 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n17934) );
  OAI222_X1 U19998 ( .A1(n17939), .A2(n14238), .B1(n17934), .B2(n17942), .C1(
        n17933), .C2(n17936), .ZN(P2_U3234) );
  INV_X1 U19999 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20437) );
  OAI222_X1 U20000 ( .A1(n17939), .A2(n19043), .B1(n20437), .B2(n17942), .C1(
        n14238), .C2(n17936), .ZN(P2_U3235) );
  INV_X1 U20001 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20439) );
  OAI222_X1 U20002 ( .A1(n17936), .A2(n19043), .B1(n20439), .B2(n17942), .C1(
        n17246), .C2(n17939), .ZN(P2_U3236) );
  INV_X1 U20003 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20441) );
  OAI222_X1 U20004 ( .A1(n17939), .A2(n17935), .B1(n20441), .B2(n17942), .C1(
        n17246), .C2(n17936), .ZN(P2_U3237) );
  INV_X1 U20005 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20443) );
  OAI222_X1 U20006 ( .A1(n17936), .A2(n17935), .B1(n20443), .B2(n17942), .C1(
        n17219), .C2(n17939), .ZN(P2_U3238) );
  INV_X1 U20007 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20445) );
  OAI222_X1 U20008 ( .A1(n17936), .A2(n17219), .B1(n20445), .B2(n17942), .C1(
        n19060), .C2(n17939), .ZN(P2_U3239) );
  INV_X1 U20009 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20447) );
  OAI222_X1 U20010 ( .A1(n17936), .A2(n19060), .B1(n20447), .B2(n17942), .C1(
        n17937), .C2(n17939), .ZN(P2_U3240) );
  INV_X1 U20011 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20450) );
  OAI222_X1 U20012 ( .A1(n17939), .A2(n17938), .B1(n20450), .B2(n17942), .C1(
        n17937), .C2(n17936), .ZN(P2_U3241) );
  OAI22_X1 U20013 ( .A1(n22262), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17942), .ZN(n17940) );
  INV_X1 U20014 ( .A(n17940), .ZN(P2_U3588) );
  OAI22_X1 U20015 ( .A1(n22262), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17942), .ZN(n17941) );
  INV_X1 U20016 ( .A(n17941), .ZN(P2_U3587) );
  MUX2_X1 U20017 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n22262), .Z(P2_U3586) );
  OAI22_X1 U20018 ( .A1(n22262), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17942), .ZN(n17943) );
  INV_X1 U20019 ( .A(n17943), .ZN(P2_U3585) );
  INV_X1 U20020 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17944) );
  NOR3_X1 U20021 ( .A1(n17944), .A2(n18218), .A3(n17945), .ZN(n17972) );
  NOR2_X1 U20022 ( .A1(n18218), .A2(n17945), .ZN(n17946) );
  OAI21_X1 U20023 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17946), .A(n18214), .ZN(
        n17947) );
  OAI22_X1 U20024 ( .A1(n17972), .A2(n17947), .B1(n18159), .B2(n18214), .ZN(
        P3_U2699) );
  NOR2_X1 U20025 ( .A1(n21290), .A2(n18218), .ZN(n18215) );
  NAND4_X1 U20026 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n18215), .ZN(n17951) );
  INV_X1 U20027 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17949) );
  NAND3_X1 U20028 ( .A1(n17951), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n18214), .ZN(
        n17948) );
  OAI221_X1 U20029 ( .B1(n17951), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n18214), 
        .C2(n17949), .A(n17948), .ZN(P3_U2700) );
  NAND2_X1 U20030 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17950) );
  INV_X1 U20031 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20792) );
  OAI21_X1 U20032 ( .B1(n18218), .B2(n17950), .A(n20792), .ZN(n17952) );
  NAND3_X1 U20033 ( .A1(n18214), .A2(n17952), .A3(n17951), .ZN(n17953) );
  OAI21_X1 U20034 ( .B1(n18214), .B2(n18062), .A(n17953), .ZN(P3_U2701) );
  AOI22_X1 U20035 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17957) );
  AOI22_X1 U20036 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U20037 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U20038 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17954) );
  NAND4_X1 U20039 ( .A1(n17957), .A2(n17956), .A3(n17955), .A4(n17954), .ZN(
        n17963) );
  AOI22_X1 U20040 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17961) );
  AOI22_X1 U20041 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17960) );
  AOI22_X1 U20042 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U20043 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17958) );
  NAND4_X1 U20044 ( .A1(n17961), .A2(n17960), .A3(n17959), .A4(n17958), .ZN(
        n17962) );
  NOR2_X1 U20045 ( .A1(n17963), .A2(n17962), .ZN(n21364) );
  NAND2_X1 U20046 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17972), .ZN(n17971) );
  NOR2_X1 U20047 ( .A1(n17964), .A2(n17971), .ZN(n17965) );
  NAND2_X1 U20048 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17965), .ZN(n18087) );
  OAI21_X1 U20049 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17965), .A(n18087), .ZN(
        n17966) );
  AOI22_X1 U20050 ( .A1(n18219), .A2(n21364), .B1(n17966), .B2(n18214), .ZN(
        P3_U2695) );
  NOR2_X1 U20051 ( .A1(n21290), .A2(n17971), .ZN(n17969) );
  NAND2_X1 U20052 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17969), .ZN(n17968) );
  NAND3_X1 U20053 ( .A1(n17968), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n18214), .ZN(
        n17967) );
  OAI221_X1 U20054 ( .B1(n17968), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n18214), 
        .C2(n18233), .A(n17967), .ZN(P3_U2696) );
  OAI211_X1 U20055 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17969), .A(n17968), .B(
        n18214), .ZN(n17970) );
  OAI21_X1 U20056 ( .B1(n18214), .B2(n18267), .A(n17970), .ZN(P3_U2697) );
  INV_X1 U20057 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17974) );
  OAI21_X1 U20058 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17972), .A(n17971), .ZN(
        n17973) );
  AOI22_X1 U20059 ( .A1(n18219), .A2(n17974), .B1(n17973), .B2(n18214), .ZN(
        P3_U2698) );
  NAND2_X1 U20060 ( .A1(n18002), .A2(n18215), .ZN(n18059) );
  INV_X1 U20061 ( .A(n18059), .ZN(n17975) );
  NAND2_X1 U20062 ( .A1(n17976), .A2(n17975), .ZN(n17999) );
  AOI22_X1 U20063 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17980) );
  AOI22_X1 U20064 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17979) );
  AOI22_X1 U20065 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U20066 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17977) );
  NAND4_X1 U20067 ( .A1(n17980), .A2(n17979), .A3(n17978), .A4(n17977), .ZN(
        n17986) );
  AOI22_X1 U20068 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U20069 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U20070 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U20071 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17981) );
  NAND4_X1 U20072 ( .A1(n17984), .A2(n17983), .A3(n17982), .A4(n17981), .ZN(
        n17985) );
  NOR2_X1 U20073 ( .A1(n17986), .A2(n17985), .ZN(n21343) );
  NAND3_X1 U20074 ( .A1(n17999), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n18214), 
        .ZN(n17987) );
  OAI221_X1 U20075 ( .B1(n17999), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n18214), 
        .C2(n21343), .A(n17987), .ZN(P3_U2687) );
  AOI22_X1 U20076 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U20077 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17990) );
  AOI22_X1 U20078 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17989) );
  AOI22_X1 U20079 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17988) );
  NAND4_X1 U20080 ( .A1(n17991), .A2(n17990), .A3(n17989), .A4(n17988), .ZN(
        n17997) );
  AOI22_X1 U20081 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U20082 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U20083 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17993) );
  AOI22_X1 U20084 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17992) );
  NAND4_X1 U20085 ( .A1(n17995), .A2(n17994), .A3(n17993), .A4(n17992), .ZN(
        n17996) );
  NOR2_X1 U20086 ( .A1(n17997), .A2(n17996), .ZN(n21356) );
  NAND2_X1 U20087 ( .A1(n18217), .A2(n18002), .ZN(n18043) );
  OAI21_X1 U20088 ( .B1(n17998), .B2(n18043), .A(n20971), .ZN(n18000) );
  NAND3_X1 U20089 ( .A1(n18000), .A2(n17999), .A3(n18214), .ZN(n18001) );
  OAI21_X1 U20090 ( .B1(n21356), .B2(n18214), .A(n18001), .ZN(P3_U2688) );
  NAND3_X1 U20091 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18217), .A3(n18002), 
        .ZN(n18016) );
  NAND2_X1 U20092 ( .A1(n18214), .A2(n18016), .ZN(n18045) );
  AOI22_X1 U20093 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U20094 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18014) );
  INV_X1 U20095 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U20096 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18003), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18004) );
  OAI21_X1 U20097 ( .B1(n18006), .B2(n18005), .A(n18004), .ZN(n18012) );
  AOI22_X1 U20098 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U20099 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18051), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U20100 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U20101 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18007) );
  NAND4_X1 U20102 ( .A1(n18010), .A2(n18009), .A3(n18008), .A4(n18007), .ZN(
        n18011) );
  AOI211_X1 U20103 ( .C1(n18244), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n18012), .B(n18011), .ZN(n18013) );
  NAND3_X1 U20104 ( .A1(n18015), .A2(n18014), .A3(n18013), .ZN(n21196) );
  NOR2_X1 U20105 ( .A1(n21290), .A2(n18016), .ZN(n18018) );
  AOI22_X1 U20106 ( .A1(n18219), .A2(n21196), .B1(n18018), .B2(n20948), .ZN(
        n18017) );
  OAI21_X1 U20107 ( .B1(n20948), .B2(n18045), .A(n18017), .ZN(P3_U2690) );
  NAND2_X1 U20108 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18018), .ZN(n18031) );
  AOI22_X1 U20109 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U20110 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18027) );
  AOI22_X1 U20111 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18019) );
  OAI21_X1 U20112 ( .B1(n18063), .B2(n18267), .A(n18019), .ZN(n18025) );
  AOI22_X1 U20113 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U20114 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U20115 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U20116 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18020) );
  NAND4_X1 U20117 ( .A1(n18023), .A2(n18022), .A3(n18021), .A4(n18020), .ZN(
        n18024) );
  AOI211_X1 U20118 ( .C1(n18253), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n18025), .B(n18024), .ZN(n18026) );
  NAND3_X1 U20119 ( .A1(n18028), .A2(n18027), .A3(n18026), .ZN(n21345) );
  INV_X1 U20120 ( .A(n21345), .ZN(n18030) );
  NAND3_X1 U20121 ( .A1(n18031), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n18214), 
        .ZN(n18029) );
  OAI221_X1 U20122 ( .B1(n18031), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n18214), 
        .C2(n18030), .A(n18029), .ZN(P3_U2689) );
  AOI22_X1 U20123 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14064), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U20124 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18035) );
  AOI22_X1 U20125 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18032), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U20126 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18033) );
  NAND4_X1 U20127 ( .A1(n18036), .A2(n18035), .A3(n18034), .A4(n18033), .ZN(
        n18042) );
  AOI22_X1 U20128 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18040) );
  AOI22_X1 U20129 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18039) );
  AOI22_X1 U20130 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U20131 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18037) );
  NAND4_X1 U20132 ( .A1(n18040), .A2(n18039), .A3(n18038), .A4(n18037), .ZN(
        n18041) );
  NOR2_X1 U20133 ( .A1(n18042), .A2(n18041), .ZN(n21200) );
  INV_X1 U20134 ( .A(n18043), .ZN(n18044) );
  NOR2_X1 U20135 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18044), .ZN(n18046) );
  OAI22_X1 U20136 ( .A1(n21200), .A2(n18214), .B1(n18046), .B2(n18045), .ZN(
        P3_U2691) );
  AOI22_X1 U20137 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U20138 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U20139 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U20140 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18047) );
  NAND4_X1 U20141 ( .A1(n18050), .A2(n18049), .A3(n18048), .A4(n18047), .ZN(
        n18057) );
  AOI22_X1 U20142 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18051), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18055) );
  AOI22_X1 U20143 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U20144 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18053) );
  AOI22_X1 U20145 ( .A1(n18245), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18052) );
  NAND4_X1 U20146 ( .A1(n18055), .A2(n18054), .A3(n18053), .A4(n18052), .ZN(
        n18056) );
  NOR2_X1 U20147 ( .A1(n18057), .A2(n18056), .ZN(n21205) );
  OAI21_X1 U20148 ( .B1(n18058), .B2(n18087), .A(n18214), .ZN(n18073) );
  OAI21_X1 U20149 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18073), .A(n18059), .ZN(
        n18060) );
  AOI21_X1 U20150 ( .B1(n18219), .B2(n21205), .A(n18060), .ZN(P3_U2692) );
  AOI22_X1 U20151 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18072) );
  AOI22_X1 U20152 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18071) );
  AOI22_X1 U20153 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18061) );
  OAI21_X1 U20154 ( .B1(n18063), .B2(n18062), .A(n18061), .ZN(n18069) );
  AOI22_X1 U20155 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U20156 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U20157 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U20158 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18064) );
  NAND4_X1 U20159 ( .A1(n18067), .A2(n18066), .A3(n18065), .A4(n18064), .ZN(
        n18068) );
  AOI211_X1 U20160 ( .C1(n18246), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n18069), .B(n18068), .ZN(n18070) );
  NAND3_X1 U20161 ( .A1(n18072), .A2(n18071), .A3(n18070), .ZN(n21209) );
  INV_X1 U20162 ( .A(n21209), .ZN(n18075) );
  NOR2_X1 U20163 ( .A1(n20895), .A2(n18087), .ZN(n18090) );
  NOR2_X1 U20164 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18090), .ZN(n18074) );
  OAI22_X1 U20165 ( .A1(n18075), .A2(n18214), .B1(n18074), .B2(n18073), .ZN(
        P3_U2693) );
  AOI22_X1 U20166 ( .A1(n14064), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U20167 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18271), .B1(
        n18076), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U20168 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20821), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18247), .ZN(n18078) );
  AOI22_X1 U20169 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20808), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18265), .ZN(n18077) );
  NAND4_X1 U20170 ( .A1(n18080), .A2(n18079), .A3(n18078), .A4(n18077), .ZN(
        n18086) );
  AOI22_X1 U20171 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18263), .ZN(n18084) );
  AOI22_X1 U20172 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18245), .ZN(n18083) );
  AOI22_X1 U20173 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18255), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18082) );
  AOI22_X1 U20174 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n11171), .ZN(n18081) );
  NAND4_X1 U20175 ( .A1(n18084), .A2(n18083), .A3(n18082), .A4(n18081), .ZN(
        n18085) );
  NOR2_X1 U20176 ( .A1(n18086), .A2(n18085), .ZN(n21215) );
  AOI21_X1 U20177 ( .B1(n20895), .B2(n18087), .A(n18219), .ZN(n18088) );
  INV_X1 U20178 ( .A(n18088), .ZN(n18089) );
  OAI22_X1 U20179 ( .A1(n21215), .A2(n18214), .B1(n18090), .B2(n18089), .ZN(
        P3_U2694) );
  OAI33_X1 U20180 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21290), .A3(n18092), 
        .B1(n21169), .B2(n18219), .B3(n18091), .ZN(P3_U2672) );
  NAND2_X1 U20181 ( .A1(n21366), .A2(n18093), .ZN(n18106) );
  NAND2_X1 U20182 ( .A1(n18214), .A2(n18094), .ZN(n18172) );
  AOI22_X1 U20183 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U20184 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18097) );
  AOI22_X1 U20185 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U20186 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18095) );
  NAND4_X1 U20187 ( .A1(n18098), .A2(n18097), .A3(n18096), .A4(n18095), .ZN(
        n18104) );
  AOI22_X1 U20188 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18102) );
  AOI22_X1 U20189 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U20190 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18100) );
  AOI22_X1 U20191 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18262), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18099) );
  NAND4_X1 U20192 ( .A1(n18102), .A2(n18101), .A3(n18100), .A4(n18099), .ZN(
        n18103) );
  NOR2_X1 U20193 ( .A1(n18104), .A2(n18103), .ZN(n21255) );
  OR2_X1 U20194 ( .A1(n21255), .A2(n18214), .ZN(n18105) );
  OAI221_X1 U20195 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18106), .C1(n21046), 
        .C2(n18172), .A(n18105), .ZN(P3_U2682) );
  NOR2_X1 U20196 ( .A1(n21046), .A2(n18106), .ZN(n18144) );
  NAND2_X1 U20197 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18144), .ZN(n18138) );
  NAND2_X1 U20198 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18143), .ZN(n18128) );
  NAND2_X1 U20199 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18132), .ZN(n18126) );
  OAI21_X1 U20200 ( .B1(n18123), .B2(n18107), .A(n18116), .ZN(n21325) );
  NAND3_X1 U20201 ( .A1(n18126), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18214), 
        .ZN(n18108) );
  OAI221_X1 U20202 ( .B1(n18126), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18214), 
        .C2(n21325), .A(n18108), .ZN(P3_U2676) );
  OAI21_X1 U20203 ( .B1(n18115), .B2(n18110), .A(n18109), .ZN(n21313) );
  INV_X1 U20204 ( .A(n18215), .ZN(n18221) );
  NAND2_X1 U20205 ( .A1(n18214), .A2(n18126), .ZN(n18111) );
  OAI21_X1 U20206 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18221), .A(n18111), .ZN(
        n18118) );
  OAI221_X1 U20207 ( .B1(n18118), .B2(n18215), .C1(n18118), .C2(n18119), .A(
        P3_EBX_REG_29__SCAN_IN), .ZN(n18114) );
  INV_X1 U20208 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21140) );
  NAND3_X1 U20209 ( .A1(n21366), .A2(n18112), .A3(n21140), .ZN(n18113) );
  OAI211_X1 U20210 ( .C1(n18214), .C2(n21313), .A(n18114), .B(n18113), .ZN(
        P3_U2674) );
  AOI21_X1 U20211 ( .B1(n18117), .B2(n18116), .A(n18115), .ZN(n21314) );
  AOI22_X1 U20212 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18118), .B1(n21314), 
        .B2(n18219), .ZN(n18121) );
  NAND4_X1 U20213 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n18132), .A4(n18119), .ZN(n18120) );
  NAND2_X1 U20214 ( .A1(n18121), .A2(n18120), .ZN(P3_U2675) );
  AOI21_X1 U20215 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18214), .A(n18132), .ZN(
        n18122) );
  INV_X1 U20216 ( .A(n18122), .ZN(n18125) );
  AOI21_X1 U20217 ( .B1(n18124), .B2(n18129), .A(n18123), .ZN(n21295) );
  AOI22_X1 U20218 ( .A1(n18126), .A2(n18125), .B1(n21295), .B2(n18219), .ZN(
        n18127) );
  INV_X1 U20219 ( .A(n18127), .ZN(P3_U2677) );
  INV_X1 U20220 ( .A(n18128), .ZN(n18137) );
  AOI21_X1 U20221 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18214), .A(n18137), .ZN(
        n18131) );
  OAI21_X1 U20222 ( .B1(n18133), .B2(n18130), .A(n18129), .ZN(n21294) );
  OAI22_X1 U20223 ( .A1(n18132), .A2(n18131), .B1(n21294), .B2(n18214), .ZN(
        P3_U2678) );
  AOI21_X1 U20224 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18214), .A(n18143), .ZN(
        n18136) );
  AOI21_X1 U20225 ( .B1(n18134), .B2(n18139), .A(n18133), .ZN(n21326) );
  INV_X1 U20226 ( .A(n21326), .ZN(n18135) );
  OAI22_X1 U20227 ( .A1(n18137), .A2(n18136), .B1(n18214), .B2(n18135), .ZN(
        P3_U2679) );
  INV_X1 U20228 ( .A(n18138), .ZN(n18156) );
  AOI21_X1 U20229 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18214), .A(n18156), .ZN(
        n18142) );
  OAI21_X1 U20230 ( .B1(n18141), .B2(n18140), .A(n18139), .ZN(n21337) );
  OAI22_X1 U20231 ( .A1(n18143), .A2(n18142), .B1(n18214), .B2(n21337), .ZN(
        P3_U2680) );
  AOI21_X1 U20232 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18214), .A(n18144), .ZN(
        n18155) );
  AOI22_X1 U20233 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18148) );
  AOI22_X1 U20234 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18147) );
  AOI22_X1 U20235 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18146) );
  AOI22_X1 U20236 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18145) );
  NAND4_X1 U20237 ( .A1(n18148), .A2(n18147), .A3(n18146), .A4(n18145), .ZN(
        n18154) );
  AOI22_X1 U20238 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20239 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U20240 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20241 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18149) );
  NAND4_X1 U20242 ( .A1(n18152), .A2(n18151), .A3(n18150), .A4(n18149), .ZN(
        n18153) );
  NOR2_X1 U20243 ( .A1(n18154), .A2(n18153), .ZN(n21266) );
  OAI22_X1 U20244 ( .A1(n18156), .A2(n18155), .B1(n21266), .B2(n18214), .ZN(
        P3_U2681) );
  AOI22_X1 U20245 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18169) );
  AOI22_X1 U20246 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U20247 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18158) );
  OAI21_X1 U20248 ( .B1(n18160), .B2(n18159), .A(n18158), .ZN(n18166) );
  AOI22_X1 U20249 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18164) );
  AOI22_X1 U20250 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18245), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18163) );
  AOI22_X1 U20251 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U20252 ( .A1(n20808), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18161) );
  NAND4_X1 U20253 ( .A1(n18164), .A2(n18163), .A3(n18162), .A4(n18161), .ZN(
        n18165) );
  AOI211_X1 U20254 ( .C1(n18272), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n18166), .B(n18165), .ZN(n18167) );
  NAND3_X1 U20255 ( .A1(n18169), .A2(n18168), .A3(n18167), .ZN(n21260) );
  NAND2_X1 U20256 ( .A1(n18219), .A2(n21260), .ZN(n18170) );
  OAI221_X1 U20257 ( .B1(n18172), .B2(n18171), .C1(n18172), .C2(n18196), .A(
        n18170), .ZN(P3_U2683) );
  AOI22_X1 U20258 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U20259 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18175) );
  AOI22_X1 U20260 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U20261 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18173) );
  NAND4_X1 U20262 ( .A1(n18176), .A2(n18175), .A3(n18174), .A4(n18173), .ZN(
        n18182) );
  AOI22_X1 U20263 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18245), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U20264 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18179) );
  AOI22_X1 U20265 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18178) );
  AOI22_X1 U20266 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18177) );
  NAND4_X1 U20267 ( .A1(n18180), .A2(n18179), .A3(n18178), .A4(n18177), .ZN(
        n18181) );
  NOR2_X1 U20268 ( .A1(n18182), .A2(n18181), .ZN(n21281) );
  OAI211_X1 U20269 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18210), .A(n18215), .B(
        n18183), .ZN(n18185) );
  NAND2_X1 U20270 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18218), .ZN(n18184) );
  OAI211_X1 U20271 ( .C1(n21281), .C2(n18214), .A(n18185), .B(n18184), .ZN(
        P3_U2685) );
  AOI22_X1 U20272 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18189) );
  AOI22_X1 U20273 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U20274 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n20808), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U20275 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18199), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18186) );
  NAND4_X1 U20276 ( .A1(n18189), .A2(n18188), .A3(n18187), .A4(n18186), .ZN(
        n18195) );
  AOI22_X1 U20277 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18193) );
  AOI22_X1 U20278 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U20279 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18246), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U20280 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18190) );
  NAND4_X1 U20281 ( .A1(n18193), .A2(n18192), .A3(n18191), .A4(n18190), .ZN(
        n18194) );
  NOR2_X1 U20282 ( .A1(n18195), .A2(n18194), .ZN(n21277) );
  OAI21_X1 U20283 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18197), .A(n18196), .ZN(
        n18198) );
  AOI22_X1 U20284 ( .A1(n18219), .A2(n21277), .B1(n18198), .B2(n18214), .ZN(
        P3_U2684) );
  AOI22_X1 U20285 ( .A1(n11172), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18245), .ZN(n18203) );
  AOI22_X1 U20286 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U20287 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20808), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18199), .ZN(n18201) );
  AOI22_X1 U20288 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21408), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n20821), .ZN(n18200) );
  NAND4_X1 U20289 ( .A1(n18203), .A2(n18202), .A3(n18201), .A4(n18200), .ZN(
        n18209) );
  AOI22_X1 U20290 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11171), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18254), .ZN(n18207) );
  AOI22_X1 U20291 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U20292 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18246), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U20293 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18204) );
  NAND4_X1 U20294 ( .A1(n18207), .A2(n18206), .A3(n18205), .A4(n18204), .ZN(
        n18208) );
  NOR2_X1 U20295 ( .A1(n18209), .A2(n18208), .ZN(n21287) );
  AOI211_X1 U20296 ( .C1(n21006), .C2(n18211), .A(n18210), .B(n18221), .ZN(
        n18212) );
  AOI21_X1 U20297 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18218), .A(n18212), .ZN(
        n18213) );
  OAI21_X1 U20298 ( .B1(n21287), .B2(n18214), .A(n18213), .ZN(P3_U2686) );
  INV_X1 U20299 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20780) );
  NOR2_X1 U20300 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20793) );
  AOI21_X1 U20301 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20793), .ZN(n20779) );
  AOI22_X1 U20302 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18219), .B1(
        n18215), .B2(n20779), .ZN(n18216) );
  OAI21_X1 U20303 ( .B1(n18217), .B2(n20780), .A(n18216), .ZN(P3_U2702) );
  AOI22_X1 U20304 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18219), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18218), .ZN(n18220) );
  OAI21_X1 U20305 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18221), .A(n18220), .ZN(
        P3_U2703) );
  AOI21_X1 U20306 ( .B1(n18224), .B2(n18223), .A(n18222), .ZN(n21843) );
  INV_X1 U20307 ( .A(n21843), .ZN(n18225) );
  OAI21_X1 U20308 ( .B1(n21897), .B2(n18225), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18226) );
  OAI21_X1 U20309 ( .B1(n18227), .B2(n20715), .A(n18226), .ZN(P3_U2634) );
  INV_X1 U20310 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21901) );
  AOI21_X1 U20311 ( .B1(n21901), .B2(n18229), .A(n18228), .ZN(n21891) );
  OAI21_X1 U20312 ( .B1(n21891), .B2(n19280), .A(n18231), .ZN(n18230) );
  OAI221_X1 U20313 ( .B1(n21852), .B2(n20717), .C1(n21852), .C2(n18231), .A(
        n18230), .ZN(P3_U2863) );
  INV_X1 U20314 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18602) );
  INV_X1 U20315 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18393) );
  INV_X1 U20316 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21791) );
  INV_X1 U20317 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21790) );
  INV_X1 U20318 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21825) );
  INV_X1 U20319 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18621) );
  NOR2_X1 U20320 ( .A1(n21825), .A2(n18621), .ZN(n21524) );
  NOR3_X1 U20321 ( .A1(n21791), .A2(n21790), .A3(n21525), .ZN(n18380) );
  INV_X1 U20322 ( .A(n18380), .ZN(n21543) );
  NOR2_X1 U20323 ( .A1(n18393), .A2(n21543), .ZN(n21558) );
  INV_X1 U20324 ( .A(n21558), .ZN(n21555) );
  NOR2_X1 U20325 ( .A1(n18602), .A2(n21555), .ZN(n21568) );
  NAND2_X1 U20326 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21568), .ZN(
        n21755) );
  AOI22_X1 U20327 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U20328 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U20329 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18232) );
  OAI21_X1 U20330 ( .B1(n18268), .B2(n18233), .A(n18232), .ZN(n18240) );
  AOI22_X1 U20331 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18238) );
  AOI22_X1 U20332 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U20333 ( .A1(n18234), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18236) );
  AOI22_X1 U20334 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18235) );
  NAND4_X1 U20335 ( .A1(n18238), .A2(n18237), .A3(n18236), .A4(n18235), .ZN(
        n18239) );
  AOI211_X1 U20336 ( .C1(n18279), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n18240), .B(n18239), .ZN(n18241) );
  NAND3_X1 U20337 ( .A1(n18243), .A2(n18242), .A3(n18241), .ZN(n18332) );
  AOI22_X1 U20338 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U20339 ( .A1(n18246), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18245), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U20340 ( .A1(n20821), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18250) );
  AOI22_X1 U20341 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18247), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18249) );
  NAND4_X1 U20342 ( .A1(n18252), .A2(n18251), .A3(n18250), .A4(n18249), .ZN(
        n18261) );
  AOI22_X1 U20343 ( .A1(n18051), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U20344 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18253), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U20345 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20346 ( .A1(n18255), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18256) );
  NAND4_X1 U20347 ( .A1(n18259), .A2(n18258), .A3(n18257), .A4(n18256), .ZN(
        n18260) );
  NAND3_X1 U20348 ( .A1(n18314), .A2(n18316), .A3(n18290), .ZN(n18284) );
  AOI22_X1 U20349 ( .A1(n18262), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18234), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18282) );
  AOI22_X1 U20350 ( .A1(n18264), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18263), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20351 ( .A1(n21408), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18265), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18266) );
  OAI21_X1 U20352 ( .B1(n18268), .B2(n18267), .A(n18266), .ZN(n18278) );
  AOI22_X1 U20353 ( .A1(n18270), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U20354 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14088), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U20355 ( .A1(n18272), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11171), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U20356 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11172), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18273) );
  NAND4_X1 U20357 ( .A1(n18276), .A2(n18275), .A3(n18274), .A4(n18273), .ZN(
        n18277) );
  AOI211_X1 U20358 ( .C1(n18279), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n18278), .B(n18277), .ZN(n18280) );
  NOR2_X1 U20359 ( .A1(n18284), .A2(n21225), .ZN(n18283) );
  AND2_X1 U20360 ( .A1(n18332), .A2(n18283), .ZN(n18304) );
  XOR2_X1 U20361 ( .A(n18332), .B(n18283), .Z(n18300) );
  XOR2_X1 U20362 ( .A(n21225), .B(n18284), .Z(n18296) );
  INV_X1 U20363 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21426) );
  NAND2_X1 U20364 ( .A1(n18314), .A2(n18290), .ZN(n18291) );
  XOR2_X1 U20365 ( .A(n18291), .B(n18316), .Z(n18687) );
  NAND2_X1 U20366 ( .A1(n18296), .A2(n18297), .ZN(n18298) );
  XOR2_X1 U20367 ( .A(n18297), .B(n18296), .Z(n18675) );
  NAND2_X1 U20368 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18675), .ZN(
        n18674) );
  NAND2_X1 U20369 ( .A1(n18298), .A2(n18674), .ZN(n18301) );
  NOR2_X1 U20370 ( .A1(n18300), .A2(n18301), .ZN(n18664) );
  INV_X1 U20371 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21431) );
  NAND2_X1 U20372 ( .A1(n18304), .A2(n18299), .ZN(n18305) );
  INV_X1 U20373 ( .A(n18299), .ZN(n18303) );
  AND2_X1 U20374 ( .A1(n18301), .A2(n18300), .ZN(n18665) );
  AOI21_X1 U20375 ( .B1(n18304), .B2(n18303), .A(n18665), .ZN(n18302) );
  NAND2_X1 U20376 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18648), .ZN(
        n18647) );
  NAND2_X2 U20377 ( .A1(n18305), .A2(n18647), .ZN(n21520) );
  NAND3_X1 U20378 ( .A1(n18314), .A2(n18316), .A3(n18313), .ZN(n18308) );
  INV_X1 U20379 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21492) );
  XNOR2_X1 U20380 ( .A(n21225), .B(n18308), .ZN(n18321) );
  XOR2_X1 U20381 ( .A(n21492), .B(n18321), .Z(n18680) );
  AOI22_X1 U20382 ( .A1(n18311), .A2(n18310), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18309), .ZN(n18312) );
  NAND2_X1 U20383 ( .A1(n18314), .A2(n18313), .ZN(n18315) );
  XNOR2_X1 U20384 ( .A(n18316), .B(n18315), .ZN(n18319) );
  NAND2_X1 U20385 ( .A1(n18319), .A2(n18318), .ZN(n18320) );
  NAND2_X1 U20386 ( .A1(n18680), .A2(n18679), .ZN(n18678) );
  NAND2_X2 U20387 ( .A1(n18678), .A2(n18322), .ZN(n18356) );
  AOI21_X1 U20388 ( .B1(n21439), .B2(n21705), .A(n18511), .ZN(n18324) );
  NAND2_X1 U20389 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18668), .ZN(
        n18667) );
  NAND2_X1 U20390 ( .A1(n18324), .A2(n18356), .ZN(n18325) );
  NAND2_X2 U20391 ( .A1(n18667), .A2(n18325), .ZN(n18657) );
  NOR2_X1 U20392 ( .A1(n18511), .A2(n18657), .ZN(n18357) );
  INV_X1 U20393 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21817) );
  NOR2_X4 U20394 ( .A1(n18332), .A2(n18739), .ZN(n18660) );
  INV_X1 U20395 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21770) );
  INV_X1 U20396 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21780) );
  NOR2_X1 U20397 ( .A1(n21770), .A2(n21780), .ZN(n21759) );
  INV_X1 U20398 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18349) );
  NAND2_X1 U20399 ( .A1(n21759), .A2(n18349), .ZN(n21769) );
  OAI21_X1 U20400 ( .B1(n18576), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n18327), .ZN(n21012) );
  INV_X1 U20401 ( .A(n21012), .ZN(n21015) );
  INV_X1 U20402 ( .A(n18744), .ZN(n18536) );
  INV_X1 U20403 ( .A(n18576), .ZN(n18328) );
  OAI21_X1 U20404 ( .B1(n21014), .B2(n18702), .A(n18745), .ZN(n18582) );
  AOI21_X1 U20405 ( .B1(n18536), .B2(n18328), .A(n18582), .ZN(n18344) );
  INV_X1 U20406 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18330) );
  INV_X1 U20407 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20782) );
  NAND3_X1 U20408 ( .A1(n21014), .A2(n18330), .A3(n18534), .ZN(n18343) );
  INV_X2 U20409 ( .A(n21808), .ZN(n21832) );
  NAND2_X1 U20410 ( .A1(n21832), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18329) );
  OAI211_X1 U20411 ( .C1(n18344), .C2(n18330), .A(n18343), .B(n18329), .ZN(
        n18331) );
  AOI21_X1 U20412 ( .B1(n18570), .B2(n21015), .A(n18331), .ZN(n18341) );
  INV_X1 U20413 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21577) );
  NAND2_X1 U20414 ( .A1(n21558), .A2(n21520), .ZN(n18599) );
  NOR2_X2 U20415 ( .A1(n18602), .A2(n18599), .ZN(n21572) );
  AOI22_X1 U20416 ( .A1(n18660), .A2(n11152), .B1(n18700), .B2(n21732), .ZN(
        n18373) );
  OAI21_X1 U20417 ( .B1(n21759), .B2(n18523), .A(n18373), .ZN(n18585) );
  NAND2_X1 U20418 ( .A1(n18332), .A2(n18704), .ZN(n18634) );
  NOR2_X1 U20419 ( .A1(n18511), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18432) );
  AOI21_X1 U20420 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18511), .A(
        n18432), .ZN(n18339) );
  NAND2_X1 U20421 ( .A1(n21825), .A2(n18621), .ZN(n18631) );
  NOR3_X1 U20422 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n18631), .ZN(n18390) );
  AOI22_X1 U20423 ( .A1(n18511), .A2(n21817), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18619), .ZN(n18658) );
  AOI21_X1 U20424 ( .B1(n18390), .B2(n18333), .A(n18511), .ZN(n18338) );
  INV_X1 U20425 ( .A(n18338), .ZN(n18334) );
  INV_X1 U20426 ( .A(n21755), .ZN(n21751) );
  NAND2_X1 U20427 ( .A1(n21751), .A2(n18623), .ZN(n18335) );
  NAND2_X1 U20428 ( .A1(n18334), .A2(n18335), .ZN(n18459) );
  NAND2_X1 U20429 ( .A1(n21759), .A2(n18459), .ZN(n18348) );
  NOR2_X2 U20430 ( .A1(n18338), .A2(n18337), .ZN(n18584) );
  XNOR2_X1 U20432 ( .A(n18339), .B(n18404), .ZN(n21752) );
  AOI22_X1 U20433 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18585), .B1(
        n18661), .B2(n21752), .ZN(n18340) );
  OAI211_X1 U20434 ( .C1(n18523), .C2(n21769), .A(n18341), .B(n18340), .ZN(
        P3_U2812) );
  NAND2_X1 U20435 ( .A1(n21759), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21428) );
  INV_X1 U20436 ( .A(n21428), .ZN(n21429) );
  NAND2_X1 U20437 ( .A1(n21429), .A2(n18586), .ZN(n18438) );
  NOR3_X1 U20438 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18486), .A3(
        n18399), .ZN(n18346) );
  NAND2_X1 U20439 ( .A1(n21832), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18342) );
  OAI221_X1 U20440 ( .B1(n18400), .B2(n18344), .C1(n18400), .C2(n18343), .A(
        n18342), .ZN(n18345) );
  AOI211_X1 U20441 ( .C1(n21028), .C2(n18570), .A(n18346), .B(n18345), .ZN(
        n18352) );
  NAND2_X1 U20442 ( .A1(n21429), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21731) );
  NOR2_X1 U20443 ( .A1(n11152), .A2(n21731), .ZN(n21736) );
  NOR2_X1 U20444 ( .A1(n21732), .A2(n21731), .ZN(n18347) );
  OAI22_X1 U20445 ( .A1(n21736), .A2(n18612), .B1(n18347), .B2(n18734), .ZN(
        n18435) );
  INV_X1 U20446 ( .A(n18432), .ZN(n18403) );
  NOR2_X1 U20447 ( .A1(n18403), .A2(n18404), .ZN(n18418) );
  NOR3_X1 U20448 ( .A1(n18619), .A2(n18349), .A3(n18348), .ZN(n18431) );
  NOR2_X1 U20449 ( .A1(n18418), .A2(n18431), .ZN(n18350) );
  INV_X1 U20450 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21741) );
  XOR2_X1 U20451 ( .A(n18350), .B(n21741), .Z(n21739) );
  AOI22_X1 U20452 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18435), .B1(
        n18661), .B2(n21739), .ZN(n18351) );
  OAI211_X1 U20453 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18438), .A(
        n18352), .B(n18351), .ZN(P3_U2811) );
  AOI21_X1 U20454 ( .B1(n21572), .B2(n18700), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18363) );
  INV_X1 U20455 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20976) );
  INV_X1 U20456 ( .A(n18353), .ZN(n18354) );
  NAND2_X1 U20457 ( .A1(n18354), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18592) );
  INV_X1 U20458 ( .A(n18592), .ZN(n18365) );
  XNOR2_X1 U20459 ( .A(n20976), .B(n18365), .ZN(n20981) );
  NAND2_X1 U20460 ( .A1(n18354), .A2(n18534), .ZN(n18368) );
  OAI21_X1 U20461 ( .B1(n18354), .B2(n18702), .A(n18745), .ZN(n18598) );
  AOI21_X1 U20462 ( .B1(n18536), .B2(n18592), .A(n18598), .ZN(n18369) );
  NAND2_X1 U20463 ( .A1(n21832), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21581) );
  OAI221_X1 U20464 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18368), .C1(
        n20976), .C2(n18369), .A(n21581), .ZN(n18361) );
  NOR2_X1 U20465 ( .A1(n21817), .A2(n21431), .ZN(n18355) );
  NAND3_X1 U20466 ( .A1(n18356), .A2(n18511), .A3(n18355), .ZN(n18640) );
  INV_X1 U20467 ( .A(n18640), .ZN(n18620) );
  NAND2_X1 U20468 ( .A1(n21558), .A2(n18620), .ZN(n18600) );
  NAND2_X1 U20469 ( .A1(n18357), .A2(n21817), .ZN(n18641) );
  INV_X1 U20470 ( .A(n18641), .ZN(n18389) );
  NAND3_X1 U20471 ( .A1(n18390), .A2(n18389), .A3(n18393), .ZN(n18601) );
  AOI22_X1 U20472 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18600), .B1(
        n18601), .B2(n18602), .ZN(n18358) );
  XOR2_X1 U20473 ( .A(n21577), .B(n18358), .Z(n21583) );
  NAND2_X1 U20474 ( .A1(n18660), .A2(n11152), .ZN(n18359) );
  OAI22_X1 U20475 ( .A1(n21583), .A2(n18634), .B1(n21575), .B2(n18359), .ZN(
        n18360) );
  AOI211_X1 U20476 ( .C1(n18570), .C2(n20981), .A(n18361), .B(n18360), .ZN(
        n18362) );
  OAI21_X1 U20477 ( .B1(n18373), .B2(n18363), .A(n18362), .ZN(P3_U2815) );
  AOI22_X1 U20478 ( .A1(n18511), .A2(n21780), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18619), .ZN(n18364) );
  XOR2_X1 U20479 ( .A(n18459), .B(n18364), .Z(n21785) );
  OAI221_X1 U20480 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18365), .A(n18578), .ZN(
        n20990) );
  OAI21_X1 U20481 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18366), .ZN(n18367) );
  OAI22_X1 U20482 ( .A1(n18580), .A2(n20990), .B1(n18368), .B2(n18367), .ZN(
        n18371) );
  INV_X1 U20483 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20997) );
  NAND2_X1 U20484 ( .A1(n21832), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n21786) );
  OAI21_X1 U20485 ( .B1(n18369), .B2(n20997), .A(n21786), .ZN(n18370) );
  AOI211_X1 U20486 ( .C1(n18661), .C2(n21785), .A(n18371), .B(n18370), .ZN(
        n18372) );
  OAI221_X1 U20487 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18523), 
        .C1(n21780), .C2(n18373), .A(n18372), .ZN(P3_U2814) );
  NOR2_X1 U20488 ( .A1(n18631), .A2(n18641), .ZN(n18613) );
  NOR2_X1 U20489 ( .A1(n21791), .A2(n21525), .ZN(n21546) );
  INV_X1 U20490 ( .A(n21546), .ZN(n18379) );
  NOR3_X1 U20491 ( .A1(n18619), .A2(n11145), .A3(n18379), .ZN(n18391) );
  AOI21_X1 U20492 ( .B1(n18613), .B2(n21791), .A(n18391), .ZN(n18375) );
  XOR2_X1 U20493 ( .A(n18375), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n21552) );
  CLKBUF_X1 U20494 ( .A(n18376), .Z(n18594) );
  NAND2_X1 U20495 ( .A1(n18594), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18378) );
  INV_X1 U20496 ( .A(n18378), .ZN(n18609) );
  NAND2_X1 U20497 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18609), .ZN(
        n18590) );
  OAI21_X1 U20498 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18609), .A(
        n18590), .ZN(n20937) );
  INV_X1 U20499 ( .A(n20937), .ZN(n20939) );
  NAND2_X1 U20500 ( .A1(n18594), .A2(n18534), .ZN(n18386) );
  INV_X1 U20501 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20943) );
  OAI21_X1 U20502 ( .B1(n18594), .B2(n18702), .A(n18745), .ZN(n18377) );
  AOI21_X1 U20503 ( .B1(n18536), .B2(n18378), .A(n18377), .ZN(n18398) );
  NAND2_X1 U20504 ( .A1(n21832), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21550) );
  OAI221_X1 U20505 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18386), .C1(
        n20943), .C2(n18398), .A(n21550), .ZN(n18384) );
  NOR2_X1 U20506 ( .A1(n18646), .A2(n18379), .ZN(n18382) );
  NAND2_X1 U20507 ( .A1(n21520), .A2(n18380), .ZN(n21538) );
  AOI22_X1 U20508 ( .A1(n18700), .A2(n21538), .B1(n18660), .B2(n21542), .ZN(
        n18394) );
  INV_X1 U20509 ( .A(n18394), .ZN(n18381) );
  MUX2_X1 U20510 ( .A(n18382), .B(n18381), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18383) );
  AOI211_X1 U20511 ( .C1(n18570), .C2(n20939), .A(n18384), .B(n18383), .ZN(
        n18385) );
  OAI21_X1 U20512 ( .B1(n21552), .B2(n18634), .A(n18385), .ZN(P3_U2818) );
  INV_X1 U20513 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18591) );
  INV_X1 U20514 ( .A(n18590), .ZN(n20952) );
  AOI22_X1 U20515 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20952), .B1(
        n18590), .B2(n18591), .ZN(n20951) );
  AOI211_X1 U20516 ( .C1(n20943), .C2(n18591), .A(n20975), .B(n18386), .ZN(
        n18388) );
  NOR2_X1 U20517 ( .A1(n21808), .A2(n20954), .ZN(n18387) );
  AOI211_X1 U20518 ( .C1(n18570), .C2(n20951), .A(n18388), .B(n18387), .ZN(
        n18397) );
  NOR2_X1 U20519 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21543), .ZN(
        n21789) );
  INV_X1 U20520 ( .A(n18646), .ZN(n18630) );
  AOI22_X1 U20521 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18391), .B1(
        n18390), .B2(n18389), .ZN(n18392) );
  XOR2_X1 U20522 ( .A(n18392), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n21799) );
  OAI22_X1 U20523 ( .A1(n21799), .A2(n18634), .B1(n18394), .B2(n18393), .ZN(
        n18395) );
  AOI21_X1 U20524 ( .B1(n21789), .B2(n18630), .A(n18395), .ZN(n18396) );
  OAI211_X1 U20525 ( .C1(n18398), .C2(n18591), .A(n18397), .B(n18396), .ZN(
        P3_U2817) );
  NOR2_X1 U20526 ( .A1(n18400), .A2(n18399), .ZN(n18425) );
  NAND2_X1 U20527 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18425), .ZN(
        n18439) );
  OAI21_X1 U20528 ( .B1(n18401), .B2(n18744), .A(n18745), .ZN(n18402) );
  AOI21_X1 U20529 ( .B1(n18653), .B2(n18439), .A(n18402), .ZN(n18427) );
  OAI21_X1 U20530 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18579), .A(
        n18427), .ZN(n18415) );
  AOI22_X1 U20531 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18415), .B1(
        n18570), .B2(n21056), .ZN(n18412) );
  INV_X1 U20532 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21588) );
  NOR4_X1 U20533 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n18403), .ZN(n18448) );
  INV_X1 U20534 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18434) );
  NOR2_X1 U20535 ( .A1(n18434), .A2(n21741), .ZN(n21437) );
  NAND2_X1 U20536 ( .A1(n21437), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21589) );
  INV_X1 U20537 ( .A(n21589), .ZN(n18406) );
  NAND3_X1 U20538 ( .A1(n18406), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18404), .ZN(n18467) );
  INV_X1 U20539 ( .A(n18467), .ZN(n18405) );
  OAI21_X1 U20540 ( .B1(n18448), .B2(n18405), .A(n18466), .ZN(n18449) );
  XOR2_X1 U20541 ( .A(n21588), .B(n18449), .Z(n21584) );
  NAND2_X1 U20542 ( .A1(n21429), .A2(n18406), .ZN(n18460) );
  NOR2_X1 U20543 ( .A1(n18460), .A2(n18523), .ZN(n18408) );
  NOR2_X2 U20544 ( .A1(n18460), .A2(n11152), .ZN(n21434) );
  INV_X1 U20545 ( .A(n21434), .ZN(n18443) );
  NOR2_X2 U20546 ( .A1(n21732), .A2(n18460), .ZN(n18447) );
  INV_X1 U20547 ( .A(n18447), .ZN(n21436) );
  AOI22_X1 U20548 ( .A1(n18660), .A2(n18443), .B1(n18700), .B2(n21436), .ZN(
        n18424) );
  INV_X1 U20549 ( .A(n18424), .ZN(n18407) );
  MUX2_X1 U20550 ( .A(n18408), .B(n18407), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18409) );
  AOI21_X1 U20551 ( .B1(n18661), .B2(n21584), .A(n18409), .ZN(n18411) );
  NAND2_X1 U20552 ( .A1(n21832), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21594) );
  NOR2_X1 U20553 ( .A1(n18486), .A2(n18439), .ZN(n18417) );
  OAI211_X1 U20554 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18417), .B(n18440), .ZN(n18410) );
  NAND4_X1 U20555 ( .A1(n18412), .A2(n18411), .A3(n21594), .A4(n18410), .ZN(
        P3_U2808) );
  INV_X1 U20556 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18423) );
  INV_X1 U20557 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21445) );
  OAI22_X1 U20558 ( .A1(n21808), .A2(n21445), .B1(n18580), .B2(n18413), .ZN(
        n18414) );
  AOI221_X1 U20559 ( .B1(n18417), .B2(n18416), .C1(n18415), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18414), .ZN(n18422) );
  NOR2_X1 U20560 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18419) );
  AOI22_X1 U20561 ( .A1(n21437), .A2(n18431), .B1(n18419), .B2(n18418), .ZN(
        n18420) );
  XOR2_X1 U20562 ( .A(n18423), .B(n18420), .Z(n21443) );
  AND2_X1 U20563 ( .A1(n18423), .A2(n21437), .ZN(n21442) );
  INV_X1 U20564 ( .A(n18438), .ZN(n18480) );
  AOI22_X1 U20565 ( .A1(n18661), .A2(n21443), .B1(n21442), .B2(n18480), .ZN(
        n18421) );
  OAI211_X1 U20566 ( .C1(n18424), .C2(n18423), .A(n18422), .B(n18421), .ZN(
        P3_U2809) );
  NAND2_X1 U20567 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18434), .ZN(
        n21750) );
  INV_X1 U20568 ( .A(n18579), .ZN(n18429) );
  AOI21_X1 U20569 ( .B1(n18425), .B2(n19606), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18426) );
  NAND2_X1 U20570 ( .A1(n21832), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21747) );
  OAI21_X1 U20571 ( .B1(n18427), .B2(n18426), .A(n21747), .ZN(n18428) );
  AOI221_X1 U20572 ( .B1(n18570), .B2(n18430), .C1(n18429), .C2(n18430), .A(
        n18428), .ZN(n18437) );
  OAI221_X1 U20573 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18432), 
        .C1(n21741), .C2(n18431), .A(n18466), .ZN(n18433) );
  XOR2_X1 U20574 ( .A(n18434), .B(n18433), .Z(n21745) );
  AOI22_X1 U20575 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18435), .B1(
        n18661), .B2(n21745), .ZN(n18436) );
  OAI211_X1 U20576 ( .C1(n18438), .C2(n21750), .A(n18437), .B(n18436), .ZN(
        P3_U2810) );
  NOR2_X1 U20577 ( .A1(n18440), .A2(n18439), .ZN(n18453) );
  NAND2_X1 U20578 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18453), .ZN(
        n18484) );
  INV_X1 U20579 ( .A(n18745), .ZN(n18728) );
  AOI21_X1 U20580 ( .B1(n19606), .B2(n18484), .A(n18728), .ZN(n18457) );
  OAI21_X1 U20581 ( .B1(n18441), .B2(n18744), .A(n18457), .ZN(n18442) );
  AOI22_X1 U20582 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18442), .B1(
        n18570), .B2(n21072), .ZN(n18456) );
  NAND2_X1 U20583 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18479) );
  NOR2_X2 U20584 ( .A1(n18479), .A2(n18443), .ZN(n21716) );
  INV_X1 U20585 ( .A(n18479), .ZN(n18462) );
  NAND2_X1 U20586 ( .A1(n18462), .A2(n18447), .ZN(n21714) );
  NAND2_X1 U20587 ( .A1(n18700), .A2(n21714), .ZN(n18444) );
  OAI21_X1 U20588 ( .B1(n21716), .B2(n18612), .A(n18444), .ZN(n18481) );
  INV_X1 U20589 ( .A(n18444), .ZN(n18446) );
  NOR2_X1 U20590 ( .A1(n21716), .A2(n18612), .ZN(n18445) );
  AOI22_X1 U20591 ( .A1(n18447), .A2(n18446), .B1(n21434), .B2(n18445), .ZN(
        n18451) );
  NAND2_X1 U20592 ( .A1(n18448), .A2(n21588), .ZN(n18463) );
  AOI221_X1 U20593 ( .B1(n21588), .B2(n18463), .C1(n18619), .C2(n18463), .A(
        n18449), .ZN(n18450) );
  XNOR2_X1 U20594 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18450), .ZN(
        n21722) );
  OAI22_X1 U20595 ( .A1(n18451), .A2(n21588), .B1(n18634), .B2(n21722), .ZN(
        n18452) );
  AOI21_X1 U20596 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18481), .A(
        n18452), .ZN(n18455) );
  NAND2_X1 U20597 ( .A1(n21832), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21720) );
  NAND3_X1 U20598 ( .A1(n18453), .A2(n21073), .A3(n18534), .ZN(n18454) );
  NAND4_X1 U20599 ( .A1(n18456), .A2(n18455), .A3(n21720), .A4(n18454), .ZN(
        P3_U2807) );
  OAI21_X1 U20600 ( .B1(n18458), .B2(n18744), .A(n18457), .ZN(n18477) );
  AOI22_X1 U20601 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18477), .B1(
        n18570), .B2(n21095), .ZN(n18472) );
  INV_X1 U20602 ( .A(n18459), .ZN(n18464) );
  INV_X1 U20603 ( .A(n18460), .ZN(n18461) );
  NAND2_X1 U20604 ( .A1(n18462), .A2(n18461), .ZN(n18524) );
  OAI22_X1 U20605 ( .A1(n18464), .A2(n18524), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18463), .ZN(n18465) );
  NOR2_X2 U20606 ( .A1(n18474), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18473) );
  INV_X1 U20607 ( .A(n18501), .ZN(n18496) );
  NOR2_X1 U20608 ( .A1(n18511), .A2(n18473), .ZN(n18498) );
  AOI21_X1 U20609 ( .B1(n18511), .B2(n18496), .A(n18498), .ZN(n18468) );
  XOR2_X1 U20610 ( .A(n18468), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21606) );
  NAND2_X1 U20611 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21716), .ZN(
        n18493) );
  XOR2_X1 U20612 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18493), .Z(
        n21602) );
  INV_X1 U20613 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21611) );
  INV_X1 U20614 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18525) );
  XOR2_X1 U20615 ( .A(n21611), .B(n18494), .Z(n21596) );
  OAI22_X1 U20616 ( .A1(n18612), .A2(n21602), .B1(n18734), .B2(n21596), .ZN(
        n18469) );
  AOI21_X1 U20617 ( .B1(n18661), .B2(n21606), .A(n18469), .ZN(n18471) );
  NAND2_X1 U20618 ( .A1(n21832), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21607) );
  NOR2_X1 U20619 ( .A1(n18486), .A2(n18484), .ZN(n18478) );
  OAI211_X1 U20620 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18478), .B(n18485), .ZN(n18470) );
  NAND4_X1 U20621 ( .A1(n18472), .A2(n18471), .A3(n21607), .A4(n18470), .ZN(
        P3_U2805) );
  AOI21_X1 U20622 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18474), .A(
        n18473), .ZN(n21730) );
  OAI22_X1 U20623 ( .A1(n21808), .A2(n18838), .B1(n18580), .B2(n18475), .ZN(
        n18476) );
  AOI221_X1 U20624 ( .B1(n18478), .B2(n21091), .C1(n18477), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18476), .ZN(n18483) );
  NOR3_X1 U20625 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18479), .A3(
        n21589), .ZN(n21723) );
  AOI22_X1 U20626 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18481), .B1(
        n21723), .B2(n18480), .ZN(n18482) );
  OAI211_X1 U20627 ( .C1(n21730), .C2(n18634), .A(n18483), .B(n18482), .ZN(
        P3_U2806) );
  NOR2_X1 U20628 ( .A1(n18485), .A2(n18484), .ZN(n18517) );
  NAND2_X1 U20629 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18517), .ZN(
        n18488) );
  NOR3_X1 U20630 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18486), .A3(
        n18488), .ZN(n18508) );
  OAI21_X1 U20631 ( .B1(n14158), .B2(n18744), .A(n18745), .ZN(n18487) );
  AOI21_X1 U20632 ( .B1(n18653), .B2(n18488), .A(n18487), .ZN(n18519) );
  OAI21_X1 U20633 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18579), .A(
        n18519), .ZN(n18512) );
  NAND2_X1 U20634 ( .A1(n21832), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21709) );
  NOR2_X1 U20635 ( .A1(n21125), .A2(n18488), .ZN(n18533) );
  NAND3_X1 U20636 ( .A1(n18533), .A2(n18489), .A3(n18534), .ZN(n18490) );
  OAI211_X1 U20637 ( .C1(n18580), .C2(n18491), .A(n21709), .B(n18490), .ZN(
        n18492) );
  AOI221_X1 U20638 ( .B1(n18508), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n18512), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18492), .ZN(
        n18507) );
  INV_X1 U20639 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18529) );
  NOR2_X1 U20640 ( .A1(n18529), .A2(n21611), .ZN(n21627) );
  INV_X1 U20641 ( .A(n21627), .ZN(n18495) );
  NOR2_X2 U20642 ( .A1(n18493), .A2(n18495), .ZN(n21629) );
  AOI22_X1 U20643 ( .A1(n18660), .A2(n21641), .B1(n18700), .B2(n21612), .ZN(
        n18530) );
  NAND2_X1 U20644 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18530), .ZN(
        n18513) );
  OAI211_X1 U20645 ( .C1(n18660), .C2(n18700), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18513), .ZN(n18506) );
  NOR4_X2 U20646 ( .A1(n18525), .A2(n18524), .A3(n18495), .A4(n18523), .ZN(
        n18557) );
  INV_X1 U20647 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21645) );
  NAND3_X1 U20648 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18557), .A3(
        n21645), .ZN(n18505) );
  NOR2_X1 U20649 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18511), .ZN(
        n18542) );
  AOI21_X1 U20650 ( .B1(n18511), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18542), .ZN(n21707) );
  NAND2_X1 U20651 ( .A1(n18496), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18500) );
  AND2_X1 U20652 ( .A1(n18511), .A2(n21611), .ZN(n18497) );
  INV_X1 U20653 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21631) );
  NAND2_X1 U20654 ( .A1(n18502), .A2(n21631), .ZN(n21708) );
  INV_X1 U20655 ( .A(n21708), .ZN(n18543) );
  NAND2_X1 U20656 ( .A1(n18503), .A2(n21707), .ZN(n21687) );
  OAI211_X1 U20657 ( .C1(n21707), .C2(n18503), .A(n18661), .B(n21687), .ZN(
        n18504) );
  NAND4_X1 U20658 ( .A1(n18507), .A2(n18506), .A3(n18505), .A4(n18504), .ZN(
        P3_U2802) );
  AOI21_X1 U20659 ( .B1(n18570), .B2(n21122), .A(n18508), .ZN(n18516) );
  OAI21_X1 U20660 ( .B1(n18511), .B2(n18510), .A(n18509), .ZN(n21625) );
  AOI22_X1 U20661 ( .A1(n18661), .A2(n21625), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18512), .ZN(n18515) );
  OAI21_X1 U20662 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18557), .A(
        n18513), .ZN(n18514) );
  NAND2_X1 U20663 ( .A1(n21832), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21637) );
  NAND4_X1 U20664 ( .A1(n18516), .A2(n18515), .A3(n18514), .A4(n21637), .ZN(
        P3_U2803) );
  AOI21_X1 U20665 ( .B1(n18517), .B2(n19606), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18518) );
  INV_X1 U20666 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21624) );
  OAI22_X1 U20667 ( .A1(n18519), .A2(n18518), .B1(n21808), .B2(n21624), .ZN(
        n18520) );
  AOI221_X1 U20668 ( .B1(n18570), .B2(n21113), .C1(n18429), .C2(n21113), .A(
        n18520), .ZN(n18528) );
  OAI21_X1 U20669 ( .B1(n18522), .B2(n18529), .A(n18521), .ZN(n21616) );
  NOR3_X1 U20670 ( .A1(n18525), .A2(n18524), .A3(n18523), .ZN(n18526) );
  NOR2_X1 U20671 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21611), .ZN(
        n21621) );
  AOI22_X1 U20672 ( .A1(n18661), .A2(n21616), .B1(n18526), .B2(n21621), .ZN(
        n18527) );
  OAI211_X1 U20673 ( .C1(n18530), .C2(n18529), .A(n18528), .B(n18527), .ZN(
        P3_U2804) );
  INV_X1 U20674 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21665) );
  INV_X1 U20675 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21664) );
  NOR2_X1 U20676 ( .A1(n21665), .A2(n21664), .ZN(n21675) );
  NAND2_X1 U20677 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21650) );
  AND2_X1 U20678 ( .A1(n21675), .A2(n21649), .ZN(n18531) );
  INV_X1 U20679 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21674) );
  XOR2_X1 U20680 ( .A(n18531), .B(n21674), .Z(n21678) );
  NAND2_X1 U20681 ( .A1(n21832), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n21683) );
  INV_X1 U20682 ( .A(n21683), .ZN(n18541) );
  NAND2_X1 U20683 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18533), .ZN(
        n18560) );
  NOR2_X1 U20684 ( .A1(n21150), .A2(n18560), .ZN(n18535) );
  NAND2_X1 U20685 ( .A1(n18535), .A2(n18534), .ZN(n18554) );
  XNOR2_X1 U20686 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18539) );
  NOR2_X1 U20687 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18579), .ZN(
        n18569) );
  INV_X1 U20688 ( .A(n18535), .ZN(n18537) );
  AOI22_X1 U20689 ( .A1(n19606), .A2(n18537), .B1(n18536), .B2(n18568), .ZN(
        n18538) );
  NAND2_X1 U20690 ( .A1(n18538), .A2(n18745), .ZN(n18562) );
  NOR2_X1 U20691 ( .A1(n18569), .A2(n18562), .ZN(n18553) );
  OAI22_X1 U20692 ( .A1(n18554), .A2(n18539), .B1(n18553), .B2(n21171), .ZN(
        n18540) );
  AOI211_X1 U20693 ( .C1(n21018), .C2(n18570), .A(n18541), .B(n18540), .ZN(
        n18549) );
  NAND2_X1 U20694 ( .A1(n18543), .A2(n18542), .ZN(n18563) );
  NOR2_X1 U20695 ( .A1(n21645), .A2(n18619), .ZN(n18544) );
  NAND2_X1 U20696 ( .A1(n18545), .A2(n18544), .ZN(n21689) );
  OAI33_X1 U20697 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18563), .B1(n21664), .B2(
        n21689), .B3(n21665), .ZN(n18546) );
  XNOR2_X1 U20698 ( .A(n18546), .B(n21674), .ZN(n21682) );
  NOR2_X1 U20699 ( .A1(n21650), .A2(n21612), .ZN(n21696) );
  NAND2_X1 U20700 ( .A1(n21675), .A2(n21696), .ZN(n18547) );
  XOR2_X1 U20701 ( .A(n18547), .B(n21674), .Z(n21681) );
  AOI22_X1 U20702 ( .A1(n18661), .A2(n21682), .B1(n18700), .B2(n21681), .ZN(
        n18548) );
  OAI211_X1 U20703 ( .C1(n21678), .C2(n18612), .A(n18549), .B(n18548), .ZN(
        P3_U2799) );
  OAI22_X1 U20704 ( .A1(n21665), .A2(n21689), .B1(n18563), .B2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18550) );
  XOR2_X1 U20705 ( .A(n18550), .B(n21664), .Z(n21672) );
  NOR2_X1 U20706 ( .A1(n21650), .A2(n21665), .ZN(n21663) );
  INV_X1 U20707 ( .A(n21663), .ZN(n21640) );
  NOR2_X1 U20708 ( .A1(n21612), .A2(n21640), .ZN(n21642) );
  AOI21_X1 U20709 ( .B1(n21629), .B2(n21663), .A(n18612), .ZN(n18565) );
  INV_X1 U20710 ( .A(n18565), .ZN(n18551) );
  OAI21_X1 U20711 ( .B1(n21642), .B2(n18734), .A(n18551), .ZN(n18566) );
  INV_X1 U20712 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21155) );
  OAI21_X1 U20713 ( .B1(n18567), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n18552), .ZN(n21165) );
  OAI22_X1 U20714 ( .A1(n18553), .A2(n21155), .B1(n18580), .B2(n21165), .ZN(
        n18556) );
  INV_X1 U20715 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21167) );
  OAI22_X1 U20716 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18554), .B1(
        n21808), .B2(n21167), .ZN(n18555) );
  AOI211_X1 U20717 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18566), .A(
        n18556), .B(n18555), .ZN(n18559) );
  NAND3_X1 U20718 ( .A1(n21663), .A2(n18557), .A3(n21664), .ZN(n18558) );
  OAI211_X1 U20719 ( .C1(n21672), .C2(n18634), .A(n18559), .B(n18558), .ZN(
        P3_U2800) );
  OAI21_X1 U20720 ( .B1(n18560), .B2(n19516), .A(n21150), .ZN(n18561) );
  AOI22_X1 U20721 ( .A1(n21801), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18562), 
        .B2(n18561), .ZN(n18574) );
  NAND2_X1 U20722 ( .A1(n18563), .A2(n21689), .ZN(n18564) );
  XOR2_X1 U20723 ( .A(n18564), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21656) );
  AOI22_X1 U20724 ( .A1(n21649), .A2(n18565), .B1(n18661), .B2(n21656), .ZN(
        n18573) );
  OAI221_X1 U20725 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21696), 
        .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n18700), .A(n18566), .ZN(
        n18572) );
  AOI21_X1 U20726 ( .B1(n18568), .B2(n21150), .A(n18567), .ZN(n21145) );
  OAI21_X1 U20727 ( .B1(n18570), .B2(n18569), .A(n21145), .ZN(n18571) );
  NAND4_X1 U20728 ( .A1(n18574), .A2(n18573), .A3(n18572), .A4(n18571), .ZN(
        P3_U2801) );
  OAI21_X1 U20729 ( .B1(n18575), .B2(n19516), .A(n18577), .ZN(n18581) );
  AOI21_X1 U20730 ( .B1(n18578), .B2(n18577), .A(n18576), .ZN(n21003) );
  NAND2_X1 U20731 ( .A1(n18580), .A2(n18579), .ZN(n18736) );
  AOI22_X1 U20732 ( .A1(n18582), .A2(n18581), .B1(n21003), .B2(n18736), .ZN(
        n18589) );
  OAI21_X1 U20733 ( .B1(n18584), .B2(n21770), .A(n18583), .ZN(n21776) );
  AOI22_X1 U20734 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18585), .B1(
        n18661), .B2(n21776), .ZN(n18588) );
  NAND3_X1 U20735 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18586), .A3(
        n21770), .ZN(n18587) );
  NAND2_X1 U20736 ( .A1(n21832), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21777) );
  NAND4_X1 U20737 ( .A1(n18589), .A2(n18588), .A3(n18587), .A4(n21777), .ZN(
        P3_U2813) );
  NOR2_X1 U20738 ( .A1(n18591), .A2(n18590), .ZN(n18593) );
  OAI21_X1 U20739 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18593), .A(
        n18592), .ZN(n20959) );
  NAND2_X1 U20740 ( .A1(n18594), .A2(n19606), .ZN(n18611) );
  INV_X1 U20741 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18595) );
  OAI21_X1 U20742 ( .B1(n18596), .B2(n18611), .A(n18595), .ZN(n18597) );
  AOI22_X1 U20743 ( .A1(n21832), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18598), 
        .B2(n18597), .ZN(n18607) );
  AOI21_X1 U20744 ( .B1(n18602), .B2(n18599), .A(n21572), .ZN(n21562) );
  NAND2_X1 U20745 ( .A1(n18601), .A2(n18600), .ZN(n18603) );
  XOR2_X1 U20746 ( .A(n18603), .B(n18602), .Z(n21566) );
  OAI21_X1 U20747 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18604), .A(
        n21575), .ZN(n21561) );
  OAI22_X1 U20748 ( .A1(n21566), .A2(n18634), .B1(n18612), .B2(n21561), .ZN(
        n18605) );
  AOI21_X1 U20749 ( .B1(n18700), .B2(n21562), .A(n18605), .ZN(n18606) );
  OAI211_X1 U20750 ( .C1(n18726), .C2(n20959), .A(n18607), .B(n18606), .ZN(
        P3_U2816) );
  INV_X1 U20751 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20929) );
  INV_X1 U20752 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20900) );
  INV_X1 U20753 ( .A(n18608), .ZN(n20855) );
  NAND3_X1 U20754 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20855), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20881) );
  INV_X1 U20755 ( .A(n20881), .ZN(n18652) );
  NAND2_X1 U20756 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18652), .ZN(
        n18651) );
  NOR2_X1 U20757 ( .A1(n20900), .A2(n18651), .ZN(n20891) );
  NAND2_X1 U20758 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20891), .ZN(
        n18625) );
  AOI21_X1 U20759 ( .B1(n20929), .B2(n18625), .A(n18609), .ZN(n20925) );
  NAND2_X1 U20760 ( .A1(n18745), .A2(n18702), .ZN(n18737) );
  INV_X1 U20761 ( .A(n18737), .ZN(n18636) );
  NAND3_X1 U20762 ( .A1(n18649), .A2(n20855), .A3(n19606), .ZN(n18637) );
  NOR2_X1 U20763 ( .A1(n20900), .A2(n18637), .ZN(n18635) );
  NAND2_X1 U20764 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18635), .ZN(
        n18626) );
  OAI21_X1 U20765 ( .B1(n18636), .B2(n20929), .A(n18626), .ZN(n18610) );
  AOI22_X1 U20766 ( .A1(n20925), .A2(n18736), .B1(n18611), .B2(n18610), .ZN(
        n18618) );
  OAI22_X1 U20767 ( .A1(n21521), .A2(n18612), .B1(n18734), .B2(n21520), .ZN(
        n18643) );
  AOI21_X1 U20768 ( .B1(n18620), .B2(n21524), .A(n18613), .ZN(n18614) );
  XOR2_X1 U20769 ( .A(n21791), .B(n18614), .Z(n21533) );
  AOI22_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18643), .B1(
        n18661), .B2(n21533), .ZN(n18617) );
  NAND2_X1 U20771 ( .A1(n21832), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18616) );
  NOR2_X1 U20772 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21525), .ZN(
        n21532) );
  OAI221_X1 U20773 ( .B1(n21532), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), 
        .C1(n21532), .C2(n21525), .A(n18630), .ZN(n18615) );
  NAND4_X1 U20774 ( .A1(n18618), .A2(n18617), .A3(n18616), .A4(n18615), .ZN(
        P3_U2819) );
  OAI221_X1 U20775 ( .B1(n18620), .B2(n18619), .C1(n18620), .C2(n21825), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18624) );
  OAI221_X1 U20776 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18641), .C1(
        n21825), .C2(n18640), .A(n18621), .ZN(n18622) );
  OAI221_X1 U20777 ( .B1(n18624), .B2(n18623), .C1(n18624), .C2(n21825), .A(
        n18622), .ZN(n21814) );
  OAI21_X1 U20778 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20891), .A(
        n18625), .ZN(n20912) );
  OAI211_X1 U20779 ( .C1(n18635), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18737), .B(n18626), .ZN(n18628) );
  NAND2_X1 U20780 ( .A1(n21832), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18627) );
  OAI211_X1 U20781 ( .C1(n18726), .C2(n20912), .A(n18628), .B(n18627), .ZN(
        n18629) );
  AOI21_X1 U20782 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18643), .A(
        n18629), .ZN(n18633) );
  NAND3_X1 U20783 ( .A1(n18631), .A2(n21525), .A3(n18630), .ZN(n18632) );
  OAI211_X1 U20784 ( .C1(n21814), .C2(n18634), .A(n18633), .B(n18632), .ZN(
        P3_U2820) );
  AOI21_X1 U20785 ( .B1(n20900), .B2(n18651), .A(n20891), .ZN(n20899) );
  AOI211_X1 U20786 ( .C1(n18637), .C2(n20900), .A(n18636), .B(n18635), .ZN(
        n18639) );
  NOR2_X1 U20787 ( .A1(n21808), .A2(n21830), .ZN(n18638) );
  AOI211_X1 U20788 ( .C1(n20899), .C2(n18736), .A(n18639), .B(n18638), .ZN(
        n18645) );
  NAND2_X1 U20789 ( .A1(n18641), .A2(n18640), .ZN(n18642) );
  XOR2_X1 U20790 ( .A(n18642), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21827) );
  AOI22_X1 U20791 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18643), .B1(
        n18661), .B2(n21827), .ZN(n18644) );
  OAI211_X1 U20792 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18646), .A(
        n18645), .B(n18644), .ZN(P3_U2821) );
  OAI21_X1 U20793 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18648), .A(
        n18647), .ZN(n21518) );
  NAND2_X1 U20794 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20855), .ZN(
        n18650) );
  AOI211_X1 U20795 ( .C1(n18654), .C2(n18650), .A(n18649), .B(n19516), .ZN(
        n18656) );
  OAI21_X1 U20796 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18652), .A(
        n18651), .ZN(n20883) );
  AOI21_X1 U20797 ( .B1(n18653), .B2(n18608), .A(n18728), .ZN(n18669) );
  OAI22_X1 U20798 ( .A1(n18726), .A2(n20883), .B1(n18654), .B2(n18669), .ZN(
        n18655) );
  AOI211_X1 U20799 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n21832), .A(n18656), .B(
        n18655), .ZN(n18663) );
  XNOR2_X1 U20800 ( .A(n18658), .B(n18657), .ZN(n18659) );
  INV_X1 U20801 ( .A(n18659), .ZN(n21514) );
  AOI22_X1 U20802 ( .A1(n21514), .A2(n18661), .B1(n18660), .B2(n18659), .ZN(
        n18662) );
  OAI211_X1 U20803 ( .C1(n18734), .C2(n21518), .A(n18663), .B(n18662), .ZN(
        P3_U2822) );
  NOR2_X1 U20804 ( .A1(n18665), .A2(n18664), .ZN(n18666) );
  XOR2_X1 U20805 ( .A(n18666), .B(n21431), .Z(n21507) );
  NOR2_X1 U20806 ( .A1(n18608), .A2(n19516), .ZN(n18672) );
  NOR2_X1 U20807 ( .A1(n18608), .A2(n20782), .ZN(n18676) );
  OAI21_X1 U20808 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18676), .A(
        n20881), .ZN(n20864) );
  OAI22_X1 U20809 ( .A1(n18726), .A2(n20864), .B1(n21808), .B2(n20877), .ZN(
        n18671) );
  OAI21_X1 U20810 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18668), .A(
        n18667), .ZN(n21506) );
  OAI22_X1 U20811 ( .A1(n18739), .A2(n21506), .B1(n20871), .B2(n18669), .ZN(
        n18670) );
  AOI211_X1 U20812 ( .C1(n18672), .C2(n20871), .A(n18671), .B(n18670), .ZN(
        n18673) );
  OAI21_X1 U20813 ( .B1(n18734), .B2(n21507), .A(n18673), .ZN(P3_U2823) );
  OAI21_X1 U20814 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18675), .A(
        n18674), .ZN(n21501) );
  INV_X1 U20815 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20853) );
  NAND2_X1 U20816 ( .A1(n18677), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18685) );
  AOI21_X1 U20817 ( .B1(n20853), .B2(n18685), .A(n18676), .ZN(n20854) );
  NAND2_X1 U20818 ( .A1(n18677), .A2(n19606), .ZN(n18681) );
  NAND2_X1 U20819 ( .A1(n21832), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21499) );
  OAI21_X1 U20820 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18681), .A(
        n21499), .ZN(n18683) );
  OAI21_X1 U20821 ( .B1(n18680), .B2(n18679), .A(n18678), .ZN(n21494) );
  NAND2_X1 U20822 ( .A1(n18737), .A2(n18681), .ZN(n18689) );
  OAI22_X1 U20823 ( .A1(n18739), .A2(n21494), .B1(n20853), .B2(n18689), .ZN(
        n18682) );
  AOI211_X1 U20824 ( .C1(n20854), .C2(n18736), .A(n18683), .B(n18682), .ZN(
        n18684) );
  OAI21_X1 U20825 ( .B1(n18734), .B2(n21501), .A(n18684), .ZN(P3_U2824) );
  NOR2_X1 U20826 ( .A1(n18690), .A2(n20782), .ZN(n18696) );
  OAI21_X1 U20827 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18696), .A(
        n18685), .ZN(n20839) );
  XOR2_X1 U20828 ( .A(n21426), .B(n18686), .Z(n18688) );
  XNOR2_X1 U20829 ( .A(n18688), .B(n18687), .ZN(n21488) );
  AOI221_X1 U20830 ( .B1(n18728), .B2(n20843), .C1(n18690), .C2(n20843), .A(
        n18689), .ZN(n18694) );
  OAI21_X1 U20831 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18692), .A(
        n18691), .ZN(n21479) );
  OAI22_X1 U20832 ( .A1(n21808), .A2(n20834), .B1(n18739), .B2(n21479), .ZN(
        n18693) );
  AOI211_X1 U20833 ( .C1(n18700), .C2(n21488), .A(n18694), .B(n18693), .ZN(
        n18695) );
  OAI21_X1 U20834 ( .B1(n18726), .B2(n20839), .A(n18695), .ZN(P3_U2825) );
  NAND2_X1 U20835 ( .A1(n18703), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18711) );
  INV_X1 U20836 ( .A(n18711), .ZN(n20828) );
  INV_X1 U20837 ( .A(n18696), .ZN(n20836) );
  OAI21_X1 U20838 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20828), .A(
        n20836), .ZN(n20829) );
  NOR3_X1 U20839 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18697), .A3(
        n19516), .ZN(n18698) );
  AOI211_X1 U20840 ( .C1(n18701), .C2(n18700), .A(n18699), .B(n18698), .ZN(
        n18707) );
  OAI21_X1 U20841 ( .B1(n18703), .B2(n18702), .A(n18745), .ZN(n18718) );
  AOI22_X1 U20842 ( .A1(n18705), .A2(n18704), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18718), .ZN(n18706) );
  OAI211_X1 U20843 ( .C1(n18726), .C2(n20829), .A(n18707), .B(n18706), .ZN(
        P3_U2826) );
  OAI21_X1 U20844 ( .B1(n18710), .B2(n18709), .A(n18708), .ZN(n21478) );
  INV_X1 U20845 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20804) );
  NOR2_X1 U20846 ( .A1(n18728), .A2(n20804), .ZN(n18717) );
  NOR2_X1 U20847 ( .A1(n20804), .A2(n20782), .ZN(n18712) );
  OAI21_X1 U20848 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18712), .A(
        n18711), .ZN(n20807) );
  OAI21_X1 U20849 ( .B1(n18715), .B2(n18714), .A(n18713), .ZN(n21472) );
  OAI22_X1 U20850 ( .A1(n18726), .A2(n20807), .B1(n18739), .B2(n21472), .ZN(
        n18716) );
  AOI221_X1 U20851 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18718), .C1(
        n18717), .C2(n18718), .A(n18716), .ZN(n18719) );
  NAND2_X1 U20852 ( .A1(n21832), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21476) );
  OAI211_X1 U20853 ( .C1(n18734), .C2(n21478), .A(n18719), .B(n21476), .ZN(
        P3_U2827) );
  OAI21_X1 U20854 ( .B1(n18722), .B2(n18721), .A(n18720), .ZN(n21461) );
  AOI22_X1 U20855 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20782), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20804), .ZN(n20800) );
  OAI21_X1 U20856 ( .B1(n18725), .B2(n18724), .A(n18723), .ZN(n21465) );
  OAI22_X1 U20857 ( .A1(n18726), .A2(n20800), .B1(n18734), .B2(n21465), .ZN(
        n18727) );
  AOI221_X1 U20858 ( .B1(n18728), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19606), .C2(n20804), .A(n18727), .ZN(n18729) );
  NAND2_X1 U20859 ( .A1(n21832), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21470) );
  OAI211_X1 U20860 ( .C1(n18739), .C2(n21461), .A(n18729), .B(n21470), .ZN(
        P3_U2828) );
  OAI21_X1 U20861 ( .B1(n18733), .B2(n18740), .A(n18730), .ZN(n21453) );
  AOI21_X1 U20862 ( .B1(n18733), .B2(n18732), .A(n18731), .ZN(n21454) );
  OAI22_X1 U20863 ( .A1(n21454), .A2(n18734), .B1(n21808), .B2(n20787), .ZN(
        n18735) );
  AOI221_X1 U20864 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18737), .C1(
        n20782), .C2(n18736), .A(n18735), .ZN(n18738) );
  OAI21_X1 U20865 ( .B1(n18739), .B2(n21453), .A(n18738), .ZN(P3_U2829) );
  NOR2_X1 U20866 ( .A1(n18741), .A2(n18740), .ZN(n18743) );
  INV_X1 U20867 ( .A(n18743), .ZN(n18742) );
  AOI22_X1 U20868 ( .A1(n18743), .A2(n21483), .B1(n21834), .B2(n18742), .ZN(
        n21447) );
  NAND3_X1 U20869 ( .A1(n18746), .A2(n18745), .A3(n18744), .ZN(n18747) );
  AOI22_X1 U20870 ( .A1(n21832), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18747), .ZN(n18748) );
  OAI21_X1 U20871 ( .B1(n21447), .B2(n21900), .A(n18748), .ZN(P3_U2830) );
  INV_X1 U20872 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21864) );
  NOR2_X1 U20873 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19277), .ZN(
        n19311) );
  NAND2_X1 U20874 ( .A1(n21861), .A2(n21864), .ZN(n19340) );
  INV_X1 U20875 ( .A(n19340), .ZN(n19342) );
  NOR2_X1 U20876 ( .A1(n21861), .A2(n21864), .ZN(n19288) );
  NOR2_X1 U20877 ( .A1(n19342), .A2(n19288), .ZN(n18749) );
  AOI22_X1 U20878 ( .A1(n18751), .A2(n19311), .B1(n18750), .B2(n18749), .ZN(
        n18752) );
  OAI21_X1 U20879 ( .B1(n18753), .B2(n21864), .A(n18752), .ZN(P3_U2866) );
  OAI21_X1 U20880 ( .B1(n18755), .B2(n18754), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18756) );
  OAI21_X1 U20881 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18757), .A(
        n18756), .ZN(P3_U2864) );
  NOR4_X1 U20882 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18761) );
  NOR4_X1 U20883 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18760) );
  NOR4_X1 U20884 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18759) );
  NOR4_X1 U20885 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18758) );
  NAND4_X1 U20886 ( .A1(n18761), .A2(n18760), .A3(n18759), .A4(n18758), .ZN(
        n18767) );
  NOR4_X1 U20887 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18765) );
  AOI211_X1 U20888 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18764) );
  NOR4_X1 U20889 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18763) );
  NOR4_X1 U20890 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18762) );
  NAND4_X1 U20891 ( .A1(n18765), .A2(n18764), .A3(n18763), .A4(n18762), .ZN(
        n18766) );
  NOR2_X1 U20892 ( .A1(n18767), .A2(n18766), .ZN(n18780) );
  INV_X1 U20893 ( .A(n18780), .ZN(n18777) );
  NOR2_X1 U20894 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18769) );
  NAND2_X1 U20895 ( .A1(n18777), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18768) );
  OAI21_X1 U20896 ( .B1(n18777), .B2(n18769), .A(n18768), .ZN(P3_U3293) );
  AOI211_X1 U20897 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18770) );
  AOI21_X1 U20898 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18770), .ZN(n18772) );
  INV_X1 U20899 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U20900 ( .A1(n18780), .A2(n18772), .B1(n18771), .B2(n18777), .ZN(
        P3_U3292) );
  INV_X1 U20901 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18774) );
  NOR3_X1 U20902 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18776) );
  NOR2_X1 U20903 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18776), .ZN(n18773) );
  MUX2_X1 U20904 ( .A(n18774), .B(n18773), .S(n18780), .Z(n18775) );
  INV_X1 U20905 ( .A(n18775), .ZN(P3_U2638) );
  INV_X1 U20906 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22235) );
  AOI21_X1 U20907 ( .B1(n20787), .B2(n22235), .A(n18776), .ZN(n18779) );
  INV_X1 U20908 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18778) );
  AOI22_X1 U20909 ( .A1(n18780), .A2(n18779), .B1(n18778), .B2(n18777), .ZN(
        P3_U2639) );
  INV_X1 U20910 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18845) );
  AOI22_X1 U20911 ( .A1(n22240), .A2(n18781), .B1(n18845), .B2(n18842), .ZN(
        P3_U3297) );
  OAI22_X1 U20912 ( .A1(n18842), .A2(n18782), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n22240), .ZN(n18783) );
  INV_X1 U20913 ( .A(n18783), .ZN(P3_U3294) );
  AOI21_X1 U20914 ( .B1(n22285), .B2(n22287), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18784) );
  AOI22_X1 U20915 ( .A1(n22240), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18784), 
        .B2(n18842), .ZN(P3_U2635) );
  INV_X1 U20916 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21376) );
  AOI22_X1 U20917 ( .A1(n21886), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18785) );
  OAI21_X1 U20918 ( .B1(n21376), .B2(n18801), .A(n18785), .ZN(P3_U2767) );
  INV_X1 U20919 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21369) );
  AOI22_X1 U20920 ( .A1(n21886), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18786) );
  OAI21_X1 U20921 ( .B1(n21369), .B2(n18801), .A(n18786), .ZN(P3_U2766) );
  INV_X1 U20922 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21219) );
  AOI22_X1 U20923 ( .A1(n21886), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18787) );
  OAI21_X1 U20924 ( .B1(n21219), .B2(n18801), .A(n18787), .ZN(P3_U2765) );
  INV_X1 U20925 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20756) );
  AOI22_X1 U20926 ( .A1(n21886), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18788) );
  OAI21_X1 U20927 ( .B1(n20756), .B2(n18801), .A(n18788), .ZN(P3_U2764) );
  INV_X1 U20928 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21220) );
  AOI22_X1 U20929 ( .A1(n21886), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18789) );
  OAI21_X1 U20930 ( .B1(n21220), .B2(n18801), .A(n18789), .ZN(P3_U2763) );
  INV_X1 U20931 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U20932 ( .A1(n21886), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18790) );
  OAI21_X1 U20933 ( .B1(n20759), .B2(n18801), .A(n18790), .ZN(P3_U2762) );
  INV_X1 U20934 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21221) );
  AOI22_X1 U20935 ( .A1(n21886), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18791) );
  OAI21_X1 U20936 ( .B1(n21221), .B2(n18801), .A(n18791), .ZN(P3_U2761) );
  INV_X1 U20937 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U20938 ( .A1(n21886), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18792) );
  OAI21_X1 U20939 ( .B1(n20762), .B2(n18801), .A(n18792), .ZN(P3_U2760) );
  INV_X1 U20940 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21360) );
  AOI22_X1 U20941 ( .A1(n20719), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18793) );
  OAI21_X1 U20942 ( .B1(n21360), .B2(n18801), .A(n18793), .ZN(P3_U2759) );
  INV_X1 U20943 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21248) );
  AOI22_X1 U20944 ( .A1(n20719), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18794) );
  OAI21_X1 U20945 ( .B1(n21248), .B2(n18801), .A(n18794), .ZN(P3_U2758) );
  INV_X1 U20946 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20767) );
  AOI22_X1 U20947 ( .A1(n20719), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18795) );
  OAI21_X1 U20948 ( .B1(n20767), .B2(n18801), .A(n18795), .ZN(P3_U2757) );
  INV_X1 U20949 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21203) );
  AOI22_X1 U20950 ( .A1(n20719), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18796) );
  OAI21_X1 U20951 ( .B1(n21203), .B2(n18801), .A(n18796), .ZN(P3_U2756) );
  INV_X1 U20952 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U20953 ( .A1(n20719), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18797) );
  OAI21_X1 U20954 ( .B1(n20770), .B2(n18801), .A(n18797), .ZN(P3_U2755) );
  INV_X1 U20955 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U20956 ( .A1(n20719), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18798) );
  OAI21_X1 U20957 ( .B1(n20772), .B2(n18801), .A(n18798), .ZN(P3_U2754) );
  INV_X1 U20958 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21348) );
  AOI22_X1 U20959 ( .A1(n20719), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18799) );
  OAI21_X1 U20960 ( .B1(n21348), .B2(n18801), .A(n18799), .ZN(P3_U2753) );
  INV_X1 U20961 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21351) );
  AOI22_X1 U20962 ( .A1(n20719), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18800) );
  OAI21_X1 U20963 ( .B1(n21351), .B2(n18801), .A(n18800), .ZN(P3_U2752) );
  INV_X1 U20964 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20729) );
  NAND2_X1 U20965 ( .A1(n18803), .A2(n18802), .ZN(n18821) );
  AOI22_X1 U20966 ( .A1(n20719), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18804) );
  OAI21_X1 U20967 ( .B1(n20729), .B2(n18821), .A(n18804), .ZN(P3_U2751) );
  INV_X1 U20968 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21251) );
  AOI22_X1 U20969 ( .A1(n20719), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18805) );
  OAI21_X1 U20970 ( .B1(n21251), .B2(n18821), .A(n18805), .ZN(P3_U2750) );
  INV_X1 U20971 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20732) );
  AOI22_X1 U20972 ( .A1(n20719), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18806) );
  OAI21_X1 U20973 ( .B1(n20732), .B2(n18821), .A(n18806), .ZN(P3_U2749) );
  INV_X1 U20974 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21273) );
  AOI22_X1 U20975 ( .A1(n20719), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18807) );
  OAI21_X1 U20976 ( .B1(n21273), .B2(n18821), .A(n18807), .ZN(P3_U2748) );
  INV_X1 U20977 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21263) );
  AOI22_X1 U20978 ( .A1(n20719), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18808) );
  OAI21_X1 U20979 ( .B1(n21263), .B2(n18821), .A(n18808), .ZN(P3_U2747) );
  INV_X1 U20980 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21258) );
  AOI22_X1 U20981 ( .A1(n20719), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18809) );
  OAI21_X1 U20982 ( .B1(n21258), .B2(n18821), .A(n18809), .ZN(P3_U2746) );
  INV_X1 U20983 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U20984 ( .A1(n20719), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18810) );
  OAI21_X1 U20985 ( .B1(n20737), .B2(n18821), .A(n18810), .ZN(P3_U2745) );
  INV_X1 U20986 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U20987 ( .A1(n20719), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18811) );
  OAI21_X1 U20988 ( .B1(n20739), .B2(n18821), .A(n18811), .ZN(P3_U2744) );
  INV_X1 U20989 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U20990 ( .A1(n20719), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18812), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18813) );
  OAI21_X1 U20991 ( .B1(n20741), .B2(n18821), .A(n18813), .ZN(P3_U2743) );
  INV_X1 U20992 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20743) );
  AOI22_X1 U20993 ( .A1(n20719), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18814) );
  OAI21_X1 U20994 ( .B1(n20743), .B2(n18821), .A(n18814), .ZN(P3_U2742) );
  INV_X1 U20995 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21297) );
  AOI22_X1 U20996 ( .A1(n20719), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18815) );
  OAI21_X1 U20997 ( .B1(n21297), .B2(n18821), .A(n18815), .ZN(P3_U2741) );
  INV_X1 U20998 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20746) );
  AOI22_X1 U20999 ( .A1(n20719), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18816) );
  OAI21_X1 U21000 ( .B1(n20746), .B2(n18821), .A(n18816), .ZN(P3_U2740) );
  INV_X1 U21001 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20748) );
  AOI22_X1 U21002 ( .A1(n20719), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18817) );
  OAI21_X1 U21003 ( .B1(n20748), .B2(n18821), .A(n18817), .ZN(P3_U2739) );
  INV_X1 U21004 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n21309) );
  AOI22_X1 U21005 ( .A1(n20719), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18818) );
  OAI21_X1 U21006 ( .B1(n21309), .B2(n18821), .A(n18818), .ZN(P3_U2738) );
  INV_X1 U21007 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U21008 ( .A1(n20719), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18819), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18820) );
  OAI21_X1 U21009 ( .B1(n20751), .B2(n18821), .A(n18820), .ZN(P3_U2737) );
  AOI21_X1 U21010 ( .B1(n18842), .B2(P3_ADS_N_REG_SCAN_IN), .A(n22236), .ZN(
        n18822) );
  INV_X1 U21011 ( .A(n18822), .ZN(P3_U2633) );
  NOR2_X1 U21012 ( .A1(n18842), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18834) );
  INV_X1 U21013 ( .A(n18839), .ZN(n18836) );
  AOI22_X1 U21014 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18842), .ZN(n18823) );
  OAI21_X1 U21015 ( .B1(n20788), .B2(n18841), .A(n18823), .ZN(P3_U3032) );
  AOI22_X1 U21016 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18842), .ZN(n18824) );
  OAI21_X1 U21017 ( .B1(n20801), .B2(n18841), .A(n18824), .ZN(P3_U3033) );
  AOI22_X1 U21018 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n18842), .ZN(n18825) );
  OAI21_X1 U21019 ( .B1(n20819), .B2(n18841), .A(n18825), .ZN(P3_U3034) );
  AOI22_X1 U21020 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n18842), .ZN(n18826) );
  OAI21_X1 U21021 ( .B1(n20834), .B2(n18841), .A(n18826), .ZN(P3_U3035) );
  INV_X1 U21022 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20849) );
  AOI22_X1 U21023 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n18842), .ZN(n18827) );
  OAI21_X1 U21024 ( .B1(n20849), .B2(n18841), .A(n18827), .ZN(P3_U3036) );
  AOI22_X1 U21025 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n18842), .ZN(n18828) );
  OAI21_X1 U21026 ( .B1(n20877), .B2(n18841), .A(n18828), .ZN(P3_U3037) );
  AOI22_X1 U21027 ( .A1(n18834), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n18842), .ZN(n18829) );
  OAI21_X1 U21028 ( .B1(n18839), .B2(n20877), .A(n18829), .ZN(P3_U3038) );
  AOI22_X1 U21029 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n18842), .ZN(n18830) );
  OAI21_X1 U21030 ( .B1(n21830), .B2(n18841), .A(n18830), .ZN(P3_U3039) );
  AOI22_X1 U21031 ( .A1(n18834), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n18842), .ZN(n18831) );
  OAI21_X1 U21032 ( .B1(n18839), .B2(n21830), .A(n18831), .ZN(P3_U3040) );
  AOI22_X1 U21033 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n18842), .ZN(n18832) );
  OAI21_X1 U21034 ( .B1(n21535), .B2(n18841), .A(n18832), .ZN(P3_U3041) );
  INV_X1 U21035 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20414) );
  OAI222_X1 U21036 ( .A1(n21535), .A2(n18839), .B1(n20414), .B2(n22240), .C1(
        n20953), .C2(n18841), .ZN(P3_U3042) );
  INV_X1 U21037 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20416) );
  OAI222_X1 U21038 ( .A1(n18841), .A2(n20954), .B1(n20416), .B2(n22240), .C1(
        n20953), .C2(n18839), .ZN(P3_U3043) );
  INV_X1 U21039 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20418) );
  OAI222_X1 U21040 ( .A1(n18841), .A2(n20962), .B1(n20418), .B2(n22240), .C1(
        n20954), .C2(n18839), .ZN(P3_U3044) );
  INV_X1 U21041 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20420) );
  OAI222_X1 U21042 ( .A1(n18841), .A2(n20986), .B1(n20420), .B2(n22240), .C1(
        n20962), .C2(n18839), .ZN(P3_U3045) );
  INV_X1 U21043 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20422) );
  OAI222_X1 U21044 ( .A1(n18841), .A2(n20993), .B1(n20422), .B2(n22240), .C1(
        n20986), .C2(n18839), .ZN(P3_U3046) );
  INV_X1 U21045 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20424) );
  OAI222_X1 U21046 ( .A1(n20993), .A2(n18839), .B1(n20424), .B2(n22240), .C1(
        n21010), .C2(n18841), .ZN(P3_U3047) );
  INV_X1 U21047 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20426) );
  INV_X1 U21048 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21025) );
  OAI222_X1 U21049 ( .A1(n21010), .A2(n18839), .B1(n20426), .B2(n22240), .C1(
        n21025), .C2(n18841), .ZN(P3_U3048) );
  INV_X1 U21050 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20428) );
  INV_X1 U21051 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21039) );
  OAI222_X1 U21052 ( .A1(n21025), .A2(n18839), .B1(n20428), .B2(n22240), .C1(
        n21039), .C2(n18841), .ZN(P3_U3049) );
  INV_X1 U21053 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20430) );
  OAI222_X1 U21054 ( .A1(n18841), .A2(n18833), .B1(n20430), .B2(n22240), .C1(
        n21039), .C2(n18839), .ZN(P3_U3050) );
  INV_X1 U21055 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20432) );
  OAI222_X1 U21056 ( .A1(n18841), .A2(n21445), .B1(n20432), .B2(n22240), .C1(
        n18833), .C2(n18839), .ZN(P3_U3051) );
  INV_X1 U21057 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20434) );
  OAI222_X1 U21058 ( .A1(n18841), .A2(n21066), .B1(n20434), .B2(n22240), .C1(
        n21445), .C2(n18839), .ZN(P3_U3052) );
  AOI22_X1 U21059 ( .A1(n18834), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n18842), .ZN(n18835) );
  OAI21_X1 U21060 ( .B1(n18839), .B2(n21066), .A(n18835), .ZN(P3_U3053) );
  AOI22_X1 U21061 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n18836), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n18842), .ZN(n18837) );
  OAI21_X1 U21062 ( .B1(n18838), .B2(n18841), .A(n18837), .ZN(P3_U3054) );
  INV_X1 U21063 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21101) );
  INV_X1 U21064 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20438) );
  OAI222_X1 U21065 ( .A1(n18841), .A2(n21101), .B1(n20438), .B2(n22240), .C1(
        n18838), .C2(n18839), .ZN(P3_U3055) );
  INV_X1 U21066 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20440) );
  OAI222_X1 U21067 ( .A1(n18841), .A2(n21624), .B1(n20440), .B2(n22240), .C1(
        n21101), .C2(n18839), .ZN(P3_U3056) );
  INV_X1 U21068 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20442) );
  OAI222_X1 U21069 ( .A1(n18841), .A2(n21133), .B1(n20442), .B2(n22240), .C1(
        n21624), .C2(n18839), .ZN(P3_U3057) );
  INV_X1 U21070 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20444) );
  OAI222_X1 U21071 ( .A1(n18841), .A2(n21136), .B1(n20444), .B2(n22240), .C1(
        n21133), .C2(n18839), .ZN(P3_U3058) );
  INV_X1 U21072 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20446) );
  INV_X1 U21073 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21661) );
  OAI222_X1 U21074 ( .A1(n21136), .A2(n18839), .B1(n20446), .B2(n22240), .C1(
        n21661), .C2(n18841), .ZN(P3_U3059) );
  INV_X1 U21075 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20448) );
  OAI222_X1 U21076 ( .A1(n18841), .A2(n21167), .B1(n20448), .B2(n22240), .C1(
        n21661), .C2(n18839), .ZN(P3_U3060) );
  INV_X1 U21077 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18840) );
  INV_X1 U21078 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20451) );
  OAI222_X1 U21079 ( .A1(n18841), .A2(n18840), .B1(n20451), .B2(n22240), .C1(
        n21167), .C2(n18839), .ZN(P3_U3061) );
  MUX2_X1 U21080 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .B(P3_BE_N_REG_0__SCAN_IN), .S(n18842), .Z(P3_U3277) );
  MUX2_X1 U21081 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n18842), .Z(P3_U3276) );
  OAI22_X1 U21082 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n22240), .ZN(n18843) );
  INV_X1 U21083 ( .A(n18843), .ZN(P3_U3275) );
  OAI22_X1 U21084 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n22240), .ZN(n18844) );
  INV_X1 U21085 ( .A(n18844), .ZN(P3_U3274) );
  NOR4_X1 U21086 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18847)
         );
  NOR4_X1 U21087 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18845), .ZN(n18846) );
  INV_X2 U21088 ( .A(n19603), .ZN(U215) );
  NAND3_X1 U21089 ( .A1(n18847), .A2(n18846), .A3(U215), .ZN(U213) );
  NAND3_X1 U21090 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18848), .A3(n22264), 
        .ZN(n18849) );
  OAI211_X1 U21091 ( .C1(n18852), .C2(n18851), .A(n18850), .B(n18849), .ZN(
        n18861) );
  INV_X1 U21092 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22271) );
  AOI211_X1 U21093 ( .C1(n22272), .C2(P2_STATEBS16_REG_SCAN_IN), .A(n18853), 
        .B(n19096), .ZN(n18859) );
  NOR2_X1 U21094 ( .A1(n22275), .A2(n19835), .ZN(n18857) );
  INV_X1 U21095 ( .A(n22272), .ZN(n18854) );
  NAND3_X1 U21096 ( .A1(n18855), .A2(n20289), .A3(n18854), .ZN(n18856) );
  OAI21_X1 U21097 ( .B1(n18857), .B2(n19235), .A(n18856), .ZN(n18858) );
  OAI21_X1 U21098 ( .B1(n18859), .B2(n18858), .A(n18861), .ZN(n18860) );
  OAI21_X1 U21099 ( .B1(n18861), .B2(n22271), .A(n18860), .ZN(P2_U3610) );
  OAI22_X1 U21100 ( .A1(n19072), .A2(n20275), .B1(n19059), .B2(n18862), .ZN(
        n18863) );
  INV_X1 U21101 ( .A(n18863), .ZN(n18868) );
  AOI22_X1 U21102 ( .A1(n19068), .A2(n18864), .B1(n11144), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n18867) );
  NAND2_X1 U21103 ( .A1(n18865), .A2(n19067), .ZN(n18866) );
  AND3_X1 U21104 ( .A1(n18868), .A2(n18867), .A3(n18866), .ZN(n18873) );
  AOI22_X1 U21105 ( .A1(n18937), .A2(n18870), .B1(n18869), .B2(n20282), .ZN(
        n18872) );
  OAI21_X1 U21106 ( .B1(n19028), .B2(n18932), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18871) );
  NAND3_X1 U21107 ( .A1(n18873), .A2(n18872), .A3(n18871), .ZN(P2_U2855) );
  INV_X1 U21108 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18874) );
  OAI21_X1 U21109 ( .B1(n18874), .B2(n19007), .A(n18958), .ZN(n18877) );
  OAI22_X1 U21110 ( .A1(n18875), .A2(n18996), .B1(n19059), .B2(n12984), .ZN(
        n18876) );
  AOI211_X1 U21111 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19028), .A(
        n18877), .B(n18876), .ZN(n18885) );
  NAND2_X1 U21112 ( .A1(n11223), .A2(n18878), .ZN(n18879) );
  XNOR2_X1 U21113 ( .A(n18880), .B(n18879), .ZN(n18883) );
  INV_X1 U21114 ( .A(n18881), .ZN(n18882) );
  AOI22_X1 U21115 ( .A1(n18883), .A2(n19055), .B1(n18882), .B2(n19067), .ZN(
        n18884) );
  OAI211_X1 U21116 ( .C1(n19072), .C2(n19969), .A(n18885), .B(n18884), .ZN(
        P2_U2849) );
  NOR2_X1 U21117 ( .A1(n19054), .A2(n18886), .ZN(n18887) );
  XOR2_X1 U21118 ( .A(n18888), .B(n18887), .Z(n18898) );
  INV_X1 U21119 ( .A(n19736), .ZN(n18896) );
  AOI22_X1 U21120 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_7__SCAN_IN), .B2(n19009), .ZN(n18889) );
  NAND2_X1 U21121 ( .A1(n18958), .A2(n18889), .ZN(n18890) );
  AOI21_X1 U21122 ( .B1(n11144), .B2(P2_EBX_REG_7__SCAN_IN), .A(n18890), .ZN(
        n18893) );
  OR2_X1 U21123 ( .A1(n19011), .A2(n18891), .ZN(n18892) );
  OAI211_X1 U21124 ( .C1(n18894), .C2(n18996), .A(n18893), .B(n18892), .ZN(
        n18895) );
  AOI21_X1 U21125 ( .B1(n18896), .B2(n18916), .A(n18895), .ZN(n18897) );
  OAI21_X1 U21126 ( .B1(n19230), .B2(n18898), .A(n18897), .ZN(P2_U2848) );
  NAND2_X1 U21127 ( .A1(n11222), .A2(n18899), .ZN(n18901) );
  XNOR2_X1 U21128 ( .A(n18901), .B(n18900), .ZN(n18910) );
  NAND2_X1 U21129 ( .A1(n18902), .A2(n19067), .ZN(n18906) );
  AOI22_X1 U21130 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19009), .ZN(n18903) );
  NAND2_X1 U21131 ( .A1(n18958), .A2(n18903), .ZN(n18904) );
  AOI21_X1 U21132 ( .B1(n11144), .B2(P2_EBX_REG_10__SCAN_IN), .A(n18904), .ZN(
        n18905) );
  OAI211_X1 U21133 ( .C1(n19072), .C2(n19727), .A(n18906), .B(n18905), .ZN(
        n18907) );
  AOI21_X1 U21134 ( .B1(n19068), .B2(n18908), .A(n18907), .ZN(n18909) );
  OAI21_X1 U21135 ( .B1(n18910), .B2(n19230), .A(n18909), .ZN(P2_U2845) );
  INV_X1 U21136 ( .A(n18911), .ZN(n18920) );
  INV_X1 U21137 ( .A(n19724), .ZN(n18915) );
  AOI22_X1 U21138 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11144), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19009), .ZN(n18912) );
  OAI211_X1 U21139 ( .C1(n19061), .C2(n18913), .A(n17323), .B(n18912), .ZN(
        n18914) );
  AOI21_X1 U21140 ( .B1(n18916), .B2(n18915), .A(n18914), .ZN(n18917) );
  OAI21_X1 U21141 ( .B1(n18918), .B2(n19011), .A(n18917), .ZN(n18919) );
  AOI21_X1 U21142 ( .B1(n18920), .B2(n19068), .A(n18919), .ZN(n18924) );
  OAI211_X1 U21143 ( .C1(n18922), .C2(n18925), .A(n18937), .B(n18921), .ZN(
        n18923) );
  OAI211_X1 U21144 ( .C1(n18926), .C2(n18925), .A(n18924), .B(n18923), .ZN(
        P2_U2844) );
  OAI21_X1 U21145 ( .B1(n18928), .B2(n18927), .A(n17502), .ZN(n19718) );
  AOI22_X1 U21146 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n11144), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19009), .ZN(n18929) );
  OAI211_X1 U21147 ( .C1(n19061), .C2(n18930), .A(n17323), .B(n18929), .ZN(
        n18931) );
  AOI21_X1 U21148 ( .B1(n18933), .B2(n18932), .A(n18931), .ZN(n18934) );
  OAI21_X1 U21149 ( .B1(n19122), .B2(n19011), .A(n18934), .ZN(n18935) );
  AOI21_X1 U21150 ( .B1(n18936), .B2(n19068), .A(n18935), .ZN(n18941) );
  OAI211_X1 U21151 ( .C1(n18939), .C2(n18938), .A(n18937), .B(n18942), .ZN(
        n18940) );
  OAI211_X1 U21152 ( .C1(n19072), .C2(n19718), .A(n18941), .B(n18940), .ZN(
        P2_U2842) );
  NAND2_X1 U21153 ( .A1(n11223), .A2(n18942), .ZN(n18943) );
  XOR2_X1 U21154 ( .A(n18944), .B(n18943), .Z(n18952) );
  AOI22_X1 U21155 ( .A1(n18945), .A2(n19068), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19028), .ZN(n18946) );
  OAI21_X1 U21156 ( .B1(n13484), .B2(n19059), .A(n18946), .ZN(n18947) );
  AOI211_X1 U21157 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n11144), .A(n19142), .B(
        n18947), .ZN(n18951) );
  OAI22_X1 U21158 ( .A1(n18948), .A2(n19011), .B1(n19715), .B2(n19072), .ZN(
        n18949) );
  INV_X1 U21159 ( .A(n18949), .ZN(n18950) );
  OAI211_X1 U21160 ( .C1(n19230), .C2(n18952), .A(n18951), .B(n18950), .ZN(
        P2_U2841) );
  NOR2_X1 U21161 ( .A1(n19054), .A2(n18953), .ZN(n18955) );
  XOR2_X1 U21162 ( .A(n18955), .B(n18954), .Z(n18965) );
  NAND2_X1 U21163 ( .A1(n18956), .A2(n19067), .ZN(n18961) );
  AOI22_X1 U21164 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19009), .ZN(n18957) );
  NAND2_X1 U21165 ( .A1(n18958), .A2(n18957), .ZN(n18959) );
  AOI21_X1 U21166 ( .B1(n11144), .B2(P2_EBX_REG_15__SCAN_IN), .A(n18959), .ZN(
        n18960) );
  OAI211_X1 U21167 ( .C1(n19072), .C2(n19712), .A(n18961), .B(n18960), .ZN(
        n18962) );
  AOI21_X1 U21168 ( .B1(n18963), .B2(n19068), .A(n18962), .ZN(n18964) );
  OAI21_X1 U21169 ( .B1(n19230), .B2(n18965), .A(n18964), .ZN(P2_U2840) );
  NOR2_X1 U21170 ( .A1(n19054), .A2(n18966), .ZN(n18967) );
  XOR2_X1 U21171 ( .A(n18968), .B(n18967), .Z(n18977) );
  AOI22_X1 U21172 ( .A1(n18969), .A2(n19068), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19028), .ZN(n18970) );
  OAI21_X1 U21173 ( .B1(n17457), .B2(n19059), .A(n18970), .ZN(n18971) );
  AOI211_X1 U21174 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n11144), .A(n19142), .B(
        n18971), .ZN(n18976) );
  OAI22_X1 U21175 ( .A1(n18973), .A2(n19011), .B1(n18972), .B2(n19072), .ZN(
        n18974) );
  INV_X1 U21176 ( .A(n18974), .ZN(n18975) );
  OAI211_X1 U21177 ( .C1(n19230), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P2_U2838) );
  NAND2_X1 U21178 ( .A1(n11222), .A2(n18978), .ZN(n18979) );
  XOR2_X1 U21179 ( .A(n18980), .B(n18979), .Z(n18991) );
  AOI22_X1 U21180 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19009), .ZN(n18981) );
  OAI21_X1 U21181 ( .B1(n18982), .B2(n18996), .A(n18981), .ZN(n18983) );
  AOI211_X1 U21182 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n11144), .A(n19142), .B(
        n18983), .ZN(n18990) );
  NAND2_X1 U21183 ( .A1(n18985), .A2(n18984), .ZN(n18987) );
  INV_X1 U21184 ( .A(n17186), .ZN(n18986) );
  NAND2_X1 U21185 ( .A1(n18987), .A2(n18986), .ZN(n20171) );
  NOR2_X1 U21186 ( .A1(n19072), .A2(n20171), .ZN(n18988) );
  AOI21_X1 U21187 ( .B1(n19148), .B2(n19067), .A(n18988), .ZN(n18989) );
  OAI211_X1 U21188 ( .C1(n19230), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P2_U2837) );
  NOR2_X1 U21189 ( .A1(n19054), .A2(n18992), .ZN(n18993) );
  XOR2_X1 U21190 ( .A(n18994), .B(n18993), .Z(n19004) );
  AOI22_X1 U21191 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19009), .ZN(n18995) );
  OAI21_X1 U21192 ( .B1(n18997), .B2(n18996), .A(n18995), .ZN(n18998) );
  AOI211_X1 U21193 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n11144), .A(n19142), .B(
        n18998), .ZN(n19003) );
  OAI22_X1 U21194 ( .A1(n19011), .A2(n19000), .B1(n19072), .B2(n18999), .ZN(
        n19001) );
  INV_X1 U21195 ( .A(n19001), .ZN(n19002) );
  OAI211_X1 U21196 ( .C1(n19230), .C2(n19004), .A(n19003), .B(n19002), .ZN(
        P2_U2836) );
  OAI22_X1 U21197 ( .A1(n19007), .A2(n19006), .B1(n19061), .B2(n19005), .ZN(
        n19008) );
  AOI21_X1 U21198 ( .B1(P2_REIP_REG_21__SCAN_IN), .B2(n19009), .A(n19008), 
        .ZN(n19010) );
  OAI21_X1 U21199 ( .B1(n19012), .B2(n19011), .A(n19010), .ZN(n19013) );
  AOI21_X1 U21200 ( .B1(n19014), .B2(n19068), .A(n19013), .ZN(n19021) );
  NOR2_X1 U21201 ( .A1(n19054), .A2(n19015), .ZN(n19018) );
  INV_X1 U21202 ( .A(n19018), .ZN(n19016) );
  OAI221_X1 U21203 ( .B1(n19019), .B2(n19018), .C1(n19017), .C2(n19016), .A(
        n19055), .ZN(n19020) );
  OAI211_X1 U21204 ( .C1(n19072), .C2(n19022), .A(n19021), .B(n19020), .ZN(
        P2_U2834) );
  NAND2_X1 U21205 ( .A1(n11223), .A2(n19023), .ZN(n19025) );
  XOR2_X1 U21206 ( .A(n19026), .B(n19025), .Z(n19036) );
  NAND2_X1 U21207 ( .A1(n19027), .A2(n19067), .ZN(n19030) );
  AOI22_X1 U21208 ( .A1(n11144), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19028), .ZN(n19029) );
  OAI211_X1 U21209 ( .C1(n19031), .C2(n19059), .A(n19030), .B(n19029), .ZN(
        n19032) );
  AOI21_X1 U21210 ( .B1(n19033), .B2(n19068), .A(n19032), .ZN(n19034) );
  INV_X1 U21211 ( .A(n19034), .ZN(n19035) );
  AOI21_X1 U21212 ( .B1(n19055), .B2(n19036), .A(n19035), .ZN(n19037) );
  OAI21_X1 U21213 ( .B1(n19038), .B2(n19072), .A(n19037), .ZN(P2_U2833) );
  NOR2_X1 U21214 ( .A1(n19054), .A2(n19039), .ZN(n19041) );
  OAI21_X1 U21215 ( .B1(n19042), .B2(n19041), .A(n19055), .ZN(n19040) );
  AOI21_X1 U21216 ( .B1(n19042), .B2(n19041), .A(n19040), .ZN(n19046) );
  OAI22_X1 U21217 ( .A1(n19044), .A2(n19061), .B1(n19043), .B2(n19059), .ZN(
        n19045) );
  AOI211_X1 U21218 ( .C1(n11144), .C2(P2_EBX_REG_25__SCAN_IN), .A(n19046), .B(
        n19045), .ZN(n19051) );
  INV_X1 U21219 ( .A(n19047), .ZN(n19048) );
  AOI22_X1 U21220 ( .A1(n19049), .A2(n19068), .B1(n19067), .B2(n19048), .ZN(
        n19050) );
  OAI211_X1 U21221 ( .C1(n19052), .C2(n19072), .A(n19051), .B(n19050), .ZN(
        P2_U2830) );
  NOR2_X1 U21222 ( .A1(n19054), .A2(n19053), .ZN(n19057) );
  OAI21_X1 U21223 ( .B1(n19058), .B2(n19057), .A(n19055), .ZN(n19056) );
  AOI21_X1 U21224 ( .B1(n19058), .B2(n19057), .A(n19056), .ZN(n19064) );
  OAI22_X1 U21225 ( .A1(n19062), .A2(n19061), .B1(n19060), .B2(n19059), .ZN(
        n19063) );
  AOI211_X1 U21226 ( .C1(n11144), .C2(P2_EBX_REG_29__SCAN_IN), .A(n19064), .B(
        n19063), .ZN(n19071) );
  AOI22_X1 U21227 ( .A1(n19069), .A2(n19068), .B1(n19067), .B2(n19066), .ZN(
        n19070) );
  OAI211_X1 U21228 ( .C1(n19073), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        P2_U2826) );
  INV_X1 U21229 ( .A(n19099), .ZN(n19102) );
  OR2_X1 U21230 ( .A1(n19075), .A2(n19074), .ZN(n19091) );
  OAI21_X1 U21231 ( .B1(n19082), .B2(n19076), .A(n17630), .ZN(n19078) );
  OAI211_X1 U21232 ( .C1(n19080), .C2(n19079), .A(n19078), .B(n19077), .ZN(
        n19088) );
  INV_X1 U21233 ( .A(n19081), .ZN(n19085) );
  NAND3_X1 U21234 ( .A1(n19082), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19083) );
  OAI211_X1 U21235 ( .C1(n19086), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        n19087) );
  MUX2_X1 U21236 ( .A(n19088), .B(n19087), .S(n12519), .Z(n19089) );
  INV_X1 U21237 ( .A(n19089), .ZN(n19090) );
  NAND2_X1 U21238 ( .A1(n19091), .A2(n19090), .ZN(n19169) );
  INV_X1 U21239 ( .A(n19169), .ZN(n19092) );
  OAI22_X1 U21240 ( .A1(n20018), .A2(n19236), .B1(n19092), .B2(n19224), .ZN(
        n19093) );
  OAI22_X1 U21241 ( .A1(n19102), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19093), .B2(n19099), .ZN(n19094) );
  INV_X1 U21242 ( .A(n19094), .ZN(P2_U3596) );
  NOR2_X1 U21243 ( .A1(n19096), .A2(n19095), .ZN(n19097) );
  NAND2_X1 U21244 ( .A1(n19098), .A2(n19097), .ZN(n19203) );
  OR3_X1 U21245 ( .A1(n19099), .A2(n19224), .A3(n19203), .ZN(n19100) );
  OAI21_X1 U21246 ( .B1(n19102), .B2(n19101), .A(n19100), .ZN(P2_U3595) );
  OAI22_X1 U21247 ( .A1(n19104), .A2(n19112), .B1(n19134), .B2(n19103), .ZN(
        n19105) );
  INV_X1 U21248 ( .A(n19105), .ZN(n19118) );
  NAND2_X1 U21249 ( .A1(n19106), .A2(n19160), .ZN(n19109) );
  NAND2_X1 U21250 ( .A1(n19107), .A2(n19157), .ZN(n19108) );
  OAI211_X1 U21251 ( .C1(n19110), .C2(n19130), .A(n19109), .B(n19108), .ZN(
        n19111) );
  INV_X1 U21252 ( .A(n19111), .ZN(n19117) );
  NAND2_X1 U21253 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19142), .ZN(n19116) );
  NAND3_X1 U21254 ( .A1(n19114), .A2(n19113), .A3(n19112), .ZN(n19115) );
  NAND4_X1 U21255 ( .A1(n19118), .A2(n19117), .A3(n19116), .A4(n19115), .ZN(
        P2_U3022) );
  OAI22_X1 U21256 ( .A1(n19119), .A2(n13121), .B1(n19134), .B2(n19718), .ZN(
        n19120) );
  AOI21_X1 U21257 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19142), .A(n19120), 
        .ZN(n19127) );
  OAI22_X1 U21258 ( .A1(n19124), .A2(n19123), .B1(n19130), .B2(n19122), .ZN(
        n19125) );
  AOI21_X1 U21259 ( .B1(n17765), .B2(n19157), .A(n19125), .ZN(n19126) );
  OAI211_X1 U21260 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        P2_U3033) );
  NOR2_X1 U21261 ( .A1(n19131), .A2(n19130), .ZN(n19136) );
  OAI21_X1 U21262 ( .B1(n19134), .B2(n19133), .A(n19132), .ZN(n19135) );
  AOI211_X1 U21263 ( .C1(n19137), .C2(n19160), .A(n19136), .B(n19135), .ZN(
        n19138) );
  OAI221_X1 U21264 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19141), 
        .C1(n19140), .C2(n19139), .A(n19138), .ZN(P2_U3030) );
  INV_X1 U21265 ( .A(n20171), .ZN(n19147) );
  NAND2_X1 U21266 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19142), .ZN(n19143) );
  OAI211_X1 U21267 ( .C1(n19145), .C2(n13175), .A(n19144), .B(n19143), .ZN(
        n19146) );
  AOI21_X1 U21268 ( .B1(n19147), .B2(n19154), .A(n19146), .ZN(n19151) );
  AOI22_X1 U21269 ( .A1(n19149), .A2(n19160), .B1(n19159), .B2(n19148), .ZN(
        n19150) );
  OAI211_X1 U21270 ( .C1(n19153), .C2(n19152), .A(n19151), .B(n19150), .ZN(
        P2_U3028) );
  AOI22_X1 U21271 ( .A1(n19155), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19154), .B2(n19731), .ZN(n19167) );
  AOI222_X1 U21272 ( .A1(n19161), .A2(n19160), .B1(n19159), .B2(n19158), .C1(
        n19157), .C2(n19156), .ZN(n19166) );
  NAND2_X1 U21273 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19142), .ZN(n19165) );
  OAI211_X1 U21274 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n19163), .B(n19162), .ZN(n19164) );
  NAND4_X1 U21275 ( .A1(n19167), .A2(n19166), .A3(n19165), .A4(n19164), .ZN(
        P2_U3038) );
  NAND2_X1 U21276 ( .A1(n19184), .A2(n12519), .ZN(n19168) );
  OAI21_X1 U21277 ( .B1(n19169), .B2(n19184), .A(n19168), .ZN(n19183) );
  INV_X1 U21278 ( .A(n19184), .ZN(n19173) );
  MUX2_X1 U21279 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19174), .S(
        n19173), .Z(n19210) );
  NAND2_X1 U21280 ( .A1(n19170), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19171) );
  OAI21_X1 U21281 ( .B1(n19172), .B2(n19171), .A(n19910), .ZN(n19177) );
  NAND2_X1 U21282 ( .A1(n19172), .A2(n19171), .ZN(n19176) );
  OAI21_X1 U21283 ( .B1(n19906), .B2(n19174), .A(n19173), .ZN(n19175) );
  AOI21_X1 U21284 ( .B1(n19177), .B2(n19176), .A(n19175), .ZN(n19178) );
  AOI21_X1 U21285 ( .B1(n19210), .B2(n19906), .A(n19178), .ZN(n19179) );
  OAI21_X1 U21286 ( .B1(n19183), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19179), .ZN(n19182) );
  NAND2_X1 U21287 ( .A1(n19183), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19180) );
  NAND3_X1 U21288 ( .A1(n19182), .A2(n19181), .A3(n19180), .ZN(n19213) );
  INV_X1 U21289 ( .A(n19183), .ZN(n19211) );
  NAND2_X1 U21290 ( .A1(n19184), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19208) );
  INV_X1 U21291 ( .A(n19185), .ZN(n19198) );
  INV_X1 U21292 ( .A(n19186), .ZN(n19187) );
  OAI22_X1 U21293 ( .A1(n19242), .A2(n19189), .B1(n19188), .B2(n19187), .ZN(
        n19191) );
  NAND2_X1 U21294 ( .A1(n19191), .A2(n19190), .ZN(n19196) );
  AOI22_X1 U21295 ( .A1(n19197), .A2(n19194), .B1(n19193), .B2(n19192), .ZN(
        n19195) );
  OAI211_X1 U21296 ( .C1(n19198), .C2(n19197), .A(n19196), .B(n19195), .ZN(
        n19249) );
  INV_X1 U21297 ( .A(n19199), .ZN(n19200) );
  NOR3_X1 U21298 ( .A1(n19202), .A2(n19201), .A3(n19200), .ZN(n19248) );
  OAI21_X1 U21299 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19248), .ZN(n19204) );
  NAND3_X1 U21300 ( .A1(n19205), .A2(n19204), .A3(n19203), .ZN(n19206) );
  NOR2_X1 U21301 ( .A1(n19249), .A2(n19206), .ZN(n19207) );
  NAND2_X1 U21302 ( .A1(n19208), .A2(n19207), .ZN(n19209) );
  AOI21_X1 U21303 ( .B1(n19211), .B2(n19210), .A(n19209), .ZN(n19212) );
  NOR2_X1 U21304 ( .A1(n19835), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19214) );
  NAND2_X1 U21305 ( .A1(n19246), .A2(n19214), .ZN(n19216) );
  NAND2_X1 U21306 ( .A1(n19216), .A2(n19215), .ZN(n19221) );
  INV_X1 U21307 ( .A(n19217), .ZN(n19219) );
  NAND2_X1 U21308 ( .A1(n19219), .A2(n19218), .ZN(n19220) );
  NOR2_X1 U21309 ( .A1(n19233), .A2(n19222), .ZN(n19239) );
  INV_X1 U21310 ( .A(n19239), .ZN(n19229) );
  OAI21_X1 U21311 ( .B1(n19224), .B2(n19223), .A(n19247), .ZN(n19228) );
  NAND2_X1 U21312 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19835), .ZN(n19226) );
  NAND2_X1 U21313 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22275), .ZN(n19225) );
  AOI21_X1 U21314 ( .B1(n19226), .B2(n19229), .A(n19225), .ZN(n19227) );
  AOI21_X1 U21315 ( .B1(n19229), .B2(n19228), .A(n19227), .ZN(n19231) );
  NAND2_X1 U21316 ( .A1(n19231), .A2(n19230), .ZN(P2_U3177) );
  OAI221_X1 U21317 ( .B1(n19834), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19834), 
        .C2(n19233), .A(n19232), .ZN(P2_U3593) );
  OAI221_X1 U21318 ( .B1(n19234), .B2(n22275), .C1(n19234), .C2(n19835), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19245) );
  AOI21_X1 U21319 ( .B1(n19237), .B2(n19236), .A(n19235), .ZN(n19238) );
  AOI21_X1 U21320 ( .B1(n19239), .B2(n22275), .A(n19238), .ZN(n19241) );
  AOI211_X1 U21321 ( .C1(n19243), .C2(n19242), .A(n19241), .B(n19240), .ZN(
        n19244) );
  OAI211_X1 U21322 ( .C1(n19246), .C2(n19247), .A(n19245), .B(n19244), .ZN(
        P2_U3176) );
  NOR2_X1 U21323 ( .A1(n19248), .A2(n19247), .ZN(n19251) );
  MUX2_X1 U21324 ( .A(P2_MORE_REG_SCAN_IN), .B(n19249), .S(n19251), .Z(
        P2_U3609) );
  OAI21_X1 U21325 ( .B1(n19251), .B2(n12926), .A(n19250), .ZN(P2_U2819) );
  INV_X1 U21326 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20707) );
  INV_X1 U21327 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U21328 ( .A1(n19603), .A2(n20707), .B1(n19751), .B2(U215), .ZN(U282) );
  OAI22_X1 U21329 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19603), .ZN(n19252) );
  INV_X1 U21330 ( .A(n19252), .ZN(U281) );
  OAI22_X1 U21331 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19603), .ZN(n19253) );
  INV_X1 U21332 ( .A(n19253), .ZN(U280) );
  OAI22_X1 U21333 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19603), .ZN(n19254) );
  INV_X1 U21334 ( .A(n19254), .ZN(U279) );
  OAI22_X1 U21335 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19603), .ZN(n19255) );
  INV_X1 U21336 ( .A(n19255), .ZN(U278) );
  OAI22_X1 U21337 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19603), .ZN(n19256) );
  INV_X1 U21338 ( .A(n19256), .ZN(U277) );
  OAI22_X1 U21339 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19603), .ZN(n19257) );
  INV_X1 U21340 ( .A(n19257), .ZN(U276) );
  OAI22_X1 U21341 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19603), .ZN(n19258) );
  INV_X1 U21342 ( .A(n19258), .ZN(U275) );
  OAI22_X1 U21343 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19603), .ZN(n19259) );
  INV_X1 U21344 ( .A(n19259), .ZN(U274) );
  OAI22_X1 U21345 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19603), .ZN(n19260) );
  INV_X1 U21346 ( .A(n19260), .ZN(U273) );
  OAI22_X1 U21347 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19603), .ZN(n19261) );
  INV_X1 U21348 ( .A(n19261), .ZN(U272) );
  OAI22_X1 U21349 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19603), .ZN(n19262) );
  INV_X1 U21350 ( .A(n19262), .ZN(U271) );
  OAI22_X1 U21351 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19275), .ZN(n19263) );
  INV_X1 U21352 ( .A(n19263), .ZN(U270) );
  OAI22_X1 U21353 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19603), .ZN(n19264) );
  INV_X1 U21354 ( .A(n19264), .ZN(U269) );
  OAI22_X1 U21355 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19275), .ZN(n19265) );
  INV_X1 U21356 ( .A(n19265), .ZN(U268) );
  OAI22_X1 U21357 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19603), .ZN(n19266) );
  INV_X1 U21358 ( .A(n19266), .ZN(U267) );
  OAI22_X1 U21359 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19275), .ZN(n19267) );
  INV_X1 U21360 ( .A(n19267), .ZN(U266) );
  OAI22_X1 U21361 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19603), .ZN(n19268) );
  INV_X1 U21362 ( .A(n19268), .ZN(U265) );
  OAI22_X1 U21363 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19275), .ZN(n19269) );
  INV_X1 U21364 ( .A(n19269), .ZN(U264) );
  OAI22_X1 U21365 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19275), .ZN(n19270) );
  INV_X1 U21366 ( .A(n19270), .ZN(U263) );
  OAI22_X1 U21367 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19275), .ZN(n19271) );
  INV_X1 U21368 ( .A(n19271), .ZN(U262) );
  OAI22_X1 U21369 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19275), .ZN(n19272) );
  INV_X1 U21370 ( .A(n19272), .ZN(U261) );
  OAI22_X1 U21371 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19275), .ZN(n19273) );
  INV_X1 U21372 ( .A(n19273), .ZN(U260) );
  OAI22_X1 U21373 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19275), .ZN(n19274) );
  INV_X1 U21374 ( .A(n19274), .ZN(U259) );
  OAI22_X1 U21375 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19275), .ZN(n19276) );
  INV_X1 U21376 ( .A(n19276), .ZN(U258) );
  NOR2_X1 U21377 ( .A1(n21864), .A2(n19277), .ZN(n19343) );
  NAND2_X1 U21378 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19343), .ZN(
        n19695) );
  NOR2_X1 U21379 ( .A1(n19279), .A2(n19278), .ZN(n19396) );
  NAND2_X1 U21380 ( .A1(n19396), .A2(n21290), .ZN(n19356) );
  NAND2_X1 U21381 ( .A1(n19288), .A2(n21855), .ZN(n19287) );
  INV_X1 U21382 ( .A(n19287), .ZN(n19281) );
  NAND2_X1 U21383 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19281), .ZN(
        n19706) );
  INV_X1 U21384 ( .A(n19706), .ZN(n19620) );
  AND2_X1 U21385 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19606), .ZN(n19353) );
  AND2_X1 U21386 ( .A1(n21876), .A2(n19343), .ZN(n19608) );
  INV_X1 U21387 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21223) );
  NOR2_X2 U21388 ( .A1(n21223), .A2(n19518), .ZN(n19348) );
  AOI22_X1 U21389 ( .A1(n19620), .A2(n19353), .B1(n19608), .B2(n19348), .ZN(
        n19283) );
  NOR2_X1 U21390 ( .A1(n19280), .A2(n19518), .ZN(n19296) );
  AOI22_X1 U21391 ( .A1(n19606), .A2(n19281), .B1(n19343), .B2(n19296), .ZN(
        n19611) );
  NAND2_X1 U21392 ( .A1(n21852), .A2(n19281), .ZN(n19618) );
  INV_X1 U21393 ( .A(n19618), .ZN(n19626) );
  NOR2_X2 U21394 ( .A1(n19516), .A2(n19751), .ZN(n19349) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19611), .B1(
        n19626), .B2(n19349), .ZN(n19282) );
  OAI211_X1 U21396 ( .C1(n19695), .C2(n19356), .A(n19283), .B(n19282), .ZN(
        P3_U2995) );
  NAND2_X1 U21397 ( .A1(n19343), .A2(n21852), .ZN(n19602) );
  NAND2_X1 U21398 ( .A1(n21861), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19303) );
  NOR2_X1 U21399 ( .A1(n21855), .A2(n19303), .ZN(n19295) );
  NAND2_X1 U21400 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19295), .ZN(
        n19624) );
  INV_X1 U21401 ( .A(n19624), .ZN(n19632) );
  NAND2_X1 U21402 ( .A1(n19706), .A2(n19602), .ZN(n19352) );
  AND2_X1 U21403 ( .A1(n21876), .A2(n19352), .ZN(n19614) );
  AOI22_X1 U21404 ( .A1(n19349), .A2(n19632), .B1(n19348), .B2(n19614), .ZN(
        n19286) );
  NAND2_X1 U21405 ( .A1(n19618), .A2(n19624), .ZN(n19291) );
  NOR2_X1 U21406 ( .A1(n19518), .A2(n19284), .ZN(n19351) );
  AOI22_X1 U21407 ( .A1(n19606), .A2(n19291), .B1(n19351), .B2(n19352), .ZN(
        n19615) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19615), .B1(
        n19626), .B2(n19353), .ZN(n19285) );
  OAI211_X1 U21409 ( .C1(n19356), .C2(n19602), .A(n19286), .B(n19285), .ZN(
        P3_U2987) );
  NAND2_X1 U21410 ( .A1(n21852), .A2(n19295), .ZN(n19630) );
  INV_X1 U21411 ( .A(n19630), .ZN(n19637) );
  NOR2_X1 U21412 ( .A1(n19347), .A2(n19287), .ZN(n19619) );
  AOI22_X1 U21413 ( .A1(n19349), .A2(n19637), .B1(n19348), .B2(n19619), .ZN(
        n19290) );
  AND2_X1 U21414 ( .A1(n21855), .A2(n19296), .ZN(n19341) );
  AOI22_X1 U21415 ( .A1(n19606), .A2(n19295), .B1(n19288), .B2(n19341), .ZN(
        n19621) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19621), .B1(
        n19353), .B2(n19632), .ZN(n19289) );
  OAI211_X1 U21417 ( .C1(n19356), .C2(n19706), .A(n19290), .B(n19289), .ZN(
        P3_U2979) );
  AND2_X1 U21418 ( .A1(n21876), .A2(n19291), .ZN(n19625) );
  AOI22_X1 U21419 ( .A1(n19353), .A2(n19637), .B1(n19348), .B2(n19625), .ZN(
        n19293) );
  INV_X1 U21420 ( .A(n19303), .ZN(n19304) );
  NOR2_X1 U21421 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21852), .ZN(
        n19335) );
  NAND2_X1 U21422 ( .A1(n19304), .A2(n19335), .ZN(n19530) );
  NAND2_X1 U21423 ( .A1(n19630), .A2(n19530), .ZN(n19299) );
  AOI22_X1 U21424 ( .A1(n19606), .A2(n19299), .B1(n19351), .B2(n19291), .ZN(
        n19627) );
  INV_X1 U21425 ( .A(n19530), .ZN(n19643) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19627), .B1(
        n19349), .B2(n19643), .ZN(n19292) );
  OAI211_X1 U21427 ( .C1(n19618), .C2(n19356), .A(n19293), .B(n19292), .ZN(
        P3_U2971) );
  NAND2_X1 U21428 ( .A1(n21855), .A2(n21852), .ZN(n21857) );
  NOR2_X2 U21429 ( .A1(n21857), .A2(n19303), .ZN(n19648) );
  INV_X1 U21430 ( .A(n19295), .ZN(n19294) );
  NOR2_X1 U21431 ( .A1(n19347), .A2(n19294), .ZN(n19631) );
  AOI22_X1 U21432 ( .A1(n19349), .A2(n19648), .B1(n19348), .B2(n19631), .ZN(
        n19298) );
  AOI22_X1 U21433 ( .A1(n19606), .A2(n19304), .B1(n19296), .B2(n19295), .ZN(
        n19633) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19633), .B1(
        n19353), .B2(n19643), .ZN(n19297) );
  OAI211_X1 U21435 ( .C1(n19356), .C2(n19624), .A(n19298), .B(n19297), .ZN(
        P3_U2963) );
  AND2_X1 U21436 ( .A1(n21876), .A2(n19299), .ZN(n19636) );
  AOI22_X1 U21437 ( .A1(n19353), .A2(n19648), .B1(n19348), .B2(n19636), .ZN(
        n19302) );
  INV_X1 U21438 ( .A(n19648), .ZN(n19641) );
  NAND2_X1 U21439 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19311), .ZN(
        n19573) );
  NAND2_X1 U21440 ( .A1(n19641), .A2(n19573), .ZN(n19308) );
  INV_X1 U21441 ( .A(n19308), .ZN(n19307) );
  OAI22_X1 U21442 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19530), .B1(n19307), 
        .B2(n19333), .ZN(n19300) );
  OAI21_X1 U21443 ( .B1(n19637), .B2(n19300), .A(n19607), .ZN(n19638) );
  INV_X1 U21444 ( .A(n19573), .ZN(n19654) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19638), .B1(
        n19349), .B2(n19654), .ZN(n19301) );
  OAI211_X1 U21446 ( .C1(n19356), .C2(n19630), .A(n19302), .B(n19301), .ZN(
        P3_U2955) );
  NAND2_X1 U21447 ( .A1(n21852), .A2(n19311), .ZN(n19652) );
  INV_X1 U21448 ( .A(n19652), .ZN(n19660) );
  NAND2_X1 U21449 ( .A1(n21855), .A2(n21876), .ZN(n19339) );
  NOR2_X1 U21450 ( .A1(n19303), .A2(n19339), .ZN(n19642) );
  AOI22_X1 U21451 ( .A1(n19349), .A2(n19660), .B1(n19348), .B2(n19642), .ZN(
        n19306) );
  AOI22_X1 U21452 ( .A1(n19606), .A2(n19311), .B1(n19304), .B2(n19341), .ZN(
        n19644) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19644), .B1(
        n19353), .B2(n19654), .ZN(n19305) );
  OAI211_X1 U21454 ( .C1(n19356), .C2(n19530), .A(n19306), .B(n19305), .ZN(
        P3_U2947) );
  NOR2_X1 U21455 ( .A1(n19347), .A2(n19307), .ZN(n19647) );
  AOI22_X1 U21456 ( .A1(n19353), .A2(n19660), .B1(n19348), .B2(n19647), .ZN(
        n19310) );
  NAND2_X1 U21457 ( .A1(n21864), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19319) );
  INV_X1 U21458 ( .A(n19319), .ZN(n19320) );
  NAND2_X1 U21459 ( .A1(n19335), .A2(n19320), .ZN(n19658) );
  NAND2_X1 U21460 ( .A1(n19652), .A2(n19658), .ZN(n19315) );
  AOI22_X1 U21461 ( .A1(n19606), .A2(n19315), .B1(n19351), .B2(n19308), .ZN(
        n19649) );
  INV_X1 U21462 ( .A(n19658), .ZN(n19666) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19649), .B1(
        n19349), .B2(n19666), .ZN(n19309) );
  OAI211_X1 U21464 ( .C1(n19356), .C2(n19641), .A(n19310), .B(n19309), .ZN(
        P3_U2939) );
  AOI21_X1 U21465 ( .B1(n21855), .B2(n19333), .A(n19518), .ZN(n19327) );
  OAI211_X1 U21466 ( .C1(n19654), .C2(n21885), .A(n19320), .B(n19327), .ZN(
        n19655) );
  INV_X1 U21467 ( .A(n19311), .ZN(n19312) );
  NOR2_X1 U21468 ( .A1(n19347), .A2(n19312), .ZN(n19653) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19655), .B1(
        n19348), .B2(n19653), .ZN(n19314) );
  NOR2_X2 U21470 ( .A1(n21857), .A2(n19319), .ZN(n19671) );
  AOI22_X1 U21471 ( .A1(n19349), .A2(n19671), .B1(n19353), .B2(n19666), .ZN(
        n19313) );
  OAI211_X1 U21472 ( .C1(n19356), .C2(n19573), .A(n19314), .B(n19313), .ZN(
        P3_U2931) );
  AND2_X1 U21473 ( .A1(n21876), .A2(n19315), .ZN(n19659) );
  AOI22_X1 U21474 ( .A1(n19353), .A2(n19671), .B1(n19348), .B2(n19659), .ZN(
        n19318) );
  INV_X1 U21475 ( .A(n19671), .ZN(n19580) );
  NOR2_X1 U21476 ( .A1(n21855), .A2(n19340), .ZN(n19328) );
  NAND2_X1 U21477 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19328), .ZN(
        n19664) );
  NAND2_X1 U21478 ( .A1(n19580), .A2(n19664), .ZN(n19324) );
  INV_X1 U21479 ( .A(n19324), .ZN(n19323) );
  OAI22_X1 U21480 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19658), .B1(n19323), 
        .B2(n19333), .ZN(n19316) );
  OAI21_X1 U21481 ( .B1(n19660), .B2(n19316), .A(n19607), .ZN(n19661) );
  INV_X1 U21482 ( .A(n19664), .ZN(n19677) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19661), .B1(
        n19349), .B2(n19677), .ZN(n19317) );
  OAI211_X1 U21484 ( .C1(n19356), .C2(n19652), .A(n19318), .B(n19317), .ZN(
        P3_U2923) );
  NOR2_X1 U21485 ( .A1(n19339), .A2(n19319), .ZN(n19665) );
  AOI22_X1 U21486 ( .A1(n19353), .A2(n19677), .B1(n19348), .B2(n19665), .ZN(
        n19322) );
  AOI22_X1 U21487 ( .A1(n19606), .A2(n19328), .B1(n19341), .B2(n19320), .ZN(
        n19667) );
  NAND2_X1 U21488 ( .A1(n21852), .A2(n19328), .ZN(n19675) );
  INV_X1 U21489 ( .A(n19675), .ZN(n19683) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19667), .B1(
        n19349), .B2(n19683), .ZN(n19321) );
  OAI211_X1 U21491 ( .C1(n19356), .C2(n19658), .A(n19322), .B(n19321), .ZN(
        P3_U2915) );
  NOR2_X1 U21492 ( .A1(n19347), .A2(n19323), .ZN(n19670) );
  AOI22_X1 U21493 ( .A1(n19353), .A2(n19683), .B1(n19348), .B2(n19670), .ZN(
        n19326) );
  NAND2_X1 U21494 ( .A1(n19342), .A2(n19335), .ZN(n19589) );
  NAND2_X1 U21495 ( .A1(n19675), .A2(n19589), .ZN(n19332) );
  AOI22_X1 U21496 ( .A1(n19606), .A2(n19332), .B1(n19351), .B2(n19324), .ZN(
        n19672) );
  INV_X1 U21497 ( .A(n19589), .ZN(n19690) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19672), .B1(
        n19349), .B2(n19690), .ZN(n19325) );
  OAI211_X1 U21499 ( .C1(n19356), .C2(n19580), .A(n19326), .B(n19325), .ZN(
        P3_U2907) );
  NOR2_X1 U21500 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19340), .ZN(n19334) );
  OAI21_X1 U21501 ( .B1(n19677), .B2(n19334), .A(n19327), .ZN(n19678) );
  INV_X1 U21502 ( .A(n19328), .ZN(n19329) );
  NOR2_X1 U21503 ( .A1(n19347), .A2(n19329), .ZN(n19676) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19678), .B1(
        n19348), .B2(n19676), .ZN(n19331) );
  NOR2_X2 U21505 ( .A1(n21857), .A2(n19340), .ZN(n19701) );
  AOI22_X1 U21506 ( .A1(n19349), .A2(n19701), .B1(n19353), .B2(n19690), .ZN(
        n19330) );
  OAI211_X1 U21507 ( .C1(n19356), .C2(n19664), .A(n19331), .B(n19330), .ZN(
        P3_U2899) );
  INV_X1 U21508 ( .A(n19695), .ZN(n19682) );
  AND2_X1 U21509 ( .A1(n21876), .A2(n19332), .ZN(n19681) );
  AOI22_X1 U21510 ( .A1(n19349), .A2(n19682), .B1(n19348), .B2(n19681), .ZN(
        n19338) );
  INV_X1 U21511 ( .A(n19701), .ZN(n19687) );
  NAND2_X1 U21512 ( .A1(n19695), .A2(n19687), .ZN(n19350) );
  INV_X1 U21513 ( .A(n19350), .ZN(n19346) );
  OAI21_X1 U21514 ( .B1(n19346), .B2(n19333), .A(n19675), .ZN(n19336) );
  OAI221_X1 U21515 ( .B1(n19336), .B2(n19335), .C1(n19336), .C2(n19334), .A(
        n19607), .ZN(n19684) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19684), .B1(
        n19353), .B2(n19701), .ZN(n19337) );
  OAI211_X1 U21517 ( .C1(n19356), .C2(n19675), .A(n19338), .B(n19337), .ZN(
        P3_U2891) );
  NOR2_X1 U21518 ( .A1(n19340), .A2(n19339), .ZN(n19688) );
  AOI22_X1 U21519 ( .A1(n19682), .A2(n19353), .B1(n19348), .B2(n19688), .ZN(
        n19345) );
  AOI22_X1 U21520 ( .A1(n19606), .A2(n19343), .B1(n19342), .B2(n19341), .ZN(
        n19691) );
  INV_X1 U21521 ( .A(n19602), .ZN(n19699) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19691), .B1(
        n19349), .B2(n19699), .ZN(n19344) );
  OAI211_X1 U21523 ( .C1(n19356), .C2(n19589), .A(n19345), .B(n19344), .ZN(
        P3_U2883) );
  NOR2_X1 U21524 ( .A1(n19347), .A2(n19346), .ZN(n19697) );
  AOI22_X1 U21525 ( .A1(n19349), .A2(n19620), .B1(n19348), .B2(n19697), .ZN(
        n19355) );
  AOI22_X1 U21526 ( .A1(n19606), .A2(n19352), .B1(n19351), .B2(n19350), .ZN(
        n19702) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19702), .B1(
        n19353), .B2(n19699), .ZN(n19354) );
  OAI211_X1 U21528 ( .C1(n19356), .C2(n19687), .A(n19355), .B(n19354), .ZN(
        P3_U2875) );
  OAI22_X1 U21529 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19603), .ZN(n19357) );
  INV_X1 U21530 ( .A(n19357), .ZN(U257) );
  NAND2_X1 U21531 ( .A1(n19396), .A2(n19358), .ZN(n19394) );
  AND2_X1 U21532 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19606), .ZN(n19390) );
  INV_X1 U21533 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21271) );
  NOR2_X2 U21534 ( .A1(n21271), .A2(n19518), .ZN(n19389) );
  AOI22_X1 U21535 ( .A1(n19626), .A2(n19390), .B1(n19608), .B2(n19389), .ZN(
        n19360) );
  INV_X1 U21536 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n21265) );
  NOR2_X2 U21537 ( .A1(n21265), .A2(n19516), .ZN(n19391) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19611), .B1(
        n19620), .B2(n19391), .ZN(n19359) );
  OAI211_X1 U21539 ( .C1(n19695), .C2(n19394), .A(n19360), .B(n19359), .ZN(
        P3_U2994) );
  AOI22_X1 U21540 ( .A1(n19632), .A2(n19390), .B1(n19614), .B2(n19389), .ZN(
        n19362) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19615), .B1(
        n19626), .B2(n19391), .ZN(n19361) );
  OAI211_X1 U21542 ( .C1(n19602), .C2(n19394), .A(n19362), .B(n19361), .ZN(
        P3_U2986) );
  AOI22_X1 U21543 ( .A1(n19637), .A2(n19390), .B1(n19619), .B2(n19389), .ZN(
        n19364) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19621), .B1(
        n19632), .B2(n19391), .ZN(n19363) );
  OAI211_X1 U21545 ( .C1(n19706), .C2(n19394), .A(n19364), .B(n19363), .ZN(
        P3_U2978) );
  AOI22_X1 U21546 ( .A1(n19637), .A2(n19391), .B1(n19625), .B2(n19389), .ZN(
        n19366) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19627), .B1(
        n19643), .B2(n19390), .ZN(n19365) );
  OAI211_X1 U21548 ( .C1(n19618), .C2(n19394), .A(n19366), .B(n19365), .ZN(
        P3_U2970) );
  AOI22_X1 U21549 ( .A1(n19643), .A2(n19391), .B1(n19631), .B2(n19389), .ZN(
        n19368) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19633), .B1(
        n19648), .B2(n19390), .ZN(n19367) );
  OAI211_X1 U21551 ( .C1(n19624), .C2(n19394), .A(n19368), .B(n19367), .ZN(
        P3_U2962) );
  AOI22_X1 U21552 ( .A1(n19654), .A2(n19390), .B1(n19636), .B2(n19389), .ZN(
        n19370) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19638), .B1(
        n19648), .B2(n19391), .ZN(n19369) );
  OAI211_X1 U21554 ( .C1(n19630), .C2(n19394), .A(n19370), .B(n19369), .ZN(
        P3_U2954) );
  AOI22_X1 U21555 ( .A1(n19654), .A2(n19391), .B1(n19642), .B2(n19389), .ZN(
        n19372) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19644), .B1(
        n19660), .B2(n19390), .ZN(n19371) );
  OAI211_X1 U21557 ( .C1(n19530), .C2(n19394), .A(n19372), .B(n19371), .ZN(
        P3_U2946) );
  AOI22_X1 U21558 ( .A1(n19666), .A2(n19390), .B1(n19647), .B2(n19389), .ZN(
        n19374) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19649), .B1(
        n19660), .B2(n19391), .ZN(n19373) );
  OAI211_X1 U21560 ( .C1(n19641), .C2(n19394), .A(n19374), .B(n19373), .ZN(
        P3_U2938) );
  AOI22_X1 U21561 ( .A1(n19666), .A2(n19391), .B1(n19653), .B2(n19389), .ZN(
        n19376) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19655), .B1(
        n19671), .B2(n19390), .ZN(n19375) );
  OAI211_X1 U21563 ( .C1(n19573), .C2(n19394), .A(n19376), .B(n19375), .ZN(
        P3_U2930) );
  AOI22_X1 U21564 ( .A1(n19677), .A2(n19390), .B1(n19659), .B2(n19389), .ZN(
        n19378) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19661), .B1(
        n19671), .B2(n19391), .ZN(n19377) );
  OAI211_X1 U21566 ( .C1(n19652), .C2(n19394), .A(n19378), .B(n19377), .ZN(
        P3_U2922) );
  AOI22_X1 U21567 ( .A1(n19677), .A2(n19391), .B1(n19665), .B2(n19389), .ZN(
        n19380) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19667), .B1(
        n19683), .B2(n19390), .ZN(n19379) );
  OAI211_X1 U21569 ( .C1(n19658), .C2(n19394), .A(n19380), .B(n19379), .ZN(
        P3_U2914) );
  AOI22_X1 U21570 ( .A1(n19683), .A2(n19391), .B1(n19670), .B2(n19389), .ZN(
        n19382) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19672), .B1(
        n19690), .B2(n19390), .ZN(n19381) );
  OAI211_X1 U21572 ( .C1(n19580), .C2(n19394), .A(n19382), .B(n19381), .ZN(
        P3_U2906) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19678), .B1(
        n19676), .B2(n19389), .ZN(n19384) );
  AOI22_X1 U21574 ( .A1(n19690), .A2(n19391), .B1(n19701), .B2(n19390), .ZN(
        n19383) );
  OAI211_X1 U21575 ( .C1(n19664), .C2(n19394), .A(n19384), .B(n19383), .ZN(
        P3_U2898) );
  AOI22_X1 U21576 ( .A1(n19682), .A2(n19390), .B1(n19681), .B2(n19389), .ZN(
        n19386) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19684), .B1(
        n19701), .B2(n19391), .ZN(n19385) );
  OAI211_X1 U21578 ( .C1(n19675), .C2(n19394), .A(n19386), .B(n19385), .ZN(
        P3_U2890) );
  AOI22_X1 U21579 ( .A1(n19682), .A2(n19391), .B1(n19688), .B2(n19389), .ZN(
        n19388) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19691), .B1(
        n19699), .B2(n19390), .ZN(n19387) );
  OAI211_X1 U21581 ( .C1(n19589), .C2(n19394), .A(n19388), .B(n19387), .ZN(
        P3_U2882) );
  AOI22_X1 U21582 ( .A1(n19620), .A2(n19390), .B1(n19697), .B2(n19389), .ZN(
        n19393) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19702), .B1(
        n19699), .B2(n19391), .ZN(n19392) );
  OAI211_X1 U21584 ( .C1(n19687), .C2(n19394), .A(n19393), .B(n19392), .ZN(
        P3_U2874) );
  OAI22_X1 U21585 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19603), .ZN(n19395) );
  INV_X1 U21586 ( .A(n19395), .ZN(U256) );
  NAND2_X1 U21587 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19606), .ZN(n19428) );
  NAND2_X1 U21588 ( .A1(n19606), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19434) );
  INV_X1 U21589 ( .A(n19434), .ZN(n19425) );
  NOR2_X2 U21590 ( .A1(n19518), .A2(n21231), .ZN(n19429) );
  AOI22_X1 U21591 ( .A1(n19620), .A2(n19425), .B1(n19608), .B2(n19429), .ZN(
        n19398) );
  INV_X1 U21592 ( .A(n19396), .ZN(n19609) );
  NOR2_X2 U21593 ( .A1(n21252), .A2(n19609), .ZN(n19431) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19431), .ZN(n19397) );
  OAI211_X1 U21595 ( .C1(n19618), .C2(n19428), .A(n19398), .B(n19397), .ZN(
        P3_U2993) );
  AOI22_X1 U21596 ( .A1(n19626), .A2(n19425), .B1(n19614), .B2(n19429), .ZN(
        n19400) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19431), .ZN(n19399) );
  OAI211_X1 U21598 ( .C1(n19624), .C2(n19428), .A(n19400), .B(n19399), .ZN(
        P3_U2985) );
  INV_X1 U21599 ( .A(n19428), .ZN(n19430) );
  AOI22_X1 U21600 ( .A1(n19637), .A2(n19430), .B1(n19619), .B2(n19429), .ZN(
        n19402) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19431), .ZN(n19401) );
  OAI211_X1 U21602 ( .C1(n19624), .C2(n19434), .A(n19402), .B(n19401), .ZN(
        P3_U2977) );
  AOI22_X1 U21603 ( .A1(n19643), .A2(n19430), .B1(n19625), .B2(n19429), .ZN(
        n19404) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19431), .ZN(n19403) );
  OAI211_X1 U21605 ( .C1(n19630), .C2(n19434), .A(n19404), .B(n19403), .ZN(
        P3_U2969) );
  AOI22_X1 U21606 ( .A1(n19643), .A2(n19425), .B1(n19631), .B2(n19429), .ZN(
        n19406) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19431), .ZN(n19405) );
  OAI211_X1 U21608 ( .C1(n19641), .C2(n19428), .A(n19406), .B(n19405), .ZN(
        P3_U2961) );
  AOI22_X1 U21609 ( .A1(n19648), .A2(n19425), .B1(n19636), .B2(n19429), .ZN(
        n19408) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19431), .ZN(n19407) );
  OAI211_X1 U21611 ( .C1(n19573), .C2(n19428), .A(n19408), .B(n19407), .ZN(
        P3_U2953) );
  AOI22_X1 U21612 ( .A1(n19654), .A2(n19425), .B1(n19642), .B2(n19429), .ZN(
        n19410) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19431), .ZN(n19409) );
  OAI211_X1 U21614 ( .C1(n19652), .C2(n19428), .A(n19410), .B(n19409), .ZN(
        P3_U2945) );
  AOI22_X1 U21615 ( .A1(n19660), .A2(n19425), .B1(n19647), .B2(n19429), .ZN(
        n19412) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19431), .ZN(n19411) );
  OAI211_X1 U21617 ( .C1(n19658), .C2(n19428), .A(n19412), .B(n19411), .ZN(
        P3_U2937) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19655), .B1(
        n19653), .B2(n19429), .ZN(n19414) );
  AOI22_X1 U21619 ( .A1(n19654), .A2(n19431), .B1(n19666), .B2(n19425), .ZN(
        n19413) );
  OAI211_X1 U21620 ( .C1(n19580), .C2(n19428), .A(n19414), .B(n19413), .ZN(
        P3_U2929) );
  AOI22_X1 U21621 ( .A1(n19677), .A2(n19430), .B1(n19659), .B2(n19429), .ZN(
        n19416) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19431), .ZN(n19415) );
  OAI211_X1 U21623 ( .C1(n19580), .C2(n19434), .A(n19416), .B(n19415), .ZN(
        P3_U2921) );
  AOI22_X1 U21624 ( .A1(n19683), .A2(n19430), .B1(n19665), .B2(n19429), .ZN(
        n19418) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19431), .ZN(n19417) );
  OAI211_X1 U21626 ( .C1(n19664), .C2(n19434), .A(n19418), .B(n19417), .ZN(
        P3_U2913) );
  AOI22_X1 U21627 ( .A1(n19690), .A2(n19430), .B1(n19670), .B2(n19429), .ZN(
        n19420) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19431), .ZN(n19419) );
  OAI211_X1 U21629 ( .C1(n19675), .C2(n19434), .A(n19420), .B(n19419), .ZN(
        P3_U2905) );
  AOI22_X1 U21630 ( .A1(n19690), .A2(n19425), .B1(n19676), .B2(n19429), .ZN(
        n19422) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19431), .ZN(n19421) );
  OAI211_X1 U21632 ( .C1(n19687), .C2(n19428), .A(n19422), .B(n19421), .ZN(
        P3_U2897) );
  AOI22_X1 U21633 ( .A1(n19701), .A2(n19425), .B1(n19681), .B2(n19429), .ZN(
        n19424) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19431), .ZN(n19423) );
  OAI211_X1 U21635 ( .C1(n19695), .C2(n19428), .A(n19424), .B(n19423), .ZN(
        P3_U2889) );
  AOI22_X1 U21636 ( .A1(n19682), .A2(n19425), .B1(n19688), .B2(n19429), .ZN(
        n19427) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19431), .ZN(n19426) );
  OAI211_X1 U21638 ( .C1(n19602), .C2(n19428), .A(n19427), .B(n19426), .ZN(
        P3_U2881) );
  AOI22_X1 U21639 ( .A1(n19620), .A2(n19430), .B1(n19697), .B2(n19429), .ZN(
        n19433) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19431), .ZN(n19432) );
  OAI211_X1 U21641 ( .C1(n19602), .C2(n19434), .A(n19433), .B(n19432), .ZN(
        P3_U2873) );
  OAI22_X1 U21642 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19603), .ZN(n19435) );
  INV_X1 U21643 ( .A(n19435), .ZN(U255) );
  NAND2_X1 U21644 ( .A1(n19606), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19463) );
  NAND2_X1 U21645 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19606), .ZN(n19473) );
  INV_X1 U21646 ( .A(n19473), .ZN(n19460) );
  INV_X1 U21647 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21236) );
  NOR2_X2 U21648 ( .A1(n19518), .A2(n21236), .ZN(n19468) );
  AOI22_X1 U21649 ( .A1(n19626), .A2(n19460), .B1(n19608), .B2(n19468), .ZN(
        n19437) );
  NOR2_X2 U21650 ( .A1(n14120), .A2(n19609), .ZN(n19470) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19470), .ZN(n19436) );
  OAI211_X1 U21652 ( .C1(n19706), .C2(n19463), .A(n19437), .B(n19436), .ZN(
        P3_U2992) );
  INV_X1 U21653 ( .A(n19463), .ZN(n19469) );
  AOI22_X1 U21654 ( .A1(n19626), .A2(n19469), .B1(n19614), .B2(n19468), .ZN(
        n19439) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19470), .ZN(n19438) );
  OAI211_X1 U21656 ( .C1(n19624), .C2(n19473), .A(n19439), .B(n19438), .ZN(
        P3_U2984) );
  AOI22_X1 U21657 ( .A1(n19632), .A2(n19469), .B1(n19619), .B2(n19468), .ZN(
        n19441) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19470), .ZN(n19440) );
  OAI211_X1 U21659 ( .C1(n19630), .C2(n19473), .A(n19441), .B(n19440), .ZN(
        P3_U2976) );
  AOI22_X1 U21660 ( .A1(n19643), .A2(n19460), .B1(n19625), .B2(n19468), .ZN(
        n19443) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19470), .ZN(n19442) );
  OAI211_X1 U21662 ( .C1(n19630), .C2(n19463), .A(n19443), .B(n19442), .ZN(
        P3_U2968) );
  AOI22_X1 U21663 ( .A1(n19648), .A2(n19460), .B1(n19631), .B2(n19468), .ZN(
        n19445) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19470), .ZN(n19444) );
  OAI211_X1 U21665 ( .C1(n19530), .C2(n19463), .A(n19445), .B(n19444), .ZN(
        P3_U2960) );
  AOI22_X1 U21666 ( .A1(n19654), .A2(n19460), .B1(n19636), .B2(n19468), .ZN(
        n19447) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19470), .ZN(n19446) );
  OAI211_X1 U21668 ( .C1(n19641), .C2(n19463), .A(n19447), .B(n19446), .ZN(
        P3_U2952) );
  AOI22_X1 U21669 ( .A1(n19654), .A2(n19469), .B1(n19642), .B2(n19468), .ZN(
        n19449) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19470), .ZN(n19448) );
  OAI211_X1 U21671 ( .C1(n19652), .C2(n19473), .A(n19449), .B(n19448), .ZN(
        P3_U2944) );
  AOI22_X1 U21672 ( .A1(n19666), .A2(n19460), .B1(n19647), .B2(n19468), .ZN(
        n19451) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19470), .ZN(n19450) );
  OAI211_X1 U21674 ( .C1(n19652), .C2(n19463), .A(n19451), .B(n19450), .ZN(
        P3_U2936) );
  AOI22_X1 U21675 ( .A1(n19666), .A2(n19469), .B1(n19653), .B2(n19468), .ZN(
        n19453) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19470), .ZN(n19452) );
  OAI211_X1 U21677 ( .C1(n19580), .C2(n19473), .A(n19453), .B(n19452), .ZN(
        P3_U2928) );
  AOI22_X1 U21678 ( .A1(n19677), .A2(n19460), .B1(n19659), .B2(n19468), .ZN(
        n19455) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19470), .ZN(n19454) );
  OAI211_X1 U21680 ( .C1(n19580), .C2(n19463), .A(n19455), .B(n19454), .ZN(
        P3_U2920) );
  AOI22_X1 U21681 ( .A1(n19677), .A2(n19469), .B1(n19665), .B2(n19468), .ZN(
        n19457) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19470), .ZN(n19456) );
  OAI211_X1 U21683 ( .C1(n19675), .C2(n19473), .A(n19457), .B(n19456), .ZN(
        P3_U2912) );
  AOI22_X1 U21684 ( .A1(n19683), .A2(n19469), .B1(n19670), .B2(n19468), .ZN(
        n19459) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19470), .ZN(n19458) );
  OAI211_X1 U21686 ( .C1(n19589), .C2(n19473), .A(n19459), .B(n19458), .ZN(
        P3_U2904) );
  AOI22_X1 U21687 ( .A1(n19701), .A2(n19460), .B1(n19676), .B2(n19468), .ZN(
        n19462) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19470), .ZN(n19461) );
  OAI211_X1 U21689 ( .C1(n19589), .C2(n19463), .A(n19462), .B(n19461), .ZN(
        P3_U2896) );
  AOI22_X1 U21690 ( .A1(n19701), .A2(n19469), .B1(n19681), .B2(n19468), .ZN(
        n19465) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19470), .ZN(n19464) );
  OAI211_X1 U21692 ( .C1(n19695), .C2(n19473), .A(n19465), .B(n19464), .ZN(
        P3_U2888) );
  AOI22_X1 U21693 ( .A1(n19682), .A2(n19469), .B1(n19688), .B2(n19468), .ZN(
        n19467) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19470), .ZN(n19466) );
  OAI211_X1 U21695 ( .C1(n19602), .C2(n19473), .A(n19467), .B(n19466), .ZN(
        P3_U2880) );
  AOI22_X1 U21696 ( .A1(n19699), .A2(n19469), .B1(n19697), .B2(n19468), .ZN(
        n19472) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19470), .ZN(n19471) );
  OAI211_X1 U21698 ( .C1(n19706), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P3_U2872) );
  OAI22_X1 U21699 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19603), .ZN(n19474) );
  INV_X1 U21700 ( .A(n19474), .ZN(U254) );
  INV_X1 U21701 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19475) );
  NOR2_X1 U21702 ( .A1(n19475), .A2(n19516), .ZN(n19505) );
  INV_X1 U21703 ( .A(n19505), .ZN(n19514) );
  NAND2_X1 U21704 ( .A1(n19606), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19508) );
  INV_X1 U21705 ( .A(n19508), .ZN(n19510) );
  INV_X1 U21706 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21240) );
  NOR2_X2 U21707 ( .A1(n19518), .A2(n21240), .ZN(n19509) );
  AOI22_X1 U21708 ( .A1(n19620), .A2(n19510), .B1(n19608), .B2(n19509), .ZN(
        n19478) );
  NOR2_X2 U21709 ( .A1(n19476), .A2(n19609), .ZN(n19511) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19511), .ZN(n19477) );
  OAI211_X1 U21711 ( .C1(n19618), .C2(n19514), .A(n19478), .B(n19477), .ZN(
        P3_U2991) );
  AOI22_X1 U21712 ( .A1(n19632), .A2(n19505), .B1(n19614), .B2(n19509), .ZN(
        n19480) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19511), .ZN(n19479) );
  OAI211_X1 U21714 ( .C1(n19618), .C2(n19508), .A(n19480), .B(n19479), .ZN(
        P3_U2983) );
  AOI22_X1 U21715 ( .A1(n19637), .A2(n19505), .B1(n19619), .B2(n19509), .ZN(
        n19482) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19511), .ZN(n19481) );
  OAI211_X1 U21717 ( .C1(n19624), .C2(n19508), .A(n19482), .B(n19481), .ZN(
        P3_U2975) );
  AOI22_X1 U21718 ( .A1(n19637), .A2(n19510), .B1(n19625), .B2(n19509), .ZN(
        n19484) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19511), .ZN(n19483) );
  OAI211_X1 U21720 ( .C1(n19530), .C2(n19514), .A(n19484), .B(n19483), .ZN(
        P3_U2967) );
  AOI22_X1 U21721 ( .A1(n19648), .A2(n19505), .B1(n19631), .B2(n19509), .ZN(
        n19486) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19511), .ZN(n19485) );
  OAI211_X1 U21723 ( .C1(n19530), .C2(n19508), .A(n19486), .B(n19485), .ZN(
        P3_U2959) );
  AOI22_X1 U21724 ( .A1(n19648), .A2(n19510), .B1(n19636), .B2(n19509), .ZN(
        n19488) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19511), .ZN(n19487) );
  OAI211_X1 U21726 ( .C1(n19573), .C2(n19514), .A(n19488), .B(n19487), .ZN(
        P3_U2951) );
  AOI22_X1 U21727 ( .A1(n19660), .A2(n19505), .B1(n19642), .B2(n19509), .ZN(
        n19490) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19511), .ZN(n19489) );
  OAI211_X1 U21729 ( .C1(n19573), .C2(n19508), .A(n19490), .B(n19489), .ZN(
        P3_U2943) );
  AOI22_X1 U21730 ( .A1(n19666), .A2(n19505), .B1(n19647), .B2(n19509), .ZN(
        n19492) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19511), .ZN(n19491) );
  OAI211_X1 U21732 ( .C1(n19652), .C2(n19508), .A(n19492), .B(n19491), .ZN(
        P3_U2935) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19655), .B1(
        n19653), .B2(n19509), .ZN(n19494) );
  AOI22_X1 U21734 ( .A1(n19654), .A2(n19511), .B1(n19666), .B2(n19510), .ZN(
        n19493) );
  OAI211_X1 U21735 ( .C1(n19580), .C2(n19514), .A(n19494), .B(n19493), .ZN(
        P3_U2927) );
  AOI22_X1 U21736 ( .A1(n19671), .A2(n19510), .B1(n19659), .B2(n19509), .ZN(
        n19496) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19511), .ZN(n19495) );
  OAI211_X1 U21738 ( .C1(n19664), .C2(n19514), .A(n19496), .B(n19495), .ZN(
        P3_U2919) );
  AOI22_X1 U21739 ( .A1(n19677), .A2(n19510), .B1(n19665), .B2(n19509), .ZN(
        n19498) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19511), .ZN(n19497) );
  OAI211_X1 U21741 ( .C1(n19675), .C2(n19514), .A(n19498), .B(n19497), .ZN(
        P3_U2911) );
  AOI22_X1 U21742 ( .A1(n19690), .A2(n19505), .B1(n19670), .B2(n19509), .ZN(
        n19500) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19511), .ZN(n19499) );
  OAI211_X1 U21744 ( .C1(n19675), .C2(n19508), .A(n19500), .B(n19499), .ZN(
        P3_U2903) );
  AOI22_X1 U21745 ( .A1(n19701), .A2(n19505), .B1(n19676), .B2(n19509), .ZN(
        n19502) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19511), .ZN(n19501) );
  OAI211_X1 U21747 ( .C1(n19589), .C2(n19508), .A(n19502), .B(n19501), .ZN(
        P3_U2895) );
  AOI22_X1 U21748 ( .A1(n19682), .A2(n19505), .B1(n19681), .B2(n19509), .ZN(
        n19504) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19511), .ZN(n19503) );
  OAI211_X1 U21750 ( .C1(n19687), .C2(n19508), .A(n19504), .B(n19503), .ZN(
        P3_U2887) );
  AOI22_X1 U21751 ( .A1(n19699), .A2(n19505), .B1(n19688), .B2(n19509), .ZN(
        n19507) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19511), .ZN(n19506) );
  OAI211_X1 U21753 ( .C1(n19695), .C2(n19508), .A(n19507), .B(n19506), .ZN(
        P3_U2879) );
  AOI22_X1 U21754 ( .A1(n19699), .A2(n19510), .B1(n19697), .B2(n19509), .ZN(
        n19513) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19511), .ZN(n19512) );
  OAI211_X1 U21756 ( .C1(n19706), .C2(n19514), .A(n19513), .B(n19512), .ZN(
        P3_U2871) );
  OAI22_X1 U21757 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19603), .ZN(n19515) );
  INV_X1 U21758 ( .A(n19515), .ZN(U253) );
  INV_X1 U21759 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19517) );
  NOR2_X1 U21760 ( .A1(n19517), .A2(n19516), .ZN(n19554) );
  INV_X1 U21761 ( .A(n19554), .ZN(n19544) );
  NAND2_X1 U21762 ( .A1(n19606), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19558) );
  INV_X1 U21763 ( .A(n19558), .ZN(n19541) );
  INV_X1 U21764 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21246) );
  NOR2_X2 U21765 ( .A1(n19518), .A2(n21246), .ZN(n19553) );
  AOI22_X1 U21766 ( .A1(n19620), .A2(n19541), .B1(n19608), .B2(n19553), .ZN(
        n19521) );
  NOR2_X2 U21767 ( .A1(n19519), .A2(n19609), .ZN(n19555) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19555), .ZN(n19520) );
  OAI211_X1 U21769 ( .C1(n19618), .C2(n19544), .A(n19521), .B(n19520), .ZN(
        P3_U2990) );
  AOI22_X1 U21770 ( .A1(n19626), .A2(n19541), .B1(n19614), .B2(n19553), .ZN(
        n19523) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19555), .ZN(n19522) );
  OAI211_X1 U21772 ( .C1(n19624), .C2(n19544), .A(n19523), .B(n19522), .ZN(
        P3_U2982) );
  AOI22_X1 U21773 ( .A1(n19632), .A2(n19541), .B1(n19619), .B2(n19553), .ZN(
        n19525) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19555), .ZN(n19524) );
  OAI211_X1 U21775 ( .C1(n19630), .C2(n19544), .A(n19525), .B(n19524), .ZN(
        P3_U2974) );
  AOI22_X1 U21776 ( .A1(n19637), .A2(n19541), .B1(n19625), .B2(n19553), .ZN(
        n19527) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19555), .ZN(n19526) );
  OAI211_X1 U21778 ( .C1(n19530), .C2(n19544), .A(n19527), .B(n19526), .ZN(
        P3_U2966) );
  AOI22_X1 U21779 ( .A1(n19648), .A2(n19554), .B1(n19631), .B2(n19553), .ZN(
        n19529) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19555), .ZN(n19528) );
  OAI211_X1 U21781 ( .C1(n19530), .C2(n19558), .A(n19529), .B(n19528), .ZN(
        P3_U2958) );
  AOI22_X1 U21782 ( .A1(n19654), .A2(n19554), .B1(n19636), .B2(n19553), .ZN(
        n19532) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19555), .ZN(n19531) );
  OAI211_X1 U21784 ( .C1(n19641), .C2(n19558), .A(n19532), .B(n19531), .ZN(
        P3_U2950) );
  AOI22_X1 U21785 ( .A1(n19660), .A2(n19554), .B1(n19642), .B2(n19553), .ZN(
        n19534) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19555), .ZN(n19533) );
  OAI211_X1 U21787 ( .C1(n19573), .C2(n19558), .A(n19534), .B(n19533), .ZN(
        P3_U2942) );
  AOI22_X1 U21788 ( .A1(n19660), .A2(n19541), .B1(n19647), .B2(n19553), .ZN(
        n19536) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19555), .ZN(n19535) );
  OAI211_X1 U21790 ( .C1(n19658), .C2(n19544), .A(n19536), .B(n19535), .ZN(
        P3_U2934) );
  AOI22_X1 U21791 ( .A1(n19671), .A2(n19554), .B1(n19653), .B2(n19553), .ZN(
        n19538) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19555), .ZN(n19537) );
  OAI211_X1 U21793 ( .C1(n19658), .C2(n19558), .A(n19538), .B(n19537), .ZN(
        P3_U2926) );
  AOI22_X1 U21794 ( .A1(n19671), .A2(n19541), .B1(n19659), .B2(n19553), .ZN(
        n19540) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19555), .ZN(n19539) );
  OAI211_X1 U21796 ( .C1(n19664), .C2(n19544), .A(n19540), .B(n19539), .ZN(
        P3_U2918) );
  AOI22_X1 U21797 ( .A1(n19677), .A2(n19541), .B1(n19665), .B2(n19553), .ZN(
        n19543) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19555), .ZN(n19542) );
  OAI211_X1 U21799 ( .C1(n19675), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P3_U2910) );
  AOI22_X1 U21800 ( .A1(n19690), .A2(n19554), .B1(n19670), .B2(n19553), .ZN(
        n19546) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19555), .ZN(n19545) );
  OAI211_X1 U21802 ( .C1(n19675), .C2(n19558), .A(n19546), .B(n19545), .ZN(
        P3_U2902) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19678), .B1(
        n19676), .B2(n19553), .ZN(n19548) );
  AOI22_X1 U21804 ( .A1(n19677), .A2(n19555), .B1(n19701), .B2(n19554), .ZN(
        n19547) );
  OAI211_X1 U21805 ( .C1(n19589), .C2(n19558), .A(n19548), .B(n19547), .ZN(
        P3_U2894) );
  AOI22_X1 U21806 ( .A1(n19682), .A2(n19554), .B1(n19681), .B2(n19553), .ZN(
        n19550) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19555), .ZN(n19549) );
  OAI211_X1 U21808 ( .C1(n19687), .C2(n19558), .A(n19550), .B(n19549), .ZN(
        P3_U2886) );
  AOI22_X1 U21809 ( .A1(n19699), .A2(n19554), .B1(n19688), .B2(n19553), .ZN(
        n19552) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19555), .ZN(n19551) );
  OAI211_X1 U21811 ( .C1(n19695), .C2(n19558), .A(n19552), .B(n19551), .ZN(
        P3_U2878) );
  AOI22_X1 U21812 ( .A1(n19620), .A2(n19554), .B1(n19697), .B2(n19553), .ZN(
        n19557) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19555), .ZN(n19556) );
  OAI211_X1 U21814 ( .C1(n19602), .C2(n19558), .A(n19557), .B(n19556), .ZN(
        P3_U2870) );
  OAI22_X1 U21815 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19603), .ZN(n19559) );
  INV_X1 U21816 ( .A(n19559), .ZN(U252) );
  NAND2_X1 U21817 ( .A1(n19606), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19601) );
  NAND2_X1 U21818 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19606), .ZN(n19593) );
  INV_X1 U21819 ( .A(n19593), .ZN(n19597) );
  AND2_X1 U21820 ( .A1(n19607), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U21821 ( .A1(n19626), .A2(n19597), .B1(n19608), .B2(n19596), .ZN(
        n19562) );
  NOR2_X2 U21822 ( .A1(n19560), .A2(n19609), .ZN(n19598) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19598), .ZN(n19561) );
  OAI211_X1 U21824 ( .C1(n19706), .C2(n19601), .A(n19562), .B(n19561), .ZN(
        P3_U2989) );
  AOI22_X1 U21825 ( .A1(n19632), .A2(n19597), .B1(n19614), .B2(n19596), .ZN(
        n19564) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19598), .ZN(n19563) );
  OAI211_X1 U21827 ( .C1(n19618), .C2(n19601), .A(n19564), .B(n19563), .ZN(
        P3_U2981) );
  AOI22_X1 U21828 ( .A1(n19637), .A2(n19597), .B1(n19619), .B2(n19596), .ZN(
        n19566) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19598), .ZN(n19565) );
  OAI211_X1 U21830 ( .C1(n19624), .C2(n19601), .A(n19566), .B(n19565), .ZN(
        P3_U2973) );
  AOI22_X1 U21831 ( .A1(n19643), .A2(n19597), .B1(n19625), .B2(n19596), .ZN(
        n19568) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19598), .ZN(n19567) );
  OAI211_X1 U21833 ( .C1(n19630), .C2(n19601), .A(n19568), .B(n19567), .ZN(
        P3_U2965) );
  INV_X1 U21834 ( .A(n19601), .ZN(n19590) );
  AOI22_X1 U21835 ( .A1(n19643), .A2(n19590), .B1(n19631), .B2(n19596), .ZN(
        n19570) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19598), .ZN(n19569) );
  OAI211_X1 U21837 ( .C1(n19641), .C2(n19593), .A(n19570), .B(n19569), .ZN(
        P3_U2957) );
  AOI22_X1 U21838 ( .A1(n19648), .A2(n19590), .B1(n19636), .B2(n19596), .ZN(
        n19572) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19598), .ZN(n19571) );
  OAI211_X1 U21840 ( .C1(n19573), .C2(n19593), .A(n19572), .B(n19571), .ZN(
        P3_U2949) );
  AOI22_X1 U21841 ( .A1(n19654), .A2(n19590), .B1(n19642), .B2(n19596), .ZN(
        n19575) );
  AOI22_X1 U21842 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19598), .ZN(n19574) );
  OAI211_X1 U21843 ( .C1(n19652), .C2(n19593), .A(n19575), .B(n19574), .ZN(
        P3_U2941) );
  AOI22_X1 U21844 ( .A1(n19666), .A2(n19597), .B1(n19647), .B2(n19596), .ZN(
        n19577) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19598), .ZN(n19576) );
  OAI211_X1 U21846 ( .C1(n19652), .C2(n19601), .A(n19577), .B(n19576), .ZN(
        P3_U2933) );
  AOI22_X1 U21847 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19655), .B1(
        n19653), .B2(n19596), .ZN(n19579) );
  AOI22_X1 U21848 ( .A1(n19654), .A2(n19598), .B1(n19666), .B2(n19590), .ZN(
        n19578) );
  OAI211_X1 U21849 ( .C1(n19580), .C2(n19593), .A(n19579), .B(n19578), .ZN(
        P3_U2925) );
  AOI22_X1 U21850 ( .A1(n19671), .A2(n19590), .B1(n19659), .B2(n19596), .ZN(
        n19582) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19598), .ZN(n19581) );
  OAI211_X1 U21852 ( .C1(n19664), .C2(n19593), .A(n19582), .B(n19581), .ZN(
        P3_U2917) );
  AOI22_X1 U21853 ( .A1(n19683), .A2(n19597), .B1(n19665), .B2(n19596), .ZN(
        n19584) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19598), .ZN(n19583) );
  OAI211_X1 U21855 ( .C1(n19664), .C2(n19601), .A(n19584), .B(n19583), .ZN(
        P3_U2909) );
  AOI22_X1 U21856 ( .A1(n19690), .A2(n19597), .B1(n19670), .B2(n19596), .ZN(
        n19586) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19598), .ZN(n19585) );
  OAI211_X1 U21858 ( .C1(n19675), .C2(n19601), .A(n19586), .B(n19585), .ZN(
        P3_U2901) );
  AOI22_X1 U21859 ( .A1(n19701), .A2(n19597), .B1(n19676), .B2(n19596), .ZN(
        n19588) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19598), .ZN(n19587) );
  OAI211_X1 U21861 ( .C1(n19589), .C2(n19601), .A(n19588), .B(n19587), .ZN(
        P3_U2893) );
  AOI22_X1 U21862 ( .A1(n19701), .A2(n19590), .B1(n19681), .B2(n19596), .ZN(
        n19592) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19598), .ZN(n19591) );
  OAI211_X1 U21864 ( .C1(n19695), .C2(n19593), .A(n19592), .B(n19591), .ZN(
        P3_U2885) );
  AOI22_X1 U21865 ( .A1(n19699), .A2(n19597), .B1(n19688), .B2(n19596), .ZN(
        n19595) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19598), .ZN(n19594) );
  OAI211_X1 U21867 ( .C1(n19695), .C2(n19601), .A(n19595), .B(n19594), .ZN(
        P3_U2877) );
  AOI22_X1 U21868 ( .A1(n19620), .A2(n19597), .B1(n19697), .B2(n19596), .ZN(
        n19600) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19598), .ZN(n19599) );
  OAI211_X1 U21870 ( .C1(n19602), .C2(n19601), .A(n19600), .B(n19599), .ZN(
        P3_U2869) );
  OAI22_X1 U21871 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19603), .ZN(n19605) );
  INV_X1 U21872 ( .A(n19605), .ZN(U251) );
  NAND2_X1 U21873 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19606), .ZN(n19705) );
  NAND2_X1 U21874 ( .A1(n19606), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19694) );
  INV_X1 U21875 ( .A(n19694), .ZN(n19698) );
  AND2_X1 U21876 ( .A1(n19607), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19696) );
  AOI22_X1 U21877 ( .A1(n19620), .A2(n19698), .B1(n19608), .B2(n19696), .ZN(
        n19613) );
  NOR2_X2 U21878 ( .A1(n19610), .A2(n19609), .ZN(n19700) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19611), .B1(
        n19682), .B2(n19700), .ZN(n19612) );
  OAI211_X1 U21880 ( .C1(n19618), .C2(n19705), .A(n19613), .B(n19612), .ZN(
        P3_U2988) );
  INV_X1 U21881 ( .A(n19705), .ZN(n19689) );
  AOI22_X1 U21882 ( .A1(n19632), .A2(n19689), .B1(n19614), .B2(n19696), .ZN(
        n19617) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19615), .B1(
        n19699), .B2(n19700), .ZN(n19616) );
  OAI211_X1 U21884 ( .C1(n19618), .C2(n19694), .A(n19617), .B(n19616), .ZN(
        P3_U2980) );
  AOI22_X1 U21885 ( .A1(n19637), .A2(n19689), .B1(n19619), .B2(n19696), .ZN(
        n19623) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19621), .B1(
        n19620), .B2(n19700), .ZN(n19622) );
  OAI211_X1 U21887 ( .C1(n19624), .C2(n19694), .A(n19623), .B(n19622), .ZN(
        P3_U2972) );
  AOI22_X1 U21888 ( .A1(n19643), .A2(n19689), .B1(n19625), .B2(n19696), .ZN(
        n19629) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19627), .B1(
        n19626), .B2(n19700), .ZN(n19628) );
  OAI211_X1 U21890 ( .C1(n19630), .C2(n19694), .A(n19629), .B(n19628), .ZN(
        P3_U2964) );
  AOI22_X1 U21891 ( .A1(n19643), .A2(n19698), .B1(n19631), .B2(n19696), .ZN(
        n19635) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19633), .B1(
        n19632), .B2(n19700), .ZN(n19634) );
  OAI211_X1 U21893 ( .C1(n19641), .C2(n19705), .A(n19635), .B(n19634), .ZN(
        P3_U2956) );
  AOI22_X1 U21894 ( .A1(n19654), .A2(n19689), .B1(n19636), .B2(n19696), .ZN(
        n19640) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19638), .B1(
        n19637), .B2(n19700), .ZN(n19639) );
  OAI211_X1 U21896 ( .C1(n19641), .C2(n19694), .A(n19640), .B(n19639), .ZN(
        P3_U2948) );
  AOI22_X1 U21897 ( .A1(n19654), .A2(n19698), .B1(n19642), .B2(n19696), .ZN(
        n19646) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19700), .ZN(n19645) );
  OAI211_X1 U21899 ( .C1(n19652), .C2(n19705), .A(n19646), .B(n19645), .ZN(
        P3_U2940) );
  AOI22_X1 U21900 ( .A1(n19666), .A2(n19689), .B1(n19647), .B2(n19696), .ZN(
        n19651) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19649), .B1(
        n19648), .B2(n19700), .ZN(n19650) );
  OAI211_X1 U21902 ( .C1(n19652), .C2(n19694), .A(n19651), .B(n19650), .ZN(
        P3_U2932) );
  AOI22_X1 U21903 ( .A1(n19671), .A2(n19689), .B1(n19653), .B2(n19696), .ZN(
        n19657) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19700), .ZN(n19656) );
  OAI211_X1 U21905 ( .C1(n19658), .C2(n19694), .A(n19657), .B(n19656), .ZN(
        P3_U2924) );
  AOI22_X1 U21906 ( .A1(n19671), .A2(n19698), .B1(n19659), .B2(n19696), .ZN(
        n19663) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19700), .ZN(n19662) );
  OAI211_X1 U21908 ( .C1(n19664), .C2(n19705), .A(n19663), .B(n19662), .ZN(
        P3_U2916) );
  AOI22_X1 U21909 ( .A1(n19677), .A2(n19698), .B1(n19665), .B2(n19696), .ZN(
        n19669) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19700), .ZN(n19668) );
  OAI211_X1 U21911 ( .C1(n19675), .C2(n19705), .A(n19669), .B(n19668), .ZN(
        P3_U2908) );
  AOI22_X1 U21912 ( .A1(n19690), .A2(n19689), .B1(n19670), .B2(n19696), .ZN(
        n19674) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19672), .B1(
        n19671), .B2(n19700), .ZN(n19673) );
  OAI211_X1 U21914 ( .C1(n19675), .C2(n19694), .A(n19674), .B(n19673), .ZN(
        P3_U2900) );
  AOI22_X1 U21915 ( .A1(n19690), .A2(n19698), .B1(n19676), .B2(n19696), .ZN(
        n19680) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19700), .ZN(n19679) );
  OAI211_X1 U21917 ( .C1(n19687), .C2(n19705), .A(n19680), .B(n19679), .ZN(
        P3_U2892) );
  AOI22_X1 U21918 ( .A1(n19682), .A2(n19689), .B1(n19681), .B2(n19696), .ZN(
        n19686) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19700), .ZN(n19685) );
  OAI211_X1 U21920 ( .C1(n19687), .C2(n19694), .A(n19686), .B(n19685), .ZN(
        P3_U2884) );
  AOI22_X1 U21921 ( .A1(n19699), .A2(n19689), .B1(n19688), .B2(n19696), .ZN(
        n19693) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19691), .B1(
        n19690), .B2(n19700), .ZN(n19692) );
  OAI211_X1 U21923 ( .C1(n19695), .C2(n19694), .A(n19693), .B(n19692), .ZN(
        P3_U2876) );
  AOI22_X1 U21924 ( .A1(n19699), .A2(n19698), .B1(n19697), .B2(n19696), .ZN(
        n19704) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19702), .B1(
        n19701), .B2(n19700), .ZN(n19703) );
  OAI211_X1 U21926 ( .C1(n19706), .C2(n19705), .A(n19704), .B(n19703), .ZN(
        P3_U2868) );
  AOI22_X1 U21927 ( .A1(n20170), .A2(BUF2_REG_31__SCAN_IN), .B1(n20277), .B2(
        n19707), .ZN(n19709) );
  AOI22_X1 U21928 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20276), .B1(n20169), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19708) );
  NAND2_X1 U21929 ( .A1(n19709), .A2(n19708), .ZN(P2_U2888) );
  OAI222_X1 U21930 ( .A1(n19712), .A2(n20023), .B1(n19711), .B2(n20066), .C1(
        n19710), .C2(n20285), .ZN(P2_U2904) );
  OAI222_X1 U21931 ( .A1(n19715), .A2(n20023), .B1(n19714), .B2(n20066), .C1(
        n20285), .C2(n19713), .ZN(P2_U2905) );
  OAI222_X1 U21932 ( .A1(n19718), .A2(n20023), .B1(n19717), .B2(n20066), .C1(
        n20285), .C2(n19716), .ZN(P2_U2906) );
  OAI222_X1 U21933 ( .A1(n19721), .A2(n20023), .B1(n19720), .B2(n20066), .C1(
        n20285), .C2(n19719), .ZN(P2_U2907) );
  OAI222_X1 U21934 ( .A1(n19724), .A2(n20023), .B1(n19723), .B2(n20066), .C1(
        n20285), .C2(n19722), .ZN(P2_U2908) );
  AOI22_X1 U21935 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n20276), .B1(n19725), 
        .B2(n20011), .ZN(n19726) );
  OAI21_X1 U21936 ( .B1(n20023), .B2(n19727), .A(n19726), .ZN(P2_U2909) );
  OAI222_X1 U21937 ( .A1(n19730), .A2(n20023), .B1(n19729), .B2(n20066), .C1(
        n20285), .C2(n19728), .ZN(P2_U2910) );
  INV_X1 U21938 ( .A(n19731), .ZN(n19734) );
  OAI222_X1 U21939 ( .A1(n19734), .A2(n20023), .B1(n19733), .B2(n20066), .C1(
        n20285), .C2(n19732), .ZN(P2_U2911) );
  OAI222_X1 U21940 ( .A1(n19736), .A2(n20023), .B1(n19735), .B2(n20066), .C1(
        n20285), .C2(n19741), .ZN(P2_U2912) );
  AOI22_X2 U21941 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20292), .ZN(n19967) );
  NAND3_X1 U21942 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19755) );
  INV_X1 U21943 ( .A(n19746), .ZN(n19739) );
  INV_X1 U21944 ( .A(n19958), .ZN(n20290) );
  OAI21_X1 U21945 ( .B1(n19739), .B2(n20290), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19740) );
  OAI21_X1 U21946 ( .B1(n19755), .B2(n19953), .A(n19740), .ZN(n20291) );
  AOI22_X1 U21947 ( .A1(n20291), .A2(n19742), .B1(n20290), .B2(n11166), .ZN(
        n19754) );
  INV_X1 U21948 ( .A(n19776), .ZN(n19743) );
  NAND2_X1 U21949 ( .A1(n19743), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19770) );
  OAI21_X1 U21950 ( .B1(n19770), .B2(n19814), .A(n19755), .ZN(n19748) );
  NOR2_X1 U21951 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19744), .ZN(n19956) );
  INV_X1 U21952 ( .A(n19956), .ZN(n19942) );
  AOI21_X1 U21953 ( .B1(n19959), .B2(n20290), .A(n19955), .ZN(n19745) );
  OAI21_X1 U21954 ( .B1(n19746), .B2(n19942), .A(n19745), .ZN(n19747) );
  NAND2_X1 U21955 ( .A1(n19748), .A2(n19747), .ZN(n20294) );
  OAI22_X2 U21956 ( .A1(n20705), .A2(n19752), .B1(n19751), .B2(n19750), .ZN(
        n19952) );
  AOI22_X1 U21957 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n19952), .ZN(n19753) );
  OAI211_X1 U21958 ( .C1(n19967), .C2(n20399), .A(n19754), .B(n19753), .ZN(
        P2_U3175) );
  NOR2_X1 U21959 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19755), .ZN(
        n20297) );
  AOI22_X1 U21960 ( .A1(n19952), .A2(n20306), .B1(n11166), .B2(n20297), .ZN(
        n19767) );
  NAND2_X1 U21961 ( .A1(n20303), .A2(n20232), .ZN(n19756) );
  AOI21_X1 U21962 ( .B1(n19756), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19953), 
        .ZN(n19761) );
  NAND3_X1 U21963 ( .A1(n19910), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19782) );
  NOR2_X1 U21964 ( .A1(n19856), .A2(n19782), .ZN(n20304) );
  INV_X1 U21965 ( .A(n20304), .ZN(n19759) );
  NOR2_X1 U21966 ( .A1(n19762), .A2(n19942), .ZN(n19757) );
  NOR2_X1 U21967 ( .A1(n19955), .A2(n19757), .ZN(n19758) );
  AOI21_X1 U21968 ( .B1(n19761), .B2(n19759), .A(n19758), .ZN(n19760) );
  AOI21_X1 U21969 ( .B1(n20297), .B2(n19959), .A(n19760), .ZN(n20300) );
  OAI21_X1 U21970 ( .B1(n20297), .B2(n20304), .A(n19761), .ZN(n19765) );
  INV_X1 U21971 ( .A(n19762), .ZN(n19763) );
  OAI21_X1 U21972 ( .B1(n19763), .B2(n20297), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19764) );
  NAND2_X1 U21973 ( .A1(n19765), .A2(n19764), .ZN(n20299) );
  AOI22_X1 U21974 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20300), .B1(
        n19742), .B2(n20299), .ZN(n19766) );
  OAI211_X1 U21975 ( .C1(n19967), .C2(n20232), .A(n19767), .B(n19766), .ZN(
        P2_U3167) );
  INV_X1 U21976 ( .A(n19772), .ZN(n19768) );
  OAI21_X1 U21977 ( .B1(n19768), .B2(n20304), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19769) );
  OAI21_X1 U21978 ( .B1(n19782), .B2(n19953), .A(n19769), .ZN(n20305) );
  AOI22_X1 U21979 ( .A1(n20305), .A2(n19742), .B1(n20304), .B2(n11166), .ZN(
        n19778) );
  NAND2_X1 U21980 ( .A1(n19782), .A2(n19770), .ZN(n19774) );
  AOI21_X1 U21981 ( .B1(n19959), .B2(n20304), .A(n19955), .ZN(n19771) );
  OAI21_X1 U21982 ( .B1(n19772), .B2(n19942), .A(n19771), .ZN(n19773) );
  NAND2_X1 U21983 ( .A1(n19774), .A2(n19773), .ZN(n20307) );
  AOI22_X1 U21984 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20307), .B1(
        n20313), .B2(n19952), .ZN(n19777) );
  OAI211_X1 U21985 ( .C1(n19967), .C2(n20303), .A(n19778), .B(n19777), .ZN(
        P2_U3159) );
  INV_X1 U21986 ( .A(n19779), .ZN(n19780) );
  NAND2_X1 U21987 ( .A1(n19780), .A2(n19863), .ZN(n19889) );
  INV_X1 U21988 ( .A(n19781), .ZN(n19785) );
  NOR2_X1 U21989 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19782), .ZN(
        n20311) );
  OAI21_X1 U21990 ( .B1(n19783), .B2(n20311), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19784) );
  OAI21_X1 U21991 ( .B1(n19889), .B2(n19785), .A(n19784), .ZN(n20312) );
  AOI22_X1 U21992 ( .A1(n20312), .A2(n19742), .B1(n11166), .B2(n20311), .ZN(
        n19793) );
  INV_X1 U21993 ( .A(n20311), .ZN(n19786) );
  AOI21_X1 U21994 ( .B1(n19786), .B2(n19953), .A(n20286), .ZN(n19791) );
  NOR2_X1 U21995 ( .A1(n19787), .A2(n19942), .ZN(n19790) );
  NOR2_X2 U21996 ( .A1(n19821), .A2(n19884), .ZN(n20237) );
  OAI21_X1 U21997 ( .B1(n20237), .B2(n20313), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19788) );
  OAI21_X1 U21998 ( .B1(n19889), .B2(n19905), .A(n19788), .ZN(n19789) );
  AOI22_X1 U21999 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19952), .B2(n20237), .ZN(n19792) );
  OAI211_X1 U22000 ( .C1(n19967), .C2(n20310), .A(n19793), .B(n19792), .ZN(
        P2_U3151) );
  INV_X1 U22001 ( .A(n20237), .ZN(n20322) );
  NAND3_X1 U22002 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19906), .ZN(n19803) );
  INV_X1 U22003 ( .A(n19794), .ZN(n19795) );
  NOR2_X1 U22004 ( .A1(n19856), .A2(n19803), .ZN(n20317) );
  OAI21_X1 U22005 ( .B1(n19795), .B2(n20317), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19796) );
  OAI21_X1 U22006 ( .B1(n19803), .B2(n19953), .A(n19796), .ZN(n20318) );
  AOI22_X1 U22007 ( .A1(n20318), .A2(n19742), .B1(n11166), .B2(n20317), .ZN(
        n19802) );
  OAI21_X1 U22008 ( .B1(n20018), .B2(n19908), .A(n19803), .ZN(n19800) );
  AOI21_X1 U22009 ( .B1(n19959), .B2(n20317), .A(n19955), .ZN(n19797) );
  OAI21_X1 U22010 ( .B1(n19798), .B2(n19942), .A(n19797), .ZN(n19799) );
  NAND2_X1 U22011 ( .A1(n19800), .A2(n19799), .ZN(n20319) );
  AOI22_X1 U22012 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20319), .B1(
        n20324), .B2(n19952), .ZN(n19801) );
  OAI211_X1 U22013 ( .C1(n19967), .C2(n20322), .A(n19802), .B(n19801), .ZN(
        P2_U3143) );
  NOR2_X1 U22014 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19803), .ZN(
        n20323) );
  AOI22_X1 U22015 ( .A1(n19952), .A2(n20243), .B1(n11166), .B2(n20323), .ZN(
        n19813) );
  OAI21_X1 U22016 ( .B1(n20324), .B2(n20243), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19804) );
  NAND2_X1 U22017 ( .A1(n19804), .A2(n19939), .ZN(n19811) );
  NAND3_X1 U22018 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19910), .A3(
        n19906), .ZN(n19831) );
  NOR2_X1 U22019 ( .A1(n19856), .A2(n19831), .ZN(n20329) );
  NOR2_X1 U22020 ( .A1(n20329), .A2(n20323), .ZN(n19810) );
  INV_X1 U22021 ( .A(n19810), .ZN(n19807) );
  AOI21_X1 U22022 ( .B1(n19808), .B2(n19834), .A(n20323), .ZN(n19805) );
  NOR2_X1 U22023 ( .A1(n19805), .A2(n20286), .ZN(n19806) );
  OAI22_X1 U22024 ( .A1(n19811), .A2(n19807), .B1(n19955), .B2(n19806), .ZN(
        n20326) );
  OAI21_X1 U22025 ( .B1(n19808), .B2(n20323), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19809) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20326), .B1(
        n19742), .B2(n20325), .ZN(n19812) );
  OAI211_X1 U22027 ( .C1(n19967), .C2(n20240), .A(n19813), .B(n19812), .ZN(
        P2_U3135) );
  NAND2_X1 U22028 ( .A1(n19814), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19871) );
  INV_X1 U22029 ( .A(n19871), .ZN(n19815) );
  AND2_X1 U22030 ( .A1(n20015), .A2(n19815), .ZN(n19938) );
  NAND2_X1 U22031 ( .A1(n19909), .A2(n19938), .ZN(n19823) );
  INV_X1 U22032 ( .A(n19831), .ZN(n19822) );
  NAND2_X1 U22033 ( .A1(n19823), .A2(n19831), .ZN(n19820) );
  INV_X1 U22034 ( .A(n20329), .ZN(n19816) );
  NAND2_X1 U22035 ( .A1(n19953), .A2(n19816), .ZN(n19817) );
  NAND2_X1 U22036 ( .A1(n19959), .A2(n19817), .ZN(n19818) );
  OAI21_X1 U22037 ( .B1(n19942), .B2(n19824), .A(n19818), .ZN(n19819) );
  INV_X1 U22038 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U22039 ( .A1(n19952), .A2(n20336), .B1(n11166), .B2(n20329), .ZN(
        n19829) );
  NAND3_X1 U22040 ( .A1(n19823), .A2(n19939), .A3(n19822), .ZN(n19827) );
  INV_X1 U22041 ( .A(n19824), .ZN(n19825) );
  OAI21_X1 U22042 ( .B1(n19825), .B2(n20329), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19826) );
  NAND2_X1 U22043 ( .A1(n19827), .A2(n19826), .ZN(n20330) );
  INV_X1 U22044 ( .A(n19967), .ZN(n19895) );
  AOI22_X1 U22045 ( .A1(n19742), .A2(n20330), .B1(n20243), .B2(n19895), .ZN(
        n19828) );
  OAI211_X1 U22046 ( .C1(n19984), .C2(n19830), .A(n19829), .B(n19828), .ZN(
        P2_U3127) );
  NOR2_X1 U22047 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n20335) );
  AOI22_X1 U22048 ( .A1(n19952), .A2(n20246), .B1(n11166), .B2(n20335), .ZN(
        n19844) );
  AOI21_X1 U22049 ( .B1(n20346), .B2(n20249), .A(n22228), .ZN(n19832) );
  NOR2_X1 U22050 ( .A1(n19832), .A2(n19953), .ZN(n19839) );
  NAND2_X1 U22051 ( .A1(n19905), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19890) );
  INV_X1 U22052 ( .A(n19890), .ZN(n19873) );
  NAND2_X1 U22053 ( .A1(n19833), .A2(n19873), .ZN(n19838) );
  OAI21_X1 U22054 ( .B1(n19840), .B2(n19835), .A(n19834), .ZN(n19836) );
  AOI21_X1 U22055 ( .B1(n19839), .B2(n19838), .A(n19836), .ZN(n19837) );
  OAI21_X1 U22056 ( .B1(n20335), .B2(n19837), .A(n19959), .ZN(n20338) );
  INV_X1 U22057 ( .A(n19838), .ZN(n20341) );
  OAI21_X1 U22058 ( .B1(n20341), .B2(n20335), .A(n19839), .ZN(n19842) );
  OAI21_X1 U22059 ( .B1(n19840), .B2(n20335), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19841) );
  NAND2_X1 U22060 ( .A1(n19842), .A2(n19841), .ZN(n20337) );
  AOI22_X1 U22061 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n19742), .ZN(n19843) );
  OAI211_X1 U22062 ( .C1(n19967), .C2(n20249), .A(n19844), .B(n19843), .ZN(
        P2_U3119) );
  NAND2_X1 U22063 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19873), .ZN(
        n19852) );
  OAI21_X1 U22064 ( .B1(n19872), .B2(n19845), .A(n19852), .ZN(n19849) );
  AOI21_X1 U22065 ( .B1(n19850), .B2(n19956), .A(n20341), .ZN(n19847) );
  INV_X1 U22066 ( .A(n19955), .ZN(n19846) );
  OAI21_X1 U22067 ( .B1(n19847), .B2(n20286), .A(n19846), .ZN(n19848) );
  INV_X1 U22068 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U22069 ( .B1(n19850), .B2(n20341), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19851) );
  OAI21_X1 U22070 ( .B1(n19852), .B2(n19953), .A(n19851), .ZN(n20342) );
  AOI22_X1 U22071 ( .A1(n20342), .A2(n19742), .B1(n20341), .B2(n11166), .ZN(
        n19854) );
  AOI22_X1 U22072 ( .A1(n20246), .A2(n19895), .B1(n20350), .B2(n19952), .ZN(
        n19853) );
  OAI211_X1 U22073 ( .C1(n19989), .C2(n19855), .A(n19854), .B(n19853), .ZN(
        P2_U3111) );
  INV_X1 U22074 ( .A(n19923), .ZN(n19858) );
  NAND2_X1 U22075 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19856), .ZN(
        n19921) );
  NOR2_X1 U22076 ( .A1(n19921), .A2(n19890), .ZN(n20347) );
  OAI21_X1 U22077 ( .B1(n19860), .B2(n20347), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19857) );
  OAI21_X1 U22078 ( .B1(n19890), .B2(n19858), .A(n19857), .ZN(n20348) );
  AOI22_X1 U22079 ( .A1(n20348), .A2(n19742), .B1(n11166), .B2(n20347), .ZN(
        n19868) );
  INV_X1 U22080 ( .A(n20347), .ZN(n19859) );
  AOI21_X1 U22081 ( .B1(n19859), .B2(n19953), .A(n20286), .ZN(n19866) );
  INV_X1 U22082 ( .A(n19860), .ZN(n19861) );
  NOR2_X1 U22083 ( .A1(n19861), .A2(n19942), .ZN(n19865) );
  OAI21_X1 U22084 ( .B1(n20355), .B2(n20350), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19862) );
  OAI21_X1 U22085 ( .B1(n19863), .B2(n19890), .A(n19862), .ZN(n19864) );
  AOI22_X1 U22086 ( .A1(n19952), .A2(n20355), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n20349), .ZN(n19867) );
  OAI211_X1 U22087 ( .C1(n19967), .C2(n20200), .A(n19868), .B(n19867), .ZN(
        P2_U3103) );
  INV_X1 U22088 ( .A(n19872), .ZN(n19870) );
  INV_X1 U22089 ( .A(n19946), .ZN(n19869) );
  NAND2_X1 U22090 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19910), .ZN(
        n19936) );
  NOR2_X1 U22091 ( .A1(n19936), .A2(n19890), .ZN(n20354) );
  AOI22_X1 U22092 ( .A1(n20362), .A2(n19952), .B1(n11166), .B2(n20354), .ZN(
        n19882) );
  OAI21_X1 U22093 ( .B1(n19872), .B2(n19871), .A(n19939), .ZN(n19880) );
  NAND2_X1 U22094 ( .A1(n19910), .A2(n19873), .ZN(n19879) );
  INV_X1 U22095 ( .A(n19879), .ZN(n19876) );
  OAI21_X1 U22096 ( .B1(n19939), .B2(n20354), .A(n19959), .ZN(n19874) );
  OAI21_X1 U22097 ( .B1(n11190), .B2(n19942), .A(n19874), .ZN(n19875) );
  OAI21_X1 U22098 ( .B1(n19880), .B2(n19876), .A(n19875), .ZN(n20357) );
  OAI21_X1 U22099 ( .B1(n11191), .B2(n20354), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19878) );
  OAI21_X1 U22100 ( .B1(n19880), .B2(n19879), .A(n19878), .ZN(n20356) );
  AOI22_X1 U22101 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20357), .B1(
        n19742), .B2(n20356), .ZN(n19881) );
  OAI211_X1 U22102 ( .C1(n19967), .C2(n20353), .A(n19882), .B(n19881), .ZN(
        P2_U3095) );
  INV_X1 U22103 ( .A(n19947), .ZN(n19886) );
  INV_X1 U22104 ( .A(n19884), .ZN(n19885) );
  NAND2_X1 U22105 ( .A1(n20368), .A2(n20360), .ZN(n19887) );
  NAND2_X1 U22106 ( .A1(n19887), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19888) );
  NAND2_X1 U22107 ( .A1(n19888), .A2(n19939), .ZN(n19900) );
  NOR2_X1 U22108 ( .A1(n19889), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19896) );
  NOR3_X2 U22109 ( .A1(n19890), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20361) );
  OAI21_X1 U22110 ( .B1(n19939), .B2(n20361), .A(n19959), .ZN(n19891) );
  OAI21_X1 U22111 ( .B1(n19942), .B2(n19892), .A(n19891), .ZN(n19893) );
  INV_X1 U22112 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U22113 ( .A1(n19895), .A2(n20362), .B1(n11166), .B2(n20361), .ZN(
        n19902) );
  INV_X1 U22114 ( .A(n19896), .ZN(n19899) );
  OAI21_X1 U22115 ( .B1(n19897), .B2(n20361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19898) );
  AOI22_X1 U22116 ( .A1(n19742), .A2(n20364), .B1(n20370), .B2(n19952), .ZN(
        n19901) );
  OAI211_X1 U22117 ( .C1(n20363), .C2(n19903), .A(n19902), .B(n19901), .ZN(
        P2_U3087) );
  NAND2_X1 U22118 ( .A1(n19906), .A2(n19905), .ZN(n19935) );
  NOR2_X1 U22119 ( .A1(n19907), .A2(n19935), .ZN(n20369) );
  AOI22_X1 U22120 ( .A1(n19952), .A2(n20378), .B1(n20369), .B2(n11166), .ZN(
        n19920) );
  OAI21_X1 U22121 ( .B1(n19909), .B2(n19908), .A(n19939), .ZN(n19918) );
  NOR2_X1 U22122 ( .A1(n19910), .A2(n19935), .ZN(n19914) );
  INV_X1 U22123 ( .A(n19915), .ZN(n19912) );
  OAI21_X1 U22124 ( .B1(n19939), .B2(n20369), .A(n19959), .ZN(n19911) );
  OAI21_X1 U22125 ( .B1(n19912), .B2(n19942), .A(n19911), .ZN(n19913) );
  OAI21_X1 U22126 ( .B1(n19918), .B2(n19914), .A(n19913), .ZN(n20372) );
  INV_X1 U22127 ( .A(n19914), .ZN(n19917) );
  OAI21_X1 U22128 ( .B1(n19915), .B2(n20369), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19916) );
  OAI21_X1 U22129 ( .B1(n19918), .B2(n19917), .A(n19916), .ZN(n20371) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20372), .B1(
        n19742), .B2(n20371), .ZN(n19919) );
  OAI211_X1 U22131 ( .C1(n19967), .C2(n20368), .A(n19920), .B(n19919), .ZN(
        P2_U3079) );
  NOR2_X1 U22132 ( .A1(n19921), .A2(n19935), .ZN(n20376) );
  OAI21_X1 U22133 ( .B1(n19927), .B2(n20376), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19924) );
  INV_X1 U22134 ( .A(n19935), .ZN(n19922) );
  NAND2_X1 U22135 ( .A1(n19923), .A2(n19922), .ZN(n19926) );
  NAND2_X1 U22136 ( .A1(n19924), .A2(n19926), .ZN(n20377) );
  AOI22_X1 U22137 ( .A1(n20377), .A2(n19742), .B1(n11166), .B2(n20376), .ZN(
        n19934) );
  OAI221_X1 U22138 ( .B1(n22228), .B2(n20388), .C1(n22228), .C2(n20375), .A(
        n19926), .ZN(n19931) );
  INV_X1 U22139 ( .A(n19927), .ZN(n19929) );
  INV_X1 U22140 ( .A(n20376), .ZN(n19928) );
  OAI21_X1 U22141 ( .B1(n19929), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19928), 
        .ZN(n19930) );
  MUX2_X1 U22142 ( .A(n19931), .B(n19930), .S(n19953), .Z(n19932) );
  NAND2_X1 U22143 ( .A1(n19932), .A2(n19959), .ZN(n20379) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n19952), .ZN(n19933) );
  OAI211_X1 U22145 ( .C1(n19967), .C2(n20375), .A(n19934), .B(n19933), .ZN(
        P2_U3071) );
  NOR2_X1 U22146 ( .A1(n19935), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19944) );
  INV_X1 U22147 ( .A(n19944), .ZN(n19950) );
  NOR2_X1 U22148 ( .A1(n19936), .A2(n19935), .ZN(n20382) );
  OAI21_X1 U22149 ( .B1(n12825), .B2(n20382), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19937) );
  OAI21_X1 U22150 ( .B1(n19950), .B2(n19953), .A(n19937), .ZN(n20383) );
  AOI22_X1 U22151 ( .A1(n20383), .A2(n19742), .B1(n11166), .B2(n20382), .ZN(
        n19949) );
  AND2_X1 U22152 ( .A1(n20018), .A2(n19938), .ZN(n19945) );
  OAI21_X1 U22153 ( .B1(n19939), .B2(n20382), .A(n19959), .ZN(n19940) );
  OAI21_X1 U22154 ( .B1(n19942), .B2(n19941), .A(n19940), .ZN(n19943) );
  OAI21_X1 U22155 ( .B1(n19945), .B2(n19944), .A(n19943), .ZN(n20385) );
  NOR2_X2 U22156 ( .A1(n19947), .A2(n19946), .ZN(n20392) );
  AOI22_X1 U22157 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n19952), .ZN(n19948) );
  OAI211_X1 U22158 ( .C1(n19967), .C2(n20388), .A(n19949), .B(n19948), .ZN(
        P2_U3063) );
  INV_X1 U22159 ( .A(n20399), .ZN(n20268) );
  NOR2_X1 U22160 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19950), .ZN(
        n20391) );
  AOI22_X1 U22161 ( .A1(n19952), .A2(n20268), .B1(n11166), .B2(n20391), .ZN(
        n19966) );
  AOI21_X1 U22162 ( .B1(n20273), .B2(n20399), .A(n22228), .ZN(n19954) );
  NOR2_X1 U22163 ( .A1(n19954), .A2(n19953), .ZN(n19961) );
  AOI21_X1 U22164 ( .B1(n19956), .B2(n19962), .A(n19955), .ZN(n19957) );
  AOI21_X1 U22165 ( .B1(n19961), .B2(n19958), .A(n19957), .ZN(n19960) );
  OAI21_X1 U22166 ( .B1(n20391), .B2(n19960), .A(n19959), .ZN(n20396) );
  OAI21_X1 U22167 ( .B1(n20290), .B2(n20391), .A(n19961), .ZN(n19964) );
  OAI21_X1 U22168 ( .B1(n19962), .B2(n20391), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19963) );
  NAND2_X1 U22169 ( .A1(n19964), .A2(n19963), .ZN(n20395) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20396), .B1(
        n19742), .B2(n20395), .ZN(n19965) );
  OAI211_X1 U22171 ( .C1(n19967), .C2(n20273), .A(n19966), .B(n19965), .ZN(
        P2_U3055) );
  OAI222_X1 U22172 ( .A1(n19969), .A2(n20023), .B1(n19968), .B2(n20066), .C1(
        n20285), .C2(n19970), .ZN(P2_U2913) );
  AOI22_X1 U22173 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20292), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20293), .ZN(n20010) );
  NOR2_X2 U22174 ( .A1(n13736), .A2(n20288), .ZN(n20006) );
  AOI22_X1 U22175 ( .A1(n20291), .A2(n19971), .B1(n20290), .B2(n20006), .ZN(
        n19973) );
  AOI22_X1 U22176 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20292), .ZN(n20005) );
  INV_X1 U22177 ( .A(n20005), .ZN(n20007) );
  AOI22_X1 U22178 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20294), .B1(
        n20268), .B2(n20007), .ZN(n19972) );
  OAI211_X1 U22179 ( .C1(n20010), .C2(n20232), .A(n19973), .B(n19972), .ZN(
        P2_U3174) );
  AOI22_X1 U22180 ( .A1(n20007), .A2(n20298), .B1(n20006), .B2(n20297), .ZN(
        n19975) );
  AOI22_X1 U22181 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20300), .B1(
        n19971), .B2(n20299), .ZN(n19974) );
  OAI211_X1 U22182 ( .C1(n20010), .C2(n20303), .A(n19975), .B(n19974), .ZN(
        P2_U3166) );
  AOI22_X1 U22183 ( .A1(n20305), .A2(n19971), .B1(n20304), .B2(n20006), .ZN(
        n19977) );
  AOI22_X1 U22184 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20307), .B1(
        n20306), .B2(n20007), .ZN(n19976) );
  OAI211_X1 U22185 ( .C1(n20010), .C2(n20310), .A(n19977), .B(n19976), .ZN(
        P2_U3158) );
  AOI22_X1 U22186 ( .A1(n20312), .A2(n19971), .B1(n20006), .B2(n20311), .ZN(
        n19979) );
  INV_X1 U22187 ( .A(n20010), .ZN(n20002) );
  AOI22_X1 U22188 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20237), .B2(n20002), .ZN(n19978) );
  OAI211_X1 U22189 ( .C1(n20005), .C2(n20310), .A(n19979), .B(n19978), .ZN(
        P2_U3150) );
  AOI22_X1 U22190 ( .A1(n20318), .A2(n19971), .B1(n20006), .B2(n20317), .ZN(
        n19981) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20319), .B1(
        n20237), .B2(n20007), .ZN(n19980) );
  OAI211_X1 U22192 ( .C1(n20010), .C2(n20240), .A(n19981), .B(n19980), .ZN(
        P2_U3142) );
  AOI22_X1 U22193 ( .A1(n20002), .A2(n20243), .B1(n20006), .B2(n20323), .ZN(
        n19983) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20326), .B1(
        n19971), .B2(n20325), .ZN(n19982) );
  OAI211_X1 U22195 ( .C1(n20005), .C2(n20240), .A(n19983), .B(n19982), .ZN(
        P2_U3134) );
  AOI22_X1 U22196 ( .A1(n20002), .A2(n20336), .B1(n20006), .B2(n20329), .ZN(
        n19986) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20331), .B1(
        n19971), .B2(n20330), .ZN(n19985) );
  OAI211_X1 U22198 ( .C1(n20005), .C2(n20334), .A(n19986), .B(n19985), .ZN(
        P2_U3126) );
  AOI22_X1 U22199 ( .A1(n20007), .A2(n20336), .B1(n20006), .B2(n20335), .ZN(
        n19988) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n19971), .ZN(n19987) );
  OAI211_X1 U22201 ( .C1(n20010), .C2(n20346), .A(n19988), .B(n19987), .ZN(
        P2_U3118) );
  AOI22_X1 U22202 ( .A1(n20342), .A2(n19971), .B1(n20341), .B2(n20006), .ZN(
        n19991) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20343), .B1(
        n20246), .B2(n20007), .ZN(n19990) );
  OAI211_X1 U22204 ( .C1(n20010), .C2(n20200), .A(n19991), .B(n19990), .ZN(
        P2_U3110) );
  AOI22_X1 U22205 ( .A1(n20348), .A2(n19971), .B1(n20006), .B2(n20347), .ZN(
        n19993) );
  AOI22_X1 U22206 ( .A1(n20002), .A2(n20355), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n20349), .ZN(n19992) );
  OAI211_X1 U22207 ( .C1(n20005), .C2(n20200), .A(n19993), .B(n19992), .ZN(
        P2_U3102) );
  AOI22_X1 U22208 ( .A1(n20007), .A2(n20355), .B1(n20006), .B2(n20354), .ZN(
        n19995) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20357), .B1(
        n19971), .B2(n20356), .ZN(n19994) );
  OAI211_X1 U22210 ( .C1(n20010), .C2(n20360), .A(n19995), .B(n19994), .ZN(
        P2_U3094) );
  AOI22_X1 U22211 ( .A1(n20007), .A2(n20362), .B1(n20006), .B2(n20361), .ZN(
        n19997) );
  AOI22_X1 U22212 ( .A1(n19971), .A2(n20364), .B1(n20370), .B2(n20002), .ZN(
        n19996) );
  OAI211_X1 U22213 ( .C1(n20363), .C2(n12856), .A(n19997), .B(n19996), .ZN(
        P2_U3086) );
  AOI22_X1 U22214 ( .A1(n20002), .A2(n20378), .B1(n20369), .B2(n20006), .ZN(
        n19999) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20372), .B1(
        n19971), .B2(n20371), .ZN(n19998) );
  OAI211_X1 U22216 ( .C1(n20005), .C2(n20368), .A(n19999), .B(n19998), .ZN(
        P2_U3078) );
  AOI22_X1 U22217 ( .A1(n20377), .A2(n19971), .B1(n20006), .B2(n20376), .ZN(
        n20001) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20002), .ZN(n20000) );
  OAI211_X1 U22219 ( .C1(n20005), .C2(n20375), .A(n20001), .B(n20000), .ZN(
        P2_U3070) );
  AOI22_X1 U22220 ( .A1(n20383), .A2(n19971), .B1(n20006), .B2(n20382), .ZN(
        n20004) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20002), .ZN(n20003) );
  OAI211_X1 U22222 ( .C1(n20005), .C2(n20388), .A(n20004), .B(n20003), .ZN(
        P2_U3062) );
  AOI22_X1 U22223 ( .A1(n20007), .A2(n20392), .B1(n20006), .B2(n20391), .ZN(
        n20009) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n19971), .ZN(n20008) );
  OAI211_X1 U22225 ( .C1(n20010), .C2(n20399), .A(n20009), .B(n20008), .ZN(
        P2_U3054) );
  AOI22_X1 U22226 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20276), .B1(n20024), .B2(
        n20011), .ZN(n20021) );
  NAND2_X1 U22227 ( .A1(n20013), .A2(n20012), .ZN(n20014) );
  OAI21_X1 U22228 ( .B1(n20016), .B2(n20015), .A(n20014), .ZN(n20122) );
  XNOR2_X1 U22229 ( .A(n20018), .B(n20017), .ZN(n20123) );
  NOR2_X1 U22230 ( .A1(n20122), .A2(n20123), .ZN(n20121) );
  AOI21_X1 U22231 ( .B1(n20018), .B2(n20017), .A(n20121), .ZN(n20019) );
  NOR2_X1 U22232 ( .A1(n20019), .A2(n20074), .ZN(n20075) );
  OR3_X1 U22233 ( .A1(n20075), .A2(n20076), .A3(n20222), .ZN(n20020) );
  OAI211_X1 U22234 ( .C1(n20023), .C2(n20022), .A(n20021), .B(n20020), .ZN(
        P2_U2914) );
  AOI22_X1 U22235 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20292), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20293), .ZN(n20064) );
  INV_X1 U22236 ( .A(n20024), .ZN(n20025) );
  NOR2_X2 U22237 ( .A1(n20025), .A2(n20286), .ZN(n20061) );
  AOI22_X1 U22238 ( .A1(n20291), .A2(n20061), .B1(n20290), .B2(n20027), .ZN(
        n20029) );
  AOI22_X1 U22239 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20292), .ZN(n20059) );
  INV_X1 U22240 ( .A(n20059), .ZN(n20060) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20294), .B1(
        n20268), .B2(n20060), .ZN(n20028) );
  OAI211_X1 U22242 ( .C1(n20064), .C2(n20232), .A(n20029), .B(n20028), .ZN(
        P2_U3173) );
  AOI22_X1 U22243 ( .A1(n20056), .A2(n20306), .B1(n20027), .B2(n20297), .ZN(
        n20031) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20300), .B1(
        n20061), .B2(n20299), .ZN(n20030) );
  OAI211_X1 U22245 ( .C1(n20059), .C2(n20232), .A(n20031), .B(n20030), .ZN(
        P2_U3165) );
  AOI22_X1 U22246 ( .A1(n20305), .A2(n20061), .B1(n20304), .B2(n20027), .ZN(
        n20033) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20307), .B1(
        n20313), .B2(n20056), .ZN(n20032) );
  OAI211_X1 U22248 ( .C1(n20059), .C2(n20303), .A(n20033), .B(n20032), .ZN(
        P2_U3157) );
  AOI22_X1 U22249 ( .A1(n20312), .A2(n20061), .B1(n20027), .B2(n20311), .ZN(
        n20035) );
  AOI22_X1 U22250 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20237), .B2(n20056), .ZN(n20034) );
  OAI211_X1 U22251 ( .C1(n20059), .C2(n20310), .A(n20035), .B(n20034), .ZN(
        P2_U3149) );
  AOI22_X1 U22252 ( .A1(n20318), .A2(n20061), .B1(n20027), .B2(n20317), .ZN(
        n20037) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20319), .B1(
        n20237), .B2(n20060), .ZN(n20036) );
  OAI211_X1 U22254 ( .C1(n20064), .C2(n20240), .A(n20037), .B(n20036), .ZN(
        P2_U3141) );
  AOI22_X1 U22255 ( .A1(n20056), .A2(n20243), .B1(n20027), .B2(n20323), .ZN(
        n20039) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20326), .B1(
        n20061), .B2(n20325), .ZN(n20038) );
  OAI211_X1 U22257 ( .C1(n20059), .C2(n20240), .A(n20039), .B(n20038), .ZN(
        P2_U3133) );
  AOI22_X1 U22258 ( .A1(n20060), .A2(n20243), .B1(n20027), .B2(n20329), .ZN(
        n20041) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20331), .B1(
        n20061), .B2(n20330), .ZN(n20040) );
  OAI211_X1 U22260 ( .C1(n20064), .C2(n20249), .A(n20041), .B(n20040), .ZN(
        P2_U3125) );
  AOI22_X1 U22261 ( .A1(n20060), .A2(n20336), .B1(n20027), .B2(n20335), .ZN(
        n20043) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20061), .ZN(n20042) );
  OAI211_X1 U22263 ( .C1(n20064), .C2(n20346), .A(n20043), .B(n20042), .ZN(
        P2_U3117) );
  AOI22_X1 U22264 ( .A1(n20342), .A2(n20061), .B1(n20341), .B2(n20027), .ZN(
        n20045) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20343), .B1(
        n20350), .B2(n20056), .ZN(n20044) );
  OAI211_X1 U22266 ( .C1(n20059), .C2(n20346), .A(n20045), .B(n20044), .ZN(
        P2_U3109) );
  AOI22_X1 U22267 ( .A1(n20348), .A2(n20061), .B1(n20027), .B2(n20347), .ZN(
        n20047) );
  AOI22_X1 U22268 ( .A1(n20060), .A2(n20350), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n20349), .ZN(n20046) );
  OAI211_X1 U22269 ( .C1(n20064), .C2(n20353), .A(n20047), .B(n20046), .ZN(
        P2_U3101) );
  AOI22_X1 U22270 ( .A1(n20056), .A2(n20362), .B1(n20027), .B2(n20354), .ZN(
        n20049) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20357), .B1(
        n20061), .B2(n20356), .ZN(n20048) );
  OAI211_X1 U22272 ( .C1(n20059), .C2(n20353), .A(n20049), .B(n20048), .ZN(
        P2_U3093) );
  AOI22_X1 U22273 ( .A1(n20060), .A2(n20362), .B1(n20027), .B2(n20361), .ZN(
        n20051) );
  AOI22_X1 U22274 ( .A1(n20061), .A2(n20364), .B1(n20370), .B2(n20056), .ZN(
        n20050) );
  OAI211_X1 U22275 ( .C1(n20363), .C2(n13719), .A(n20051), .B(n20050), .ZN(
        P2_U3085) );
  AOI22_X1 U22276 ( .A1(n20056), .A2(n20378), .B1(n20369), .B2(n20027), .ZN(
        n20053) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20372), .B1(
        n20061), .B2(n20371), .ZN(n20052) );
  OAI211_X1 U22278 ( .C1(n20059), .C2(n20368), .A(n20053), .B(n20052), .ZN(
        P2_U3077) );
  AOI22_X1 U22279 ( .A1(n20377), .A2(n20061), .B1(n20027), .B2(n20376), .ZN(
        n20055) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20056), .ZN(n20054) );
  OAI211_X1 U22281 ( .C1(n20059), .C2(n20375), .A(n20055), .B(n20054), .ZN(
        P2_U3069) );
  AOI22_X1 U22282 ( .A1(n20383), .A2(n20061), .B1(n20027), .B2(n20382), .ZN(
        n20058) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20056), .ZN(n20057) );
  OAI211_X1 U22284 ( .C1(n20059), .C2(n20388), .A(n20058), .B(n20057), .ZN(
        P2_U3061) );
  AOI22_X1 U22285 ( .A1(n20060), .A2(n20392), .B1(n20027), .B2(n20391), .ZN(
        n20063) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20061), .ZN(n20062) );
  OAI211_X1 U22287 ( .C1(n20064), .C2(n20399), .A(n20063), .B(n20062), .ZN(
        P2_U3053) );
  OAI22_X1 U22288 ( .A1(n20067), .A2(n20080), .B1(n20066), .B2(n20065), .ZN(
        n20068) );
  INV_X1 U22289 ( .A(n20068), .ZN(n20073) );
  AOI22_X1 U22290 ( .A1(n20170), .A2(BUF2_REG_20__SCAN_IN), .B1(n20169), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n20072) );
  AOI22_X1 U22291 ( .A1(n20070), .A2(n20279), .B1(n20277), .B2(n20069), .ZN(
        n20071) );
  NAND3_X1 U22292 ( .A1(n20073), .A2(n20072), .A3(n20071), .ZN(P2_U2899) );
  AOI22_X1 U22293 ( .A1(n20277), .A2(n20074), .B1(n20276), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n20079) );
  XOR2_X1 U22294 ( .A(n20076), .B(n20075), .Z(n20077) );
  NAND2_X1 U22295 ( .A1(n20077), .A2(n20279), .ZN(n20078) );
  OAI211_X1 U22296 ( .C1(n20080), .C2(n20285), .A(n20079), .B(n20078), .ZN(
        P2_U2915) );
  AOI22_X1 U22297 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20292), .ZN(n20119) );
  NOR2_X2 U22298 ( .A1(n20080), .A2(n20286), .ZN(n20116) );
  NOR2_X2 U22299 ( .A1(n20081), .A2(n20288), .ZN(n20114) );
  AOI22_X1 U22300 ( .A1(n20291), .A2(n20116), .B1(n20290), .B2(n20114), .ZN(
        n20083) );
  AOI22_X1 U22301 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20292), .ZN(n20109) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n20115), .ZN(n20082) );
  OAI211_X1 U22303 ( .C1(n20119), .C2(n20399), .A(n20083), .B(n20082), .ZN(
        P2_U3172) );
  INV_X1 U22304 ( .A(n20119), .ZN(n20106) );
  AOI22_X1 U22305 ( .A1(n20106), .A2(n20298), .B1(n20114), .B2(n20297), .ZN(
        n20085) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20300), .B1(
        n20116), .B2(n20299), .ZN(n20084) );
  OAI211_X1 U22307 ( .C1(n20109), .C2(n20303), .A(n20085), .B(n20084), .ZN(
        P2_U3164) );
  AOI22_X1 U22308 ( .A1(n20305), .A2(n20116), .B1(n20304), .B2(n20114), .ZN(
        n20087) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20307), .B1(
        n20306), .B2(n20106), .ZN(n20086) );
  OAI211_X1 U22310 ( .C1(n20109), .C2(n20310), .A(n20087), .B(n20086), .ZN(
        P2_U3156) );
  AOI22_X1 U22311 ( .A1(n20312), .A2(n20116), .B1(n20114), .B2(n20311), .ZN(
        n20089) );
  AOI22_X1 U22312 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20237), .B2(n20115), .ZN(n20088) );
  OAI211_X1 U22313 ( .C1(n20119), .C2(n20310), .A(n20089), .B(n20088), .ZN(
        P2_U3148) );
  AOI22_X1 U22314 ( .A1(n20318), .A2(n20116), .B1(n20114), .B2(n20317), .ZN(
        n20091) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20319), .B1(
        n20237), .B2(n20106), .ZN(n20090) );
  OAI211_X1 U22316 ( .C1(n20109), .C2(n20240), .A(n20091), .B(n20090), .ZN(
        P2_U3140) );
  AOI22_X1 U22317 ( .A1(n20106), .A2(n20324), .B1(n20114), .B2(n20323), .ZN(
        n20093) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20326), .B1(
        n20116), .B2(n20325), .ZN(n20092) );
  OAI211_X1 U22319 ( .C1(n20109), .C2(n20334), .A(n20093), .B(n20092), .ZN(
        P2_U3132) );
  AOI22_X1 U22320 ( .A1(n20115), .A2(n20336), .B1(n20114), .B2(n20329), .ZN(
        n20095) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20331), .B1(
        n20116), .B2(n20330), .ZN(n20094) );
  OAI211_X1 U22322 ( .C1(n20119), .C2(n20334), .A(n20095), .B(n20094), .ZN(
        P2_U3124) );
  AOI22_X1 U22323 ( .A1(n20115), .A2(n20246), .B1(n20114), .B2(n20335), .ZN(
        n20097) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20116), .ZN(n20096) );
  OAI211_X1 U22325 ( .C1(n20119), .C2(n20249), .A(n20097), .B(n20096), .ZN(
        P2_U3116) );
  AOI22_X1 U22326 ( .A1(n20342), .A2(n20116), .B1(n20341), .B2(n20114), .ZN(
        n20099) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20343), .B1(
        n20350), .B2(n20115), .ZN(n20098) );
  OAI211_X1 U22328 ( .C1(n20119), .C2(n20346), .A(n20099), .B(n20098), .ZN(
        P2_U3108) );
  AOI22_X1 U22329 ( .A1(n20348), .A2(n20116), .B1(n20114), .B2(n20347), .ZN(
        n20101) );
  AOI22_X1 U22330 ( .A1(n20115), .A2(n20355), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n20349), .ZN(n20100) );
  OAI211_X1 U22331 ( .C1(n20119), .C2(n20200), .A(n20101), .B(n20100), .ZN(
        P2_U3100) );
  AOI22_X1 U22332 ( .A1(n20106), .A2(n20355), .B1(n20114), .B2(n20354), .ZN(
        n20103) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20357), .B1(
        n20116), .B2(n20356), .ZN(n20102) );
  OAI211_X1 U22334 ( .C1(n20109), .C2(n20360), .A(n20103), .B(n20102), .ZN(
        P2_U3092) );
  AOI22_X1 U22335 ( .A1(n20106), .A2(n20362), .B1(n20114), .B2(n20361), .ZN(
        n20105) );
  AOI22_X1 U22336 ( .A1(n20116), .A2(n20364), .B1(n20370), .B2(n20115), .ZN(
        n20104) );
  OAI211_X1 U22337 ( .C1(n20363), .C2(n13688), .A(n20105), .B(n20104), .ZN(
        P2_U3084) );
  AOI22_X1 U22338 ( .A1(n20106), .A2(n20370), .B1(n20369), .B2(n20114), .ZN(
        n20108) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20372), .B1(
        n20116), .B2(n20371), .ZN(n20107) );
  OAI211_X1 U22340 ( .C1(n20109), .C2(n20375), .A(n20108), .B(n20107), .ZN(
        P2_U3076) );
  AOI22_X1 U22341 ( .A1(n20377), .A2(n20116), .B1(n20114), .B2(n20376), .ZN(
        n20111) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20115), .ZN(n20110) );
  OAI211_X1 U22343 ( .C1(n20119), .C2(n20375), .A(n20111), .B(n20110), .ZN(
        P2_U3068) );
  AOI22_X1 U22344 ( .A1(n20383), .A2(n20116), .B1(n20114), .B2(n20382), .ZN(
        n20113) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20115), .ZN(n20112) );
  OAI211_X1 U22346 ( .C1(n20119), .C2(n20388), .A(n20113), .B(n20112), .ZN(
        P2_U3060) );
  AOI22_X1 U22347 ( .A1(n20115), .A2(n20268), .B1(n20391), .B2(n20114), .ZN(
        n20118) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20116), .ZN(n20117) );
  OAI211_X1 U22349 ( .C1(n20119), .C2(n20273), .A(n20118), .B(n20117), .ZN(
        P2_U3052) );
  AOI22_X1 U22350 ( .A1(n20120), .A2(n20277), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20276), .ZN(n20126) );
  AOI21_X1 U22351 ( .B1(n20123), .B2(n20122), .A(n20121), .ZN(n20124) );
  OR2_X1 U22352 ( .A1(n20124), .A2(n20222), .ZN(n20125) );
  OAI211_X1 U22353 ( .C1(n20127), .C2(n20285), .A(n20126), .B(n20125), .ZN(
        P2_U2916) );
  AOI22_X1 U22354 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20292), .ZN(n20158) );
  NOR2_X2 U22355 ( .A1(n20127), .A2(n20286), .ZN(n20163) );
  NOR2_X2 U22356 ( .A1(n12531), .A2(n20288), .ZN(n20161) );
  AOI22_X1 U22357 ( .A1(n20291), .A2(n20163), .B1(n20290), .B2(n20161), .ZN(
        n20129) );
  AOI22_X1 U22358 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20292), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20293), .ZN(n20166) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n20155), .ZN(n20128) );
  OAI211_X1 U22360 ( .C1(n20158), .C2(n20399), .A(n20129), .B(n20128), .ZN(
        P2_U3171) );
  AOI22_X1 U22361 ( .A1(n20155), .A2(n20306), .B1(n20161), .B2(n20297), .ZN(
        n20131) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20300), .B1(
        n20163), .B2(n20299), .ZN(n20130) );
  OAI211_X1 U22363 ( .C1(n20158), .C2(n20232), .A(n20131), .B(n20130), .ZN(
        P2_U3163) );
  AOI22_X1 U22364 ( .A1(n20305), .A2(n20163), .B1(n20304), .B2(n20161), .ZN(
        n20133) );
  INV_X1 U22365 ( .A(n20158), .ZN(n20162) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20307), .B1(
        n20306), .B2(n20162), .ZN(n20132) );
  OAI211_X1 U22367 ( .C1(n20166), .C2(n20310), .A(n20133), .B(n20132), .ZN(
        P2_U3155) );
  AOI22_X1 U22368 ( .A1(n20312), .A2(n20163), .B1(n20161), .B2(n20311), .ZN(
        n20135) );
  AOI22_X1 U22369 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20237), .B2(n20155), .ZN(n20134) );
  OAI211_X1 U22370 ( .C1(n20158), .C2(n20310), .A(n20135), .B(n20134), .ZN(
        P2_U3147) );
  AOI22_X1 U22371 ( .A1(n20318), .A2(n20163), .B1(n20161), .B2(n20317), .ZN(
        n20137) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20319), .B1(
        n20324), .B2(n20155), .ZN(n20136) );
  OAI211_X1 U22373 ( .C1(n20158), .C2(n20322), .A(n20137), .B(n20136), .ZN(
        P2_U3139) );
  AOI22_X1 U22374 ( .A1(n20162), .A2(n20324), .B1(n20161), .B2(n20323), .ZN(
        n20139) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20326), .B1(
        n20163), .B2(n20325), .ZN(n20138) );
  OAI211_X1 U22376 ( .C1(n20166), .C2(n20334), .A(n20139), .B(n20138), .ZN(
        P2_U3131) );
  AOI22_X1 U22377 ( .A1(n20155), .A2(n20336), .B1(n20161), .B2(n20329), .ZN(
        n20141) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20331), .B1(
        n20163), .B2(n20330), .ZN(n20140) );
  OAI211_X1 U22379 ( .C1(n20158), .C2(n20334), .A(n20141), .B(n20140), .ZN(
        P2_U3123) );
  AOI22_X1 U22380 ( .A1(n20155), .A2(n20246), .B1(n20161), .B2(n20335), .ZN(
        n20143) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20163), .ZN(n20142) );
  OAI211_X1 U22382 ( .C1(n20158), .C2(n20249), .A(n20143), .B(n20142), .ZN(
        P2_U3115) );
  AOI22_X1 U22383 ( .A1(n20342), .A2(n20163), .B1(n20341), .B2(n20161), .ZN(
        n20145) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20343), .B1(
        n20246), .B2(n20162), .ZN(n20144) );
  OAI211_X1 U22385 ( .C1(n20166), .C2(n20200), .A(n20145), .B(n20144), .ZN(
        P2_U3107) );
  AOI22_X1 U22386 ( .A1(n20348), .A2(n20163), .B1(n20161), .B2(n20347), .ZN(
        n20147) );
  AOI22_X1 U22387 ( .A1(n20155), .A2(n20355), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n20349), .ZN(n20146) );
  OAI211_X1 U22388 ( .C1(n20158), .C2(n20200), .A(n20147), .B(n20146), .ZN(
        P2_U3099) );
  AOI22_X1 U22389 ( .A1(n20155), .A2(n20362), .B1(n20161), .B2(n20354), .ZN(
        n20149) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20357), .B1(
        n20163), .B2(n20356), .ZN(n20148) );
  OAI211_X1 U22391 ( .C1(n20158), .C2(n20353), .A(n20149), .B(n20148), .ZN(
        P2_U3091) );
  AOI22_X1 U22392 ( .A1(n20162), .A2(n20362), .B1(n20161), .B2(n20361), .ZN(
        n20151) );
  AOI22_X1 U22393 ( .A1(n20163), .A2(n20364), .B1(n20370), .B2(n20155), .ZN(
        n20150) );
  OAI211_X1 U22394 ( .C1(n20363), .C2(n20152), .A(n20151), .B(n20150), .ZN(
        P2_U3083) );
  AOI22_X1 U22395 ( .A1(n20155), .A2(n20378), .B1(n20369), .B2(n20161), .ZN(
        n20154) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20372), .B1(
        n20163), .B2(n20371), .ZN(n20153) );
  OAI211_X1 U22397 ( .C1(n20158), .C2(n20368), .A(n20154), .B(n20153), .ZN(
        P2_U3075) );
  AOI22_X1 U22398 ( .A1(n20377), .A2(n20163), .B1(n20161), .B2(n20376), .ZN(
        n20157) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20155), .ZN(n20156) );
  OAI211_X1 U22400 ( .C1(n20158), .C2(n20375), .A(n20157), .B(n20156), .ZN(
        P2_U3067) );
  AOI22_X1 U22401 ( .A1(n20383), .A2(n20163), .B1(n20161), .B2(n20382), .ZN(
        n20160) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20385), .B1(
        n20262), .B2(n20162), .ZN(n20159) );
  OAI211_X1 U22403 ( .C1(n20166), .C2(n20273), .A(n20160), .B(n20159), .ZN(
        P2_U3059) );
  AOI22_X1 U22404 ( .A1(n20162), .A2(n20392), .B1(n20161), .B2(n20391), .ZN(
        n20165) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20163), .ZN(n20164) );
  OAI211_X1 U22406 ( .C1(n20166), .C2(n20399), .A(n20165), .B(n20164), .ZN(
        P2_U3051) );
  AOI22_X1 U22407 ( .A1(n20168), .A2(n20167), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n20276), .ZN(n20177) );
  AOI22_X1 U22408 ( .A1(n20170), .A2(BUF2_REG_18__SCAN_IN), .B1(n20169), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n20176) );
  OAI22_X1 U22409 ( .A1(n20173), .A2(n20222), .B1(n20172), .B2(n20171), .ZN(
        n20174) );
  INV_X1 U22410 ( .A(n20174), .ZN(n20175) );
  NAND3_X1 U22411 ( .A1(n20177), .A2(n20176), .A3(n20175), .ZN(P2_U2901) );
  AOI22_X1 U22412 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20292), .ZN(n20212) );
  NOR2_X2 U22413 ( .A1(n20178), .A2(n20286), .ZN(n20215) );
  NOR2_X2 U22414 ( .A1(n20179), .A2(n20288), .ZN(n20213) );
  AOI22_X1 U22415 ( .A1(n20291), .A2(n20215), .B1(n20290), .B2(n20213), .ZN(
        n20181) );
  AOI22_X1 U22416 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20292), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20293), .ZN(n20218) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n20209), .ZN(n20180) );
  OAI211_X1 U22418 ( .C1(n20212), .C2(n20399), .A(n20181), .B(n20180), .ZN(
        P2_U3170) );
  INV_X1 U22419 ( .A(n20212), .ZN(n20214) );
  AOI22_X1 U22420 ( .A1(n20214), .A2(n20298), .B1(n20213), .B2(n20297), .ZN(
        n20183) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20300), .B1(
        n20215), .B2(n20299), .ZN(n20182) );
  OAI211_X1 U22422 ( .C1(n20218), .C2(n20303), .A(n20183), .B(n20182), .ZN(
        P2_U3162) );
  AOI22_X1 U22423 ( .A1(n20305), .A2(n20215), .B1(n20304), .B2(n20213), .ZN(
        n20185) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20307), .B1(
        n20313), .B2(n20209), .ZN(n20184) );
  OAI211_X1 U22425 ( .C1(n20212), .C2(n20303), .A(n20185), .B(n20184), .ZN(
        P2_U3154) );
  AOI22_X1 U22426 ( .A1(n20312), .A2(n20215), .B1(n20213), .B2(n20311), .ZN(
        n20187) );
  AOI22_X1 U22427 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20237), .B2(n20209), .ZN(n20186) );
  OAI211_X1 U22428 ( .C1(n20212), .C2(n20310), .A(n20187), .B(n20186), .ZN(
        P2_U3146) );
  AOI22_X1 U22429 ( .A1(n20318), .A2(n20215), .B1(n20213), .B2(n20317), .ZN(
        n20189) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20319), .B1(
        n20237), .B2(n20214), .ZN(n20188) );
  OAI211_X1 U22431 ( .C1(n20218), .C2(n20240), .A(n20189), .B(n20188), .ZN(
        P2_U3138) );
  AOI22_X1 U22432 ( .A1(n20214), .A2(n20324), .B1(n20213), .B2(n20323), .ZN(
        n20191) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20326), .B1(
        n20215), .B2(n20325), .ZN(n20190) );
  OAI211_X1 U22434 ( .C1(n20218), .C2(n20334), .A(n20191), .B(n20190), .ZN(
        P2_U3130) );
  AOI22_X1 U22435 ( .A1(n20214), .A2(n20243), .B1(n20213), .B2(n20329), .ZN(
        n20193) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20331), .B1(
        n20215), .B2(n20330), .ZN(n20192) );
  OAI211_X1 U22437 ( .C1(n20218), .C2(n20249), .A(n20193), .B(n20192), .ZN(
        P2_U3122) );
  AOI22_X1 U22438 ( .A1(n20209), .A2(n20246), .B1(n20213), .B2(n20335), .ZN(
        n20195) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20215), .ZN(n20194) );
  OAI211_X1 U22440 ( .C1(n20212), .C2(n20249), .A(n20195), .B(n20194), .ZN(
        P2_U3114) );
  AOI22_X1 U22441 ( .A1(n20342), .A2(n20215), .B1(n20341), .B2(n20213), .ZN(
        n20197) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20343), .B1(
        n20246), .B2(n20214), .ZN(n20196) );
  OAI211_X1 U22443 ( .C1(n20218), .C2(n20200), .A(n20197), .B(n20196), .ZN(
        P2_U3106) );
  AOI22_X1 U22444 ( .A1(n20348), .A2(n20215), .B1(n20213), .B2(n20347), .ZN(
        n20199) );
  AOI22_X1 U22445 ( .A1(n20209), .A2(n20355), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n20349), .ZN(n20198) );
  OAI211_X1 U22446 ( .C1(n20212), .C2(n20200), .A(n20199), .B(n20198), .ZN(
        P2_U3098) );
  AOI22_X1 U22447 ( .A1(n20214), .A2(n20355), .B1(n20213), .B2(n20354), .ZN(
        n20202) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20357), .B1(
        n20215), .B2(n20356), .ZN(n20201) );
  OAI211_X1 U22449 ( .C1(n20218), .C2(n20360), .A(n20202), .B(n20201), .ZN(
        P2_U3090) );
  AOI22_X1 U22450 ( .A1(n20214), .A2(n20362), .B1(n20213), .B2(n20361), .ZN(
        n20204) );
  AOI22_X1 U22451 ( .A1(n20215), .A2(n20364), .B1(n20370), .B2(n20209), .ZN(
        n20203) );
  OAI211_X1 U22452 ( .C1(n20363), .C2(n13655), .A(n20204), .B(n20203), .ZN(
        P2_U3082) );
  AOI22_X1 U22453 ( .A1(n20209), .A2(n20378), .B1(n20369), .B2(n20213), .ZN(
        n20206) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20372), .B1(
        n20215), .B2(n20371), .ZN(n20205) );
  OAI211_X1 U22455 ( .C1(n20212), .C2(n20368), .A(n20206), .B(n20205), .ZN(
        P2_U3074) );
  AOI22_X1 U22456 ( .A1(n20377), .A2(n20215), .B1(n20213), .B2(n20376), .ZN(
        n20208) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20209), .ZN(n20207) );
  OAI211_X1 U22458 ( .C1(n20212), .C2(n20375), .A(n20208), .B(n20207), .ZN(
        P2_U3066) );
  AOI22_X1 U22459 ( .A1(n20383), .A2(n20215), .B1(n20213), .B2(n20382), .ZN(
        n20211) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20209), .ZN(n20210) );
  OAI211_X1 U22461 ( .C1(n20212), .C2(n20388), .A(n20211), .B(n20210), .ZN(
        P2_U3058) );
  AOI22_X1 U22462 ( .A1(n20214), .A2(n20392), .B1(n20213), .B2(n20391), .ZN(
        n20217) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20215), .ZN(n20216) );
  OAI211_X1 U22464 ( .C1(n20218), .C2(n20399), .A(n20217), .B(n20216), .ZN(
        P2_U3050) );
  AOI22_X1 U22465 ( .A1(n20277), .A2(n20219), .B1(n20276), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n20225) );
  AOI21_X1 U22466 ( .B1(n20278), .B2(n20221), .A(n20220), .ZN(n20223) );
  OR2_X1 U22467 ( .A1(n20223), .A2(n20222), .ZN(n20224) );
  OAI211_X1 U22468 ( .C1(n20226), .C2(n20285), .A(n20225), .B(n20224), .ZN(
        P2_U2918) );
  AOI22_X1 U22469 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20292), .ZN(n20274) );
  NOR2_X2 U22470 ( .A1(n20226), .A2(n20286), .ZN(n20270) );
  NOR2_X2 U22471 ( .A1(n20227), .A2(n20288), .ZN(n20267) );
  AOI22_X1 U22472 ( .A1(n20291), .A2(n20270), .B1(n20290), .B2(n20267), .ZN(
        n20229) );
  AOI22_X1 U22473 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20292), .ZN(n20261) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n20269), .ZN(n20228) );
  OAI211_X1 U22475 ( .C1(n20274), .C2(n20399), .A(n20229), .B(n20228), .ZN(
        P2_U3169) );
  AOI22_X1 U22476 ( .A1(n20269), .A2(n20306), .B1(n20267), .B2(n20297), .ZN(
        n20231) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20300), .B1(
        n20270), .B2(n20299), .ZN(n20230) );
  OAI211_X1 U22478 ( .C1(n20274), .C2(n20232), .A(n20231), .B(n20230), .ZN(
        P2_U3161) );
  AOI22_X1 U22479 ( .A1(n20305), .A2(n20270), .B1(n20304), .B2(n20267), .ZN(
        n20234) );
  INV_X1 U22480 ( .A(n20274), .ZN(n20258) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20307), .B1(
        n20306), .B2(n20258), .ZN(n20233) );
  OAI211_X1 U22482 ( .C1(n20261), .C2(n20310), .A(n20234), .B(n20233), .ZN(
        P2_U3153) );
  AOI22_X1 U22483 ( .A1(n20312), .A2(n20270), .B1(n20267), .B2(n20311), .ZN(
        n20236) );
  AOI22_X1 U22484 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20237), .B2(n20269), .ZN(n20235) );
  OAI211_X1 U22485 ( .C1(n20274), .C2(n20310), .A(n20236), .B(n20235), .ZN(
        P2_U3145) );
  AOI22_X1 U22486 ( .A1(n20318), .A2(n20270), .B1(n20267), .B2(n20317), .ZN(
        n20239) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20319), .B1(
        n20237), .B2(n20258), .ZN(n20238) );
  OAI211_X1 U22488 ( .C1(n20261), .C2(n20240), .A(n20239), .B(n20238), .ZN(
        P2_U3137) );
  AOI22_X1 U22489 ( .A1(n20258), .A2(n20324), .B1(n20267), .B2(n20323), .ZN(
        n20242) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20326), .B1(
        n20270), .B2(n20325), .ZN(n20241) );
  OAI211_X1 U22491 ( .C1(n20261), .C2(n20334), .A(n20242), .B(n20241), .ZN(
        P2_U3129) );
  AOI22_X1 U22492 ( .A1(n20258), .A2(n20243), .B1(n20267), .B2(n20329), .ZN(
        n20245) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20331), .B1(
        n20270), .B2(n20330), .ZN(n20244) );
  OAI211_X1 U22494 ( .C1(n20261), .C2(n20249), .A(n20245), .B(n20244), .ZN(
        P2_U3121) );
  AOI22_X1 U22495 ( .A1(n20269), .A2(n20246), .B1(n20267), .B2(n20335), .ZN(
        n20248) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20270), .ZN(n20247) );
  OAI211_X1 U22497 ( .C1(n20274), .C2(n20249), .A(n20248), .B(n20247), .ZN(
        P2_U3113) );
  AOI22_X1 U22498 ( .A1(n20342), .A2(n20270), .B1(n20341), .B2(n20267), .ZN(
        n20251) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20343), .B1(
        n20350), .B2(n20269), .ZN(n20250) );
  OAI211_X1 U22500 ( .C1(n20274), .C2(n20346), .A(n20251), .B(n20250), .ZN(
        P2_U3105) );
  AOI22_X1 U22501 ( .A1(n20348), .A2(n20270), .B1(n20267), .B2(n20347), .ZN(
        n20253) );
  AOI22_X1 U22502 ( .A1(n20258), .A2(n20350), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n20349), .ZN(n20252) );
  OAI211_X1 U22503 ( .C1(n20261), .C2(n20353), .A(n20253), .B(n20252), .ZN(
        P2_U3097) );
  AOI22_X1 U22504 ( .A1(n20258), .A2(n20355), .B1(n20267), .B2(n20354), .ZN(
        n20255) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20357), .B1(
        n20270), .B2(n20356), .ZN(n20254) );
  OAI211_X1 U22506 ( .C1(n20261), .C2(n20360), .A(n20255), .B(n20254), .ZN(
        P2_U3089) );
  AOI22_X1 U22507 ( .A1(n20258), .A2(n20362), .B1(n20267), .B2(n20361), .ZN(
        n20257) );
  AOI22_X1 U22508 ( .A1(n20270), .A2(n20364), .B1(n20370), .B2(n20269), .ZN(
        n20256) );
  OAI211_X1 U22509 ( .C1(n20363), .C2(n12687), .A(n20257), .B(n20256), .ZN(
        P2_U3081) );
  AOI22_X1 U22510 ( .A1(n20258), .A2(n20370), .B1(n20369), .B2(n20267), .ZN(
        n20260) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20372), .B1(
        n20270), .B2(n20371), .ZN(n20259) );
  OAI211_X1 U22512 ( .C1(n20261), .C2(n20375), .A(n20260), .B(n20259), .ZN(
        P2_U3073) );
  AOI22_X1 U22513 ( .A1(n20377), .A2(n20270), .B1(n20267), .B2(n20376), .ZN(
        n20264) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20379), .B1(
        n20262), .B2(n20269), .ZN(n20263) );
  OAI211_X1 U22515 ( .C1(n20274), .C2(n20375), .A(n20264), .B(n20263), .ZN(
        P2_U3065) );
  AOI22_X1 U22516 ( .A1(n20383), .A2(n20270), .B1(n20267), .B2(n20382), .ZN(
        n20266) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20269), .ZN(n20265) );
  OAI211_X1 U22518 ( .C1(n20274), .C2(n20388), .A(n20266), .B(n20265), .ZN(
        P2_U3057) );
  AOI22_X1 U22519 ( .A1(n20269), .A2(n20268), .B1(n20391), .B2(n20267), .ZN(
        n20272) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20270), .ZN(n20271) );
  OAI211_X1 U22521 ( .C1(n20274), .C2(n20273), .A(n20272), .B(n20271), .ZN(
        P2_U3049) );
  INV_X1 U22522 ( .A(n20275), .ZN(n20281) );
  AOI22_X1 U22523 ( .A1(n20277), .A2(n20281), .B1(n20276), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n20284) );
  INV_X1 U22524 ( .A(n20278), .ZN(n20280) );
  OAI211_X1 U22525 ( .C1(n20282), .C2(n20281), .A(n20280), .B(n20279), .ZN(
        n20283) );
  OAI211_X1 U22526 ( .C1(n20287), .C2(n20285), .A(n20284), .B(n20283), .ZN(
        P2_U2919) );
  AOI22_X1 U22527 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20292), .ZN(n20389) );
  NOR2_X2 U22528 ( .A1(n20287), .A2(n20286), .ZN(n20394) );
  NOR2_X2 U22529 ( .A1(n20289), .A2(n20288), .ZN(n20390) );
  AOI22_X1 U22530 ( .A1(n20291), .A2(n20394), .B1(n20290), .B2(n20390), .ZN(
        n20296) );
  AOI22_X2 U22531 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20293), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20292), .ZN(n20400) );
  INV_X1 U22532 ( .A(n20400), .ZN(n20384) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20294), .B1(
        n20298), .B2(n20384), .ZN(n20295) );
  OAI211_X1 U22534 ( .C1(n20389), .C2(n20399), .A(n20296), .B(n20295), .ZN(
        P2_U3168) );
  AOI22_X1 U22535 ( .A1(n20393), .A2(n20298), .B1(n20390), .B2(n20297), .ZN(
        n20302) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20300), .B1(
        n20394), .B2(n20299), .ZN(n20301) );
  OAI211_X1 U22537 ( .C1(n20400), .C2(n20303), .A(n20302), .B(n20301), .ZN(
        P2_U3160) );
  AOI22_X1 U22538 ( .A1(n20305), .A2(n20394), .B1(n20304), .B2(n20390), .ZN(
        n20309) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20307), .B1(
        n20306), .B2(n20393), .ZN(n20308) );
  OAI211_X1 U22540 ( .C1(n20400), .C2(n20310), .A(n20309), .B(n20308), .ZN(
        P2_U3152) );
  AOI22_X1 U22541 ( .A1(n20312), .A2(n20394), .B1(n20390), .B2(n20311), .ZN(
        n20316) );
  AOI22_X1 U22542 ( .A1(n20314), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20393), .B2(n20313), .ZN(n20315) );
  OAI211_X1 U22543 ( .C1(n20400), .C2(n20322), .A(n20316), .B(n20315), .ZN(
        P2_U3144) );
  AOI22_X1 U22544 ( .A1(n20318), .A2(n20394), .B1(n20390), .B2(n20317), .ZN(
        n20321) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20319), .B1(
        n20324), .B2(n20384), .ZN(n20320) );
  OAI211_X1 U22546 ( .C1(n20389), .C2(n20322), .A(n20321), .B(n20320), .ZN(
        P2_U3136) );
  AOI22_X1 U22547 ( .A1(n20393), .A2(n20324), .B1(n20390), .B2(n20323), .ZN(
        n20328) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20326), .B1(
        n20394), .B2(n20325), .ZN(n20327) );
  OAI211_X1 U22549 ( .C1(n20400), .C2(n20334), .A(n20328), .B(n20327), .ZN(
        P2_U3128) );
  AOI22_X1 U22550 ( .A1(n20384), .A2(n20336), .B1(n20390), .B2(n20329), .ZN(
        n20333) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20331), .B1(
        n20394), .B2(n20330), .ZN(n20332) );
  OAI211_X1 U22552 ( .C1(n20389), .C2(n20334), .A(n20333), .B(n20332), .ZN(
        P2_U3120) );
  AOI22_X1 U22553 ( .A1(n20393), .A2(n20336), .B1(n20390), .B2(n20335), .ZN(
        n20340) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20338), .B1(
        n20337), .B2(n20394), .ZN(n20339) );
  OAI211_X1 U22555 ( .C1(n20400), .C2(n20346), .A(n20340), .B(n20339), .ZN(
        P2_U3112) );
  AOI22_X1 U22556 ( .A1(n20342), .A2(n20394), .B1(n20341), .B2(n20390), .ZN(
        n20345) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20343), .B1(
        n20350), .B2(n20384), .ZN(n20344) );
  OAI211_X1 U22558 ( .C1(n20389), .C2(n20346), .A(n20345), .B(n20344), .ZN(
        P2_U3104) );
  AOI22_X1 U22559 ( .A1(n20348), .A2(n20394), .B1(n20390), .B2(n20347), .ZN(
        n20352) );
  AOI22_X1 U22560 ( .A1(n20393), .A2(n20350), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n20349), .ZN(n20351) );
  OAI211_X1 U22561 ( .C1(n20400), .C2(n20353), .A(n20352), .B(n20351), .ZN(
        P2_U3096) );
  AOI22_X1 U22562 ( .A1(n20393), .A2(n20355), .B1(n20390), .B2(n20354), .ZN(
        n20359) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20357), .B1(
        n20394), .B2(n20356), .ZN(n20358) );
  OAI211_X1 U22564 ( .C1(n20400), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        P2_U3088) );
  AOI22_X1 U22565 ( .A1(n20393), .A2(n20362), .B1(n20390), .B2(n20361), .ZN(
        n20367) );
  INV_X1 U22566 ( .A(n20363), .ZN(n20365) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20365), .B1(
        n20394), .B2(n20364), .ZN(n20366) );
  OAI211_X1 U22568 ( .C1(n20400), .C2(n20368), .A(n20367), .B(n20366), .ZN(
        P2_U3080) );
  AOI22_X1 U22569 ( .A1(n20393), .A2(n20370), .B1(n20369), .B2(n20390), .ZN(
        n20374) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20372), .B1(
        n20394), .B2(n20371), .ZN(n20373) );
  OAI211_X1 U22571 ( .C1(n20400), .C2(n20375), .A(n20374), .B(n20373), .ZN(
        P2_U3072) );
  AOI22_X1 U22572 ( .A1(n20377), .A2(n20394), .B1(n20390), .B2(n20376), .ZN(
        n20381) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20379), .B1(
        n20378), .B2(n20393), .ZN(n20380) );
  OAI211_X1 U22574 ( .C1(n20400), .C2(n20388), .A(n20381), .B(n20380), .ZN(
        P2_U3064) );
  AOI22_X1 U22575 ( .A1(n20383), .A2(n20394), .B1(n20390), .B2(n20382), .ZN(
        n20387) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20385), .B1(
        n20392), .B2(n20384), .ZN(n20386) );
  OAI211_X1 U22577 ( .C1(n20389), .C2(n20388), .A(n20387), .B(n20386), .ZN(
        P2_U3056) );
  AOI22_X1 U22578 ( .A1(n20393), .A2(n20392), .B1(n20391), .B2(n20390), .ZN(
        n20398) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20394), .ZN(n20397) );
  OAI211_X1 U22580 ( .C1(n20400), .C2(n20399), .A(n20398), .B(n20397), .ZN(
        P2_U3048) );
  INV_X1 U22581 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20704) );
  INV_X1 U22582 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20401) );
  AOI222_X1 U22583 ( .A1(n20704), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20707), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20401), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20402) );
  OAI22_X1 U22584 ( .A1(n20449), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20402), .ZN(n20403) );
  INV_X1 U22585 ( .A(n20403), .ZN(U376) );
  OAI22_X1 U22586 ( .A1(n20449), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20402), .ZN(n20404) );
  INV_X1 U22587 ( .A(n20404), .ZN(U365) );
  OAI22_X1 U22588 ( .A1(n20449), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20402), .ZN(n20405) );
  INV_X1 U22589 ( .A(n20405), .ZN(U354) );
  OAI22_X1 U22590 ( .A1(n20449), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20402), .ZN(n20406) );
  INV_X1 U22591 ( .A(n20406), .ZN(U353) );
  OAI22_X1 U22592 ( .A1(n20449), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20452), .ZN(n20407) );
  INV_X1 U22593 ( .A(n20407), .ZN(U352) );
  OAI22_X1 U22594 ( .A1(n20449), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n20452), .ZN(n20408) );
  INV_X1 U22595 ( .A(n20408), .ZN(U351) );
  INV_X2 U22596 ( .A(n20449), .ZN(n20452) );
  OAI22_X1 U22597 ( .A1(n20449), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20452), .ZN(n20409) );
  INV_X1 U22598 ( .A(n20409), .ZN(U350) );
  OAI22_X1 U22599 ( .A1(n20449), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n20452), .ZN(n20410) );
  INV_X1 U22600 ( .A(n20410), .ZN(U349) );
  OAI22_X1 U22601 ( .A1(n20449), .A2(P3_ADDRESS_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_8__SCAN_IN), .B2(n20452), .ZN(n20411) );
  INV_X1 U22602 ( .A(n20411), .ZN(U348) );
  OAI22_X1 U22603 ( .A1(n20449), .A2(P3_ADDRESS_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n20452), .ZN(n20412) );
  INV_X1 U22604 ( .A(n20412), .ZN(U347) );
  AOI22_X1 U22605 ( .A1(n20452), .A2(n20414), .B1(n20413), .B2(n20449), .ZN(
        U375) );
  AOI22_X1 U22606 ( .A1(n20452), .A2(n20416), .B1(n20415), .B2(n20449), .ZN(
        U374) );
  AOI22_X1 U22607 ( .A1(n20452), .A2(n20418), .B1(n20417), .B2(n20449), .ZN(
        U373) );
  AOI22_X1 U22608 ( .A1(n20452), .A2(n20420), .B1(n20419), .B2(n20449), .ZN(
        U372) );
  AOI22_X1 U22609 ( .A1(n20452), .A2(n20422), .B1(n20421), .B2(n20449), .ZN(
        U371) );
  AOI22_X1 U22610 ( .A1(n20452), .A2(n20424), .B1(n20423), .B2(n20449), .ZN(
        U370) );
  AOI22_X1 U22611 ( .A1(n20452), .A2(n20426), .B1(n20425), .B2(n20449), .ZN(
        U369) );
  AOI22_X1 U22612 ( .A1(n20452), .A2(n20428), .B1(n20427), .B2(n20449), .ZN(
        U368) );
  AOI22_X1 U22613 ( .A1(n20452), .A2(n20430), .B1(n20429), .B2(n20449), .ZN(
        U367) );
  AOI22_X1 U22614 ( .A1(n20452), .A2(n20432), .B1(n20431), .B2(n20449), .ZN(
        U366) );
  AOI22_X1 U22615 ( .A1(n20452), .A2(n20434), .B1(n20433), .B2(n20449), .ZN(
        U364) );
  OAI22_X1 U22616 ( .A1(n20449), .A2(P3_ADDRESS_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n20452), .ZN(n20435) );
  INV_X1 U22617 ( .A(n20435), .ZN(U363) );
  OAI22_X1 U22618 ( .A1(n20449), .A2(P3_ADDRESS_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n20452), .ZN(n20436) );
  INV_X1 U22619 ( .A(n20436), .ZN(U362) );
  AOI22_X1 U22620 ( .A1(n20452), .A2(n20438), .B1(n20437), .B2(n20449), .ZN(
        U361) );
  AOI22_X1 U22621 ( .A1(n20452), .A2(n20440), .B1(n20439), .B2(n20449), .ZN(
        U360) );
  AOI22_X1 U22622 ( .A1(n20452), .A2(n20442), .B1(n20441), .B2(n20449), .ZN(
        U359) );
  AOI22_X1 U22623 ( .A1(n20452), .A2(n20444), .B1(n20443), .B2(n20449), .ZN(
        U358) );
  AOI22_X1 U22624 ( .A1(n20452), .A2(n20446), .B1(n20445), .B2(n20449), .ZN(
        U357) );
  AOI22_X1 U22625 ( .A1(n20452), .A2(n20448), .B1(n20447), .B2(n20449), .ZN(
        U356) );
  AOI22_X1 U22626 ( .A1(n20452), .A2(n20451), .B1(n20450), .B2(n20449), .ZN(
        U355) );
  AOI22_X1 U22627 ( .A1(n21905), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20454) );
  OAI21_X1 U22628 ( .B1(n22304), .B2(n20473), .A(n20454), .ZN(P1_U2936) );
  AOI22_X1 U22629 ( .A1(n20464), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20455) );
  OAI21_X1 U22630 ( .B1(n12070), .B2(n20473), .A(n20455), .ZN(P1_U2935) );
  AOI22_X1 U22631 ( .A1(n20464), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20456) );
  OAI21_X1 U22632 ( .B1(n12060), .B2(n20473), .A(n20456), .ZN(P1_U2934) );
  AOI22_X1 U22633 ( .A1(n20464), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20457) );
  OAI21_X1 U22634 ( .B1(n12090), .B2(n20473), .A(n20457), .ZN(P1_U2933) );
  AOI22_X1 U22635 ( .A1(n20464), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20458) );
  OAI21_X1 U22636 ( .B1(n22324), .B2(n20473), .A(n20458), .ZN(P1_U2932) );
  AOI22_X1 U22637 ( .A1(n20464), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20459) );
  OAI21_X1 U22638 ( .B1(n14869), .B2(n20473), .A(n20459), .ZN(P1_U2931) );
  AOI22_X1 U22639 ( .A1(n20464), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20460) );
  OAI21_X1 U22640 ( .B1(n12122), .B2(n20473), .A(n20460), .ZN(P1_U2930) );
  AOI22_X1 U22641 ( .A1(n20464), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20461) );
  OAI21_X1 U22642 ( .B1(n12052), .B2(n20473), .A(n20461), .ZN(P1_U2929) );
  INV_X1 U22643 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n22346) );
  AOI22_X1 U22644 ( .A1(n20464), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20462) );
  OAI21_X1 U22645 ( .B1(n22346), .B2(n20473), .A(n20462), .ZN(P1_U2928) );
  INV_X1 U22646 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n22353) );
  AOI22_X1 U22647 ( .A1(n21905), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20463) );
  OAI21_X1 U22648 ( .B1(n22353), .B2(n20473), .A(n20463), .ZN(P1_U2927) );
  AOI22_X1 U22649 ( .A1(n20464), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20465) );
  OAI21_X1 U22650 ( .B1(n15134), .B2(n20473), .A(n20465), .ZN(P1_U2926) );
  AOI22_X1 U22651 ( .A1(n21905), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20466) );
  OAI21_X1 U22652 ( .B1(n15696), .B2(n20473), .A(n20466), .ZN(P1_U2925) );
  INV_X1 U22653 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n22371) );
  AOI22_X1 U22654 ( .A1(n21905), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20467) );
  OAI21_X1 U22655 ( .B1(n22371), .B2(n20473), .A(n20467), .ZN(P1_U2924) );
  INV_X1 U22656 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n22378) );
  AOI22_X1 U22657 ( .A1(n21905), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20468) );
  OAI21_X1 U22658 ( .B1(n22378), .B2(n20473), .A(n20468), .ZN(P1_U2923) );
  INV_X1 U22659 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n22388) );
  AOI22_X1 U22660 ( .A1(n21905), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20469), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20470) );
  OAI21_X1 U22661 ( .B1(n22388), .B2(n20473), .A(n20470), .ZN(P1_U2922) );
  AOI22_X1 U22662 ( .A1(n21905), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20471), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20472) );
  OAI21_X1 U22663 ( .B1(n20474), .B2(n20473), .A(n20472), .ZN(P1_U2921) );
  INV_X2 U22664 ( .A(n22727), .ZN(n20637) );
  OR2_X1 U22665 ( .A1(n20637), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20500) );
  NOR2_X1 U22666 ( .A1(n22251), .A2(n20637), .ZN(n20511) );
  INV_X1 U22667 ( .A(n20511), .ZN(n20497) );
  OAI222_X1 U22668 ( .A1(n20500), .A2(n20476), .B1(n20475), .B2(n22727), .C1(
        n20527), .C2(n20497), .ZN(P1_U3197) );
  AOI222_X1 U22669 ( .A1(n11178), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n20509), .ZN(n20477) );
  INV_X1 U22670 ( .A(n20477), .ZN(P1_U3198) );
  AOI222_X1 U22671 ( .A1(n20509), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n11178), .ZN(n20478) );
  INV_X1 U22672 ( .A(n20478), .ZN(P1_U3199) );
  AOI222_X1 U22673 ( .A1(n20509), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n11178), .ZN(n20479) );
  INV_X1 U22674 ( .A(n20479), .ZN(P1_U3200) );
  AOI222_X1 U22675 ( .A1(n20509), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n11178), .ZN(n20480) );
  INV_X1 U22676 ( .A(n20480), .ZN(P1_U3201) );
  AOI222_X1 U22677 ( .A1(n20509), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n11178), .ZN(n20481) );
  INV_X1 U22678 ( .A(n20481), .ZN(P1_U3202) );
  AOI222_X1 U22679 ( .A1(n20511), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n11178), .ZN(n20482) );
  INV_X1 U22680 ( .A(n20482), .ZN(P1_U3203) );
  AOI222_X1 U22681 ( .A1(n20509), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n11178), .ZN(n20483) );
  INV_X1 U22682 ( .A(n20483), .ZN(P1_U3204) );
  AOI222_X1 U22683 ( .A1(n20509), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n11178), .ZN(n20484) );
  INV_X1 U22684 ( .A(n20484), .ZN(P1_U3205) );
  AOI222_X1 U22685 ( .A1(n20511), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n11178), .ZN(n20485) );
  INV_X1 U22686 ( .A(n20485), .ZN(P1_U3206) );
  AOI222_X1 U22687 ( .A1(n11178), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20509), .ZN(n20486) );
  INV_X1 U22688 ( .A(n20486), .ZN(P1_U3207) );
  AOI222_X1 U22689 ( .A1(n20511), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n11178), .ZN(n20487) );
  INV_X1 U22690 ( .A(n20487), .ZN(P1_U3208) );
  AOI222_X1 U22691 ( .A1(n11178), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20509), .ZN(n20488) );
  INV_X1 U22692 ( .A(n20488), .ZN(P1_U3209) );
  AOI222_X1 U22693 ( .A1(n20511), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n11178), .ZN(n20489) );
  INV_X1 U22694 ( .A(n20489), .ZN(P1_U3210) );
  AOI22_X1 U22695 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n11178), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20637), .ZN(n20490) );
  OAI21_X1 U22696 ( .B1(n20491), .B2(n20497), .A(n20490), .ZN(P1_U3211) );
  AOI22_X1 U22697 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20509), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20637), .ZN(n20492) );
  OAI21_X1 U22698 ( .B1(n20493), .B2(n20500), .A(n20492), .ZN(P1_U3212) );
  AOI222_X1 U22699 ( .A1(n11178), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20509), .ZN(n20494) );
  INV_X1 U22700 ( .A(n20494), .ZN(P1_U3213) );
  AOI222_X1 U22701 ( .A1(n11178), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20509), .ZN(n20495) );
  INV_X1 U22702 ( .A(n20495), .ZN(P1_U3214) );
  AOI22_X1 U22703 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n11178), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20637), .ZN(n20496) );
  OAI21_X1 U22704 ( .B1(n20498), .B2(n20497), .A(n20496), .ZN(P1_U3215) );
  AOI22_X1 U22705 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20509), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20637), .ZN(n20499) );
  OAI21_X1 U22706 ( .B1(n22166), .B2(n20500), .A(n20499), .ZN(P1_U3216) );
  AOI222_X1 U22707 ( .A1(n20511), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n11178), .ZN(n20501) );
  INV_X1 U22708 ( .A(n20501), .ZN(P1_U3217) );
  AOI222_X1 U22709 ( .A1(n11178), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20509), .ZN(n20502) );
  INV_X1 U22710 ( .A(n20502), .ZN(P1_U3218) );
  AOI222_X1 U22711 ( .A1(n20509), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n11178), .ZN(n20503) );
  INV_X1 U22712 ( .A(n20503), .ZN(P1_U3219) );
  AOI222_X1 U22713 ( .A1(n20511), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n11178), .ZN(n20504) );
  INV_X1 U22714 ( .A(n20504), .ZN(P1_U3220) );
  AOI222_X1 U22715 ( .A1(n20511), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n11178), .ZN(n20505) );
  INV_X1 U22716 ( .A(n20505), .ZN(P1_U3221) );
  AOI222_X1 U22717 ( .A1(n20509), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n11178), .ZN(n20506) );
  INV_X1 U22718 ( .A(n20506), .ZN(P1_U3222) );
  AOI222_X1 U22719 ( .A1(n11178), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20509), .ZN(n20507) );
  INV_X1 U22720 ( .A(n20507), .ZN(P1_U3223) );
  AOI222_X1 U22721 ( .A1(n11178), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20511), .ZN(n20508) );
  INV_X1 U22722 ( .A(n20508), .ZN(P1_U3224) );
  AOI222_X1 U22723 ( .A1(n11178), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20509), .ZN(n20510) );
  INV_X1 U22724 ( .A(n20510), .ZN(P1_U3225) );
  AOI222_X1 U22725 ( .A1(n20511), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20637), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n11178), .ZN(n20512) );
  INV_X1 U22726 ( .A(n20512), .ZN(P1_U3226) );
  OAI22_X1 U22727 ( .A1(n20637), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22727), .ZN(n20513) );
  INV_X1 U22728 ( .A(n20513), .ZN(P1_U3458) );
  NOR4_X1 U22729 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20523) );
  NOR4_X1 U22730 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20522) );
  INV_X1 U22731 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22225) );
  NOR4_X1 U22732 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20514) );
  OAI21_X1 U22733 ( .B1(n20530), .B2(n22225), .A(n20514), .ZN(n20520) );
  NOR4_X1 U22734 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20518) );
  NOR4_X1 U22735 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20517) );
  NOR4_X1 U22736 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20516) );
  NOR4_X1 U22737 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20515) );
  NAND4_X1 U22738 ( .A1(n20518), .A2(n20517), .A3(n20516), .A4(n20515), .ZN(
        n20519) );
  NOR4_X1 U22739 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_30__SCAN_IN), .A3(n20520), .A4(n20519), .ZN(n20521)
         );
  NAND3_X1 U22740 ( .A1(n20523), .A2(n20522), .A3(n20521), .ZN(n20534) );
  INV_X1 U22741 ( .A(n20534), .ZN(n20539) );
  INV_X1 U22742 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20524) );
  NOR2_X1 U22743 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20534), .ZN(n20536) );
  NAND2_X1 U22744 ( .A1(n20536), .A2(n22225), .ZN(n20531) );
  NAND4_X1 U22745 ( .A1(n20539), .A2(n20526), .A3(n20530), .A4(n22225), .ZN(
        n20533) );
  OAI211_X1 U22746 ( .C1(n20539), .C2(n20524), .A(n20531), .B(n20533), .ZN(
        P1_U2808) );
  OAI22_X1 U22747 ( .A1(n20637), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22727), .ZN(n20525) );
  INV_X1 U22748 ( .A(n20525), .ZN(P1_U3459) );
  NAND2_X1 U22749 ( .A1(n20536), .A2(n20526), .ZN(n20538) );
  OAI21_X1 U22750 ( .B1(n20527), .B2(n20526), .A(n20539), .ZN(n20528) );
  OAI21_X1 U22751 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20539), .A(n20528), 
        .ZN(n20529) );
  OAI221_X1 U22752 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20531), .C1(n20530), .C2(n20538), .A(n20529), .ZN(P1_U3481) );
  OAI22_X1 U22753 ( .A1(n20637), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22727), .ZN(n20532) );
  INV_X1 U22754 ( .A(n20532), .ZN(P1_U3460) );
  OAI221_X1 U22755 ( .B1(n20536), .B2(n20535), .C1(n20536), .C2(n20534), .A(
        n20533), .ZN(P1_U2807) );
  OAI22_X1 U22756 ( .A1(n20637), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22727), .ZN(n20537) );
  INV_X1 U22757 ( .A(n20537), .ZN(P1_U3461) );
  OAI21_X1 U22758 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n20539), .A(n20538), 
        .ZN(n20540) );
  INV_X1 U22759 ( .A(n20540), .ZN(P1_U3482) );
  NOR2_X1 U22760 ( .A1(n22027), .A2(n20551), .ZN(n20541) );
  AOI21_X1 U22761 ( .B1(n20624), .B2(n13591), .A(n20541), .ZN(n20542) );
  OAI21_X1 U22762 ( .B1(n20556), .B2(n20543), .A(n20542), .ZN(P1_U2855) );
  AOI22_X1 U22763 ( .A1(n20611), .A2(n13591), .B1(n20544), .B2(n22008), .ZN(
        n20545) );
  OAI21_X1 U22764 ( .B1(n20556), .B2(n15801), .A(n20545), .ZN(P1_U2857) );
  INV_X1 U22765 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n22177) );
  OAI22_X1 U22766 ( .A1(n22182), .A2(n16572), .B1(n20551), .B2(n22180), .ZN(
        n20546) );
  INV_X1 U22767 ( .A(n20546), .ZN(n20547) );
  OAI21_X1 U22768 ( .B1(n20556), .B2(n22177), .A(n20547), .ZN(P1_U2849) );
  INV_X1 U22769 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n20550) );
  NOR2_X1 U22770 ( .A1(n22169), .A2(n20551), .ZN(n20548) );
  AOI21_X1 U22771 ( .B1(n22171), .B2(n13591), .A(n20548), .ZN(n20549) );
  OAI21_X1 U22772 ( .B1(n20556), .B2(n20550), .A(n20549), .ZN(P1_U2851) );
  OAI22_X1 U22773 ( .A1(n20552), .A2(n16572), .B1(n20551), .B2(n21955), .ZN(
        n20553) );
  INV_X1 U22774 ( .A(n20553), .ZN(n20554) );
  OAI21_X1 U22775 ( .B1(n20556), .B2(n20555), .A(n20554), .ZN(P1_U2867) );
  AOI22_X1 U22776 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20564) );
  OR2_X1 U22777 ( .A1(n20558), .A2(n20557), .ZN(n20559) );
  NAND2_X1 U22778 ( .A1(n20560), .A2(n20559), .ZN(n21928) );
  INV_X1 U22779 ( .A(n21928), .ZN(n20562) );
  INV_X1 U22780 ( .A(n20561), .ZN(n22065) );
  AOI22_X1 U22781 ( .A1(n20562), .A2(n20629), .B1(n20628), .B2(n22065), .ZN(
        n20563) );
  OAI211_X1 U22782 ( .C1(n20633), .C2(n22067), .A(n20564), .B(n20563), .ZN(
        P1_U2995) );
  AOI22_X1 U22783 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20572) );
  OAI21_X1 U22784 ( .B1(n20568), .B2(n20567), .A(n20566), .ZN(n20569) );
  INV_X1 U22785 ( .A(n20569), .ZN(n21961) );
  AOI22_X1 U22786 ( .A1(n21961), .A2(n20629), .B1(n20628), .B2(n20570), .ZN(
        n20571) );
  OAI211_X1 U22787 ( .C1(n20633), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P1_U2994) );
  AOI22_X1 U22788 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20581) );
  OAI21_X1 U22789 ( .B1(n20576), .B2(n20575), .A(n20574), .ZN(n20577) );
  INV_X1 U22790 ( .A(n20577), .ZN(n21947) );
  INV_X1 U22791 ( .A(n20578), .ZN(n20579) );
  AOI22_X1 U22792 ( .A1(n21947), .A2(n20629), .B1(n20628), .B2(n20579), .ZN(
        n20580) );
  OAI211_X1 U22793 ( .C1(n20633), .C2(n20582), .A(n20581), .B(n20580), .ZN(
        P1_U2993) );
  AOI22_X1 U22794 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20588) );
  OAI21_X1 U22795 ( .B1(n20585), .B2(n20584), .A(n20583), .ZN(n20586) );
  INV_X1 U22796 ( .A(n20586), .ZN(n21966) );
  AOI22_X1 U22797 ( .A1(n21966), .A2(n20629), .B1(n20628), .B2(n22077), .ZN(
        n20587) );
  OAI211_X1 U22798 ( .C1(n20633), .C2(n22079), .A(n20588), .B(n20587), .ZN(
        P1_U2992) );
  NOR2_X1 U22799 ( .A1(n22016), .A2(n20589), .ZN(n21995) );
  NOR2_X1 U22800 ( .A1(n20590), .A2(n20593), .ZN(n20592) );
  MUX2_X1 U22801 ( .A(n20593), .B(n20592), .S(n20591), .Z(n20594) );
  XNOR2_X1 U22802 ( .A(n20594), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n21994) );
  OAI22_X1 U22803 ( .A1(n21994), .A2(n22203), .B1(n20633), .B2(n20595), .ZN(
        n20596) );
  AOI211_X1 U22804 ( .C1(n20627), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21995), .B(n20596), .ZN(n20597) );
  OAI21_X1 U22805 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(P1_U2988) );
  OAI21_X1 U22806 ( .B1(n20602), .B2(n20601), .A(n20600), .ZN(n20603) );
  INV_X1 U22807 ( .A(n20603), .ZN(n21988) );
  AOI22_X1 U22808 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20605) );
  AOI22_X1 U22809 ( .A1(n20623), .A2(n22099), .B1(n20628), .B2(n22098), .ZN(
        n20604) );
  OAI211_X1 U22810 ( .C1(n21988), .C2(n22203), .A(n20605), .B(n20604), .ZN(
        P1_U2987) );
  OAI21_X1 U22811 ( .B1(n20608), .B2(n20607), .A(n20606), .ZN(n20609) );
  INV_X1 U22812 ( .A(n20609), .ZN(n22010) );
  AOI22_X1 U22813 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n20613) );
  AOI22_X1 U22814 ( .A1(n20611), .A2(n20628), .B1(n20623), .B2(n20610), .ZN(
        n20612) );
  OAI211_X1 U22815 ( .C1(n22010), .C2(n22203), .A(n20613), .B(n20612), .ZN(
        P1_U2984) );
  NAND2_X1 U22816 ( .A1(n11595), .A2(n20614), .ZN(n20620) );
  INV_X1 U22817 ( .A(n20615), .ZN(n20616) );
  OAI21_X1 U22818 ( .B1(n20618), .B2(n20617), .A(n20616), .ZN(n20619) );
  MUX2_X1 U22819 ( .A(n11595), .B(n20620), .S(n20619), .Z(n20621) );
  XNOR2_X1 U22820 ( .A(n20621), .B(n22024), .ZN(n22034) );
  AOI22_X1 U22821 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20626) );
  AOI22_X1 U22822 ( .A1(n20624), .A2(n20628), .B1(n20623), .B2(n20622), .ZN(
        n20625) );
  OAI211_X1 U22823 ( .C1(n22203), .C2(n22034), .A(n20626), .B(n20625), .ZN(
        P1_U2982) );
  AOI22_X1 U22824 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20627), .B1(
        n22040), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n20632) );
  AOI22_X1 U22825 ( .A1(n20630), .A2(n20629), .B1(n22145), .B2(n20628), .ZN(
        n20631) );
  OAI211_X1 U22826 ( .C1(n20633), .C2(n22142), .A(n20632), .B(n20631), .ZN(
        P1_U2980) );
  OAI21_X1 U22827 ( .B1(n20634), .B2(n22220), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20635) );
  OAI21_X1 U22828 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20636), .A(n20635), 
        .ZN(P1_U2803) );
  OAI222_X1 U22829 ( .A1(n22727), .A2(n20639), .B1(n22727), .B2(n20638), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(n20637), .ZN(P1_U2804) );
  INV_X1 U22830 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20642) );
  AOI22_X1 U22831 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n11177), .ZN(n20641) );
  OAI21_X1 U22832 ( .B1(n20642), .B2(n20706), .A(n20641), .ZN(U247) );
  INV_X1 U22833 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U22834 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n11177), .ZN(n20643) );
  OAI21_X1 U22835 ( .B1(n20644), .B2(n20706), .A(n20643), .ZN(U246) );
  INV_X1 U22836 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U22837 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n11177), .ZN(n20645) );
  OAI21_X1 U22838 ( .B1(n20646), .B2(n20706), .A(n20645), .ZN(U245) );
  INV_X1 U22839 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20648) );
  AOI22_X1 U22840 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n11177), .ZN(n20647) );
  OAI21_X1 U22841 ( .B1(n20648), .B2(n20706), .A(n20647), .ZN(U244) );
  INV_X1 U22842 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U22843 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n11177), .ZN(n20649) );
  OAI21_X1 U22844 ( .B1(n20650), .B2(n20706), .A(n20649), .ZN(U243) );
  AOI22_X1 U22845 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n11177), .ZN(n20651) );
  OAI21_X1 U22846 ( .B1(n20652), .B2(n20706), .A(n20651), .ZN(U242) );
  INV_X1 U22847 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20654) );
  AOI22_X1 U22848 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n11177), .ZN(n20653) );
  OAI21_X1 U22849 ( .B1(n20654), .B2(n20706), .A(n20653), .ZN(U241) );
  INV_X1 U22850 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20656) );
  AOI22_X1 U22851 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11177), .ZN(n20655) );
  OAI21_X1 U22852 ( .B1(n20656), .B2(n20706), .A(n20655), .ZN(U240) );
  INV_X1 U22853 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20658) );
  AOI22_X1 U22854 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n11177), .ZN(n20657) );
  OAI21_X1 U22855 ( .B1(n20658), .B2(n20706), .A(n20657), .ZN(U239) );
  INV_X1 U22856 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20660) );
  AOI22_X1 U22857 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n11177), .ZN(n20659) );
  OAI21_X1 U22858 ( .B1(n20660), .B2(n20706), .A(n20659), .ZN(U238) );
  AOI22_X1 U22859 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11177), .ZN(n20661) );
  OAI21_X1 U22860 ( .B1(n20662), .B2(n20706), .A(n20661), .ZN(U237) );
  INV_X1 U22861 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20664) );
  AOI22_X1 U22862 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11177), .ZN(n20663) );
  OAI21_X1 U22863 ( .B1(n20664), .B2(n20706), .A(n20663), .ZN(U236) );
  INV_X1 U22864 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20666) );
  AOI22_X1 U22865 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11177), .ZN(n20665) );
  OAI21_X1 U22866 ( .B1(n20666), .B2(n20706), .A(n20665), .ZN(U235) );
  INV_X1 U22867 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20668) );
  AOI22_X1 U22868 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11177), .ZN(n20667) );
  OAI21_X1 U22869 ( .B1(n20668), .B2(n20706), .A(n20667), .ZN(U234) );
  INV_X1 U22870 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20670) );
  AOI22_X1 U22871 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11177), .ZN(n20669) );
  OAI21_X1 U22872 ( .B1(n20670), .B2(n20706), .A(n20669), .ZN(U233) );
  INV_X1 U22873 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20672) );
  AOI22_X1 U22874 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11177), .ZN(n20671) );
  OAI21_X1 U22875 ( .B1(n20672), .B2(n20706), .A(n20671), .ZN(U232) );
  AOI22_X1 U22876 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11177), .ZN(n20673) );
  OAI21_X1 U22877 ( .B1(n20674), .B2(n20706), .A(n20673), .ZN(U231) );
  AOI22_X1 U22878 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11177), .ZN(n20675) );
  OAI21_X1 U22879 ( .B1(n20676), .B2(n20706), .A(n20675), .ZN(U230) );
  AOI22_X1 U22880 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11177), .ZN(n20677) );
  OAI21_X1 U22881 ( .B1(n20678), .B2(n20706), .A(n20677), .ZN(U229) );
  AOI22_X1 U22882 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n11177), .ZN(n20679) );
  OAI21_X1 U22883 ( .B1(n20680), .B2(n20706), .A(n20679), .ZN(U228) );
  AOI22_X1 U22884 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n11177), .ZN(n20681) );
  OAI21_X1 U22885 ( .B1(n20682), .B2(n20706), .A(n20681), .ZN(U227) );
  AOI22_X1 U22886 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11177), .ZN(n20683) );
  OAI21_X1 U22887 ( .B1(n20684), .B2(n20706), .A(n20683), .ZN(U226) );
  AOI22_X1 U22888 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n11177), .ZN(n20685) );
  OAI21_X1 U22889 ( .B1(n20686), .B2(n20706), .A(n20685), .ZN(U225) );
  AOI22_X1 U22890 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n11177), .ZN(n20687) );
  OAI21_X1 U22891 ( .B1(n20688), .B2(n20706), .A(n20687), .ZN(U224) );
  AOI22_X1 U22892 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11177), .ZN(n20689) );
  OAI21_X1 U22893 ( .B1(n20690), .B2(n20706), .A(n20689), .ZN(U223) );
  AOI22_X1 U22894 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11177), .ZN(n20691) );
  OAI21_X1 U22895 ( .B1(n20692), .B2(n20706), .A(n20691), .ZN(U222) );
  AOI22_X1 U22896 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n11177), .ZN(n20694) );
  OAI21_X1 U22897 ( .B1(n20695), .B2(n20706), .A(n20694), .ZN(U221) );
  AOI22_X1 U22898 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n11177), .ZN(n20696) );
  OAI21_X1 U22899 ( .B1(n20697), .B2(n20706), .A(n20696), .ZN(U220) );
  AOI22_X1 U22900 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n11177), .ZN(n20698) );
  OAI21_X1 U22901 ( .B1(n20699), .B2(n20706), .A(n20698), .ZN(U219) );
  AOI22_X1 U22902 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n11177), .ZN(n20700) );
  OAI21_X1 U22903 ( .B1(n20701), .B2(n20706), .A(n20700), .ZN(U218) );
  AOI22_X1 U22904 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20693), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n11177), .ZN(n20702) );
  OAI21_X1 U22905 ( .B1(n20703), .B2(n20706), .A(n20702), .ZN(U217) );
  OAI222_X1 U22906 ( .A1(U212), .A2(n20707), .B1(n20706), .B2(n20705), .C1(
        U214), .C2(n20704), .ZN(U216) );
  AOI22_X1 U22907 ( .A1(n22727), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20708), 
        .B2(n20637), .ZN(P1_U3483) );
  OAI21_X1 U22908 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20710), .A(n20709), 
        .ZN(n20712) );
  AOI211_X1 U22909 ( .C1(n20713), .C2(n20712), .A(n22292), .B(n20711), .ZN(
        n20716) );
  OAI21_X1 U22910 ( .B1(n20716), .B2(n20715), .A(n20714), .ZN(n20723) );
  INV_X1 U22911 ( .A(n20717), .ZN(n20718) );
  AOI22_X1 U22912 ( .A1(n20719), .A2(n21875), .B1(n20718), .B2(n21897), .ZN(
        n20721) );
  NAND2_X1 U22913 ( .A1(n20721), .A2(n20720), .ZN(n20722) );
  MUX2_X1 U22914 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20723), .S(n20722), 
        .Z(P3_U3296) );
  AND3_X2 U22915 ( .A1(n21875), .A2(n20726), .A3(n20725), .ZN(n20775) );
  AOI22_X1 U22916 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20774), .ZN(n20728) );
  OAI21_X1 U22917 ( .B1(n20729), .B2(n20777), .A(n20728), .ZN(P3_U2768) );
  AOI22_X1 U22918 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20774), .ZN(n20730) );
  OAI21_X1 U22919 ( .B1(n21251), .B2(n20777), .A(n20730), .ZN(P3_U2769) );
  AOI22_X1 U22920 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20774), .ZN(n20731) );
  OAI21_X1 U22921 ( .B1(n20732), .B2(n20777), .A(n20731), .ZN(P3_U2770) );
  AOI22_X1 U22922 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20765), .ZN(n20733) );
  OAI21_X1 U22923 ( .B1(n21273), .B2(n20777), .A(n20733), .ZN(P3_U2771) );
  AOI22_X1 U22924 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20765), .ZN(n20734) );
  OAI21_X1 U22925 ( .B1(n21263), .B2(n20777), .A(n20734), .ZN(P3_U2772) );
  AOI22_X1 U22926 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20765), .ZN(n20735) );
  OAI21_X1 U22927 ( .B1(n21258), .B2(n20777), .A(n20735), .ZN(P3_U2773) );
  AOI22_X1 U22928 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20765), .ZN(n20736) );
  OAI21_X1 U22929 ( .B1(n20737), .B2(n20777), .A(n20736), .ZN(P3_U2774) );
  AOI22_X1 U22930 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20765), .ZN(n20738) );
  OAI21_X1 U22931 ( .B1(n20739), .B2(n20777), .A(n20738), .ZN(P3_U2775) );
  AOI22_X1 U22932 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20765), .ZN(n20740) );
  OAI21_X1 U22933 ( .B1(n20741), .B2(n20777), .A(n20740), .ZN(P3_U2776) );
  AOI22_X1 U22934 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20765), .ZN(n20742) );
  OAI21_X1 U22935 ( .B1(n20743), .B2(n20777), .A(n20742), .ZN(P3_U2777) );
  AOI22_X1 U22936 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20765), .ZN(n20744) );
  OAI21_X1 U22937 ( .B1(n21297), .B2(n20777), .A(n20744), .ZN(P3_U2778) );
  AOI22_X1 U22938 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20765), .ZN(n20745) );
  OAI21_X1 U22939 ( .B1(n20746), .B2(n20777), .A(n20745), .ZN(P3_U2779) );
  AOI22_X1 U22940 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20774), .ZN(n20747) );
  OAI21_X1 U22941 ( .B1(n20748), .B2(n20777), .A(n20747), .ZN(P3_U2780) );
  AOI22_X1 U22942 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20774), .ZN(n20749) );
  OAI21_X1 U22943 ( .B1(n21309), .B2(n20777), .A(n20749), .ZN(P3_U2781) );
  AOI22_X1 U22944 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20775), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20774), .ZN(n20750) );
  OAI21_X1 U22945 ( .B1(n20751), .B2(n20777), .A(n20750), .ZN(P3_U2782) );
  AOI22_X1 U22946 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20774), .ZN(n20752) );
  OAI21_X1 U22947 ( .B1(n21376), .B2(n20777), .A(n20752), .ZN(P3_U2783) );
  AOI22_X1 U22948 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20774), .ZN(n20753) );
  OAI21_X1 U22949 ( .B1(n21369), .B2(n20777), .A(n20753), .ZN(P3_U2784) );
  AOI22_X1 U22950 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20774), .ZN(n20754) );
  OAI21_X1 U22951 ( .B1(n21219), .B2(n20777), .A(n20754), .ZN(P3_U2785) );
  AOI22_X1 U22952 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20774), .ZN(n20755) );
  OAI21_X1 U22953 ( .B1(n20756), .B2(n20777), .A(n20755), .ZN(P3_U2786) );
  AOI22_X1 U22954 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20774), .ZN(n20757) );
  OAI21_X1 U22955 ( .B1(n21220), .B2(n20777), .A(n20757), .ZN(P3_U2787) );
  AOI22_X1 U22956 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20774), .ZN(n20758) );
  OAI21_X1 U22957 ( .B1(n20759), .B2(n20777), .A(n20758), .ZN(P3_U2788) );
  AOI22_X1 U22958 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20774), .ZN(n20760) );
  OAI21_X1 U22959 ( .B1(n21221), .B2(n20777), .A(n20760), .ZN(P3_U2789) );
  AOI22_X1 U22960 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20774), .ZN(n20761) );
  OAI21_X1 U22961 ( .B1(n20762), .B2(n20777), .A(n20761), .ZN(P3_U2790) );
  AOI22_X1 U22962 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20774), .ZN(n20763) );
  OAI21_X1 U22963 ( .B1(n21360), .B2(n20777), .A(n20763), .ZN(P3_U2791) );
  AOI22_X1 U22964 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20765), .ZN(n20764) );
  OAI21_X1 U22965 ( .B1(n21248), .B2(n20777), .A(n20764), .ZN(P3_U2792) );
  AOI22_X1 U22966 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20765), .ZN(n20766) );
  OAI21_X1 U22967 ( .B1(n20767), .B2(n20777), .A(n20766), .ZN(P3_U2793) );
  AOI22_X1 U22968 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20774), .ZN(n20768) );
  OAI21_X1 U22969 ( .B1(n21203), .B2(n20777), .A(n20768), .ZN(P3_U2794) );
  AOI22_X1 U22970 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20774), .ZN(n20769) );
  OAI21_X1 U22971 ( .B1(n20770), .B2(n20777), .A(n20769), .ZN(P3_U2795) );
  AOI22_X1 U22972 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20774), .ZN(n20771) );
  OAI21_X1 U22973 ( .B1(n20772), .B2(n20777), .A(n20771), .ZN(P3_U2796) );
  AOI22_X1 U22974 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20774), .ZN(n20773) );
  OAI21_X1 U22975 ( .B1(n21348), .B2(n20777), .A(n20773), .ZN(P3_U2797) );
  AOI22_X1 U22976 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20775), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20774), .ZN(n20776) );
  OAI21_X1 U22977 ( .B1(n21351), .B2(n20777), .A(n20776), .ZN(P3_U2798) );
  NAND2_X1 U22978 ( .A1(n20778), .A2(n20789), .ZN(n21381) );
  AOI22_X1 U22979 ( .A1(n21185), .A2(n20779), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n20879), .ZN(n20785) );
  NOR2_X1 U22980 ( .A1(n21151), .A2(n21882), .ZN(n20857) );
  INV_X1 U22981 ( .A(n20857), .ZN(n21180) );
  OAI21_X1 U22982 ( .B1(n20892), .B2(n21180), .A(n21170), .ZN(n20783) );
  AOI21_X1 U22983 ( .B1(n21018), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21882), .ZN(n20950) );
  OAI22_X1 U22984 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n21081), .B1(n21168), 
        .B2(n20780), .ZN(n20781) );
  AOI221_X1 U22985 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20783), .C1(
        n20782), .C2(n20950), .A(n20781), .ZN(n20784) );
  OAI211_X1 U22986 ( .C1(n21381), .C2(n20809), .A(n20785), .B(n20784), .ZN(
        P3_U2670) );
  INV_X1 U22987 ( .A(n21882), .ZN(n21157) );
  NAND2_X1 U22988 ( .A1(n21151), .A2(n21157), .ZN(n20911) );
  AOI211_X1 U22989 ( .C1(n20788), .C2(n20787), .A(n20786), .B(n21081), .ZN(
        n20797) );
  INV_X1 U22990 ( .A(n20789), .ZN(n21406) );
  NOR2_X1 U22991 ( .A1(n21406), .A2(n21851), .ZN(n21400) );
  NOR2_X1 U22992 ( .A1(n20790), .A2(n21400), .ZN(n21395) );
  AOI22_X1 U22993 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n21092), .B1(
        P3_REIP_REG_2__SCAN_IN), .B2(n20879), .ZN(n20795) );
  INV_X1 U22994 ( .A(n20814), .ZN(n20791) );
  OAI211_X1 U22995 ( .C1(n20793), .C2(n20792), .A(n21185), .B(n20791), .ZN(
        n20794) );
  OAI211_X1 U22996 ( .C1(n21395), .C2(n20809), .A(n20795), .B(n20794), .ZN(
        n20796) );
  AOI211_X1 U22997 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n21186), .A(n20797), .B(
        n20796), .ZN(n20799) );
  INV_X1 U22998 ( .A(n20803), .ZN(n21013) );
  OAI221_X1 U22999 ( .B1(n21013), .B2(n20800), .C1(n20803), .C2(n20804), .A(
        n20857), .ZN(n20798) );
  OAI211_X1 U23000 ( .C1(n20800), .C2(n20911), .A(n20799), .B(n20798), .ZN(
        P3_U2669) );
  INV_X1 U23001 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20817) );
  OAI21_X1 U23002 ( .B1(n20820), .B2(n21081), .A(n21184), .ZN(n20826) );
  OAI21_X1 U23003 ( .B1(n21081), .B2(n20802), .A(n20801), .ZN(n20812) );
  OAI21_X1 U23004 ( .B1(n20804), .B2(n20803), .A(n21018), .ZN(n20806) );
  OAI21_X1 U23005 ( .B1(n20807), .B2(n20806), .A(n21157), .ZN(n20805) );
  AOI21_X1 U23006 ( .B1(n20807), .B2(n20806), .A(n20805), .ZN(n20811) );
  AOI21_X1 U23007 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21391), .A(
        n21848), .ZN(n21411) );
  NOR2_X1 U23008 ( .A1(n20808), .A2(n21411), .ZN(n21422) );
  OAI22_X1 U23009 ( .A1(n21422), .A2(n20809), .B1(n21168), .B2(n20813), .ZN(
        n20810) );
  AOI211_X1 U23010 ( .C1(n20826), .C2(n20812), .A(n20811), .B(n20810), .ZN(
        n20816) );
  OAI211_X1 U23011 ( .C1(n20814), .C2(n20813), .A(n21185), .B(n20818), .ZN(
        n20815) );
  OAI211_X1 U23012 ( .C1(n21170), .C2(n20817), .A(n20816), .B(n20815), .ZN(
        P3_U2668) );
  AOI22_X1 U23013 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n21092), .B1(
        n21186), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n20833) );
  AOI211_X1 U23014 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20818), .A(n20840), .B(
        n21160), .ZN(n20825) );
  NAND3_X1 U23015 ( .A1(n21103), .A2(n20820), .A3(n20819), .ZN(n20823) );
  OAI21_X1 U23016 ( .B1(n20821), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n21182), .ZN(n20822) );
  NAND3_X1 U23017 ( .A1(n21808), .A2(n20823), .A3(n20822), .ZN(n20824) );
  AOI211_X1 U23018 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n20826), .A(n20825), .B(
        n20824), .ZN(n20832) );
  INV_X1 U23019 ( .A(n20911), .ZN(n20979) );
  INV_X1 U23020 ( .A(n20829), .ZN(n20827) );
  OAI211_X1 U23021 ( .C1(n20979), .C2(n20828), .A(n20827), .B(n20950), .ZN(
        n20831) );
  OAI211_X1 U23022 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20836), .A(
        n20857), .B(n20829), .ZN(n20830) );
  NAND4_X1 U23023 ( .A1(n20833), .A2(n20832), .A3(n20831), .A4(n20830), .ZN(
        P3_U2667) );
  OAI21_X1 U23024 ( .B1(n20850), .B2(n21081), .A(n21184), .ZN(n20862) );
  OAI21_X1 U23025 ( .B1(n21081), .B2(n20835), .A(n20834), .ZN(n20845) );
  OAI21_X1 U23026 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20836), .A(
        n21018), .ZN(n20838) );
  AOI21_X1 U23027 ( .B1(n20839), .B2(n20838), .A(n21882), .ZN(n20837) );
  OAI21_X1 U23028 ( .B1(n20839), .B2(n20838), .A(n20837), .ZN(n20842) );
  OAI211_X1 U23029 ( .C1(n20840), .C2(n20847), .A(n21185), .B(n20848), .ZN(
        n20841) );
  OAI211_X1 U23030 ( .C1(n21170), .C2(n20843), .A(n20842), .B(n20841), .ZN(
        n20844) );
  AOI21_X1 U23031 ( .B1(n20862), .B2(n20845), .A(n20844), .ZN(n20846) );
  OAI211_X1 U23032 ( .C1(n21168), .C2(n20847), .A(n20846), .B(n21808), .ZN(
        P3_U2666) );
  AOI22_X1 U23033 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21092), .B1(
        n21186), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n20861) );
  AOI211_X1 U23034 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20848), .A(n20868), .B(
        n21160), .ZN(n20852) );
  NAND3_X1 U23035 ( .A1(n21103), .A2(n20850), .A3(n20849), .ZN(n20875) );
  NAND2_X1 U23036 ( .A1(n21808), .A2(n20875), .ZN(n20851) );
  AOI211_X1 U23037 ( .C1(n20862), .C2(P3_REIP_REG_6__SCAN_IN), .A(n20852), .B(
        n20851), .ZN(n20860) );
  OAI211_X1 U23038 ( .C1(n20979), .C2(n20853), .A(n20854), .B(n20950), .ZN(
        n20859) );
  INV_X1 U23039 ( .A(n20854), .ZN(n20856) );
  NAND2_X1 U23040 ( .A1(n20855), .A2(n21013), .ZN(n20921) );
  NAND3_X1 U23041 ( .A1(n20857), .A2(n20856), .A3(n20921), .ZN(n20858) );
  NAND4_X1 U23042 ( .A1(n20861), .A2(n20860), .A3(n20859), .A4(n20858), .ZN(
        P3_U2665) );
  INV_X1 U23043 ( .A(n20862), .ZN(n20876) );
  NAND2_X1 U23044 ( .A1(n21018), .A2(n20921), .ZN(n20863) );
  XOR2_X1 U23045 ( .A(n20864), .B(n20863), .Z(n20873) );
  NOR3_X1 U23046 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21081), .A3(n20865), .ZN(
        n20866) );
  AOI211_X1 U23047 ( .C1(n21186), .C2(P3_EBX_REG_7__SCAN_IN), .A(n21832), .B(
        n20866), .ZN(n20870) );
  OAI211_X1 U23048 ( .C1(n20868), .C2(n20867), .A(n21185), .B(n20878), .ZN(
        n20869) );
  OAI211_X1 U23049 ( .C1(n21170), .C2(n20871), .A(n20870), .B(n20869), .ZN(
        n20872) );
  AOI21_X1 U23050 ( .B1(n21157), .B2(n20873), .A(n20872), .ZN(n20874) );
  OAI221_X1 U23051 ( .B1(n20877), .B2(n20876), .C1(n20877), .C2(n20875), .A(
        n20874), .ZN(P3_U2664) );
  INV_X1 U23052 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20889) );
  AOI211_X1 U23053 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20878), .A(n20893), .B(
        n21160), .ZN(n20887) );
  AOI21_X1 U23054 ( .B1(n21103), .B2(n20890), .A(n20879), .ZN(n20907) );
  AOI21_X1 U23055 ( .B1(n21103), .B2(n20880), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n20885) );
  OAI21_X1 U23056 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20881), .A(
        n21018), .ZN(n20882) );
  XNOR2_X1 U23057 ( .A(n20883), .B(n20882), .ZN(n20884) );
  OAI22_X1 U23058 ( .A1(n20907), .A2(n20885), .B1(n21882), .B2(n20884), .ZN(
        n20886) );
  AOI211_X1 U23059 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20887), .B(n20886), .ZN(n20888) );
  OAI211_X1 U23060 ( .C1(n21168), .C2(n20889), .A(n20888), .B(n21808), .ZN(
        P3_U2663) );
  NOR3_X1 U23061 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n21081), .A3(n20890), .ZN(
        n20915) );
  AND2_X1 U23062 ( .A1(n20892), .A2(n20891), .ZN(n20909) );
  NOR3_X1 U23063 ( .A1(n20899), .A2(n20909), .A3(n21180), .ZN(n20898) );
  OAI211_X1 U23064 ( .C1(n20893), .C2(n20895), .A(n21185), .B(n20905), .ZN(
        n20894) );
  NAND2_X1 U23065 ( .A1(n21808), .A2(n20894), .ZN(n20897) );
  OAI22_X1 U23066 ( .A1(n20900), .A2(n21170), .B1(n21168), .B2(n20895), .ZN(
        n20896) );
  NOR4_X1 U23067 ( .A1(n20915), .A2(n20898), .A3(n20897), .A4(n20896), .ZN(
        n20902) );
  OAI211_X1 U23068 ( .C1(n20979), .C2(n20900), .A(n20899), .B(n20950), .ZN(
        n20901) );
  OAI211_X1 U23069 ( .C1(n20907), .C2(n21830), .A(n20902), .B(n20901), .ZN(
        P3_U2662) );
  NOR2_X1 U23070 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n21081), .ZN(n20903) );
  AOI22_X1 U23071 ( .A1(n21186), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n20904), 
        .B2(n20903), .ZN(n20918) );
  AOI211_X1 U23072 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20905), .A(n20926), .B(
        n21160), .ZN(n20906) );
  AOI211_X1 U23073 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n21092), .A(
        n21832), .B(n20906), .ZN(n20917) );
  INV_X1 U23074 ( .A(n20907), .ZN(n20914) );
  AOI21_X1 U23075 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20909), .A(
        n21151), .ZN(n20908) );
  INV_X1 U23076 ( .A(n20908), .ZN(n20923) );
  OAI21_X1 U23077 ( .B1(n20909), .B2(n20912), .A(n21157), .ZN(n20910) );
  AOI22_X1 U23078 ( .A1(n20912), .A2(n20923), .B1(n20911), .B2(n20910), .ZN(
        n20913) );
  AOI221_X1 U23079 ( .B1(n20915), .B2(P3_REIP_REG_10__SCAN_IN), .C1(n20914), 
        .C2(P3_REIP_REG_10__SCAN_IN), .A(n20913), .ZN(n20916) );
  NAND3_X1 U23080 ( .A1(n20918), .A2(n20917), .A3(n20916), .ZN(P3_U2661) );
  OAI21_X1 U23081 ( .B1(n20919), .B2(n21081), .A(n21184), .ZN(n20945) );
  NOR2_X1 U23082 ( .A1(n21081), .A2(n20920), .ZN(n20931) );
  NOR2_X1 U23083 ( .A1(n20922), .A2(n20921), .ZN(n20974) );
  NOR2_X1 U23084 ( .A1(n20974), .A2(n21151), .ZN(n20938) );
  INV_X1 U23085 ( .A(n20925), .ZN(n20924) );
  OAI221_X1 U23086 ( .B1(n20925), .B2(n20938), .C1(n20924), .C2(n20923), .A(
        n21157), .ZN(n20928) );
  OAI211_X1 U23087 ( .C1(n20926), .C2(n20933), .A(n21185), .B(n20934), .ZN(
        n20927) );
  OAI211_X1 U23088 ( .C1(n21170), .C2(n20929), .A(n20928), .B(n20927), .ZN(
        n20930) );
  AOI221_X1 U23089 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n20945), .C1(n20931), 
        .C2(n20945), .A(n20930), .ZN(n20932) );
  OAI211_X1 U23090 ( .C1(n21168), .C2(n20933), .A(n20932), .B(n21808), .ZN(
        P3_U2660) );
  AOI211_X1 U23091 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20934), .A(n20946), .B(
        n21160), .ZN(n20935) );
  AOI211_X1 U23092 ( .C1(n21186), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21832), .B(
        n20935), .ZN(n20942) );
  INV_X1 U23093 ( .A(n20938), .ZN(n20936) );
  AOI221_X1 U23094 ( .B1(n20939), .B2(n20938), .C1(n20937), .C2(n20936), .A(
        n21882), .ZN(n20940) );
  AOI221_X1 U23095 ( .B1(n20945), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n21067), 
        .C2(n20953), .A(n20940), .ZN(n20941) );
  OAI211_X1 U23096 ( .C1(n20943), .C2(n21170), .A(n20942), .B(n20941), .ZN(
        P3_U2659) );
  AOI21_X1 U23097 ( .B1(n20975), .B2(n20974), .A(n21151), .ZN(n20960) );
  NOR2_X1 U23098 ( .A1(n20951), .A2(n21882), .ZN(n20944) );
  AOI22_X1 U23099 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n20945), .B1(n20960), 
        .B2(n20944), .ZN(n20958) );
  OAI211_X1 U23100 ( .C1(n20946), .C2(n20948), .A(n21185), .B(n20963), .ZN(
        n20947) );
  OAI211_X1 U23101 ( .C1(n21168), .C2(n20948), .A(n21808), .B(n20947), .ZN(
        n20949) );
  AOI21_X1 U23102 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n21092), .A(
        n20949), .ZN(n20957) );
  OAI211_X1 U23103 ( .C1(n20952), .C2(n21151), .A(n20951), .B(n20950), .ZN(
        n20956) );
  OAI221_X1 U23104 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n20954), .C2(n20953), .A(n21067), .ZN(n20955) );
  NAND4_X1 U23105 ( .A1(n20958), .A2(n20957), .A3(n20956), .A4(n20955), .ZN(
        P3_U2658) );
  XOR2_X1 U23106 ( .A(n20960), .B(n20959), .Z(n20968) );
  AOI21_X1 U23107 ( .B1(n21186), .B2(P3_EBX_REG_14__SCAN_IN), .A(n21832), .ZN(
        n20967) );
  NAND2_X1 U23108 ( .A1(n21183), .A2(n20998), .ZN(n20987) );
  AOI21_X1 U23109 ( .B1(n20962), .B2(n20961), .A(n20987), .ZN(n20965) );
  AOI211_X1 U23110 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20963), .A(n20969), .B(
        n21160), .ZN(n20964) );
  AOI211_X1 U23111 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20965), .B(n20964), .ZN(n20966) );
  OAI211_X1 U23112 ( .C1(n21882), .C2(n20968), .A(n20967), .B(n20966), .ZN(
        P3_U2657) );
  NOR2_X1 U23113 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n21052), .ZN(n20973) );
  OAI211_X1 U23114 ( .C1(n20969), .C2(n20971), .A(n21185), .B(n20984), .ZN(
        n20970) );
  OAI211_X1 U23115 ( .C1(n21168), .C2(n20971), .A(n21808), .B(n20970), .ZN(
        n20972) );
  AOI211_X1 U23116 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20973), .B(n20972), .ZN(n20983) );
  NAND3_X1 U23117 ( .A1(n20975), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n20974), .ZN(n20977) );
  OAI21_X1 U23118 ( .B1(n20976), .B2(n20977), .A(n21018), .ZN(n20989) );
  INV_X1 U23119 ( .A(n20989), .ZN(n20980) );
  AOI21_X1 U23120 ( .B1(n20981), .B2(n20977), .A(n21882), .ZN(n20978) );
  OAI22_X1 U23121 ( .A1(n20981), .A2(n20980), .B1(n20979), .B2(n20978), .ZN(
        n20982) );
  OAI211_X1 U23122 ( .C1(n20987), .C2(n20986), .A(n20983), .B(n20982), .ZN(
        P3_U2656) );
  AOI211_X1 U23123 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20984), .A(n21004), .B(
        n21160), .ZN(n20985) );
  AOI211_X1 U23124 ( .C1(n21186), .C2(P3_EBX_REG_16__SCAN_IN), .A(n21832), .B(
        n20985), .ZN(n20996) );
  NOR2_X1 U23125 ( .A1(n20986), .A2(n21052), .ZN(n20994) );
  OAI21_X1 U23126 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n21052), .A(n20987), 
        .ZN(n20992) );
  OAI21_X1 U23127 ( .B1(n20990), .B2(n20989), .A(n21157), .ZN(n20988) );
  AOI21_X1 U23128 ( .B1(n20990), .B2(n20989), .A(n20988), .ZN(n20991) );
  AOI221_X1 U23129 ( .B1(n20994), .B2(n20993), .C1(n20992), .C2(
        P3_REIP_REG_16__SCAN_IN), .A(n20991), .ZN(n20995) );
  OAI211_X1 U23130 ( .C1(n20997), .C2(n21170), .A(n20996), .B(n20995), .ZN(
        P3_U2655) );
  NAND3_X1 U23131 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n21049), .ZN(n21011) );
  OAI21_X1 U23132 ( .B1(n20999), .B2(n20998), .A(n21183), .ZN(n21040) );
  AOI21_X1 U23133 ( .B1(n21000), .B2(n21013), .A(n21151), .ZN(n21002) );
  OAI21_X1 U23134 ( .B1(n21003), .B2(n21002), .A(n21157), .ZN(n21001) );
  AOI21_X1 U23135 ( .B1(n21003), .B2(n21002), .A(n21001), .ZN(n21008) );
  OAI211_X1 U23136 ( .C1(n21004), .C2(n21006), .A(n21185), .B(n21019), .ZN(
        n21005) );
  OAI211_X1 U23137 ( .C1(n21168), .C2(n21006), .A(n21808), .B(n21005), .ZN(
        n21007) );
  AOI211_X1 U23138 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n21008), .B(n21007), .ZN(n21009) );
  OAI221_X1 U23139 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n21011), .C1(n21010), 
        .C2(n21040), .A(n21009), .ZN(P3_U2654) );
  AOI21_X1 U23140 ( .B1(n21014), .B2(n21013), .A(n21012), .ZN(n21017) );
  NOR2_X1 U23141 ( .A1(n11293), .A2(n21015), .ZN(n21016) );
  AOI211_X1 U23142 ( .C1(n21018), .C2(n21017), .A(n21016), .B(n21882), .ZN(
        n21023) );
  AOI211_X1 U23143 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n21019), .A(n21030), .B(
        n21160), .ZN(n21022) );
  AOI22_X1 U23144 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n21092), .B1(
        n21186), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n21020) );
  INV_X1 U23145 ( .A(n21020), .ZN(n21021) );
  NOR4_X1 U23146 ( .A1(n21832), .A2(n21023), .A3(n21022), .A4(n21021), .ZN(
        n21024) );
  OAI221_X1 U23147 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n21026), .C1(n21025), 
        .C2(n21040), .A(n21024), .ZN(P3_U2653) );
  AOI211_X1 U23148 ( .C1(n21028), .C2(n11293), .A(n21027), .B(n21882), .ZN(
        n21034) );
  OAI211_X1 U23149 ( .C1(n21030), .C2(n21032), .A(n21185), .B(n21029), .ZN(
        n21031) );
  OAI211_X1 U23150 ( .C1(n21168), .C2(n21032), .A(n21808), .B(n21031), .ZN(
        n21033) );
  AOI211_X1 U23151 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21034), .B(n21033), .ZN(n21038) );
  OAI211_X1 U23152 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n21036), .B(n21035), .ZN(n21037) );
  OAI211_X1 U23153 ( .C1(n21040), .C2(n21039), .A(n21038), .B(n21037), .ZN(
        P3_U2652) );
  AOI211_X1 U23154 ( .C1(n21043), .C2(n21042), .A(n21041), .B(n21882), .ZN(
        n21048) );
  OAI211_X1 U23155 ( .C1(n21044), .C2(n21046), .A(n21185), .B(n21057), .ZN(
        n21045) );
  OAI21_X1 U23156 ( .B1(n21046), .B2(n21168), .A(n21045), .ZN(n21047) );
  AOI211_X1 U23157 ( .C1(n21092), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n21048), .B(n21047), .ZN(n21051) );
  NAND3_X1 U23158 ( .A1(n21050), .A2(n21049), .A3(n21445), .ZN(n21065) );
  OAI211_X1 U23159 ( .C1(n21445), .C2(n21064), .A(n21051), .B(n21065), .ZN(
        P3_U2650) );
  NOR3_X1 U23160 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n21053), .A3(n21052), 
        .ZN(n21062) );
  AOI211_X1 U23161 ( .C1(n21056), .C2(n21055), .A(n21054), .B(n21882), .ZN(
        n21061) );
  AOI211_X1 U23162 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21057), .A(n21077), .B(
        n21160), .ZN(n21060) );
  AOI22_X1 U23163 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21092), .B1(
        n21186), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n21058) );
  INV_X1 U23164 ( .A(n21058), .ZN(n21059) );
  NOR4_X1 U23165 ( .A1(n21062), .A2(n21061), .A3(n21060), .A4(n21059), .ZN(
        n21063) );
  OAI221_X1 U23166 ( .B1(n21066), .B2(n21065), .C1(n21066), .C2(n21064), .A(
        n21063), .ZN(P3_U2649) );
  NAND2_X1 U23167 ( .A1(n21068), .A2(n21067), .ZN(n21080) );
  INV_X1 U23168 ( .A(n21069), .ZN(n21082) );
  OAI21_X1 U23169 ( .B1(n21082), .B2(n21081), .A(n21184), .ZN(n21097) );
  AOI211_X1 U23170 ( .C1(n21072), .C2(n21071), .A(n21070), .B(n21882), .ZN(
        n21075) );
  OAI22_X1 U23171 ( .A1(n21073), .A2(n21170), .B1(n21168), .B2(n21076), .ZN(
        n21074) );
  AOI211_X1 U23172 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n21097), .A(n21075), 
        .B(n21074), .ZN(n21079) );
  OAI211_X1 U23173 ( .C1(n21077), .C2(n21076), .A(n21185), .B(n21083), .ZN(
        n21078) );
  OAI211_X1 U23174 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n21080), .A(n21079), 
        .B(n21078), .ZN(P3_U2648) );
  NOR2_X1 U23175 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21081), .ZN(n21098) );
  AOI22_X1 U23176 ( .A1(n21186), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n21082), 
        .B2(n21098), .ZN(n21090) );
  AOI211_X1 U23177 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n21083), .A(n21100), .B(
        n21160), .ZN(n21088) );
  AOI211_X1 U23178 ( .C1(n21086), .C2(n21085), .A(n21084), .B(n21882), .ZN(
        n21087) );
  AOI211_X1 U23179 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n21097), .A(n21088), 
        .B(n21087), .ZN(n21089) );
  OAI211_X1 U23180 ( .C1(n21091), .C2(n21170), .A(n21090), .B(n21089), .ZN(
        P3_U2647) );
  AOI22_X1 U23181 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21092), .B1(
        n21186), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n21107) );
  AOI211_X1 U23182 ( .C1(n21095), .C2(n21094), .A(n21093), .B(n21882), .ZN(
        n21096) );
  AOI221_X1 U23183 ( .B1(n21098), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n21097), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n21096), .ZN(n21106) );
  OAI211_X1 U23184 ( .C1(n21100), .C2(n21099), .A(n21185), .B(n21110), .ZN(
        n21105) );
  NAND3_X1 U23185 ( .A1(n21103), .A2(n21102), .A3(n21101), .ZN(n21104) );
  NAND4_X1 U23186 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        P3_U2646) );
  INV_X1 U23187 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U23188 ( .A1(n21186), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n21109), 
        .B2(n21108), .ZN(n21118) );
  AOI211_X1 U23189 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21110), .A(n21130), .B(
        n21160), .ZN(n21115) );
  AOI211_X1 U23190 ( .C1(n21113), .C2(n21112), .A(n21111), .B(n21882), .ZN(
        n21114) );
  AOI211_X1 U23191 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n21116), .A(n21115), 
        .B(n21114), .ZN(n21117) );
  OAI211_X1 U23192 ( .C1(n21119), .C2(n21170), .A(n21118), .B(n21117), .ZN(
        P3_U2645) );
  AOI211_X1 U23193 ( .C1(n21122), .C2(n21121), .A(n21120), .B(n21882), .ZN(
        n21127) );
  OAI22_X1 U23194 ( .A1(n21125), .A2(n21170), .B1(n21124), .B2(n21123), .ZN(
        n21126) );
  AOI211_X1 U23195 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n21186), .A(n21127), .B(
        n21126), .ZN(n21132) );
  OAI211_X1 U23196 ( .C1(n21130), .C2(n21129), .A(n21185), .B(n21128), .ZN(
        n21131) );
  OAI211_X1 U23197 ( .C1(n21134), .C2(n21133), .A(n21132), .B(n21131), .ZN(
        P3_U2644) );
  NOR2_X1 U23198 ( .A1(n21136), .A2(n21135), .ZN(n21153) );
  AOI22_X1 U23199 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n21186), .B1(n21153), 
        .B2(n21661), .ZN(n21149) );
  INV_X1 U23200 ( .A(n21137), .ZN(n21139) );
  NAND2_X1 U23201 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n21138) );
  OAI21_X1 U23202 ( .B1(n21139), .B2(n21138), .A(n21183), .ZN(n21154) );
  INV_X1 U23203 ( .A(n21154), .ZN(n21176) );
  INV_X1 U23204 ( .A(n21141), .ZN(n21142) );
  NAND2_X1 U23205 ( .A1(n21141), .A2(n21140), .ZN(n21159) );
  NAND2_X1 U23206 ( .A1(n21185), .A2(n21159), .ZN(n21163) );
  AOI21_X1 U23207 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21142), .A(n21163), .ZN(
        n21147) );
  NOR2_X1 U23208 ( .A1(n21143), .A2(n21151), .ZN(n21144) );
  AOI211_X1 U23209 ( .C1(n21145), .C2(n21144), .A(n21152), .B(n21882), .ZN(
        n21146) );
  OAI211_X1 U23210 ( .C1(n21150), .C2(n21170), .A(n21149), .B(n21148), .ZN(
        P3_U2642) );
  XOR2_X1 U23211 ( .A(n21164), .B(n21165), .Z(n21158) );
  NAND2_X1 U23212 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21153), .ZN(n21166) );
  NOR2_X1 U23213 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21166), .ZN(n21177) );
  OAI22_X1 U23214 ( .A1(n21155), .A2(n21170), .B1(n21167), .B2(n21154), .ZN(
        n21156) );
  NOR2_X1 U23215 ( .A1(n21160), .A2(n21159), .ZN(n21175) );
  OAI21_X1 U23216 ( .B1(n21186), .B2(n21175), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n21161) );
  OAI211_X1 U23217 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n21163), .A(n21162), .B(
        n21161), .ZN(P3_U2641) );
  NAND2_X1 U23218 ( .A1(n21165), .A2(n21164), .ZN(n21181) );
  INV_X1 U23219 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21174) );
  NOR3_X1 U23220 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21167), .A3(n21166), 
        .ZN(n21173) );
  OAI22_X1 U23221 ( .A1(n21171), .A2(n21170), .B1(n21169), .B2(n21168), .ZN(
        n21172) );
  AOI211_X1 U23222 ( .C1(n21175), .C2(n21174), .A(n21173), .B(n21172), .ZN(
        n21179) );
  OAI21_X1 U23223 ( .B1(n21177), .B2(n21176), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n21178) );
  OAI211_X1 U23224 ( .C1(n21181), .C2(n21180), .A(n21179), .B(n21178), .ZN(
        P3_U2640) );
  AOI22_X1 U23225 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n21183), .B1(n21182), 
        .B2(n21403), .ZN(n21189) );
  NAND3_X1 U23226 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21184), .A3(
        n21423), .ZN(n21188) );
  OAI21_X1 U23227 ( .B1(n21186), .B2(n21185), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n21187) );
  NAND3_X1 U23228 ( .A1(n21189), .A2(n21188), .A3(n21187), .ZN(P3_U2671) );
  NAND2_X1 U23229 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n21249) );
  NAND4_X1 U23230 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n21190) );
  NOR3_X1 U23231 ( .A1(n21376), .A2(n21369), .A3(n21190), .ZN(n21191) );
  NAND3_X1 U23232 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(n21191), .ZN(n21247) );
  NAND2_X1 U23233 ( .A1(n21366), .A2(n21375), .ZN(n21377) );
  NOR2_X1 U23234 ( .A1(n21247), .A2(n21377), .ZN(n21357) );
  NAND2_X1 U23235 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21357), .ZN(n21213) );
  NOR2_X1 U23236 ( .A1(n21248), .A2(n21213), .ZN(n21217) );
  NAND2_X1 U23237 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21217), .ZN(n21210) );
  NOR2_X1 U23238 ( .A1(n21249), .A2(n21210), .ZN(n21344) );
  INV_X1 U23239 ( .A(n21344), .ZN(n21199) );
  NAND3_X1 U23240 ( .A1(n21353), .A2(P3_EAX_REG_13__SCAN_IN), .A3(n21199), 
        .ZN(n21198) );
  NAND2_X1 U23241 ( .A1(n21195), .A2(n21375), .ZN(n21245) );
  AOI22_X1 U23242 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21373), .B1(n21372), .B2(
        n21196), .ZN(n21197) );
  OAI211_X1 U23243 ( .C1(P3_EAX_REG_13__SCAN_IN), .C2(n21199), .A(n21198), .B(
        n21197), .ZN(P3_U2722) );
  INV_X1 U23244 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21202) );
  INV_X1 U23245 ( .A(n21210), .ZN(n21204) );
  AOI22_X1 U23246 ( .A1(n21204), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n21353), .ZN(n21201) );
  OAI222_X1 U23247 ( .A1(n21245), .A2(n21202), .B1(n21344), .B2(n21201), .C1(
        n21363), .C2(n21200), .ZN(P3_U2723) );
  INV_X1 U23248 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21208) );
  NOR2_X1 U23249 ( .A1(n21203), .A2(n21210), .ZN(n21207) );
  AOI21_X1 U23250 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n21353), .A(n21204), .ZN(
        n21206) );
  OAI222_X1 U23251 ( .A1(n21245), .A2(n21208), .B1(n21207), .B2(n21206), .C1(
        n21363), .C2(n21205), .ZN(P3_U2724) );
  AOI22_X1 U23252 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21373), .B1(n21372), .B2(
        n21209), .ZN(n21212) );
  OAI211_X1 U23253 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21217), .A(n21353), .B(
        n21210), .ZN(n21211) );
  NAND2_X1 U23254 ( .A1(n21212), .A2(n21211), .ZN(P3_U2725) );
  INV_X1 U23255 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21218) );
  OAI21_X1 U23256 ( .B1(n21248), .B2(n21359), .A(n21213), .ZN(n21214) );
  INV_X1 U23257 ( .A(n21214), .ZN(n21216) );
  OAI222_X1 U23258 ( .A1(n21245), .A2(n21218), .B1(n21217), .B2(n21216), .C1(
        n21363), .C2(n21215), .ZN(P3_U2726) );
  NOR4_X1 U23259 ( .A1(n21376), .A2(n21369), .A3(n21219), .A4(n21377), .ZN(
        n21244) );
  NAND2_X1 U23260 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21244), .ZN(n21232) );
  NOR2_X1 U23261 ( .A1(n21220), .A2(n21232), .ZN(n21235) );
  NAND2_X1 U23262 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21235), .ZN(n21224) );
  NOR2_X1 U23263 ( .A1(n21221), .A2(n21224), .ZN(n21227) );
  AOI21_X1 U23264 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21353), .A(n21227), .ZN(
        n21222) );
  OAI222_X1 U23265 ( .A1(n21223), .A2(n21245), .B1(n21357), .B2(n21222), .C1(
        n21363), .C2(n21439), .ZN(P3_U2728) );
  INV_X1 U23266 ( .A(n21224), .ZN(n21230) );
  AOI21_X1 U23267 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21353), .A(n21230), .ZN(
        n21226) );
  OAI222_X1 U23268 ( .A1(n21271), .A2(n21245), .B1(n21227), .B2(n21226), .C1(
        n21363), .C2(n21225), .ZN(P3_U2729) );
  AOI21_X1 U23269 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21353), .A(n21235), .ZN(
        n21229) );
  OAI222_X1 U23270 ( .A1(n21231), .A2(n21245), .B1(n21230), .B2(n21229), .C1(
        n21363), .C2(n21228), .ZN(P3_U2730) );
  INV_X1 U23271 ( .A(n21232), .ZN(n21239) );
  AOI21_X1 U23272 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21353), .A(n21239), .ZN(
        n21234) );
  OAI222_X1 U23273 ( .A1(n21236), .A2(n21245), .B1(n21235), .B2(n21234), .C1(
        n21363), .C2(n21233), .ZN(P3_U2731) );
  AOI21_X1 U23274 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21353), .A(n21244), .ZN(
        n21238) );
  OAI222_X1 U23275 ( .A1(n21240), .A2(n21245), .B1(n21239), .B2(n21238), .C1(
        n21363), .C2(n21237), .ZN(P3_U2732) );
  NOR3_X1 U23276 ( .A1(n21376), .A2(n21369), .A3(n21377), .ZN(n21241) );
  AOI21_X1 U23277 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21353), .A(n21241), .ZN(
        n21243) );
  OAI222_X1 U23278 ( .A1(n21246), .A2(n21245), .B1(n21244), .B2(n21243), .C1(
        n21363), .C2(n21242), .ZN(P3_U2733) );
  NOR4_X1 U23279 ( .A1(n21360), .A2(n21348), .A3(n21249), .A4(n21248), .ZN(
        n21250) );
  NOR3_X1 U23280 ( .A1(n21290), .A2(n21340), .A3(n21251), .ZN(n21282) );
  NAND2_X1 U23281 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n21282), .ZN(n21278) );
  NOR2_X1 U23282 ( .A1(n21273), .A2(n21278), .ZN(n21272) );
  NAND2_X1 U23283 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21272), .ZN(n21259) );
  NAND2_X1 U23284 ( .A1(n21353), .A2(n21259), .ZN(n21264) );
  NAND2_X1 U23285 ( .A1(n21252), .A2(n21359), .ZN(n21332) );
  INV_X1 U23286 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21254) );
  NOR2_X2 U23287 ( .A1(n21253), .A2(n21353), .ZN(n21338) );
  INV_X1 U23288 ( .A(n21338), .ZN(n21320) );
  OAI22_X1 U23289 ( .A1(n21255), .A2(n21363), .B1(n21254), .B2(n21320), .ZN(
        n21256) );
  AOI21_X1 U23290 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21339), .A(n21256), .ZN(
        n21257) );
  OAI221_X1 U23291 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21259), .C1(n21258), 
        .C2(n21264), .A(n21257), .ZN(P3_U2714) );
  AOI22_X1 U23292 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n21338), .B1(n21372), .B2(
        n21260), .ZN(n21262) );
  AOI22_X1 U23293 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21339), .B1(n21272), .B2(
        n21263), .ZN(n21261) );
  OAI211_X1 U23294 ( .C1(n21263), .C2(n21264), .A(n21262), .B(n21261), .ZN(
        P3_U2715) );
  OAI21_X1 U23295 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21377), .A(n21264), .ZN(
        n21269) );
  NAND3_X1 U23296 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .ZN(n21289) );
  NOR3_X1 U23297 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n21289), .A3(n21278), .ZN(
        n21268) );
  OAI22_X1 U23298 ( .A1(n21266), .A2(n21363), .B1(n21265), .B2(n21320), .ZN(
        n21267) );
  AOI211_X1 U23299 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n21269), .A(n21268), .B(
        n21267), .ZN(n21270) );
  OAI21_X1 U23300 ( .B1(n21271), .B2(n21332), .A(n21270), .ZN(P3_U2713) );
  AOI22_X1 U23301 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21338), .ZN(n21276) );
  AOI211_X1 U23302 ( .C1(n21273), .C2(n21278), .A(n21272), .B(n21359), .ZN(
        n21274) );
  INV_X1 U23303 ( .A(n21274), .ZN(n21275) );
  OAI211_X1 U23304 ( .C1(n21277), .C2(n21363), .A(n21276), .B(n21275), .ZN(
        P3_U2716) );
  AOI22_X1 U23305 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21338), .ZN(n21280) );
  OAI211_X1 U23306 ( .C1(n21282), .C2(P3_EAX_REG_18__SCAN_IN), .A(n21353), .B(
        n21278), .ZN(n21279) );
  OAI211_X1 U23307 ( .C1(n21281), .C2(n21363), .A(n21280), .B(n21279), .ZN(
        P3_U2717) );
  AOI22_X1 U23308 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21338), .ZN(n21286) );
  INV_X1 U23309 ( .A(n21340), .ZN(n21284) );
  INV_X1 U23310 ( .A(n21282), .ZN(n21283) );
  OAI211_X1 U23311 ( .C1(n21284), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21353), .B(
        n21283), .ZN(n21285) );
  OAI211_X1 U23312 ( .C1(n21287), .C2(n21363), .A(n21286), .B(n21285), .ZN(
        P3_U2718) );
  AOI22_X1 U23313 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21338), .ZN(n21293) );
  NAND3_X1 U23314 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n21288) );
  NAND2_X1 U23315 ( .A1(n21334), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21333) );
  NAND2_X1 U23316 ( .A1(n21328), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21327) );
  OAI211_X1 U23317 ( .C1(n21291), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21353), .B(
        n21296), .ZN(n21292) );
  OAI211_X1 U23318 ( .C1(n21294), .C2(n21363), .A(n21293), .B(n21292), .ZN(
        P3_U2710) );
  INV_X1 U23319 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n21301) );
  AOI22_X1 U23320 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n21338), .B1(n21372), .B2(
        n21295), .ZN(n21300) );
  AOI211_X1 U23321 ( .C1(n21297), .C2(n21296), .A(n21322), .B(n21359), .ZN(
        n21298) );
  INV_X1 U23322 ( .A(n21298), .ZN(n21299) );
  OAI211_X1 U23323 ( .C1(n21332), .C2(n21301), .A(n21300), .B(n21299), .ZN(
        P3_U2709) );
  NAND2_X1 U23324 ( .A1(n21322), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21321) );
  NAND2_X1 U23325 ( .A1(n21308), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21304) );
  NAND3_X1 U23326 ( .A1(n21353), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n21304), 
        .ZN(n21303) );
  NAND2_X1 U23327 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21338), .ZN(n21302) );
  OAI211_X1 U23328 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n21304), .A(n21303), .B(
        n21302), .ZN(P3_U2704) );
  AOI22_X1 U23329 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n21338), .ZN(n21306) );
  OAI211_X1 U23330 ( .C1(n21308), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21353), .B(
        n21304), .ZN(n21305) );
  OAI211_X1 U23331 ( .C1(n21307), .C2(n21363), .A(n21306), .B(n21305), .ZN(
        P3_U2705) );
  AOI22_X1 U23332 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21338), .ZN(n21312) );
  AOI211_X1 U23333 ( .C1(n21309), .C2(n21315), .A(n21308), .B(n21359), .ZN(
        n21310) );
  INV_X1 U23334 ( .A(n21310), .ZN(n21311) );
  OAI211_X1 U23335 ( .C1(n21313), .C2(n21363), .A(n21312), .B(n21311), .ZN(
        P3_U2706) );
  INV_X1 U23336 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21319) );
  AOI22_X1 U23337 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21339), .B1(n21372), .B2(
        n21314), .ZN(n21318) );
  OAI211_X1 U23338 ( .C1(n21316), .C2(P3_EAX_REG_28__SCAN_IN), .A(n21353), .B(
        n21315), .ZN(n21317) );
  OAI211_X1 U23339 ( .C1(n21320), .C2(n21319), .A(n21318), .B(n21317), .ZN(
        P3_U2707) );
  AOI22_X1 U23340 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21338), .ZN(n21324) );
  OAI211_X1 U23341 ( .C1(n21322), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21353), .B(
        n21321), .ZN(n21323) );
  OAI211_X1 U23342 ( .C1(n21325), .C2(n21363), .A(n21324), .B(n21323), .ZN(
        P3_U2708) );
  INV_X1 U23343 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21331) );
  AOI22_X1 U23344 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n21338), .B1(n21372), .B2(
        n21326), .ZN(n21330) );
  OAI211_X1 U23345 ( .C1(n21328), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21353), .B(
        n21327), .ZN(n21329) );
  OAI211_X1 U23346 ( .C1(n21332), .C2(n21331), .A(n21330), .B(n21329), .ZN(
        P3_U2711) );
  AOI22_X1 U23347 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21338), .ZN(n21336) );
  OAI211_X1 U23348 ( .C1(n21334), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21353), .B(
        n21333), .ZN(n21335) );
  OAI211_X1 U23349 ( .C1(n21337), .C2(n21363), .A(n21336), .B(n21335), .ZN(
        P3_U2712) );
  AOI22_X1 U23350 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21339), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21338), .ZN(n21342) );
  OAI211_X1 U23351 ( .C1(n21350), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21353), .B(
        n21340), .ZN(n21341) );
  OAI211_X1 U23352 ( .C1(n21343), .C2(n21363), .A(n21342), .B(n21341), .ZN(
        P3_U2719) );
  NAND2_X1 U23353 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21344), .ZN(n21349) );
  NAND2_X1 U23354 ( .A1(n21353), .A2(n21352), .ZN(n21347) );
  AOI22_X1 U23355 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21373), .B1(n21372), .B2(
        n21345), .ZN(n21346) );
  OAI221_X1 U23356 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n21349), .C1(n21348), 
        .C2(n21347), .A(n21346), .ZN(P3_U2721) );
  AOI21_X1 U23357 ( .B1(n21352), .B2(n21351), .A(n21350), .ZN(n21354) );
  AOI22_X1 U23358 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n21373), .B1(n21354), .B2(
        n21353), .ZN(n21355) );
  OAI21_X1 U23359 ( .B1(n21356), .B2(n21363), .A(n21355), .ZN(P3_U2720) );
  AOI22_X1 U23360 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21373), .B1(n21357), .B2(
        n21360), .ZN(n21362) );
  OR3_X1 U23361 ( .A1(n21360), .A2(n21359), .A3(n21358), .ZN(n21361) );
  OAI211_X1 U23362 ( .C1(n21364), .C2(n21363), .A(n21362), .B(n21361), .ZN(
        P3_U2727) );
  OR2_X1 U23363 ( .A1(n21376), .A2(n21377), .ZN(n21370) );
  AOI21_X1 U23364 ( .B1(n21366), .B2(n21376), .A(n21365), .ZN(n21368) );
  AOI22_X1 U23365 ( .A1(n21373), .A2(BUF2_REG_1__SCAN_IN), .B1(n21372), .B2(
        n15581), .ZN(n21367) );
  OAI221_X1 U23366 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n21370), .C1(n21369), 
        .C2(n21368), .A(n21367), .ZN(P3_U2734) );
  AOI22_X1 U23367 ( .A1(n21373), .A2(BUF2_REG_0__SCAN_IN), .B1(n21372), .B2(
        n21371), .ZN(n21374) );
  OAI221_X1 U23368 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21377), .C1(n21376), 
        .C2(n21375), .A(n21374), .ZN(P3_U2735) );
  INV_X1 U23369 ( .A(n21424), .ZN(n21386) );
  NOR2_X1 U23370 ( .A1(n21378), .A2(n21818), .ZN(n21380) );
  AOI22_X1 U23371 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21822), .B1(
        n21380), .B2(n21403), .ZN(n21856) );
  INV_X1 U23372 ( .A(n21423), .ZN(n21384) );
  AOI222_X1 U23373 ( .A1(n21522), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21856), 
        .B2(n21384), .C1(n21403), .C2(n21887), .ZN(n21379) );
  AOI22_X1 U23374 ( .A1(n21386), .A2(n21403), .B1(n21379), .B2(n21424), .ZN(
        P3_U3290) );
  OAI21_X1 U23375 ( .B1(n21805), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21816), .ZN(n21402) );
  OAI22_X1 U23376 ( .A1(n21380), .A2(n21381), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21402), .ZN(n21854) );
  INV_X1 U23377 ( .A(n21381), .ZN(n21383) );
  AOI22_X1 U23378 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21674), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21462), .ZN(n21397) );
  NAND2_X1 U23379 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21398) );
  INV_X1 U23380 ( .A(n21398), .ZN(n21382) );
  AOI222_X1 U23381 ( .A1(n21854), .A2(n21384), .B1(n21383), .B2(n21887), .C1(
        n21397), .C2(n21382), .ZN(n21385) );
  AOI22_X1 U23382 ( .A1(n21386), .A2(n21392), .B1(n21385), .B2(n21424), .ZN(
        P3_U3289) );
  AOI22_X1 U23383 ( .A1(n21390), .A2(n21389), .B1(n21388), .B2(n21387), .ZN(
        n21416) );
  AOI211_X1 U23384 ( .C1(n21410), .C2(n21416), .A(n21406), .B(n21851), .ZN(
        n21394) );
  AOI211_X1 U23385 ( .C1(n21851), .C2(n21392), .A(n21391), .B(n21402), .ZN(
        n21393) );
  AOI211_X1 U23386 ( .C1(n21835), .C2(n21395), .A(n21394), .B(n21393), .ZN(
        n21850) );
  OAI222_X1 U23387 ( .A1(n21398), .A2(n21397), .B1(n21423), .B2(n21850), .C1(
        n21396), .C2(n21421), .ZN(n21399) );
  AOI22_X1 U23388 ( .A1(n21887), .A2(n21400), .B1(n21424), .B2(n21399), .ZN(
        n21401) );
  OAI21_X1 U23389 ( .B1(n21851), .B2(n21424), .A(n21401), .ZN(P3_U3288) );
  NOR2_X1 U23390 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21412), .ZN(
        n21420) );
  INV_X1 U23391 ( .A(n21402), .ZN(n21419) );
  NAND2_X1 U23392 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21403), .ZN(
        n21409) );
  OAI211_X1 U23393 ( .C1(n21406), .C2(n21405), .A(n21835), .B(n21404), .ZN(
        n21407) );
  OAI22_X1 U23394 ( .A1(n21410), .A2(n21409), .B1(n21408), .B2(n21407), .ZN(
        n21418) );
  INV_X1 U23395 ( .A(n21411), .ZN(n21415) );
  NAND2_X1 U23396 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21412), .ZN(
        n21413) );
  OAI22_X1 U23397 ( .A1(n21416), .A2(n21415), .B1(n21414), .B2(n21413), .ZN(
        n21417) );
  AOI211_X1 U23398 ( .C1(n21420), .C2(n21419), .A(n21418), .B(n21417), .ZN(
        n21847) );
  OAI22_X1 U23399 ( .A1(n21847), .A2(n21423), .B1(n21422), .B2(n21421), .ZN(
        n21425) );
  MUX2_X1 U23400 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21425), .S(
        n21424), .Z(P3_U3285) );
  INV_X1 U23401 ( .A(n21818), .ZN(n21601) );
  NOR3_X1 U23402 ( .A1(n21480), .A2(n21481), .A3(n21426), .ZN(n21493) );
  NAND2_X1 U23403 ( .A1(n21427), .A2(n21493), .ZN(n21485) );
  OR2_X1 U23404 ( .A1(n21492), .A2(n21485), .ZN(n21503) );
  NOR2_X1 U23405 ( .A1(n21431), .A2(n21503), .ZN(n21821) );
  NAND2_X1 U23406 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21821), .ZN(
        n21804) );
  NOR2_X1 U23407 ( .A1(n21755), .A2(n21804), .ZN(n21753) );
  INV_X1 U23408 ( .A(n21753), .ZN(n21432) );
  NOR2_X1 U23409 ( .A1(n21428), .A2(n21432), .ZN(n21440) );
  INV_X1 U23410 ( .A(n21440), .ZN(n21585) );
  AOI211_X1 U23411 ( .C1(n21818), .C2(n21585), .A(n21763), .B(n21685), .ZN(
        n21734) );
  NAND2_X1 U23412 ( .A1(n21751), .A2(n21429), .ZN(n21441) );
  NAND2_X1 U23413 ( .A1(n21493), .A2(n21430), .ZN(n21486) );
  OR2_X1 U23414 ( .A1(n21492), .A2(n21486), .ZN(n21505) );
  OR3_X1 U23415 ( .A1(n21817), .A2(n21431), .A3(n21505), .ZN(n21754) );
  NOR2_X1 U23416 ( .A1(n21441), .A2(n21754), .ZN(n21599) );
  OAI21_X1 U23417 ( .B1(n21432), .B2(n21731), .A(n21805), .ZN(n21433) );
  OAI21_X1 U23418 ( .B1(n21599), .B2(n21756), .A(n21433), .ZN(n21738) );
  NOR2_X1 U23419 ( .A1(n21835), .A2(n21805), .ZN(n21807) );
  NAND2_X1 U23420 ( .A1(n21483), .A2(n21439), .ZN(n21735) );
  OAI22_X1 U23421 ( .A1(n21437), .A2(n21807), .B1(n21434), .B2(n21735), .ZN(
        n21435) );
  AOI211_X1 U23422 ( .C1(n21834), .C2(n21436), .A(n21738), .B(n21435), .ZN(
        n21586) );
  OAI211_X1 U23423 ( .C1(n21601), .C2(n21437), .A(n21734), .B(n21586), .ZN(
        n21438) );
  NAND2_X1 U23424 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21438), .ZN(
        n21446) );
  NOR2_X1 U23425 ( .A1(n21439), .A2(n21841), .ZN(n21688) );
  AOI22_X1 U23426 ( .A1(n21834), .A2(n21520), .B1(n21700), .B2(n21521), .ZN(
        n21544) );
  AOI22_X1 U23427 ( .A1(n21835), .A2(n21599), .B1(n21654), .B2(n21440), .ZN(
        n21597) );
  OAI21_X1 U23428 ( .B1(n21544), .B2(n21441), .A(n21597), .ZN(n21587) );
  NAND2_X1 U23429 ( .A1(n21587), .A2(n21773), .ZN(n21749) );
  INV_X1 U23430 ( .A(n21749), .ZN(n21724) );
  AOI22_X1 U23431 ( .A1(n21828), .A2(n21443), .B1(n21724), .B2(n21442), .ZN(
        n21444) );
  OAI221_X1 U23432 ( .B1(n21832), .B2(n21446), .C1(n21808), .C2(n21445), .A(
        n21444), .ZN(P3_U2841) );
  NOR2_X1 U23433 ( .A1(n21835), .A2(n21818), .ZN(n21744) );
  OAI221_X1 U23434 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21744), .C1(
        n21522), .C2(n21822), .A(n21447), .ZN(n21448) );
  AOI22_X1 U23435 ( .A1(n21801), .A2(P3_REIP_REG_0__SCAN_IN), .B1(n21773), 
        .B2(n21448), .ZN(n21449) );
  OAI21_X1 U23436 ( .B1(n21522), .B2(n21793), .A(n21449), .ZN(P3_U2862) );
  NAND2_X1 U23437 ( .A1(n21832), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21458) );
  NOR2_X1 U23438 ( .A1(n21783), .A2(n21450), .ZN(n21452) );
  NOR2_X1 U23439 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21744), .ZN(
        n21451) );
  MUX2_X1 U23440 ( .A(n21452), .B(n21451), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21456) );
  OAI22_X1 U23441 ( .A1(n21454), .A2(n21695), .B1(n21841), .B2(n21453), .ZN(
        n21455) );
  OAI21_X1 U23442 ( .B1(n21456), .B2(n21455), .A(n21668), .ZN(n21457) );
  OAI211_X1 U23443 ( .C1(n21793), .C2(n21462), .A(n21458), .B(n21457), .ZN(
        P3_U2861) );
  NAND3_X1 U23444 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21654), .A3(
        n21471), .ZN(n21459) );
  OAI211_X1 U23445 ( .C1(n21841), .C2(n21461), .A(n21460), .B(n21459), .ZN(
        n21468) );
  NOR2_X1 U23446 ( .A1(n21522), .A2(n21462), .ZN(n21464) );
  AOI21_X1 U23447 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21600), .A(
        n21764), .ZN(n21463) );
  AOI21_X1 U23448 ( .B1(n21464), .B2(n21835), .A(n21463), .ZN(n21466) );
  OAI22_X1 U23449 ( .A1(n21466), .A2(n21471), .B1(n21695), .B2(n21465), .ZN(
        n21467) );
  OAI21_X1 U23450 ( .B1(n21468), .B2(n21467), .A(n21668), .ZN(n21469) );
  OAI211_X1 U23451 ( .C1(n21793), .C2(n21471), .A(n21470), .B(n21469), .ZN(
        P3_U2860) );
  NAND2_X1 U23452 ( .A1(n21668), .A2(n21834), .ZN(n21519) );
  AND2_X1 U23453 ( .A1(n21481), .A2(n21496), .ZN(n21473) );
  OAI22_X1 U23454 ( .A1(n21474), .A2(n21473), .B1(n21472), .B2(n21841), .ZN(
        n21475) );
  AOI22_X1 U23455 ( .A1(n21773), .A2(n21475), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21803), .ZN(n21477) );
  OAI211_X1 U23456 ( .C1(n21519), .C2(n21478), .A(n21477), .B(n21476), .ZN(
        P3_U2859) );
  INV_X1 U23457 ( .A(n21479), .ZN(n21484) );
  NOR4_X1 U23458 ( .A1(n21496), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n21481), .A4(n21480), .ZN(n21482) );
  AOI21_X1 U23459 ( .B1(n21484), .B2(n21483), .A(n21482), .ZN(n21491) );
  AOI22_X1 U23460 ( .A1(n21835), .A2(n21486), .B1(n21816), .B2(n21485), .ZN(
        n21487) );
  OAI221_X1 U23461 ( .B1(n21685), .B2(n21487), .C1(n21685), .C2(n21600), .A(
        n21793), .ZN(n21497) );
  INV_X1 U23462 ( .A(n21519), .ZN(n21613) );
  AOI22_X1 U23463 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21497), .B1(
        n21613), .B2(n21488), .ZN(n21490) );
  NAND2_X1 U23464 ( .A1(n21832), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21489) );
  OAI211_X1 U23465 ( .C1(n21491), .C2(n21685), .A(n21490), .B(n21489), .ZN(
        P3_U2857) );
  NAND2_X1 U23466 ( .A1(n21493), .A2(n21492), .ZN(n21495) );
  OAI22_X1 U23467 ( .A1(n21496), .A2(n21495), .B1(n21494), .B2(n21841), .ZN(
        n21498) );
  AOI22_X1 U23468 ( .A1(n21668), .A2(n21498), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21497), .ZN(n21500) );
  OAI211_X1 U23469 ( .C1(n21519), .C2(n21501), .A(n21500), .B(n21499), .ZN(
        P3_U2856) );
  AOI22_X1 U23470 ( .A1(n21835), .A2(n21505), .B1(n21816), .B2(n21503), .ZN(
        n21502) );
  NAND3_X1 U23471 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21502), .A3(
        n21600), .ZN(n21511) );
  INV_X1 U23472 ( .A(n21654), .ZN(n21504) );
  OAI22_X1 U23473 ( .A1(n21756), .A2(n21505), .B1(n21504), .B2(n21503), .ZN(
        n21531) );
  OAI22_X1 U23474 ( .A1(n21695), .A2(n21507), .B1(n21841), .B2(n21506), .ZN(
        n21508) );
  AOI221_X1 U23475 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21511), .C1(
        n21531), .C2(n21511), .A(n21508), .ZN(n21510) );
  AOI22_X1 U23476 ( .A1(n21801), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n21803), 
        .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21509) );
  OAI21_X1 U23477 ( .B1(n21510), .B2(n21685), .A(n21509), .ZN(P3_U2855) );
  AOI22_X1 U23478 ( .A1(n21801), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n21803), 
        .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21517) );
  NAND3_X1 U23479 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21727), .A3(
        n21511), .ZN(n21513) );
  NAND3_X1 U23480 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21817), .A3(
        n21531), .ZN(n21512) );
  OAI211_X1 U23481 ( .C1(n21514), .C2(n21735), .A(n21513), .B(n21512), .ZN(
        n21515) );
  AOI22_X1 U23482 ( .A1(n21668), .A2(n21515), .B1(n21828), .B2(n21514), .ZN(
        n21516) );
  OAI211_X1 U23483 ( .C1(n21519), .C2(n21518), .A(n21517), .B(n21516), .ZN(
        P3_U2854) );
  OAI22_X1 U23484 ( .A1(n21521), .A2(n21735), .B1(n21695), .B2(n21520), .ZN(
        n21802) );
  INV_X1 U23485 ( .A(n21802), .ZN(n21529) );
  NOR2_X1 U23486 ( .A1(n21834), .A2(n21700), .ZN(n21757) );
  OR2_X1 U23487 ( .A1(n21522), .A2(n21804), .ZN(n21815) );
  OAI21_X1 U23488 ( .B1(n21825), .B2(n21815), .A(n21818), .ZN(n21523) );
  NAND2_X1 U23489 ( .A1(n21754), .A2(n21835), .ZN(n21537) );
  OAI211_X1 U23490 ( .C1(n21524), .C2(n21757), .A(n21523), .B(n21537), .ZN(
        n21810) );
  INV_X1 U23491 ( .A(n21810), .ZN(n21528) );
  NOR2_X1 U23492 ( .A1(n21546), .A2(n21756), .ZN(n21554) );
  AOI221_X1 U23493 ( .B1(n21525), .B2(n21805), .C1(n21804), .C2(n21805), .A(
        n21554), .ZN(n21539) );
  OAI211_X1 U23494 ( .C1(n21601), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21668), .B(n21539), .ZN(n21526) );
  INV_X1 U23495 ( .A(n21526), .ZN(n21527) );
  NAND3_X1 U23496 ( .A1(n21529), .A2(n21528), .A3(n21527), .ZN(n21530) );
  NAND2_X1 U23497 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21530), .ZN(
        n21536) );
  NAND3_X1 U23498 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n21531), .ZN(n21571) );
  AOI21_X1 U23499 ( .B1(n21544), .B2(n21571), .A(n21685), .ZN(n21826) );
  AOI22_X1 U23500 ( .A1(n21828), .A2(n21533), .B1(n21826), .B2(n21532), .ZN(
        n21534) );
  OAI221_X1 U23501 ( .B1(n21832), .B2(n21536), .C1(n21808), .C2(n21535), .A(
        n21534), .ZN(P3_U2851) );
  INV_X1 U23502 ( .A(n21537), .ZN(n21824) );
  INV_X1 U23503 ( .A(n21538), .ZN(n21540) );
  OAI21_X1 U23504 ( .B1(n21540), .B2(n21695), .A(n21539), .ZN(n21541) );
  AOI211_X1 U23505 ( .C1(n21700), .C2(n21542), .A(n21824), .B(n21541), .ZN(
        n21794) );
  AOI211_X1 U23506 ( .C1(n21805), .C2(n21791), .A(n21818), .B(n21790), .ZN(
        n21548) );
  NOR2_X1 U23507 ( .A1(n21543), .A2(n21815), .ZN(n21553) );
  NAND2_X1 U23508 ( .A1(n21544), .A2(n21571), .ZN(n21545) );
  AOI21_X1 U23509 ( .B1(n21546), .B2(n21545), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21547) );
  AOI211_X1 U23510 ( .C1(n21794), .C2(n21548), .A(n21553), .B(n21547), .ZN(
        n21549) );
  AOI22_X1 U23511 ( .A1(n21773), .A2(n21549), .B1(n21803), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21551) );
  OAI211_X1 U23512 ( .C1(n21552), .C2(n21813), .A(n21551), .B(n21550), .ZN(
        P3_U2850) );
  AOI22_X1 U23513 ( .A1(n21801), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n21803), 
        .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21565) );
  AOI21_X1 U23514 ( .B1(n21805), .B2(n21804), .A(n21824), .ZN(n21567) );
  OAI22_X1 U23515 ( .A1(n21601), .A2(n21553), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21756), .ZN(n21796) );
  AOI211_X1 U23516 ( .C1(n21805), .C2(n21555), .A(n21554), .B(n21796), .ZN(
        n21556) );
  OAI211_X1 U23517 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21744), .A(
        n21567), .B(n21556), .ZN(n21559) );
  NOR2_X1 U23518 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21571), .ZN(
        n21557) );
  AOI22_X1 U23519 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21559), .B1(
        n21558), .B2(n21557), .ZN(n21560) );
  OAI21_X1 U23520 ( .B1(n21735), .B2(n21561), .A(n21560), .ZN(n21563) );
  AOI22_X1 U23521 ( .A1(n21773), .A2(n21563), .B1(n21613), .B2(n21562), .ZN(
        n21564) );
  OAI211_X1 U23522 ( .C1(n21566), .C2(n21813), .A(n21565), .B(n21564), .ZN(
        P3_U2848) );
  INV_X1 U23523 ( .A(n21568), .ZN(n21570) );
  OAI211_X1 U23524 ( .C1(n21568), .C2(n21807), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21567), .ZN(n21569) );
  AOI221_X1 U23525 ( .B1(n21570), .B2(n21818), .C1(n21815), .C2(n21818), .A(
        n21569), .ZN(n21781) );
  NOR3_X1 U23526 ( .A1(n21781), .A2(n21571), .A3(n21570), .ZN(n21580) );
  INV_X1 U23527 ( .A(n21572), .ZN(n21576) );
  NAND2_X1 U23528 ( .A1(n21834), .A2(n21732), .ZN(n21771) );
  NOR2_X1 U23529 ( .A1(n21735), .A2(n21573), .ZN(n21762) );
  INV_X1 U23530 ( .A(n21762), .ZN(n21574) );
  OAI22_X1 U23531 ( .A1(n21576), .A2(n21771), .B1(n21575), .B2(n21574), .ZN(
        n21579) );
  NAND2_X1 U23532 ( .A1(n21793), .A2(n21771), .ZN(n21766) );
  NOR2_X1 U23533 ( .A1(n21762), .A2(n21766), .ZN(n21782) );
  AOI211_X1 U23534 ( .C1(n21781), .C2(n21782), .A(n21832), .B(n21577), .ZN(
        n21578) );
  AOI221_X1 U23535 ( .B1(n21580), .B2(n21668), .C1(n21579), .C2(n21773), .A(
        n21578), .ZN(n21582) );
  OAI211_X1 U23536 ( .C1(n21583), .C2(n21813), .A(n21582), .B(n21581), .ZN(
        P3_U2847) );
  AOI22_X1 U23537 ( .A1(n21803), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n21828), .B2(n21584), .ZN(n21595) );
  NOR2_X1 U23538 ( .A1(n21588), .A2(n21589), .ZN(n21598) );
  INV_X1 U23539 ( .A(n21598), .ZN(n21619) );
  NOR2_X1 U23540 ( .A1(n21585), .A2(n21619), .ZN(n21644) );
  AOI21_X1 U23541 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21644), .A(
        n21601), .ZN(n21592) );
  OAI211_X1 U23542 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21807), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n21586), .ZN(n21591) );
  INV_X1 U23543 ( .A(n21587), .ZN(n21618) );
  OAI21_X1 U23544 ( .B1(n21618), .B2(n21589), .A(n21588), .ZN(n21590) );
  OAI211_X1 U23545 ( .C1(n21592), .C2(n21591), .A(n21668), .B(n21590), .ZN(
        n21593) );
  NAND3_X1 U23546 ( .A1(n21595), .A2(n21594), .A3(n21593), .ZN(P3_U2840) );
  INV_X1 U23547 ( .A(n21596), .ZN(n21605) );
  NAND2_X1 U23548 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21620) );
  NOR4_X1 U23549 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21597), .A3(
        n21619), .A4(n21620), .ZN(n21604) );
  NAND2_X1 U23550 ( .A1(n21599), .A2(n21598), .ZN(n21628) );
  AND2_X1 U23551 ( .A1(n21835), .A2(n21628), .ZN(n21717) );
  OAI221_X1 U23552 ( .B1(n21644), .B2(n21601), .C1(n21644), .C2(n21822), .A(
        n21600), .ZN(n21713) );
  AOI211_X1 U23553 ( .C1(n21727), .C2(n21620), .A(n21717), .B(n21713), .ZN(
        n21615) );
  OAI22_X1 U23554 ( .A1(n21615), .A2(n21611), .B1(n21735), .B2(n21602), .ZN(
        n21603) );
  AOI211_X1 U23555 ( .C1(n21605), .C2(n21834), .A(n21604), .B(n21603), .ZN(
        n21609) );
  AOI22_X1 U23556 ( .A1(n21803), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n21828), .B2(n21606), .ZN(n21608) );
  OAI211_X1 U23557 ( .C1(n21609), .C2(n21685), .A(n21608), .B(n21607), .ZN(
        P3_U2837) );
  NOR2_X1 U23558 ( .A1(n21629), .A2(n21735), .ZN(n21610) );
  AOI211_X1 U23559 ( .C1(n21727), .C2(n21611), .A(n21610), .B(n21685), .ZN(
        n21614) );
  NAND2_X1 U23560 ( .A1(n21613), .A2(n21612), .ZN(n21632) );
  OAI221_X1 U23561 ( .B1(n21832), .B2(n21615), .C1(n21832), .C2(n21614), .A(
        n21632), .ZN(n21617) );
  AOI22_X1 U23562 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21617), .B1(
        n21828), .B2(n21616), .ZN(n21623) );
  NOR2_X1 U23563 ( .A1(n21619), .A2(n21618), .ZN(n21719) );
  INV_X1 U23564 ( .A(n21620), .ZN(n21626) );
  NAND4_X1 U23565 ( .A1(n21668), .A2(n21719), .A3(n21626), .A4(n21621), .ZN(
        n21622) );
  OAI211_X1 U23566 ( .C1(n21624), .C2(n21808), .A(n21623), .B(n21622), .ZN(
        P3_U2836) );
  INV_X1 U23567 ( .A(n21625), .ZN(n21639) );
  NAND2_X1 U23568 ( .A1(n21627), .A2(n21626), .ZN(n21634) );
  NOR2_X1 U23569 ( .A1(n21634), .A2(n21628), .ZN(n21652) );
  NOR2_X1 U23570 ( .A1(n21652), .A2(n21756), .ZN(n21646) );
  INV_X1 U23571 ( .A(n21634), .ZN(n21701) );
  OAI22_X1 U23572 ( .A1(n21764), .A2(n21701), .B1(n21629), .B2(n21735), .ZN(
        n21630) );
  NOR4_X1 U23573 ( .A1(n21646), .A2(n21631), .A3(n21713), .A4(n21630), .ZN(
        n21633) );
  OAI21_X1 U23574 ( .B1(n21633), .B2(n21685), .A(n21632), .ZN(n21636) );
  INV_X1 U23575 ( .A(n21719), .ZN(n21703) );
  NOR2_X1 U23576 ( .A1(n21703), .A2(n21634), .ZN(n21635) );
  AOI222_X1 U23577 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21636), 
        .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21803), .C1(n21636), 
        .C2(n21635), .ZN(n21638) );
  OAI211_X1 U23578 ( .C1(n21639), .C2(n21813), .A(n21638), .B(n21637), .ZN(
        P3_U2835) );
  NOR2_X1 U23579 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21756), .ZN(
        n21691) );
  NOR2_X1 U23580 ( .A1(n21641), .A2(n21640), .ZN(n21643) );
  OAI22_X1 U23581 ( .A1(n21643), .A2(n21735), .B1(n21642), .B2(n21695), .ZN(
        n21669) );
  NOR4_X1 U23582 ( .A1(n21691), .A2(n21685), .A3(n21665), .A4(n21669), .ZN(
        n21648) );
  NAND3_X1 U23583 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21701), .A3(
        n21644), .ZN(n21692) );
  NOR2_X1 U23584 ( .A1(n21645), .A2(n21692), .ZN(n21653) );
  AOI211_X1 U23585 ( .C1(n21818), .C2(n21692), .A(n21646), .B(n21763), .ZN(
        n21694) );
  OAI21_X1 U23586 ( .B1(n21822), .B2(n21653), .A(n21694), .ZN(n21647) );
  INV_X1 U23587 ( .A(n21647), .ZN(n21662) );
  NAND3_X1 U23588 ( .A1(n21648), .A2(n21662), .A3(n11270), .ZN(n21659) );
  INV_X1 U23589 ( .A(n21649), .ZN(n21699) );
  NOR2_X1 U23590 ( .A1(n21756), .A2(n21650), .ZN(n21651) );
  AOI22_X1 U23591 ( .A1(n21654), .A2(n21653), .B1(n21652), .B2(n21651), .ZN(
        n21677) );
  OAI21_X1 U23592 ( .B1(n21735), .B2(n21699), .A(n21677), .ZN(n21655) );
  AOI21_X1 U23593 ( .B1(n21834), .B2(n21696), .A(n21655), .ZN(n21666) );
  OAI22_X1 U23594 ( .A1(n21832), .A2(n21665), .B1(n21666), .B2(n21685), .ZN(
        n21658) );
  OAI21_X1 U23595 ( .B1(n21808), .B2(n21661), .A(n21660), .ZN(P3_U2833) );
  AOI22_X1 U23596 ( .A1(n21801), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21803), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21671) );
  OAI211_X1 U23597 ( .C1(n21783), .C2(n21663), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n21662), .ZN(n21673) );
  OAI21_X1 U23598 ( .B1(n21666), .B2(n21665), .A(n21664), .ZN(n21667) );
  OAI211_X1 U23599 ( .C1(n21669), .C2(n21673), .A(n21668), .B(n21667), .ZN(
        n21670) );
  OAI211_X1 U23600 ( .C1(n21672), .C2(n21813), .A(n21671), .B(n21670), .ZN(
        P3_U2832) );
  AND3_X1 U23601 ( .A1(n21727), .A2(n21673), .A3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21680) );
  NAND2_X1 U23602 ( .A1(n21675), .A2(n21674), .ZN(n21676) );
  OAI22_X1 U23603 ( .A1(n21678), .A2(n21735), .B1(n21677), .B2(n21676), .ZN(
        n21679) );
  AOI211_X1 U23604 ( .C1(n21834), .C2(n21681), .A(n21680), .B(n21679), .ZN(
        n21686) );
  AOI21_X1 U23605 ( .B1(n21682), .B2(n21828), .A(n11287), .ZN(n21684) );
  OAI211_X1 U23606 ( .C1(n21686), .C2(n21685), .A(n21684), .B(n21683), .ZN(
        P3_U2831) );
  NAND2_X1 U23607 ( .A1(n21687), .A2(n21688), .ZN(n21704) );
  INV_X1 U23608 ( .A(n21689), .ZN(n21690) );
  AOI21_X1 U23609 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21704), .A(
        n21690), .ZN(n21698) );
  AOI211_X1 U23610 ( .C1(n21805), .C2(n21692), .A(n21691), .B(n21803), .ZN(
        n21693) );
  OAI211_X1 U23611 ( .C1(n21696), .C2(n21695), .A(n21694), .B(n21693), .ZN(
        n21697) );
  NAND2_X1 U23612 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21701), .ZN(
        n21702) );
  OAI22_X1 U23613 ( .A1(n21705), .A2(n21704), .B1(n21703), .B2(n21702), .ZN(
        n21706) );
  OAI221_X1 U23614 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21773), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21706), .A(n21808), .ZN(
        n21711) );
  OR3_X1 U23615 ( .A1(n21708), .A2(n21813), .A3(n21707), .ZN(n21710) );
  OAI211_X1 U23616 ( .C1(n21712), .C2(n21711), .A(n21710), .B(n21709), .ZN(
        P3_U2834) );
  AOI211_X1 U23617 ( .C1(n21834), .C2(n21714), .A(n21803), .B(n21713), .ZN(
        n21715) );
  OAI21_X1 U23618 ( .B1(n21716), .B2(n21735), .A(n21715), .ZN(n21726) );
  NOR2_X1 U23619 ( .A1(n21726), .A2(n21717), .ZN(n21718) );
  AOI21_X1 U23620 ( .B1(n21718), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n21832), .ZN(n21725) );
  OAI221_X1 U23621 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21719), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21793), .A(n21725), .ZN(
        n21721) );
  OAI211_X1 U23622 ( .C1(n21813), .C2(n21722), .A(n21721), .B(n21720), .ZN(
        P3_U2839) );
  AOI22_X1 U23623 ( .A1(n21801), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n21724), 
        .B2(n21723), .ZN(n21729) );
  OAI211_X1 U23624 ( .C1(n21727), .C2(n21726), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21725), .ZN(n21728) );
  OAI211_X1 U23625 ( .C1(n21730), .C2(n21813), .A(n21729), .B(n21728), .ZN(
        P3_U2838) );
  OAI21_X1 U23626 ( .B1(n21732), .B2(n21731), .A(n21834), .ZN(n21733) );
  OAI211_X1 U23627 ( .C1(n21736), .C2(n21735), .A(n21734), .B(n21733), .ZN(
        n21737) );
  OAI21_X1 U23628 ( .B1(n21738), .B2(n21737), .A(n21808), .ZN(n21742) );
  AOI22_X1 U23629 ( .A1(n21801), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21828), 
        .B2(n21739), .ZN(n21740) );
  OAI221_X1 U23630 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21749), 
        .C1(n21741), .C2(n21742), .A(n21740), .ZN(P3_U2843) );
  NAND2_X1 U23631 ( .A1(n21741), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21743) );
  OAI21_X1 U23632 ( .B1(n21744), .B2(n21743), .A(n21742), .ZN(n21746) );
  AOI22_X1 U23633 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21746), .B1(
        n21828), .B2(n21745), .ZN(n21748) );
  OAI211_X1 U23634 ( .C1(n21750), .C2(n21749), .A(n21748), .B(n21747), .ZN(
        P3_U2842) );
  NAND2_X1 U23635 ( .A1(n21751), .A2(n21826), .ZN(n21788) );
  AOI22_X1 U23636 ( .A1(n21801), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n21828), 
        .B2(n21752), .ZN(n21768) );
  AOI21_X1 U23637 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21753), .A(
        n21764), .ZN(n21761) );
  OAI21_X1 U23638 ( .B1(n21755), .B2(n21754), .A(n21835), .ZN(n21758) );
  AOI22_X1 U23639 ( .A1(n21759), .A2(n21758), .B1(n21757), .B2(n21756), .ZN(
        n21760) );
  NOR4_X1 U23640 ( .A1(n21763), .A2(n21762), .A3(n21761), .A4(n21760), .ZN(
        n21772) );
  OAI21_X1 U23641 ( .B1(n21764), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n21772), .ZN(n21765) );
  OAI211_X1 U23642 ( .C1(n21766), .C2(n21765), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n21808), .ZN(n21767) );
  OAI211_X1 U23643 ( .C1(n21769), .C2(n21788), .A(n21768), .B(n21767), .ZN(
        P3_U2844) );
  NAND2_X1 U23644 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21770), .ZN(
        n21779) );
  NOR2_X1 U23645 ( .A1(n21832), .A2(n21770), .ZN(n21775) );
  NAND3_X1 U23646 ( .A1(n21773), .A2(n21772), .A3(n21771), .ZN(n21774) );
  AOI22_X1 U23647 ( .A1(n21828), .A2(n21776), .B1(n21775), .B2(n21774), .ZN(
        n21778) );
  OAI211_X1 U23648 ( .C1(n21779), .C2(n21788), .A(n21778), .B(n21777), .ZN(
        P3_U2845) );
  AOI221_X1 U23649 ( .B1(n21783), .B2(n21782), .C1(n21781), .C2(n21782), .A(
        n21780), .ZN(n21784) );
  AOI22_X1 U23650 ( .A1(n21785), .A2(n21828), .B1(n21784), .B2(n21808), .ZN(
        n21787) );
  OAI211_X1 U23651 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n21788), .A(
        n21787), .B(n21786), .ZN(P3_U2846) );
  AOI22_X1 U23652 ( .A1(n21801), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21826), 
        .B2(n21789), .ZN(n21798) );
  OAI21_X1 U23653 ( .B1(n21791), .B2(n21790), .A(n21805), .ZN(n21792) );
  NAND3_X1 U23654 ( .A1(n21794), .A2(n21793), .A3(n21792), .ZN(n21795) );
  OAI211_X1 U23655 ( .C1(n21796), .C2(n21795), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21808), .ZN(n21797) );
  OAI211_X1 U23656 ( .C1(n21799), .C2(n21813), .A(n21798), .B(n21797), .ZN(
        P3_U2849) );
  NOR2_X1 U23657 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21825), .ZN(
        n21800) );
  AOI22_X1 U23658 ( .A1(n21801), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21826), 
        .B2(n21800), .ZN(n21812) );
  NOR2_X1 U23659 ( .A1(n21803), .A2(n21802), .ZN(n21820) );
  NAND2_X1 U23660 ( .A1(n21805), .A2(n21804), .ZN(n21806) );
  OAI211_X1 U23661 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21807), .A(
        n21820), .B(n21806), .ZN(n21809) );
  OAI211_X1 U23662 ( .C1(n21810), .C2(n21809), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21808), .ZN(n21811) );
  OAI211_X1 U23663 ( .C1(n21814), .C2(n21813), .A(n21812), .B(n21811), .ZN(
        P3_U2852) );
  OAI211_X1 U23664 ( .C1(n21818), .C2(n21817), .A(n21816), .B(n21815), .ZN(
        n21819) );
  OAI211_X1 U23665 ( .C1(n21822), .C2(n21821), .A(n21820), .B(n21819), .ZN(
        n21823) );
  OAI21_X1 U23666 ( .B1(n21824), .B2(n21823), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21831) );
  AOI22_X1 U23667 ( .A1(n21828), .A2(n21827), .B1(n21826), .B2(n21825), .ZN(
        n21829) );
  OAI221_X1 U23668 ( .B1(n21832), .B2(n21831), .C1(n21808), .C2(n21830), .A(
        n21829), .ZN(P3_U2853) );
  NAND2_X1 U23669 ( .A1(n22292), .A2(n21886), .ZN(n21881) );
  INV_X1 U23670 ( .A(n21833), .ZN(n21880) );
  NOR2_X1 U23671 ( .A1(n21835), .A2(n21834), .ZN(n21837) );
  OAI222_X1 U23672 ( .A1(n21841), .A2(n21840), .B1(n21839), .B2(n21838), .C1(
        n21837), .C2(n21836), .ZN(n21899) );
  AND2_X1 U23673 ( .A1(n21843), .A2(n21842), .ZN(n21898) );
  OAI21_X1 U23674 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21898), .ZN(n21844) );
  OAI211_X1 U23675 ( .C1(n21849), .C2(n21846), .A(n21845), .B(n21844), .ZN(
        n21870) );
  MUX2_X1 U23676 ( .A(n21848), .B(n21847), .S(n21849), .Z(n21868) );
  INV_X1 U23677 ( .A(n21849), .ZN(n21859) );
  AOI22_X1 U23678 ( .A1(n21859), .A2(n21851), .B1(n21850), .B2(n21849), .ZN(
        n21863) );
  OR3_X1 U23679 ( .A1(n21856), .A2(n21855), .A3(n21852), .ZN(n21853) );
  AOI22_X1 U23680 ( .A1(n21856), .A2(n21855), .B1(n21854), .B2(n21853), .ZN(
        n21858) );
  OAI21_X1 U23681 ( .B1(n21859), .B2(n21858), .A(n21857), .ZN(n21862) );
  AND2_X1 U23682 ( .A1(n21863), .A2(n21862), .ZN(n21860) );
  OAI221_X1 U23683 ( .B1(n21863), .B2(n21862), .C1(n21861), .C2(n21860), .A(
        n21865), .ZN(n21867) );
  AOI21_X1 U23684 ( .B1(n21865), .B2(n21864), .A(n21863), .ZN(n21866) );
  AOI222_X1 U23685 ( .A1(n21868), .A2(n21867), .B1(n21868), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21867), .C2(n21866), .ZN(
        n21869) );
  NOR4_X1 U23686 ( .A1(n21871), .A2(n21899), .A3(n21870), .A4(n21869), .ZN(
        n21896) );
  OAI211_X1 U23687 ( .C1(n21874), .C2(n21873), .A(n21872), .B(n21896), .ZN(
        n21884) );
  OAI21_X1 U23688 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21875), .A(n21884), 
        .ZN(n21890) );
  INV_X1 U23689 ( .A(n21890), .ZN(n21877) );
  NAND3_X1 U23690 ( .A1(n21878), .A2(n21877), .A3(n21876), .ZN(n21879) );
  NAND4_X1 U23691 ( .A1(n21882), .A2(n21881), .A3(n21880), .A4(n21879), .ZN(
        P3_U2997) );
  OAI221_X1 U23692 ( .B1(n21885), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21885), 
        .C2(n21884), .A(n21883), .ZN(P3_U3282) );
  AOI22_X1 U23693 ( .A1(n21888), .A2(n21887), .B1(n22292), .B2(n21886), .ZN(
        n21889) );
  INV_X1 U23694 ( .A(n21889), .ZN(n21893) );
  NOR2_X1 U23695 ( .A1(n21891), .A2(n21890), .ZN(n21892) );
  MUX2_X1 U23696 ( .A(n21893), .B(n21892), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21895) );
  OAI211_X1 U23697 ( .C1(n21896), .C2(n21897), .A(n21895), .B(n21894), .ZN(
        P3_U2996) );
  NOR2_X1 U23698 ( .A1(n21898), .A2(n21897), .ZN(n21902) );
  MUX2_X1 U23699 ( .A(P3_MORE_REG_SCAN_IN), .B(n21899), .S(n21902), .Z(
        P3_U3295) );
  OAI21_X1 U23700 ( .B1(n21902), .B2(n21901), .A(n21900), .ZN(P3_U2637) );
  AOI211_X1 U23701 ( .C1(n21905), .C2(n22243), .A(n21904), .B(n21903), .ZN(
        n21911) );
  OAI211_X1 U23702 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21907), .A(n21906), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21908) );
  AOI21_X1 U23703 ( .B1(n21908), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n22214), 
        .ZN(n21910) );
  NAND2_X1 U23704 ( .A1(n21911), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21909) );
  OAI21_X1 U23705 ( .B1(n21911), .B2(n21910), .A(n21909), .ZN(P1_U3485) );
  NOR2_X1 U23706 ( .A1(n22016), .A2(n15977), .ZN(n21914) );
  INV_X1 U23707 ( .A(n21912), .ZN(n21913) );
  AOI211_X1 U23708 ( .C1(n21916), .C2(n21915), .A(n21914), .B(n21913), .ZN(
        n21920) );
  AOI22_X1 U23709 ( .A1(n21918), .A2(n22038), .B1(n22037), .B2(n21917), .ZN(
        n21919) );
  OAI211_X1 U23710 ( .C1(n21922), .C2(n21921), .A(n21920), .B(n21919), .ZN(
        P1_U3018) );
  NAND2_X1 U23711 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21924) );
  AOI211_X1 U23712 ( .C1(n21981), .C2(n21924), .A(n21923), .B(n21979), .ZN(
        n21939) );
  AOI22_X1 U23713 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21926), .B1(
        n21985), .B2(n21925), .ZN(n21941) );
  AOI211_X1 U23714 ( .C1(n21933), .C2(n21940), .A(n21941), .B(n21927), .ZN(
        n21931) );
  NOR2_X1 U23715 ( .A1(n21928), .A2(n22033), .ZN(n21930) );
  INV_X1 U23716 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n22053) );
  OAI22_X1 U23717 ( .A1(n22062), .A2(n22017), .B1(n22016), .B2(n22053), .ZN(
        n21929) );
  NOR3_X1 U23718 ( .A1(n21931), .A2(n21930), .A3(n21929), .ZN(n21932) );
  OAI21_X1 U23719 ( .B1(n21939), .B2(n21933), .A(n21932), .ZN(P1_U3027) );
  NOR2_X1 U23720 ( .A1(n21934), .A2(n22033), .ZN(n21935) );
  AOI211_X1 U23721 ( .C1(n22037), .C2(n21937), .A(n21936), .B(n21935), .ZN(
        n21938) );
  OAI221_X1 U23722 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21941), .C1(
        n21940), .C2(n21939), .A(n21938), .ZN(P1_U3028) );
  INV_X1 U23723 ( .A(n21965), .ZN(n21943) );
  OAI21_X1 U23724 ( .B1(n21944), .B2(n21943), .A(n21942), .ZN(n21960) );
  AOI21_X1 U23725 ( .B1(n21953), .B2(n21952), .A(n21960), .ZN(n21949) );
  INV_X1 U23726 ( .A(n21945), .ZN(n21946) );
  AOI222_X1 U23727 ( .A1(n21947), .A2(n22038), .B1(n22037), .B2(n21946), .C1(
        n22040), .C2(P1_REIP_REG_6__SCAN_IN), .ZN(n21948) );
  OAI221_X1 U23728 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21951), .C1(
        n21950), .C2(n21949), .A(n21948), .ZN(P1_U3025) );
  NAND2_X1 U23729 ( .A1(n21953), .A2(n21952), .ZN(n21964) );
  NAND2_X1 U23730 ( .A1(n21985), .A2(n21954), .ZN(n21957) );
  OAI222_X1 U23731 ( .A1(n21958), .A2(n22016), .B1(n21957), .B2(n21956), .C1(
        n22017), .C2(n21955), .ZN(n21959) );
  INV_X1 U23732 ( .A(n21959), .ZN(n21963) );
  AOI22_X1 U23733 ( .A1(n21961), .A2(n22038), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21960), .ZN(n21962) );
  OAI211_X1 U23734 ( .C1(n21965), .C2(n21964), .A(n21963), .B(n21962), .ZN(
        P1_U3026) );
  AOI222_X1 U23735 ( .A1(n21966), .A2(n22038), .B1(n22037), .B2(n22068), .C1(
        n22040), .C2(P1_REIP_REG_7__SCAN_IN), .ZN(n21968) );
  OAI211_X1 U23736 ( .C1(n21970), .C2(n21969), .A(n21968), .B(n21967), .ZN(
        P1_U3024) );
  NOR2_X1 U23737 ( .A1(n21971), .A2(n22033), .ZN(n21972) );
  AOI211_X1 U23738 ( .C1(n22037), .C2(n21974), .A(n21973), .B(n21972), .ZN(
        n21975) );
  OAI221_X1 U23739 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21978), .C1(
        n21977), .C2(n21976), .A(n21975), .ZN(P1_U3022) );
  AOI21_X1 U23740 ( .B1(n21981), .B2(n21980), .A(n21979), .ZN(n21982) );
  INV_X1 U23741 ( .A(n21982), .ZN(n21983) );
  AOI21_X1 U23742 ( .B1(n21985), .B2(n21984), .A(n21983), .ZN(n22004) );
  NAND2_X1 U23743 ( .A1(n21986), .A2(n22003), .ZN(n21992) );
  NOR3_X1 U23744 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21987), .A3(
        n22003), .ZN(n21990) );
  OAI22_X1 U23745 ( .A1(n21988), .A2(n22033), .B1(n22017), .B2(n22102), .ZN(
        n21989) );
  AOI211_X1 U23746 ( .C1(P1_REIP_REG_12__SCAN_IN), .C2(n22040), .A(n21990), 
        .B(n21989), .ZN(n21991) );
  OAI221_X1 U23747 ( .B1(n21993), .B2(n22004), .C1(n21993), .C2(n21992), .A(
        n21991), .ZN(P1_U3019) );
  OR2_X1 U23748 ( .A1(n21994), .A2(n22033), .ZN(n22001) );
  INV_X1 U23749 ( .A(n21995), .ZN(n21996) );
  OAI21_X1 U23750 ( .B1(n21997), .B2(n22017), .A(n21996), .ZN(n21998) );
  AOI21_X1 U23751 ( .B1(n21999), .B2(n22003), .A(n21998), .ZN(n22000) );
  AND2_X1 U23752 ( .A1(n22001), .A2(n22000), .ZN(n22002) );
  OAI21_X1 U23753 ( .B1(n22004), .B2(n22003), .A(n22002), .ZN(P1_U3020) );
  NAND2_X1 U23754 ( .A1(n22040), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n22005) );
  OAI221_X1 U23755 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n22025), 
        .C1(n22006), .C2(n22013), .A(n22005), .ZN(n22007) );
  AOI21_X1 U23756 ( .B1(n22008), .B2(n22037), .A(n22007), .ZN(n22009) );
  OAI21_X1 U23757 ( .B1(n22010), .B2(n22033), .A(n22009), .ZN(P1_U3016) );
  NAND2_X1 U23758 ( .A1(n22012), .A2(n22011), .ZN(n22022) );
  OAI21_X1 U23759 ( .B1(n22015), .B2(n22014), .A(n22013), .ZN(n22029) );
  NOR2_X1 U23760 ( .A1(n22016), .A2(n22131), .ZN(n22020) );
  OAI22_X1 U23761 ( .A1(n22018), .A2(n22033), .B1(n22017), .B2(n22136), .ZN(
        n22019) );
  AOI211_X1 U23762 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n22029), .A(
        n22020), .B(n22019), .ZN(n22021) );
  OAI21_X1 U23763 ( .B1(n22023), .B2(n22022), .A(n22021), .ZN(P1_U3013) );
  OAI21_X1 U23764 ( .B1(n22026), .B2(n22025), .A(n22024), .ZN(n22030) );
  INV_X1 U23765 ( .A(n22027), .ZN(n22028) );
  AOI22_X1 U23766 ( .A1(n22030), .A2(n22029), .B1(n22037), .B2(n22028), .ZN(
        n22032) );
  NAND2_X1 U23767 ( .A1(n22040), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n22031) );
  OAI211_X1 U23768 ( .C1(n22034), .C2(n22033), .A(n22032), .B(n22031), .ZN(
        P1_U3014) );
  INV_X1 U23769 ( .A(n22035), .ZN(n22039) );
  AOI22_X1 U23770 ( .A1(n22039), .A2(n22038), .B1(n22037), .B2(n22036), .ZN(
        n22049) );
  NAND2_X1 U23771 ( .A1(n22040), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n22048) );
  OAI21_X1 U23772 ( .B1(n22042), .B2(n22041), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22047) );
  NAND3_X1 U23773 ( .A1(n22045), .A2(n22044), .A3(n22043), .ZN(n22046) );
  NAND4_X1 U23774 ( .A1(n22049), .A2(n22048), .A3(n22047), .A4(n22046), .ZN(
        P1_U3009) );
  NAND2_X1 U23775 ( .A1(n22051), .A2(n22050), .ZN(n22061) );
  INV_X1 U23776 ( .A(n22052), .ZN(n22054) );
  OAI21_X1 U23777 ( .B1(n22138), .B2(n22054), .A(n22053), .ZN(n22058) );
  AOI21_X1 U23778 ( .B1(n22151), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22139), .ZN(n22055) );
  OAI21_X1 U23779 ( .B1(n22191), .B2(n22056), .A(n22055), .ZN(n22057) );
  AOI21_X1 U23780 ( .B1(n22059), .B2(n22058), .A(n22057), .ZN(n22060) );
  OAI211_X1 U23781 ( .C1(n22062), .C2(n22202), .A(n22061), .B(n22060), .ZN(
        n22063) );
  AOI21_X1 U23782 ( .B1(n22065), .B2(n22064), .A(n22063), .ZN(n22066) );
  OAI21_X1 U23783 ( .B1(n22067), .B2(n22186), .A(n22066), .ZN(P1_U2836) );
  INV_X1 U23784 ( .A(n22068), .ZN(n22070) );
  INV_X1 U23785 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n22069) );
  OAI22_X1 U23786 ( .A1(n22070), .A2(n22202), .B1(n22191), .B2(n22069), .ZN(
        n22071) );
  AOI211_X1 U23787 ( .C1(n22151), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22139), .B(n22071), .ZN(n22072) );
  OAI221_X1 U23788 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n22075), .C1(n22074), 
        .C2(n22073), .A(n22072), .ZN(n22076) );
  AOI21_X1 U23789 ( .B1(n22077), .B2(n22197), .A(n22076), .ZN(n22078) );
  OAI21_X1 U23790 ( .B1(n22079), .B2(n22186), .A(n22078), .ZN(P1_U2833) );
  AOI21_X1 U23791 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n22119), .A(n22080), .ZN(
        n22088) );
  OAI22_X1 U23792 ( .A1(n22082), .A2(n22202), .B1(n22081), .B2(n22191), .ZN(
        n22083) );
  AOI211_X1 U23793 ( .C1(n22151), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n22139), .B(n22083), .ZN(n22087) );
  AOI22_X1 U23794 ( .A1(n22085), .A2(n22197), .B1(n22195), .B2(n22084), .ZN(
        n22086) );
  OAI211_X1 U23795 ( .C1(n22089), .C2(n22088), .A(n22087), .B(n22086), .ZN(
        P1_U2831) );
  AOI211_X1 U23796 ( .C1(n22091), .C2(n22094), .A(n22090), .B(n22138), .ZN(
        n22097) );
  AOI22_X1 U23797 ( .A1(n11143), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n22151), .ZN(n22093) );
  OAI211_X1 U23798 ( .C1(n22095), .C2(n22094), .A(n22093), .B(n22122), .ZN(
        n22096) );
  AOI211_X1 U23799 ( .C1(n22098), .C2(n22197), .A(n22097), .B(n22096), .ZN(
        n22101) );
  NAND2_X1 U23800 ( .A1(n22099), .A2(n22195), .ZN(n22100) );
  OAI211_X1 U23801 ( .C1(n22102), .C2(n22202), .A(n22101), .B(n22100), .ZN(
        P1_U2828) );
  NOR2_X1 U23802 ( .A1(n22103), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n22106) );
  OAI22_X1 U23803 ( .A1(n22106), .A2(n22105), .B1(n22191), .B2(n22104), .ZN(
        n22107) );
  AOI211_X1 U23804 ( .C1(n22151), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n22139), .B(n22107), .ZN(n22112) );
  INV_X1 U23805 ( .A(n22108), .ZN(n22109) );
  AOI22_X1 U23806 ( .A1(n22110), .A2(n22197), .B1(n22109), .B2(n22195), .ZN(
        n22111) );
  OAI211_X1 U23807 ( .C1(n22202), .C2(n22113), .A(n22112), .B(n22111), .ZN(
        P1_U2826) );
  AOI22_X1 U23808 ( .A1(n11143), .A2(P1_EBX_REG_16__SCAN_IN), .B1(n22151), 
        .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n22124) );
  OAI22_X1 U23809 ( .A1(n22115), .A2(n22181), .B1(n22202), .B2(n22114), .ZN(
        n22116) );
  AOI21_X1 U23810 ( .B1(n22117), .B2(n22195), .A(n22116), .ZN(n22123) );
  OAI211_X1 U23811 ( .C1(n22120), .C2(P1_REIP_REG_16__SCAN_IN), .A(n22119), 
        .B(n22118), .ZN(n22121) );
  NAND4_X1 U23812 ( .A1(n22124), .A2(n22123), .A3(n22122), .A4(n22121), .ZN(
        P1_U2824) );
  AND2_X1 U23813 ( .A1(n22131), .A2(n22125), .ZN(n22146) );
  AOI21_X1 U23814 ( .B1(n22151), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n22139), .ZN(n22126) );
  OAI21_X1 U23815 ( .B1(n22191), .B2(n22127), .A(n22126), .ZN(n22128) );
  AOI211_X1 U23816 ( .C1(n22195), .C2(n22129), .A(n22146), .B(n22128), .ZN(
        n22135) );
  OAI22_X1 U23817 ( .A1(n22132), .A2(n22181), .B1(n22131), .B2(n22130), .ZN(
        n22133) );
  INV_X1 U23818 ( .A(n22133), .ZN(n22134) );
  OAI211_X1 U23819 ( .C1(n22202), .C2(n22136), .A(n22135), .B(n22134), .ZN(
        P1_U2822) );
  NOR3_X1 U23820 ( .A1(n22138), .A2(n22137), .A3(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n22144) );
  NAND2_X1 U23821 ( .A1(n11143), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n22141) );
  AOI21_X1 U23822 ( .B1(n22151), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22139), .ZN(n22140) );
  OAI211_X1 U23823 ( .C1(n22186), .C2(n22142), .A(n22141), .B(n22140), .ZN(
        n22143) );
  AOI211_X1 U23824 ( .C1(n22145), .C2(n22197), .A(n22144), .B(n22143), .ZN(
        n22149) );
  OAI21_X1 U23825 ( .B1(n22147), .B2(n22146), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n22148) );
  OAI211_X1 U23826 ( .C1(n22150), .C2(n22202), .A(n22149), .B(n22148), .ZN(
        P1_U2821) );
  AOI22_X1 U23827 ( .A1(n11143), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n22151), .ZN(n22158) );
  AND2_X1 U23828 ( .A1(n22153), .A2(n22152), .ZN(n22156) );
  NOR2_X1 U23829 ( .A1(n22155), .A2(n22154), .ZN(n22168) );
  OAI21_X1 U23830 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n22156), .A(n22168), 
        .ZN(n22157) );
  OAI211_X1 U23831 ( .C1(n22159), .C2(n22181), .A(n22158), .B(n22157), .ZN(
        n22160) );
  AOI21_X1 U23832 ( .B1(n22161), .B2(n22195), .A(n22160), .ZN(n22162) );
  OAI21_X1 U23833 ( .B1(n22202), .B2(n22163), .A(n22162), .ZN(P1_U2820) );
  INV_X1 U23834 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n22164) );
  OAI22_X1 U23835 ( .A1(n22191), .A2(n20550), .B1(n22164), .B2(n22188), .ZN(
        n22165) );
  AOI221_X1 U23836 ( .B1(n22168), .B2(P1_REIP_REG_21__SCAN_IN), .C1(n22167), 
        .C2(n22166), .A(n22165), .ZN(n22173) );
  NOR2_X1 U23837 ( .A1(n22169), .A2(n22202), .ZN(n22170) );
  AOI21_X1 U23838 ( .B1(n22171), .B2(n22197), .A(n22170), .ZN(n22172) );
  OAI211_X1 U23839 ( .C1(n22174), .C2(n22186), .A(n22173), .B(n22172), .ZN(
        P1_U2819) );
  INV_X1 U23840 ( .A(n22175), .ZN(n22194) );
  OAI22_X1 U23841 ( .A1(n22191), .A2(n22177), .B1(n22176), .B2(n22188), .ZN(
        n22178) );
  AOI221_X1 U23842 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n22194), .C1(n22179), 
        .C2(n22194), .A(n22178), .ZN(n22185) );
  OAI22_X1 U23843 ( .A1(n22182), .A2(n22181), .B1(n22202), .B2(n22180), .ZN(
        n22183) );
  INV_X1 U23844 ( .A(n22183), .ZN(n22184) );
  OAI211_X1 U23845 ( .C1(n22187), .C2(n22186), .A(n22185), .B(n22184), .ZN(
        P1_U2817) );
  INV_X1 U23846 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n22189) );
  OAI22_X1 U23847 ( .A1(n22191), .A2(n22190), .B1(n22189), .B2(n22188), .ZN(
        n22192) );
  AOI211_X1 U23848 ( .C1(n22194), .C2(P1_REIP_REG_24__SCAN_IN), .A(n22193), 
        .B(n22192), .ZN(n22200) );
  AOI22_X1 U23849 ( .A1(n22198), .A2(n22197), .B1(n22196), .B2(n22195), .ZN(
        n22199) );
  OAI211_X1 U23850 ( .C1(n22202), .C2(n22201), .A(n22200), .B(n22199), .ZN(
        P1_U2816) );
  OAI21_X1 U23851 ( .B1(n22205), .B2(n22204), .A(n22203), .ZN(P1_U2806) );
  INV_X1 U23852 ( .A(n22206), .ZN(n22213) );
  NOR2_X1 U23853 ( .A1(n22213), .A2(n22210), .ZN(n22212) );
  OAI211_X1 U23854 ( .C1(n22212), .C2(n22476), .A(n22208), .B(n22207), .ZN(
        P1_U3163) );
  OAI22_X1 U23855 ( .A1(n22212), .A2(n22211), .B1(n22210), .B2(n22209), .ZN(
        P1_U3466) );
  AOI21_X1 U23856 ( .B1(n22215), .B2(n22214), .A(n22213), .ZN(n22216) );
  OAI22_X1 U23857 ( .A1(n22218), .A2(n22217), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22216), .ZN(n22219) );
  OAI21_X1 U23858 ( .B1(n22221), .B2(n22220), .A(n22219), .ZN(P1_U3161) );
  INV_X1 U23859 ( .A(n22222), .ZN(n22224) );
  OAI21_X1 U23860 ( .B1(n22226), .B2(n22223), .A(n22224), .ZN(P1_U2805) );
  OAI21_X1 U23861 ( .B1(n22226), .B2(n22225), .A(n22224), .ZN(P1_U3465) );
  INV_X1 U23862 ( .A(n22227), .ZN(n22229) );
  OAI21_X1 U23863 ( .B1(n22231), .B2(n22228), .A(n22229), .ZN(P2_U2818) );
  OAI21_X1 U23864 ( .B1(n22231), .B2(n22230), .A(n22229), .ZN(P2_U3592) );
  INV_X1 U23865 ( .A(n22232), .ZN(n22234) );
  OAI21_X1 U23866 ( .B1(n22236), .B2(n22233), .A(n22234), .ZN(P3_U2636) );
  OAI21_X1 U23867 ( .B1(n22236), .B2(n22235), .A(n22234), .ZN(P3_U3281) );
  INV_X1 U23868 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22237) );
  AOI21_X1 U23869 ( .B1(HOLD), .B2(n22238), .A(n22237), .ZN(n22239) );
  AOI21_X1 U23870 ( .B1(n22292), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22287), 
        .ZN(n22298) );
  AOI21_X1 U23871 ( .B1(n22288), .B2(NA), .A(n22285), .ZN(n22291) );
  OAI22_X1 U23872 ( .A1(n22240), .A2(n22239), .B1(n22298), .B2(n22291), .ZN(
        P3_U3029) );
  INV_X1 U23873 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22244) );
  OAI21_X1 U23874 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n22244), .A(HOLD), .ZN(
        n22249) );
  INV_X1 U23875 ( .A(n22241), .ZN(n22248) );
  INV_X1 U23876 ( .A(NA), .ZN(n22265) );
  NAND2_X1 U23877 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22242), .ZN(n22253) );
  NAND2_X1 U23878 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22253), .ZN(n22256) );
  OAI211_X1 U23879 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n22265), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n22256), .ZN(n22247) );
  AOI211_X1 U23880 ( .C1(n22249), .C2(n22244), .A(n22250), .B(n22243), .ZN(
        n22245) );
  NAND3_X1 U23881 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22265), .A3(n22245), 
        .ZN(n22246) );
  OAI211_X1 U23882 ( .C1(n22249), .C2(n22248), .A(n22247), .B(n22246), .ZN(
        P1_U3196) );
  INV_X1 U23883 ( .A(HOLD), .ZN(n22269) );
  OAI21_X1 U23884 ( .B1(n22251), .B2(n22269), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22257) );
  INV_X1 U23885 ( .A(n22257), .ZN(n22252) );
  NOR2_X1 U23886 ( .A1(n22250), .A2(n22269), .ZN(n22258) );
  AOI22_X1 U23887 ( .A1(n22252), .A2(P1_STATE_REG_0__SCAN_IN), .B1(n22258), 
        .B2(n22251), .ZN(n22255) );
  NAND3_X1 U23888 ( .A1(n22255), .A2(n22254), .A3(n22253), .ZN(P1_U3195) );
  INV_X1 U23889 ( .A(n22256), .ZN(n22260) );
  AOI211_X1 U23890 ( .C1(NA), .C2(n11714), .A(n22258), .B(n22257), .ZN(n22259)
         );
  OAI22_X1 U23891 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22260), .B1(n22727), 
        .B2(n22259), .ZN(P1_U3194) );
  NAND3_X1 U23892 ( .A1(n22262), .A2(HOLD), .A3(n22261), .ZN(n22268) );
  OAI21_X1 U23893 ( .B1(n22264), .B2(n22263), .A(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n22277) );
  OAI21_X1 U23894 ( .B1(n22266), .B2(n22265), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n22283) );
  AOI22_X1 U23895 ( .A1(n22271), .A2(n17936), .B1(n22277), .B2(n22283), .ZN(
        n22267) );
  NAND2_X1 U23896 ( .A1(n22268), .A2(n22267), .ZN(P2_U3209) );
  NOR2_X1 U23897 ( .A1(n22270), .A2(n22269), .ZN(n22280) );
  NOR3_X1 U23898 ( .A1(n22280), .A2(n22271), .A3(n22282), .ZN(n22273) );
  AOI211_X1 U23899 ( .C1(n22274), .C2(HOLD), .A(n22273), .B(n22272), .ZN(
        n22276) );
  NAND2_X1 U23900 ( .A1(n22275), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22278) );
  NAND2_X1 U23901 ( .A1(n22276), .A2(n22278), .ZN(P2_U3210) );
  INV_X1 U23902 ( .A(n22277), .ZN(n22284) );
  OAI22_X1 U23903 ( .A1(NA), .A2(n22278), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22279) );
  OAI22_X1 U23904 ( .A1(n22280), .A2(n22279), .B1(HOLD), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22281) );
  OAI22_X1 U23905 ( .A1(n22284), .A2(n22283), .B1(n22282), .B2(n22281), .ZN(
        P2_U3211) );
  OAI21_X1 U23906 ( .B1(HOLD), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22295) );
  AOI21_X1 U23907 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n22295), .ZN(
        n22286) );
  AOI211_X1 U23908 ( .C1(n22285), .C2(n22287), .A(n22292), .B(n22286), .ZN(
        n22290) );
  AOI22_X1 U23909 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22287), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(n22286), .ZN(n22289) );
  AOI22_X1 U23910 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22290), .B1(n22289), 
        .B2(n22288), .ZN(P3_U3030) );
  INV_X1 U23911 ( .A(n22291), .ZN(n22297) );
  NAND2_X1 U23912 ( .A1(n22292), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n22293) );
  OAI22_X1 U23913 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n22293), .ZN(n22294) );
  AOI21_X1 U23914 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n22294), .ZN(
        n22296) );
  OAI22_X1 U23915 ( .A1(n22298), .A2(n22297), .B1(n22296), .B2(n22295), .ZN(
        P3_U3031) );
  NOR2_X1 U23916 ( .A1(n22381), .A2(n22300), .ZN(n22302) );
  AOI21_X1 U23917 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n22385), .A(n22302), 
        .ZN(n22301) );
  OAI21_X1 U23918 ( .B1(n12191), .B2(n22387), .A(n22301), .ZN(P1_U2937) );
  AOI21_X1 U23919 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n22385), .A(n22302), 
        .ZN(n22303) );
  OAI21_X1 U23920 ( .B1(n22304), .B2(n22387), .A(n22303), .ZN(P1_U2952) );
  NOR2_X1 U23921 ( .A1(n22381), .A2(n22305), .ZN(n22307) );
  AOI21_X1 U23922 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n22385), .A(n22307), 
        .ZN(n22306) );
  OAI21_X1 U23923 ( .B1(n15743), .B2(n22387), .A(n22306), .ZN(P1_U2938) );
  AOI21_X1 U23924 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n22385), .A(n22307), 
        .ZN(n22308) );
  OAI21_X1 U23925 ( .B1(n12070), .B2(n22387), .A(n22308), .ZN(P1_U2953) );
  NOR2_X1 U23926 ( .A1(n22381), .A2(n22309), .ZN(n22312) );
  AOI21_X1 U23927 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n22363), .A(n22312), 
        .ZN(n22310) );
  OAI21_X1 U23928 ( .B1(n22311), .B2(n22387), .A(n22310), .ZN(P1_U2939) );
  AOI21_X1 U23929 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n22363), .A(n22312), 
        .ZN(n22313) );
  OAI21_X1 U23930 ( .B1(n12060), .B2(n22387), .A(n22313), .ZN(P1_U2954) );
  NOR2_X1 U23931 ( .A1(n22381), .A2(n22314), .ZN(n22317) );
  AOI21_X1 U23932 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n22363), .A(n22317), 
        .ZN(n22315) );
  OAI21_X1 U23933 ( .B1(n22316), .B2(n22387), .A(n22315), .ZN(P1_U2940) );
  AOI21_X1 U23934 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n22363), .A(n22317), 
        .ZN(n22318) );
  OAI21_X1 U23935 ( .B1(n12090), .B2(n22387), .A(n22318), .ZN(P1_U2955) );
  NOR2_X1 U23936 ( .A1(n22381), .A2(n22319), .ZN(n22322) );
  AOI21_X1 U23937 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n22363), .A(n22322), 
        .ZN(n22320) );
  OAI21_X1 U23938 ( .B1(n22321), .B2(n22387), .A(n22320), .ZN(P1_U2941) );
  AOI21_X1 U23939 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n22363), .A(n22322), 
        .ZN(n22323) );
  OAI21_X1 U23940 ( .B1(n22324), .B2(n22387), .A(n22323), .ZN(P1_U2956) );
  NOR2_X1 U23941 ( .A1(n22381), .A2(n22325), .ZN(n22328) );
  AOI21_X1 U23942 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n22363), .A(n22328), 
        .ZN(n22326) );
  OAI21_X1 U23943 ( .B1(n22327), .B2(n22387), .A(n22326), .ZN(P1_U2942) );
  AOI21_X1 U23944 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n22363), .A(n22328), 
        .ZN(n22329) );
  OAI21_X1 U23945 ( .B1(n14869), .B2(n22387), .A(n22329), .ZN(P1_U2957) );
  NOR2_X1 U23946 ( .A1(n22381), .A2(n22330), .ZN(n22333) );
  AOI21_X1 U23947 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n22363), .A(n22333), 
        .ZN(n22331) );
  OAI21_X1 U23948 ( .B1(n22332), .B2(n22387), .A(n22331), .ZN(P1_U2943) );
  AOI21_X1 U23949 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n22363), .A(n22333), 
        .ZN(n22334) );
  OAI21_X1 U23950 ( .B1(n12122), .B2(n22387), .A(n22334), .ZN(P1_U2958) );
  NOR2_X1 U23951 ( .A1(n22381), .A2(n22335), .ZN(n22338) );
  AOI21_X1 U23952 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n22363), .A(n22338), 
        .ZN(n22336) );
  OAI21_X1 U23953 ( .B1(n22337), .B2(n22387), .A(n22336), .ZN(P1_U2944) );
  AOI21_X1 U23954 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n22363), .A(n22338), 
        .ZN(n22339) );
  OAI21_X1 U23955 ( .B1(n12052), .B2(n22387), .A(n22339), .ZN(P1_U2959) );
  INV_X1 U23956 ( .A(n22340), .ZN(n22341) );
  NOR2_X1 U23957 ( .A1(n22381), .A2(n22341), .ZN(n22344) );
  AOI21_X1 U23958 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n22363), .A(n22344), 
        .ZN(n22342) );
  OAI21_X1 U23959 ( .B1(n22343), .B2(n22387), .A(n22342), .ZN(P1_U2945) );
  AOI21_X1 U23960 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n22363), .A(n22344), 
        .ZN(n22345) );
  OAI21_X1 U23961 ( .B1(n22346), .B2(n22387), .A(n22345), .ZN(P1_U2960) );
  INV_X1 U23962 ( .A(n22347), .ZN(n22348) );
  NOR2_X1 U23963 ( .A1(n22381), .A2(n22348), .ZN(n22351) );
  AOI21_X1 U23964 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n22363), .A(n22351), 
        .ZN(n22349) );
  OAI21_X1 U23965 ( .B1(n22350), .B2(n22387), .A(n22349), .ZN(P1_U2946) );
  AOI21_X1 U23966 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n22363), .A(n22351), 
        .ZN(n22352) );
  OAI21_X1 U23967 ( .B1(n22353), .B2(n22387), .A(n22352), .ZN(P1_U2961) );
  NOR2_X1 U23968 ( .A1(n22381), .A2(n22354), .ZN(n22357) );
  AOI21_X1 U23969 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n22363), .A(n22357), 
        .ZN(n22355) );
  OAI21_X1 U23970 ( .B1(n22356), .B2(n22387), .A(n22355), .ZN(P1_U2947) );
  AOI21_X1 U23971 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n22363), .A(n22357), 
        .ZN(n22358) );
  OAI21_X1 U23972 ( .B1(n15134), .B2(n22387), .A(n22358), .ZN(P1_U2962) );
  NOR2_X1 U23973 ( .A1(n22381), .A2(n22359), .ZN(n22362) );
  AOI21_X1 U23974 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n22363), .A(n22362), 
        .ZN(n22360) );
  OAI21_X1 U23975 ( .B1(n22361), .B2(n22387), .A(n22360), .ZN(P1_U2948) );
  AOI21_X1 U23976 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n22363), .A(n22362), 
        .ZN(n22364) );
  OAI21_X1 U23977 ( .B1(n15696), .B2(n22387), .A(n22364), .ZN(P1_U2963) );
  INV_X1 U23978 ( .A(n22365), .ZN(n22366) );
  NOR2_X1 U23979 ( .A1(n22381), .A2(n22366), .ZN(n22369) );
  AOI21_X1 U23980 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n22385), .A(n22369), 
        .ZN(n22367) );
  OAI21_X1 U23981 ( .B1(n22368), .B2(n22387), .A(n22367), .ZN(P1_U2949) );
  AOI21_X1 U23982 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n22385), .A(n22369), 
        .ZN(n22370) );
  OAI21_X1 U23983 ( .B1(n22371), .B2(n22387), .A(n22370), .ZN(P1_U2964) );
  INV_X1 U23984 ( .A(n22372), .ZN(n22373) );
  NOR2_X1 U23985 ( .A1(n22381), .A2(n22373), .ZN(n22376) );
  AOI21_X1 U23986 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n22385), .A(n22376), 
        .ZN(n22374) );
  OAI21_X1 U23987 ( .B1(n22375), .B2(n22387), .A(n22374), .ZN(P1_U2950) );
  AOI21_X1 U23988 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n22385), .A(n22376), 
        .ZN(n22377) );
  OAI21_X1 U23989 ( .B1(n22378), .B2(n22387), .A(n22377), .ZN(P1_U2965) );
  INV_X1 U23990 ( .A(n22379), .ZN(n22380) );
  NOR2_X1 U23991 ( .A1(n22381), .A2(n22380), .ZN(n22384) );
  AOI21_X1 U23992 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n22385), .A(n22384), 
        .ZN(n22382) );
  OAI21_X1 U23993 ( .B1(n22383), .B2(n22387), .A(n22382), .ZN(P1_U2951) );
  AOI21_X1 U23994 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n22385), .A(n22384), 
        .ZN(n22386) );
  OAI21_X1 U23995 ( .B1(n22388), .B2(n22387), .A(n22386), .ZN(P1_U2966) );
  NOR3_X1 U23996 ( .A1(n22654), .A2(n22721), .A3(n22465), .ZN(n22389) );
  NOR2_X1 U23997 ( .A1(n22465), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22466) );
  NOR2_X1 U23998 ( .A1(n22389), .A2(n22466), .ZN(n22398) );
  INV_X1 U23999 ( .A(n22398), .ZN(n22391) );
  NOR2_X1 U24000 ( .A1(n22406), .A2(n22468), .ZN(n22397) );
  INV_X1 U24001 ( .A(n22394), .ZN(n22390) );
  NOR2_X1 U24002 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22392), .ZN(
        n22653) );
  AOI22_X1 U24003 ( .A1(n22721), .A2(n22490), .B1(n22653), .B2(n22489), .ZN(
        n22400) );
  INV_X1 U24004 ( .A(n22653), .ZN(n22393) );
  INV_X1 U24005 ( .A(n22411), .ZN(n22458) );
  AOI21_X1 U24006 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22393), .A(n22458), 
        .ZN(n22396) );
  NAND2_X1 U24007 ( .A1(n22394), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22395) );
  OAI211_X1 U24008 ( .C1(n22398), .C2(n22397), .A(n22396), .B(n22395), .ZN(
        n22655) );
  AOI22_X1 U24009 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22655), .B1(
        n22654), .B2(n22475), .ZN(n22399) );
  OAI211_X1 U24010 ( .C1(n22658), .C2(n22487), .A(n22400), .B(n22399), .ZN(
        P1_U3033) );
  INV_X1 U24011 ( .A(n22660), .ZN(n22551) );
  AOI22_X1 U24012 ( .A1(n22489), .A2(n22547), .B1(n22546), .B2(n22488), .ZN(
        n22402) );
  AOI22_X1 U24013 ( .A1(n22548), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n22654), .B2(n22490), .ZN(n22401) );
  OAI211_X1 U24014 ( .C1(n22493), .C2(n22551), .A(n22402), .B(n22401), .ZN(
        P1_U3041) );
  NOR3_X1 U24015 ( .A1(n22660), .A2(n22666), .A3(n22465), .ZN(n22405) );
  NOR2_X1 U24016 ( .A1(n22405), .A2(n22466), .ZN(n22413) );
  INV_X1 U24017 ( .A(n22413), .ZN(n22407) );
  NOR2_X1 U24018 ( .A1(n22406), .A2(n14933), .ZN(n22412) );
  NOR2_X1 U24019 ( .A1(n22477), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22434) );
  NOR3_X1 U24020 ( .A1(n22408), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22416) );
  NAND2_X1 U24021 ( .A1(n22454), .A2(n22416), .ZN(n22409) );
  INV_X1 U24022 ( .A(n22409), .ZN(n22659) );
  AOI22_X1 U24023 ( .A1(n22660), .A2(n22490), .B1(n22659), .B2(n22489), .ZN(
        n22415) );
  NOR2_X1 U24024 ( .A1(n22434), .A2(n22476), .ZN(n22438) );
  AOI21_X1 U24025 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22409), .A(n22438), 
        .ZN(n22410) );
  OAI211_X1 U24026 ( .C1(n22413), .C2(n22412), .A(n22411), .B(n22410), .ZN(
        n22661) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22661), .B1(
        n22666), .B2(n22475), .ZN(n22414) );
  OAI211_X1 U24028 ( .C1(n22664), .C2(n22487), .A(n22415), .B(n22414), .ZN(
        P1_U3049) );
  INV_X1 U24029 ( .A(n22416), .ZN(n22425) );
  OAI21_X1 U24030 ( .B1(n22419), .B2(n22418), .A(n22417), .ZN(n22428) );
  NOR2_X1 U24031 ( .A1(n22454), .A2(n22425), .ZN(n22665) );
  AOI21_X1 U24032 ( .B1(n22421), .B2(n22420), .A(n22665), .ZN(n22423) );
  OAI22_X1 U24033 ( .A1(n22476), .A2(n22425), .B1(n22428), .B2(n22423), .ZN(
        n22422) );
  AOI22_X1 U24034 ( .A1(n22667), .A2(n22475), .B1(n22489), .B2(n22665), .ZN(
        n22430) );
  INV_X1 U24035 ( .A(n22423), .ZN(n22427) );
  AOI21_X1 U24036 ( .B1(n22465), .B2(n22425), .A(n22424), .ZN(n22426) );
  OAI21_X1 U24037 ( .B1(n22428), .B2(n22427), .A(n22426), .ZN(n22668) );
  AOI22_X1 U24038 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22666), .B2(n22490), .ZN(n22429) );
  OAI211_X1 U24039 ( .C1(n22671), .C2(n22487), .A(n22430), .B(n22429), .ZN(
        P1_U3057) );
  NOR2_X1 U24040 ( .A1(n22674), .A2(n22465), .ZN(n22432) );
  AOI21_X1 U24041 ( .B1(n22432), .B2(n22431), .A(n22466), .ZN(n22442) );
  INV_X1 U24042 ( .A(n22442), .ZN(n22436) );
  NOR2_X1 U24043 ( .A1(n22433), .A2(n14933), .ZN(n22441) );
  AOI22_X1 U24044 ( .A1(n22674), .A2(n22475), .B1(n22489), .B2(n22672), .ZN(
        n22444) );
  INV_X1 U24045 ( .A(n22672), .ZN(n22439) );
  AOI211_X1 U24046 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22439), .A(n22438), 
        .B(n22480), .ZN(n22440) );
  OAI21_X1 U24047 ( .B1(n22442), .B2(n22441), .A(n22440), .ZN(n22675) );
  AOI22_X1 U24048 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22673), .B2(n22490), .ZN(n22443) );
  OAI211_X1 U24049 ( .C1(n22678), .C2(n22487), .A(n22444), .B(n22443), .ZN(
        P1_U3081) );
  AOI22_X1 U24050 ( .A1(n22489), .A2(n22559), .B1(n22488), .B2(n22558), .ZN(
        n22446) );
  AOI22_X1 U24051 ( .A1(n22561), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22560), .B2(n22490), .ZN(n22445) );
  OAI211_X1 U24052 ( .C1(n22493), .C2(n22684), .A(n22446), .B(n22445), .ZN(
        P1_U3097) );
  NOR3_X1 U24053 ( .A1(n22616), .A2(n22689), .A3(n22465), .ZN(n22447) );
  NOR2_X1 U24054 ( .A1(n22447), .A2(n22466), .ZN(n22462) );
  INV_X1 U24055 ( .A(n22462), .ZN(n22452) );
  AND2_X1 U24056 ( .A1(n22448), .A2(n22468), .ZN(n22461) );
  INV_X1 U24057 ( .A(n22449), .ZN(n22451) );
  NAND2_X1 U24058 ( .A1(n22454), .A2(n22453), .ZN(n22686) );
  OAI22_X1 U24059 ( .A1(n22699), .A2(n22493), .B1(n22455), .B2(n22686), .ZN(
        n22456) );
  INV_X1 U24060 ( .A(n22456), .ZN(n22464) );
  INV_X1 U24061 ( .A(n22457), .ZN(n22459) );
  AOI211_X1 U24062 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22686), .A(n22459), 
        .B(n22458), .ZN(n22460) );
  AOI22_X1 U24063 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22689), .B2(n22490), .ZN(n22463) );
  OAI211_X1 U24064 ( .C1(n22693), .C2(n22487), .A(n22464), .B(n22463), .ZN(
        P1_U3113) );
  NOR2_X1 U24065 ( .A1(n22703), .A2(n22465), .ZN(n22467) );
  AOI21_X1 U24066 ( .B1(n22467), .B2(n22715), .A(n22466), .ZN(n22484) );
  INV_X1 U24067 ( .A(n22484), .ZN(n22473) );
  NOR2_X1 U24068 ( .A1(n22469), .A2(n22468), .ZN(n22483) );
  NOR2_X1 U24069 ( .A1(n22471), .A2(n22470), .ZN(n22472) );
  NOR2_X1 U24070 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22474), .ZN(
        n22700) );
  AOI22_X1 U24071 ( .A1(n22701), .A2(n22475), .B1(n22489), .B2(n22700), .ZN(
        n22486) );
  INV_X1 U24072 ( .A(n22700), .ZN(n22481) );
  AOI21_X1 U24073 ( .B1(n22478), .B2(n22477), .A(n22476), .ZN(n22479) );
  AOI211_X1 U24074 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22481), .A(n22480), 
        .B(n22479), .ZN(n22482) );
  OAI21_X1 U24075 ( .B1(n22484), .B2(n22483), .A(n22482), .ZN(n22704) );
  AOI22_X1 U24076 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22703), .B2(n22490), .ZN(n22485) );
  OAI211_X1 U24077 ( .C1(n22708), .C2(n22487), .A(n22486), .B(n22485), .ZN(
        P1_U3129) );
  AOI22_X1 U24078 ( .A1(n22489), .A2(n22574), .B1(n22488), .B2(n22572), .ZN(
        n22492) );
  AOI22_X1 U24079 ( .A1(n22577), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n22711), .B2(n22490), .ZN(n22491) );
  OAI211_X1 U24080 ( .C1(n22493), .C2(n22725), .A(n22492), .B(n22491), .ZN(
        P1_U3145) );
  AOI22_X1 U24081 ( .A1(n22721), .A2(n22516), .B1(n22653), .B2(n22515), .ZN(
        n22495) );
  AOI22_X1 U24082 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22655), .B1(
        n22654), .B2(n11247), .ZN(n22494) );
  OAI211_X1 U24083 ( .C1(n22658), .C2(n22513), .A(n22495), .B(n22494), .ZN(
        P1_U3034) );
  AOI22_X1 U24084 ( .A1(n22515), .A2(n22547), .B1(n22546), .B2(n22514), .ZN(
        n22497) );
  AOI22_X1 U24085 ( .A1(n22548), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n22654), .B2(n22516), .ZN(n22496) );
  OAI211_X1 U24086 ( .C1(n11246), .C2(n22551), .A(n22497), .B(n22496), .ZN(
        P1_U3042) );
  AOI22_X1 U24087 ( .A1(n22666), .A2(n11247), .B1(n22515), .B2(n22659), .ZN(
        n22499) );
  AOI22_X1 U24088 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22660), .B2(n22516), .ZN(n22498) );
  OAI211_X1 U24089 ( .C1(n22664), .C2(n22513), .A(n22499), .B(n22498), .ZN(
        P1_U3050) );
  AOI22_X1 U24090 ( .A1(n22666), .A2(n22516), .B1(n22665), .B2(n22515), .ZN(
        n22501) );
  AOI22_X1 U24091 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n11247), .ZN(n22500) );
  OAI211_X1 U24092 ( .C1(n22671), .C2(n22513), .A(n22501), .B(n22500), .ZN(
        P1_U3058) );
  AOI22_X1 U24093 ( .A1(n22674), .A2(n11247), .B1(n22515), .B2(n22672), .ZN(
        n22503) );
  AOI22_X1 U24094 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22673), .B2(n22516), .ZN(n22502) );
  OAI211_X1 U24095 ( .C1(n22678), .C2(n22513), .A(n22503), .B(n22502), .ZN(
        P1_U3082) );
  AOI22_X1 U24096 ( .A1(n22515), .A2(n22559), .B1(n22514), .B2(n22558), .ZN(
        n22505) );
  AOI22_X1 U24097 ( .A1(n22561), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22560), .B2(n22516), .ZN(n22504) );
  OAI211_X1 U24098 ( .C1(n11246), .C2(n22684), .A(n22505), .B(n22504), .ZN(
        P1_U3098) );
  OAI22_X1 U24099 ( .A1(n22699), .A2(n11246), .B1(n22506), .B2(n22686), .ZN(
        n22507) );
  INV_X1 U24100 ( .A(n22507), .ZN(n22509) );
  AOI22_X1 U24101 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22689), .B2(n22516), .ZN(n22508) );
  OAI211_X1 U24102 ( .C1(n22693), .C2(n22513), .A(n22509), .B(n22508), .ZN(
        P1_U3114) );
  AOI22_X1 U24103 ( .A1(n22701), .A2(n11247), .B1(n22515), .B2(n22700), .ZN(
        n22512) );
  AOI22_X1 U24104 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22703), .B2(n22516), .ZN(n22511) );
  OAI211_X1 U24105 ( .C1(n22708), .C2(n22513), .A(n22512), .B(n22511), .ZN(
        P1_U3130) );
  AOI22_X1 U24106 ( .A1(n22515), .A2(n22574), .B1(n22514), .B2(n22572), .ZN(
        n22518) );
  AOI22_X1 U24107 ( .A1(n22577), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n22711), .B2(n22516), .ZN(n22517) );
  OAI211_X1 U24108 ( .C1(n11246), .C2(n22725), .A(n22518), .B(n22517), .ZN(
        P1_U3146) );
  AOI22_X1 U24109 ( .A1(n22721), .A2(n22541), .B1(n22653), .B2(n22540), .ZN(
        n22520) );
  AOI22_X1 U24110 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22655), .B1(
        n22654), .B2(n11249), .ZN(n22519) );
  OAI211_X1 U24111 ( .C1(n22658), .C2(n22538), .A(n22520), .B(n22519), .ZN(
        P1_U3035) );
  AOI22_X1 U24112 ( .A1(n22540), .A2(n22547), .B1(n22546), .B2(n22539), .ZN(
        n22522) );
  AOI22_X1 U24113 ( .A1(n22548), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n22654), .B2(n22541), .ZN(n22521) );
  OAI211_X1 U24114 ( .C1(n11248), .C2(n22551), .A(n22522), .B(n22521), .ZN(
        P1_U3043) );
  AOI22_X1 U24115 ( .A1(n22666), .A2(n11249), .B1(n22540), .B2(n22659), .ZN(
        n22524) );
  AOI22_X1 U24116 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22660), .B2(n22541), .ZN(n22523) );
  OAI211_X1 U24117 ( .C1(n22664), .C2(n22538), .A(n22524), .B(n22523), .ZN(
        P1_U3051) );
  AOI22_X1 U24118 ( .A1(n22666), .A2(n22541), .B1(n22665), .B2(n22540), .ZN(
        n22526) );
  AOI22_X1 U24119 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n11249), .ZN(n22525) );
  OAI211_X1 U24120 ( .C1(n22671), .C2(n22538), .A(n22526), .B(n22525), .ZN(
        P1_U3059) );
  AOI22_X1 U24121 ( .A1(n22674), .A2(n11249), .B1(n22540), .B2(n22672), .ZN(
        n22528) );
  AOI22_X1 U24122 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22673), .B2(n22541), .ZN(n22527) );
  OAI211_X1 U24123 ( .C1(n22678), .C2(n22538), .A(n22528), .B(n22527), .ZN(
        P1_U3083) );
  AOI22_X1 U24124 ( .A1(n22540), .A2(n22559), .B1(n22539), .B2(n22558), .ZN(
        n22530) );
  AOI22_X1 U24125 ( .A1(n22561), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22560), .B2(n22541), .ZN(n22529) );
  OAI211_X1 U24126 ( .C1(n11248), .C2(n22684), .A(n22530), .B(n22529), .ZN(
        P1_U3099) );
  OAI22_X1 U24127 ( .A1(n22699), .A2(n11248), .B1(n22531), .B2(n22686), .ZN(
        n22532) );
  INV_X1 U24128 ( .A(n22532), .ZN(n22534) );
  AOI22_X1 U24129 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22689), .B2(n22541), .ZN(n22533) );
  OAI211_X1 U24130 ( .C1(n22693), .C2(n22538), .A(n22534), .B(n22533), .ZN(
        P1_U3115) );
  AOI22_X1 U24131 ( .A1(n22701), .A2(n11249), .B1(n22540), .B2(n22700), .ZN(
        n22537) );
  AOI22_X1 U24132 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22703), .B2(n22541), .ZN(n22536) );
  OAI211_X1 U24133 ( .C1(n22708), .C2(n22538), .A(n22537), .B(n22536), .ZN(
        P1_U3131) );
  AOI22_X1 U24134 ( .A1(n22540), .A2(n22574), .B1(n22539), .B2(n22572), .ZN(
        n22543) );
  AOI22_X1 U24135 ( .A1(n22577), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n22711), .B2(n22541), .ZN(n22542) );
  OAI211_X1 U24136 ( .C1(n11248), .C2(n22725), .A(n22543), .B(n22542), .ZN(
        P1_U3147) );
  AOI22_X1 U24137 ( .A1(n22721), .A2(n22576), .B1(n22653), .B2(n22575), .ZN(
        n22545) );
  AOI22_X1 U24138 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22655), .B1(
        n22654), .B2(n22568), .ZN(n22544) );
  OAI211_X1 U24139 ( .C1(n22658), .C2(n22571), .A(n22545), .B(n22544), .ZN(
        P1_U3036) );
  AOI22_X1 U24140 ( .A1(n22575), .A2(n22547), .B1(n22546), .B2(n22573), .ZN(
        n22550) );
  AOI22_X1 U24141 ( .A1(n22548), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n22654), .B2(n22576), .ZN(n22549) );
  OAI211_X1 U24142 ( .C1(n22580), .C2(n22551), .A(n22550), .B(n22549), .ZN(
        P1_U3044) );
  AOI22_X1 U24143 ( .A1(n22666), .A2(n22568), .B1(n22575), .B2(n22659), .ZN(
        n22553) );
  AOI22_X1 U24144 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22660), .B2(n22576), .ZN(n22552) );
  OAI211_X1 U24145 ( .C1(n22664), .C2(n22571), .A(n22553), .B(n22552), .ZN(
        P1_U3052) );
  AOI22_X1 U24146 ( .A1(n22667), .A2(n22568), .B1(n22575), .B2(n22665), .ZN(
        n22555) );
  AOI22_X1 U24147 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22666), .B2(n22576), .ZN(n22554) );
  OAI211_X1 U24148 ( .C1(n22671), .C2(n22571), .A(n22555), .B(n22554), .ZN(
        P1_U3060) );
  AOI22_X1 U24149 ( .A1(n22673), .A2(n22576), .B1(n22672), .B2(n22575), .ZN(
        n22557) );
  AOI22_X1 U24150 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22568), .B2(n22674), .ZN(n22556) );
  OAI211_X1 U24151 ( .C1(n22678), .C2(n22571), .A(n22557), .B(n22556), .ZN(
        P1_U3084) );
  AOI22_X1 U24152 ( .A1(n22575), .A2(n22559), .B1(n22573), .B2(n22558), .ZN(
        n22563) );
  AOI22_X1 U24153 ( .A1(n22561), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22560), .B2(n22576), .ZN(n22562) );
  OAI211_X1 U24154 ( .C1(n22580), .C2(n22684), .A(n22563), .B(n22562), .ZN(
        P1_U3100) );
  OAI22_X1 U24155 ( .A1(n22699), .A2(n22580), .B1(n22564), .B2(n22686), .ZN(
        n22565) );
  INV_X1 U24156 ( .A(n22565), .ZN(n22567) );
  AOI22_X1 U24157 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22689), .B2(n22576), .ZN(n22566) );
  OAI211_X1 U24158 ( .C1(n22693), .C2(n22571), .A(n22567), .B(n22566), .ZN(
        P1_U3116) );
  AOI22_X1 U24159 ( .A1(n22701), .A2(n22568), .B1(n22575), .B2(n22700), .ZN(
        n22570) );
  AOI22_X1 U24160 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22703), .B2(n22576), .ZN(n22569) );
  OAI211_X1 U24161 ( .C1(n22708), .C2(n22571), .A(n22570), .B(n22569), .ZN(
        P1_U3132) );
  AOI22_X1 U24162 ( .A1(n22575), .A2(n22574), .B1(n22573), .B2(n22572), .ZN(
        n22579) );
  AOI22_X1 U24163 ( .A1(n22577), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n22711), .B2(n22576), .ZN(n22578) );
  OAI211_X1 U24164 ( .C1(n22580), .C2(n22725), .A(n22579), .B(n22578), .ZN(
        P1_U3148) );
  AOI22_X1 U24165 ( .A1(n22721), .A2(n22595), .B1(n22603), .B2(n22653), .ZN(
        n22582) );
  AOI22_X1 U24166 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22654), .B2(n14669), .ZN(n22581) );
  OAI211_X1 U24167 ( .C1(n22658), .C2(n22598), .A(n22582), .B(n22581), .ZN(
        P1_U3037) );
  AOI22_X1 U24168 ( .A1(n22666), .A2(n14669), .B1(n22659), .B2(n22603), .ZN(
        n22584) );
  AOI22_X1 U24169 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22661), .B1(
        n22660), .B2(n22595), .ZN(n22583) );
  OAI211_X1 U24170 ( .C1(n22664), .C2(n22598), .A(n22584), .B(n22583), .ZN(
        P1_U3053) );
  AOI22_X1 U24171 ( .A1(n22666), .A2(n22595), .B1(n22603), .B2(n22665), .ZN(
        n22586) );
  AOI22_X1 U24172 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22667), .B2(n14669), .ZN(n22585) );
  OAI211_X1 U24173 ( .C1(n22671), .C2(n22598), .A(n22586), .B(n22585), .ZN(
        P1_U3061) );
  AOI22_X1 U24174 ( .A1(n22673), .A2(n22595), .B1(n22603), .B2(n22672), .ZN(
        n22588) );
  AOI22_X1 U24175 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22674), .B2(n14669), .ZN(n22587) );
  OAI211_X1 U24176 ( .C1(n22678), .C2(n22598), .A(n22588), .B(n22587), .ZN(
        P1_U3085) );
  AOI22_X1 U24177 ( .A1(n22603), .A2(n22680), .B1(n22602), .B2(n22679), .ZN(
        n22590) );
  AOI22_X1 U24178 ( .A1(n22681), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n22689), .B2(n14669), .ZN(n22589) );
  OAI211_X1 U24179 ( .C1(n22606), .C2(n22684), .A(n22590), .B(n22589), .ZN(
        P1_U3109) );
  INV_X1 U24180 ( .A(n22686), .ZN(n22615) );
  AOI22_X1 U24181 ( .A1(n22689), .A2(n22595), .B1(n22603), .B2(n22615), .ZN(
        n22592) );
  AOI22_X1 U24182 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22616), .B2(n14669), .ZN(n22591) );
  OAI211_X1 U24183 ( .C1(n22693), .C2(n22598), .A(n22592), .B(n22591), .ZN(
        P1_U3117) );
  AOI22_X1 U24184 ( .A1(n22603), .A2(n22695), .B1(n22602), .B2(n22694), .ZN(
        n22594) );
  AOI22_X1 U24185 ( .A1(n22696), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n22703), .B2(n14669), .ZN(n22593) );
  OAI211_X1 U24186 ( .C1(n22606), .C2(n22699), .A(n22594), .B(n22593), .ZN(
        P1_U3125) );
  AOI22_X1 U24187 ( .A1(n22701), .A2(n14669), .B1(n22700), .B2(n22603), .ZN(
        n22597) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22595), .ZN(n22596) );
  OAI211_X1 U24189 ( .C1(n22708), .C2(n22598), .A(n22597), .B(n22596), .ZN(
        P1_U3133) );
  INV_X1 U24190 ( .A(n22599), .ZN(n22710) );
  AOI22_X1 U24191 ( .A1(n22602), .A2(n22710), .B1(n22603), .B2(n22709), .ZN(
        n22601) );
  AOI22_X1 U24192 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n22711), .B2(n14669), .ZN(n22600) );
  OAI211_X1 U24193 ( .C1(n22606), .C2(n22715), .A(n22601), .B(n22600), .ZN(
        P1_U3141) );
  AOI22_X1 U24194 ( .A1(n22603), .A2(n22718), .B1(n22602), .B2(n22716), .ZN(
        n22605) );
  AOI22_X1 U24195 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22721), .B2(n14669), .ZN(n22604) );
  OAI211_X1 U24196 ( .C1(n22606), .C2(n22725), .A(n22605), .B(n22604), .ZN(
        P1_U3157) );
  AOI22_X1 U24197 ( .A1(n22721), .A2(n22620), .B1(n22653), .B2(n22619), .ZN(
        n22608) );
  AOI22_X1 U24198 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22654), .B2(n14557), .ZN(n22607) );
  OAI211_X1 U24199 ( .C1(n22658), .C2(n22623), .A(n22608), .B(n22607), .ZN(
        P1_U3038) );
  AOI22_X1 U24200 ( .A1(n22666), .A2(n14557), .B1(n22659), .B2(n22619), .ZN(
        n22610) );
  AOI22_X1 U24201 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22660), .B2(n22620), .ZN(n22609) );
  OAI211_X1 U24202 ( .C1(n22664), .C2(n22623), .A(n22610), .B(n22609), .ZN(
        P1_U3054) );
  AOI22_X1 U24203 ( .A1(n22666), .A2(n22620), .B1(n22665), .B2(n22619), .ZN(
        n22612) );
  AOI22_X1 U24204 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22667), .B2(n14557), .ZN(n22611) );
  OAI211_X1 U24205 ( .C1(n22671), .C2(n22623), .A(n22612), .B(n22611), .ZN(
        P1_U3062) );
  AOI22_X1 U24206 ( .A1(n22674), .A2(n14557), .B1(n22672), .B2(n22619), .ZN(
        n22614) );
  AOI22_X1 U24207 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22673), .B2(n22620), .ZN(n22613) );
  OAI211_X1 U24208 ( .C1(n22678), .C2(n22623), .A(n22614), .B(n22613), .ZN(
        P1_U3086) );
  AOI22_X1 U24209 ( .A1(n22689), .A2(n22620), .B1(n22615), .B2(n22619), .ZN(
        n22618) );
  AOI22_X1 U24210 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22616), .B2(n14557), .ZN(n22617) );
  OAI211_X1 U24211 ( .C1(n22693), .C2(n22623), .A(n22618), .B(n22617), .ZN(
        P1_U3118) );
  AOI22_X1 U24212 ( .A1(n22701), .A2(n14557), .B1(n22700), .B2(n22619), .ZN(
        n22622) );
  AOI22_X1 U24213 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22703), .B2(n22620), .ZN(n22621) );
  OAI211_X1 U24214 ( .C1(n22708), .C2(n22623), .A(n22622), .B(n22621), .ZN(
        P1_U3134) );
  AOI22_X1 U24215 ( .A1(n22721), .A2(n22641), .B1(n22648), .B2(n22653), .ZN(
        n22625) );
  AOI22_X1 U24216 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n22654), .B2(n22649), .ZN(n22624) );
  OAI211_X1 U24217 ( .C1(n22658), .C2(n22644), .A(n22625), .B(n22624), .ZN(
        P1_U3039) );
  AOI22_X1 U24218 ( .A1(n22660), .A2(n22641), .B1(n22648), .B2(n22659), .ZN(
        n22627) );
  AOI22_X1 U24219 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22666), .B2(n22649), .ZN(n22626) );
  OAI211_X1 U24220 ( .C1(n22664), .C2(n22644), .A(n22627), .B(n22626), .ZN(
        P1_U3055) );
  AOI22_X1 U24221 ( .A1(n22666), .A2(n22641), .B1(n22648), .B2(n22665), .ZN(
        n22629) );
  AOI22_X1 U24222 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22667), .B2(n22649), .ZN(n22628) );
  OAI211_X1 U24223 ( .C1(n22671), .C2(n22644), .A(n22629), .B(n22628), .ZN(
        P1_U3063) );
  AOI22_X1 U24224 ( .A1(n22674), .A2(n22649), .B1(n22672), .B2(n22648), .ZN(
        n22631) );
  AOI22_X1 U24225 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22641), .B2(n22673), .ZN(n22630) );
  OAI211_X1 U24226 ( .C1(n22678), .C2(n22644), .A(n22631), .B(n22630), .ZN(
        P1_U3087) );
  AOI22_X1 U24227 ( .A1(n22648), .A2(n22680), .B1(n22647), .B2(n22679), .ZN(
        n22633) );
  AOI22_X1 U24228 ( .A1(n22681), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n22689), .B2(n22649), .ZN(n22632) );
  OAI211_X1 U24229 ( .C1(n22652), .C2(n22684), .A(n22633), .B(n22632), .ZN(
        P1_U3111) );
  OAI22_X1 U24230 ( .A1(n22699), .A2(n22635), .B1(n22686), .B2(n22634), .ZN(
        n22636) );
  INV_X1 U24231 ( .A(n22636), .ZN(n22638) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22690), .B1(
        n22689), .B2(n22641), .ZN(n22637) );
  OAI211_X1 U24233 ( .C1(n22693), .C2(n22644), .A(n22638), .B(n22637), .ZN(
        P1_U3119) );
  AOI22_X1 U24234 ( .A1(n22648), .A2(n22695), .B1(n22647), .B2(n22694), .ZN(
        n22640) );
  AOI22_X1 U24235 ( .A1(n22696), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n22703), .B2(n22649), .ZN(n22639) );
  OAI211_X1 U24236 ( .C1(n22652), .C2(n22699), .A(n22640), .B(n22639), .ZN(
        P1_U3127) );
  AOI22_X1 U24237 ( .A1(n22701), .A2(n22649), .B1(n22700), .B2(n22648), .ZN(
        n22643) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22641), .ZN(n22642) );
  OAI211_X1 U24239 ( .C1(n22708), .C2(n22644), .A(n22643), .B(n22642), .ZN(
        P1_U3135) );
  AOI22_X1 U24240 ( .A1(n22647), .A2(n22710), .B1(n22648), .B2(n22709), .ZN(
        n22646) );
  AOI22_X1 U24241 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n22711), .B2(n22649), .ZN(n22645) );
  OAI211_X1 U24242 ( .C1(n22652), .C2(n22715), .A(n22646), .B(n22645), .ZN(
        P1_U3143) );
  AOI22_X1 U24243 ( .A1(n22648), .A2(n22718), .B1(n22647), .B2(n22716), .ZN(
        n22651) );
  AOI22_X1 U24244 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n22721), .B2(n22649), .ZN(n22650) );
  OAI211_X1 U24245 ( .C1(n22652), .C2(n22725), .A(n22651), .B(n22650), .ZN(
        P1_U3159) );
  AOI22_X1 U24246 ( .A1(n22721), .A2(n22702), .B1(n22719), .B2(n22653), .ZN(
        n22657) );
  AOI22_X1 U24247 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22654), .B2(n22720), .ZN(n22656) );
  OAI211_X1 U24248 ( .C1(n22658), .C2(n22707), .A(n22657), .B(n22656), .ZN(
        P1_U3040) );
  AOI22_X1 U24249 ( .A1(n22666), .A2(n22720), .B1(n22659), .B2(n22719), .ZN(
        n22663) );
  AOI22_X1 U24250 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22661), .B1(
        n22660), .B2(n22702), .ZN(n22662) );
  OAI211_X1 U24251 ( .C1(n22664), .C2(n22707), .A(n22663), .B(n22662), .ZN(
        P1_U3056) );
  AOI22_X1 U24252 ( .A1(n22666), .A2(n22702), .B1(n22719), .B2(n22665), .ZN(
        n22670) );
  AOI22_X1 U24253 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22667), .B2(n22720), .ZN(n22669) );
  OAI211_X1 U24254 ( .C1(n22671), .C2(n22707), .A(n22670), .B(n22669), .ZN(
        P1_U3064) );
  AOI22_X1 U24255 ( .A1(n22673), .A2(n22702), .B1(n22719), .B2(n22672), .ZN(
        n22677) );
  AOI22_X1 U24256 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22674), .B2(n22720), .ZN(n22676) );
  OAI211_X1 U24257 ( .C1(n22678), .C2(n22707), .A(n22677), .B(n22676), .ZN(
        P1_U3088) );
  AOI22_X1 U24258 ( .A1(n22719), .A2(n22680), .B1(n22717), .B2(n22679), .ZN(
        n22683) );
  AOI22_X1 U24259 ( .A1(n22681), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n22689), .B2(n22720), .ZN(n22682) );
  OAI211_X1 U24260 ( .C1(n22726), .C2(n22684), .A(n22683), .B(n22682), .ZN(
        P1_U3112) );
  OAI22_X1 U24261 ( .A1(n22699), .A2(n22687), .B1(n22686), .B2(n22685), .ZN(
        n22688) );
  INV_X1 U24262 ( .A(n22688), .ZN(n22692) );
  AOI22_X1 U24263 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22690), .B1(
        n22689), .B2(n22702), .ZN(n22691) );
  OAI211_X1 U24264 ( .C1(n22693), .C2(n22707), .A(n22692), .B(n22691), .ZN(
        P1_U3120) );
  AOI22_X1 U24265 ( .A1(n22719), .A2(n22695), .B1(n22717), .B2(n22694), .ZN(
        n22698) );
  AOI22_X1 U24266 ( .A1(n22696), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n22703), .B2(n22720), .ZN(n22697) );
  OAI211_X1 U24267 ( .C1(n22726), .C2(n22699), .A(n22698), .B(n22697), .ZN(
        P1_U3128) );
  AOI22_X1 U24268 ( .A1(n22701), .A2(n22720), .B1(n22700), .B2(n22719), .ZN(
        n22706) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22702), .ZN(n22705) );
  OAI211_X1 U24270 ( .C1(n22708), .C2(n22707), .A(n22706), .B(n22705), .ZN(
        P1_U3136) );
  AOI22_X1 U24271 ( .A1(n22717), .A2(n22710), .B1(n22719), .B2(n22709), .ZN(
        n22714) );
  AOI22_X1 U24272 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n22711), .B2(n22720), .ZN(n22713) );
  OAI211_X1 U24273 ( .C1(n22726), .C2(n22715), .A(n22714), .B(n22713), .ZN(
        P1_U3144) );
  AOI22_X1 U24274 ( .A1(n22719), .A2(n22718), .B1(n22717), .B2(n22716), .ZN(
        n22724) );
  AOI22_X1 U24275 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22721), .B2(n22720), .ZN(n22723) );
  OAI211_X1 U24276 ( .C1(n22726), .C2(n22725), .A(n22724), .B(n22723), .ZN(
        P1_U3160) );
  OAI22_X1 U24277 ( .A1(n20637), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22727), .ZN(n22728) );
  INV_X1 U24278 ( .A(n22728), .ZN(P1_U3486) );
  AND2_X2 U11414 ( .A1(n14304), .A2(n14474), .ZN(n16824) );
  AND2_X1 U11699 ( .A1(n11313), .A2(n16829), .ZN(n11955) );
  INV_X1 U11689 ( .A(n13952), .ZN(n13720) );
  CLKBUF_X2 U12517 ( .A(n13445), .Z(n13890) );
  NAND2_X1 U11309 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21404) );
  NOR2_X2 U11496 ( .A1(n21404), .A2(n20778), .ZN(n15590) );
  CLKBUF_X3 U12592 ( .A(n11176), .Z(n20026) );
  NAND2_X1 U13341 ( .A1(n11907), .A2(n11854), .ZN(n16254) );
  INV_X1 U11463 ( .A(n18511), .ZN(n18619) );
  NAND2_X1 U11723 ( .A1(n13148), .A2(n13147), .ZN(n17785) );
  CLKBUF_X1 U11252 ( .A(n12608), .Z(n11155) );
  CLKBUF_X2 U11254 ( .A(n11444), .Z(n11227) );
  CLKBUF_X1 U11315 ( .A(n11333), .Z(n11168) );
  CLKBUF_X1 U11356 ( .A(n11506), .Z(n11507) );
  CLKBUF_X1 U11358 ( .A(n12066), .Z(n12067) );
  CLKBUF_X1 U11368 ( .A(n16360), .Z(n16401) );
  CLKBUF_X1 U11369 ( .A(n12805), .Z(n13892) );
  NOR2_X2 U11372 ( .A1(n11603), .A2(n11410), .ZN(n16825) );
  CLKBUF_X1 U11376 ( .A(n15827), .Z(n20590) );
  CLKBUF_X1 U11379 ( .A(n16360), .Z(n11221) );
  CLKBUF_X1 U11386 ( .A(n13345), .Z(n13343) );
  CLKBUF_X1 U11390 ( .A(n12565), .Z(n13230) );
  CLKBUF_X1 U11391 ( .A(n17277), .Z(n11188) );
  CLKBUF_X1 U11399 ( .A(n13083), .Z(n12889) );
  CLKBUF_X1 U11401 ( .A(n13072), .Z(n12836) );
  CLKBUF_X1 U11408 ( .A(n12813), .Z(n19860) );
  CLKBUF_X1 U11410 ( .A(n12826), .Z(n19808) );
  CLKBUF_X1 U11416 ( .A(n11588), .Z(n15726) );
  CLKBUF_X1 U11419 ( .A(n11420), .Z(n14622) );
  CLKBUF_X1 U11423 ( .A(n16531), .Z(n16571) );
  XNOR2_X1 U11450 ( .A(n11609), .B(n11608), .ZN(n12074) );
  CLKBUF_X1 U11472 ( .A(n11407), .Z(n14559) );
  CLKBUF_X1 U11494 ( .A(n11232), .Z(n11222) );
  CLKBUF_X1 U11535 ( .A(n17798), .Z(n11193) );
  CLKBUF_X1 U11536 ( .A(n13188), .Z(n17744) );
  NAND2_X1 U11578 ( .A1(n18619), .A2(n18583), .ZN(n18466) );
  CLKBUF_X1 U11611 ( .A(n13592), .Z(n16497) );
  CLKBUF_X1 U11661 ( .A(n12409), .Z(n16490) );
  CLKBUF_X1 U11719 ( .A(n20464), .Z(n21905) );
  CLKBUF_X1 U11726 ( .A(n11788), .Z(n14287) );
  CLKBUF_X1 U11756 ( .A(n15866), .Z(n11158) );
  NAND2_X1 U11759 ( .A1(n11641), .A2(n11630), .ZN(n14759) );
  CLKBUF_X1 U12036 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17687) );
  CLKBUF_X1 U12040 ( .A(n16870), .Z(n11201) );
  CLKBUF_X1 U12068 ( .A(n17876), .Z(n17912) );
  AND2_X1 U12110 ( .A1(n11255), .A2(n11254), .ZN(n17267) );
  CLKBUF_X1 U12131 ( .A(n18812), .Z(n18819) );
  CLKBUF_X1 U12182 ( .A(n20765), .Z(n20774) );
  AOI211_X1 U12233 ( .C1(n21176), .C2(P3_REIP_REG_29__SCAN_IN), .A(n21147), 
        .B(n21146), .ZN(n21148) );
  OR2_X1 U12305 ( .A1(n13313), .A2(n20288), .ZN(n22730) );
  OR2_X1 U12307 ( .A1(n16652), .A2(n16734), .ZN(n22731) );
  CLKBUF_X1 U12309 ( .A(n21886), .Z(n20719) );
endmodule

