

module b21_C_SARLock_k_64_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4244, n4245, n4246, n4249, n4250, n4251, n4252, n4253, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993;

  INV_X1 U4751 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n8588) );
  CLKBUF_X2 U4752 ( .A(n5781), .Z(n8456) );
  OAI22_X1 U4753 ( .A1(n6469), .A2(n7759), .B1(n9864), .B2(n7799), .ZN(n6064)
         );
  CLKBUF_X2 U4754 ( .A(n7649), .Z(n7674) );
  AND2_X2 U4755 ( .A1(n5768), .A2(n5774), .ZN(n5722) );
  OR2_X1 U4756 ( .A1(n5357), .A2(n4872), .ZN(n4873) );
  NAND2_X2 U4757 ( .A1(n5777), .A2(n8964), .ZN(n5798) );
  OR2_X1 U4758 ( .A1(n5672), .A2(n6206), .ZN(n5653) );
  OR2_X1 U4759 ( .A1(n5852), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9462) );
  INV_X1 U4760 ( .A(n9462), .ZN(n4244) );
  INV_X1 U4761 ( .A(n8588), .ZN(n4245) );
  INV_X1 U4762 ( .A(n4245), .ZN(n4246) );
  INV_X1 U4763 ( .A(n4245), .ZN(P1_U3084) );
  NAND3_X1 U4764 ( .A1(n4833), .A2(n4932), .A3(n4832), .ZN(n5173) );
  CLKBUF_X2 U4765 ( .A(n6269), .Z(n7384) );
  AND2_X1 U4766 ( .A1(n5798), .A2(n4619), .ZN(n7385) );
  INV_X1 U4767 ( .A(n6365), .ZN(n6257) );
  CLKBUF_X2 U4768 ( .A(n4919), .Z(n4251) );
  INV_X1 U4770 ( .A(n8013), .ZN(n9838) );
  NAND2_X1 U4771 ( .A1(n4493), .A2(n6860), .ZN(n6906) );
  INV_X1 U4772 ( .A(n6721), .ZN(n9770) );
  INV_X2 U4773 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6206) );
  NAND3_X1 U4774 ( .A1(n4871), .A2(n4594), .A3(n4813), .ZN(n7540) );
  AND4_X1 U4775 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n4927), .ZN(n6565)
         );
  INV_X1 U4776 ( .A(n5396), .ZN(n5426) );
  AND2_X1 U4777 ( .A1(n4723), .A2(n4738), .ZN(n9022) );
  XNOR2_X1 U4778 ( .A(n5652), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U4779 ( .A1(n5640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5642) );
  INV_X1 U4780 ( .A(n6480), .ZN(n7945) );
  INV_X1 U4781 ( .A(n6356), .ZN(n7946) );
  BUF_X1 U4782 ( .A(n6075), .Z(n4250) );
  NAND2_X1 U4783 ( .A1(n5655), .A2(n5654), .ZN(n7534) );
  AND2_X1 U4784 ( .A1(n4846), .A2(n4845), .ZN(n4919) );
  OAI21_X2 U4785 ( .B1(n7908), .B2(n7765), .A(n7766), .ZN(n7808) );
  XNOR2_X2 U4786 ( .A(n5022), .B(n4815), .ZN(n6908) );
  NAND2_X2 U4787 ( .A1(n8411), .A2(n7591), .ZN(n8410) );
  OAI21_X2 U4789 ( .B1(n7536), .B2(n7537), .A(n6249), .ZN(n6297) );
  NOR2_X2 U4790 ( .A1(n8343), .A2(n8034), .ZN(n8188) );
  AOI21_X2 U4791 ( .B1(n8067), .B2(n5376), .A(n5553), .ZN(n8050) );
  XNOR2_X2 U4792 ( .A(n7715), .B(n7713), .ZN(n7920) );
  NAND2_X2 U4793 ( .A1(n7711), .A2(n7710), .ZN(n7715) );
  AOI21_X2 U4794 ( .B1(n7272), .B2(n5142), .A(n4807), .ZN(n8265) );
  NAND4_X4 U4795 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n6414)
         );
  NAND2_X2 U4796 ( .A1(n5781), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5701) );
  XNOR2_X2 U4797 ( .A(n5041), .B(n4816), .ZN(n7025) );
  XNOR2_X2 U4798 ( .A(n5642), .B(n5641), .ZN(n5746) );
  OAI211_X2 U4799 ( .C1(n8664), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6591)
         );
  OR2_X2 U4800 ( .A1(n6445), .A2(n8642), .ZN(n9694) );
  OR2_X2 U4801 ( .A1(n4250), .A2(n8642), .ZN(n6584) );
  NAND2_X2 U4802 ( .A1(n4532), .A2(n4535), .ZN(n8642) );
  XNOR2_X1 U4803 ( .A(n5425), .B(n5424), .ZN(n8665) );
  NAND2_X1 U4804 ( .A1(n5577), .A2(n5576), .ZN(n9825) );
  NAND2_X1 U4805 ( .A1(n7946), .A2(n6349), .ZN(n5454) );
  NAND2_X1 U4806 ( .A1(n6563), .A2(n9829), .ZN(n5577) );
  NAND3_X1 U4807 ( .A1(n4789), .A2(n4886), .A3(n4788), .ZN(n7949) );
  INV_X1 U4808 ( .A(n7540), .ZN(n6349) );
  INV_X4 U4809 ( .A(n7798), .ZN(n7759) );
  INV_X2 U4810 ( .A(n8451), .ZN(n7614) );
  INV_X1 U4811 ( .A(n6644), .ZN(n4249) );
  CLKBUF_X3 U4812 ( .A(n7385), .Z(n8666) );
  BUF_X1 U4813 ( .A(n6112), .Z(n4334) );
  CLKBUF_X2 U4814 ( .A(n4923), .Z(n4924) );
  INV_X4 U4815 ( .A(n7680), .ZN(n8448) );
  XNOR2_X1 U4816 ( .A(n4855), .B(n4854), .ZN(n5623) );
  NOR2_X1 U4817 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5632) );
  AOI21_X1 U4818 ( .B1(n8057), .B2(n8271), .A(n8056), .ZN(n8292) );
  AOI21_X1 U4819 ( .B1(n4366), .B2(n4368), .A(n6759), .ZN(n4365) );
  NOR2_X1 U4820 ( .A1(n8794), .A2(n8793), .ZN(n8862) );
  AOI21_X1 U4821 ( .B1(n4369), .B2(n4367), .A(n5572), .ZN(n4366) );
  AND2_X1 U4822 ( .A1(n4373), .A2(n4370), .ZN(n4369) );
  NAND2_X1 U4823 ( .A1(n4698), .A2(n4699), .ZN(n4700) );
  NAND2_X1 U4824 ( .A1(n4626), .A2(n4625), .ZN(n8132) );
  OAI21_X1 U4825 ( .B1(n4545), .B2(n4544), .A(n8781), .ZN(n8788) );
  AOI22_X2 U4826 ( .A1(n8665), .A2(n5427), .B1(P1_DATAO_REG_31__SCAN_IN), .B2(
        n5426), .ZN(n8288) );
  NAND2_X1 U4827 ( .A1(n4596), .A2(n4595), .ZN(n8206) );
  XNOR2_X1 U4828 ( .A(n5417), .B(n5395), .ZN(n8663) );
  NAND2_X1 U4829 ( .A1(n7718), .A2(n7717), .ZN(n7847) );
  NAND2_X1 U4830 ( .A1(n8032), .A2(n8031), .ZN(n8215) );
  AND2_X1 U4831 ( .A1(n7752), .A2(n7753), .ZN(n4329) );
  NAND2_X1 U4832 ( .A1(n5319), .A2(n5318), .ZN(n8315) );
  NAND2_X1 U4833 ( .A1(n7292), .A2(n7291), .ZN(n7711) );
  NAND2_X1 U4834 ( .A1(n5362), .A2(n5361), .ZN(n4415) );
  XNOR2_X1 U4835 ( .A(n5313), .B(n5308), .ZN(n7313) );
  NAND2_X1 U4836 ( .A1(n6905), .A2(n6904), .ZN(n6907) );
  NAND2_X1 U4837 ( .A1(n5265), .A2(n5264), .ZN(n8327) );
  AOI211_X1 U4838 ( .C1(n4530), .C2(n8710), .A(n8709), .B(n8715), .ZN(n4529)
         );
  NAND2_X1 U4839 ( .A1(n5230), .A2(n5229), .ZN(n8338) );
  OAI21_X1 U4840 ( .B1(n8713), .B2(n8707), .A(n8706), .ZN(n4530) );
  NAND2_X1 U4841 ( .A1(n4420), .A2(n4418), .ZN(n5255) );
  NAND2_X1 U4842 ( .A1(n5112), .A2(n5111), .ZN(n7295) );
  NAND2_X1 U4843 ( .A1(n4416), .A2(n4681), .ZN(n5191) );
  NAND2_X1 U4844 ( .A1(n4417), .A2(n5106), .ZN(n5122) );
  AND2_X1 U4845 ( .A1(n5470), .A2(n5476), .ZN(n6878) );
  OAI211_X1 U4846 ( .C1(n6417), .C2(n4721), .A(n9704), .B(n4720), .ZN(n6588)
         );
  OAI22_X1 U4847 ( .A1(n5843), .A2(n5819), .B1(n9807), .B2(n5879), .ZN(n9609)
         );
  INV_X1 U4848 ( .A(n9887), .ZN(n9829) );
  AND2_X1 U4849 ( .A1(n4818), .A2(n4917), .ZN(n9887) );
  AND4_X2 U4850 ( .A1(n4852), .A2(n4851), .A3(n4850), .A4(n4849), .ZN(n6356)
         );
  NAND2_X1 U4851 ( .A1(n5288), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4851) );
  CLKBUF_X2 U4852 ( .A(n5288), .Z(n4252) );
  AND2_X1 U4853 ( .A1(n4874), .A2(n4873), .ZN(n4878) );
  INV_X1 U4854 ( .A(n5711), .ZN(n7641) );
  INV_X1 U4856 ( .A(n6076), .ZN(n9732) );
  OR2_X1 U4857 ( .A1(n4882), .A2(n5851), .ZN(n4593) );
  OAI211_X1 U4858 ( .C1(n8664), .C2(n5858), .A(n5736), .B(n5735), .ZN(n9693)
         );
  INV_X2 U4859 ( .A(n8664), .ZN(n7463) );
  XNOR2_X1 U4860 ( .A(n4467), .B(n4466), .ZN(n6272) );
  NAND2_X1 U4861 ( .A1(n4679), .A2(n4680), .ZN(n4944) );
  NAND2_X2 U4862 ( .A1(n5623), .A2(n7310), .ZN(n6112) );
  CLKBUF_X1 U4863 ( .A(n7649), .Z(n8445) );
  NAND2_X1 U4864 ( .A1(n4856), .A2(n4859), .ZN(n7310) );
  NAND2_X1 U4865 ( .A1(n4900), .A2(n4899), .ZN(n4339) );
  NAND2_X1 U4866 ( .A1(n4856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4855) );
  INV_X1 U4867 ( .A(n7050), .ZN(n6760) );
  AOI21_X1 U4868 ( .B1(n4607), .B2(n4609), .A(n4992), .ZN(n4606) );
  AND2_X1 U4869 ( .A1(n8396), .A2(n4844), .ZN(n4845) );
  NAND2_X1 U4870 ( .A1(n5677), .A2(n5675), .ZN(n8964) );
  MUX2_X1 U4871 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5653), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5655) );
  XNOR2_X1 U4872 ( .A(n5405), .B(n4836), .ZN(n6928) );
  NAND2_X1 U4873 ( .A1(n5654), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U4874 ( .A1(n5692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U4875 ( .A1(n5432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U4876 ( .A1(n4582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U4877 ( .A(n5647), .B(n5646), .ZN(n7198) );
  NAND2_X1 U4878 ( .A1(n4551), .A2(n5666), .ZN(n5916) );
  NAND2_X2 U4879 ( .A1(n5852), .A2(P1_U3084), .ZN(n9464) );
  INV_X1 U4880 ( .A(n5662), .ZN(n4551) );
  NAND4_X2 U4881 ( .A1(n5633), .A2(n5632), .A3(n6204), .A4(n5631), .ZN(n5667)
         );
  AND2_X1 U4882 ( .A1(n4276), .A2(n5213), .ZN(n4784) );
  AND4_X1 U4883 ( .A1(n4516), .A2(n4515), .A3(n5629), .A4(n4748), .ZN(n5805)
         );
  AND4_X1 U4884 ( .A1(n4830), .A2(n5065), .A3(n5091), .A4(n5153), .ZN(n4832)
         );
  AND4_X1 U4885 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4833)
         );
  INV_X1 U4886 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4834) );
  INV_X1 U4887 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5091) );
  INV_X1 U4888 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5153) );
  INV_X1 U4889 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U4890 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4515) );
  INV_X1 U4891 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5631) );
  NOR2_X1 U4892 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4516) );
  NOR2_X1 U4893 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4830) );
  NOR2_X2 U4894 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4869) );
  NOR2_X1 U4895 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4826) );
  INV_X1 U4896 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5213) );
  INV_X1 U4897 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4854) );
  NOR2_X1 U4898 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4827) );
  NOR2_X1 U4899 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5705) );
  NOR2_X1 U4900 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4828) );
  XNOR2_X1 U4901 ( .A(n5644), .B(n5643), .ZN(n7301) );
  OAI21_X1 U4902 ( .B1(n8727), .B2(n4559), .A(n4557), .ZN(n4556) );
  CLKBUF_X1 U4903 ( .A(n6373), .Z(n4328) );
  NAND2_X1 U4904 ( .A1(n5454), .A2(n6353), .ZN(n6373) );
  NAND2_X1 U4905 ( .A1(n6345), .A2(n6470), .ZN(n5579) );
  NAND4_X1 U4906 ( .A1(n5720), .A2(n5721), .A3(n5719), .A4(n4531), .ZN(n6075)
         );
  XNOR2_X1 U4907 ( .A(n6076), .B(n6414), .ZN(n8807) );
  OR2_X4 U4908 ( .A1(n9921), .A2(n9838), .ZN(n7798) );
  NAND2_X1 U4909 ( .A1(n6356), .A2(n7540), .ZN(n6353) );
  NAND2_X2 U4910 ( .A1(n8103), .A2(n5546), .ZN(n8092) );
  NAND2_X2 U4911 ( .A1(n5342), .A2(n5341), .ZN(n8103) );
  NAND2_X1 U4912 ( .A1(n6355), .A2(n5440), .ZN(n6476) );
  INV_X1 U4913 ( .A(n5357), .ZN(n5288) );
  NAND2_X2 U4914 ( .A1(n8265), .A2(n5500), .ZN(n5169) );
  OAI21_X2 U4915 ( .B1(n6476), .B2(n4918), .A(n5576), .ZN(n9839) );
  NAND2_X2 U4916 ( .A1(n4846), .A2(n8401), .ZN(n4923) );
  INV_X2 U4917 ( .A(n5711), .ZN(n4253) );
  OAI21_X1 U4920 ( .B1(n4529), .B2(n4280), .A(n4524), .ZN(n8717) );
  NAND2_X1 U4921 ( .A1(n9007), .A2(n8777), .ZN(n4544) );
  INV_X1 U4922 ( .A(n8778), .ZN(n4545) );
  AOI21_X1 U4923 ( .B1(n4687), .B2(n4689), .A(n4685), .ZN(n4684) );
  INV_X1 U4924 ( .A(n5170), .ZN(n4685) );
  OR2_X1 U4925 ( .A1(n8298), .A2(n8095), .ZN(n8046) );
  OAI21_X1 U4926 ( .B1(n8829), .B2(n8966), .A(n9199), .ZN(n8850) );
  NAND2_X1 U4927 ( .A1(n5105), .A2(n4817), .ZN(n4417) );
  NAND2_X1 U4928 ( .A1(n5798), .A2(n5852), .ZN(n8664) );
  NOR2_X1 U4929 ( .A1(n5569), .A2(n4397), .ZN(n4396) );
  INV_X1 U4930 ( .A(n5486), .ZN(n4397) );
  OAI21_X1 U4931 ( .B1(n8727), .B2(n8726), .A(n4561), .ZN(n4560) );
  NOR2_X1 U4932 ( .A1(n8730), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U4933 ( .A1(n4563), .A2(n8785), .ZN(n4562) );
  NAND2_X1 U4934 ( .A1(n5548), .A2(n5437), .ZN(n4712) );
  AND2_X1 U4935 ( .A1(n5567), .A2(n4372), .ZN(n4371) );
  NAND2_X1 U4936 ( .A1(n4300), .A2(n4374), .ZN(n4372) );
  AND2_X1 U4937 ( .A1(n4410), .A2(n4815), .ZN(n4409) );
  NAND2_X1 U4938 ( .A1(n5004), .A2(n5006), .ZN(n4410) );
  NAND2_X1 U4939 ( .A1(n4710), .A2(n5558), .ZN(n4709) );
  AOI21_X1 U4940 ( .B1(n4735), .B2(n4734), .A(n4305), .ZN(n4731) );
  AND2_X1 U4941 ( .A1(n4640), .A2(n4639), .ZN(n4638) );
  INV_X1 U4942 ( .A(n9024), .ZN(n4639) );
  OR2_X1 U4943 ( .A1(n9227), .A2(n9027), .ZN(n7527) );
  INV_X1 U4944 ( .A(n9044), .ZN(n8603) );
  NOR2_X1 U4945 ( .A1(n8814), .A2(n4758), .ZN(n4757) );
  INV_X1 U4946 ( .A(n7189), .ZN(n4758) );
  AND2_X1 U4947 ( .A1(n7218), .A2(n9125), .ZN(n5767) );
  AOI21_X1 U4948 ( .B1(n5749), .B2(n5875), .A(n5876), .ZN(n6399) );
  INV_X1 U4949 ( .A(n4432), .ZN(n4431) );
  OAI21_X1 U4950 ( .B1(n4435), .B2(n4433), .A(n5325), .ZN(n4432) );
  NOR2_X2 U4951 ( .A1(n5667), .A2(n5637), .ZN(n5638) );
  AOI21_X1 U4952 ( .B1(n4422), .B2(n4424), .A(n4419), .ZN(n4418) );
  INV_X1 U4953 ( .A(n5246), .ZN(n4419) );
  AOI21_X1 U4954 ( .B1(n4684), .B2(n4686), .A(n4682), .ZN(n4681) );
  NAND2_X1 U4955 ( .A1(n5122), .A2(n4684), .ZN(n4416) );
  INV_X1 U4956 ( .A(n5172), .ZN(n4682) );
  NAND2_X1 U4957 ( .A1(n7559), .A2(n4591), .ZN(n7292) );
  AND2_X1 U4958 ( .A1(n7253), .A2(n7252), .ZN(n4591) );
  NAND2_X1 U4959 ( .A1(n6735), .A2(n4590), .ZN(n6830) );
  AND2_X1 U4960 ( .A1(n6740), .A2(n6734), .ZN(n4590) );
  OR2_X1 U4961 ( .A1(n6123), .A2(n6122), .ZN(n4451) );
  NAND2_X1 U4962 ( .A1(n4713), .A2(n8045), .ZN(n4604) );
  OR2_X1 U4963 ( .A1(n5306), .A2(n8038), .ZN(n5536) );
  NAND2_X1 U4964 ( .A1(n4623), .A2(n4620), .ZN(n8245) );
  AND2_X1 U4965 ( .A1(n8246), .A2(n4264), .ZN(n4620) );
  AND2_X1 U4966 ( .A1(n7265), .A2(n5490), .ZN(n4800) );
  NAND2_X1 U4967 ( .A1(n4610), .A2(n4612), .ZN(n7266) );
  AOI21_X1 U4968 ( .B1(n7144), .B2(n4611), .A(n4614), .ZN(n4612) );
  AND2_X1 U4969 ( .A1(n6568), .A2(n6599), .ZN(n6569) );
  NOR2_X1 U4970 ( .A1(n9831), .A2(n9897), .ZN(n6607) );
  CLKBUF_X1 U4971 ( .A(n5623), .Z(n5624) );
  INV_X1 U4972 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4783) );
  AND2_X1 U4973 ( .A1(n8504), .A2(n7609), .ZN(n4673) );
  OR2_X1 U4974 ( .A1(n7451), .A2(n7450), .ZN(n7469) );
  NOR2_X1 U4975 ( .A1(n8783), .A2(n8782), .ZN(n8794) );
  NAND2_X1 U4976 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  AOI21_X1 U4977 ( .B1(n9068), .B2(n4742), .A(n4320), .ZN(n4741) );
  NOR2_X1 U4978 ( .A1(n9120), .A2(n7485), .ZN(n9135) );
  NAND2_X1 U4979 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  INV_X1 U4980 ( .A(n7198), .ZN(n4718) );
  INV_X1 U4981 ( .A(n7301), .ZN(n4719) );
  INV_X1 U4982 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U4983 ( .A1(n4683), .A2(n4687), .ZN(n5171) );
  NAND2_X1 U4984 ( .A1(n5122), .A2(n4690), .ZN(n4683) );
  NAND2_X1 U4985 ( .A1(n8444), .A2(n8443), .ZN(n9214) );
  NAND2_X1 U4986 ( .A1(n9460), .A2(n7463), .ZN(n8444) );
  OR2_X1 U4987 ( .A1(n8465), .A2(n8596), .ZN(n4495) );
  OAI21_X1 U4988 ( .B1(n4824), .B2(n5468), .A(n5467), .ZN(n5479) );
  NOR2_X1 U4989 ( .A1(n5464), .A2(n5437), .ZN(n5468) );
  NAND2_X1 U4990 ( .A1(n4358), .A2(n5535), .ZN(n4357) );
  OAI21_X1 U4991 ( .B1(n4361), .B2(n5480), .A(n4359), .ZN(n4358) );
  NOR2_X1 U4992 ( .A1(n4360), .A2(n4317), .ZN(n4359) );
  AOI21_X1 U4993 ( .B1(n5479), .B2(n4363), .A(n4362), .ZN(n4361) );
  NAND2_X1 U4994 ( .A1(n5477), .A2(n5569), .ZN(n4356) );
  INV_X1 U4995 ( .A(n4398), .ZN(n4393) );
  NAND2_X1 U4996 ( .A1(n4396), .A2(n5485), .ZN(n4390) );
  NAND2_X1 U4997 ( .A1(n4398), .A2(n5488), .ZN(n4391) );
  NOR2_X1 U4998 ( .A1(n5495), .A2(n5494), .ZN(n4395) );
  AND2_X1 U4999 ( .A1(n4386), .A2(n4385), .ZN(n5504) );
  AND2_X1 U5000 ( .A1(n8274), .A2(n5499), .ZN(n4394) );
  OAI21_X1 U5001 ( .B1(n4528), .B2(n4526), .A(n4525), .ZN(n4524) );
  NOR2_X1 U5002 ( .A1(n8715), .A2(n8785), .ZN(n4525) );
  NAND2_X1 U5003 ( .A1(n4318), .A2(n4527), .ZN(n4526) );
  NOR2_X1 U5004 ( .A1(n8713), .A2(n8712), .ZN(n4528) );
  OR2_X1 U5005 ( .A1(n8726), .A2(n8723), .ZN(n4559) );
  NOR2_X1 U5006 ( .A1(n4668), .A2(n4558), .ZN(n4557) );
  NOR2_X1 U5007 ( .A1(n8743), .A2(n8742), .ZN(n4555) );
  AOI21_X1 U5008 ( .B1(n5528), .B2(n4347), .A(n8159), .ZN(n4346) );
  NOR2_X1 U5009 ( .A1(n5535), .A2(n4348), .ZN(n4347) );
  INV_X1 U5010 ( .A(n5527), .ZN(n4348) );
  AOI21_X1 U5011 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n5514) );
  NOR2_X1 U5012 ( .A1(n5523), .A2(n5512), .ZN(n4353) );
  NAND2_X1 U5013 ( .A1(n4711), .A2(n5546), .ZN(n4380) );
  NOR2_X1 U5014 ( .A1(n4382), .A2(n4288), .ZN(n4381) );
  NOR2_X1 U5015 ( .A1(n4274), .A2(n4383), .ZN(n4382) );
  INV_X1 U5016 ( .A(n5559), .ZN(n4377) );
  NAND2_X1 U5017 ( .A1(n4371), .A2(n4375), .ZN(n4370) );
  INV_X1 U5018 ( .A(n5566), .ZN(n4373) );
  INV_X1 U5019 ( .A(n8543), .ZN(n4513) );
  AND2_X1 U5020 ( .A1(n5649), .A2(n5646), .ZN(n4762) );
  NOR2_X1 U5021 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5649) );
  INV_X1 U5022 ( .A(n4687), .ZN(n4686) );
  INV_X1 U5023 ( .A(SI_13_), .ZN(n5087) );
  AND2_X1 U5024 ( .A1(n7829), .A2(n4581), .ZN(n4580) );
  INV_X1 U5025 ( .A(n7740), .ZN(n4578) );
  INV_X1 U5026 ( .A(n6928), .ZN(n6053) );
  OR2_X1 U5027 ( .A1(n7985), .A2(n4324), .ZN(n4448) );
  NOR2_X1 U5028 ( .A1(n8290), .A2(n8298), .ZN(n4487) );
  INV_X1 U5029 ( .A(n5536), .ZN(n4781) );
  OAI21_X1 U5030 ( .B1(n5307), .B2(n4781), .A(n8121), .ZN(n4780) );
  NOR2_X1 U5031 ( .A1(n8175), .A2(n4634), .ZN(n4633) );
  INV_X1 U5032 ( .A(n4811), .ZN(n4634) );
  OR2_X1 U5033 ( .A1(n8327), .A2(n7890), .ZN(n5525) );
  AND2_X1 U5034 ( .A1(n5272), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U5035 ( .A1(n4795), .A2(n4796), .ZN(n4794) );
  NOR2_X1 U5036 ( .A1(n4768), .A2(n4765), .ZN(n4764) );
  NOR2_X1 U5037 ( .A1(n4471), .A2(n6824), .ZN(n4470) );
  INV_X1 U5038 ( .A(n4472), .ZN(n4471) );
  NAND2_X1 U5039 ( .A1(n9887), .A2(n7944), .ZN(n5576) );
  NAND2_X1 U5040 ( .A1(n6055), .A2(n6346), .ZN(n5578) );
  OR2_X1 U5041 ( .A1(n4885), .A2(n6272), .ZN(n4916) );
  INV_X1 U5042 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4838) );
  AND2_X1 U5043 ( .A1(n7108), .A2(n4707), .ZN(n4706) );
  INV_X1 U5044 ( .A(n7067), .ZN(n4705) );
  NAND2_X1 U5045 ( .A1(n8787), .A2(n8786), .ZN(n8792) );
  NOR2_X1 U5046 ( .A1(n9203), .A2(n8988), .ZN(n8829) );
  AND2_X1 U5047 ( .A1(n9199), .A2(n8966), .ZN(n8828) );
  INV_X1 U5048 ( .A(n7534), .ZN(n5656) );
  OR2_X1 U5049 ( .A1(n9214), .A2(n9217), .ZN(n4458) );
  INV_X1 U5050 ( .A(n4663), .ZN(n4660) );
  INV_X1 U5051 ( .A(n4661), .ZN(n4659) );
  NOR2_X1 U5052 ( .A1(n8975), .A2(n4662), .ZN(n4661) );
  NOR2_X1 U5053 ( .A1(n4732), .A2(n4728), .ZN(n4727) );
  INV_X1 U5054 ( .A(n7435), .ZN(n4728) );
  AND2_X1 U5055 ( .A1(n9008), .A2(n8776), .ZN(n8826) );
  NAND2_X1 U5056 ( .A1(n4260), .A2(n4292), .ZN(n4734) );
  NAND2_X1 U5057 ( .A1(n4260), .A2(n4736), .ZN(n4735) );
  NOR2_X1 U5058 ( .A1(n9244), .A2(n4463), .ZN(n4462) );
  INV_X1 U5059 ( .A(n4464), .ZN(n4463) );
  NOR2_X1 U5060 ( .A1(n9248), .A2(n9253), .ZN(n4464) );
  NAND2_X1 U5061 ( .A1(n4653), .A2(n8711), .ZN(n4647) );
  NAND2_X1 U5062 ( .A1(n9513), .A2(n7483), .ZN(n4654) );
  NAND2_X1 U5063 ( .A1(n8808), .A2(n6622), .ZN(n4746) );
  NOR2_X1 U5064 ( .A1(n7523), .A2(n4458), .ZN(n9013) );
  INV_X1 U5065 ( .A(SI_15_), .ZN(n9321) );
  NOR2_X1 U5066 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  AND2_X1 U5067 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  NAND2_X1 U5068 ( .A1(n5386), .A2(n5385), .ZN(n5394) );
  NOR2_X1 U5069 ( .A1(n5312), .A2(n4436), .ZN(n4435) );
  INV_X1 U5070 ( .A(n5298), .ZN(n4436) );
  NOR2_X1 U5071 ( .A1(n5222), .A2(n4426), .ZN(n4425) );
  INV_X1 U5072 ( .A(n5208), .ZN(n4426) );
  AND2_X1 U5073 ( .A1(n5246), .A2(n5228), .ZN(n5244) );
  NAND2_X1 U5074 ( .A1(n5206), .A2(n5205), .ZN(n4715) );
  INV_X1 U5075 ( .A(n5120), .ZN(n4691) );
  AND2_X1 U5076 ( .A1(n6205), .A2(n6204), .ZN(n6210) );
  AOI21_X1 U5077 ( .B1(n4404), .B2(n4407), .A(n4402), .ZN(n4401) );
  AOI21_X1 U5078 ( .B1(n4409), .B2(n4406), .A(n4405), .ZN(n4404) );
  INV_X1 U5079 ( .A(n5023), .ZN(n4405) );
  INV_X1 U5080 ( .A(n5006), .ZN(n4406) );
  INV_X1 U5081 ( .A(n4409), .ZN(n4407) );
  INV_X1 U5082 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4341) );
  INV_X1 U5083 ( .A(n6843), .ZN(n4576) );
  INV_X1 U5084 ( .A(n6998), .ZN(n4574) );
  INV_X1 U5085 ( .A(n6838), .ZN(n4575) );
  AND4_X1 U5086 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n8038)
         );
  AND4_X1 U5087 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n8030)
         );
  AND4_X1 U5088 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n7275)
         );
  INV_X1 U5089 ( .A(n5398), .ZN(n5408) );
  OAI21_X1 U5090 ( .B1(n4923), .B2(n4792), .A(n4786), .ZN(n4790) );
  NAND2_X1 U5091 ( .A1(n4787), .A2(n4848), .ZN(n4786) );
  AND2_X1 U5092 ( .A1(n8401), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4787) );
  OR2_X1 U5093 ( .A1(n6146), .A2(n6145), .ZN(n4446) );
  XNOR2_X1 U5094 ( .A(n4448), .B(n8007), .ZN(n7987) );
  INV_X1 U5095 ( .A(n8288), .ZN(n4484) );
  INV_X1 U5096 ( .A(n4485), .ZN(n4481) );
  NOR2_X1 U5097 ( .A1(n8023), .A2(n4486), .ZN(n4485) );
  INV_X1 U5098 ( .A(n4487), .ZN(n4486) );
  OR2_X1 U5099 ( .A1(n5367), .A2(n7803), .ZN(n8058) );
  INV_X1 U5100 ( .A(n8046), .ZN(n4603) );
  INV_X1 U5101 ( .A(n8045), .ZN(n4605) );
  AND2_X1 U5102 ( .A1(n8046), .A2(n5375), .ZN(n8072) );
  AND2_X1 U5103 ( .A1(n8125), .A2(n8114), .ZN(n8109) );
  AND2_X1 U5104 ( .A1(n8109), .A2(n8091), .ZN(n8086) );
  OR2_X1 U5105 ( .A1(n8315), .A2(n8041), .ZN(n8042) );
  OR2_X1 U5106 ( .A1(n5320), .A2(n9346), .ZN(n5336) );
  NAND2_X1 U5107 ( .A1(n8139), .A2(n5307), .ZN(n8138) );
  INV_X1 U5108 ( .A(n4631), .ZN(n4630) );
  OAI22_X1 U5109 ( .A1(n8175), .A2(n4632), .B1(n8195), .B2(n8327), .ZN(n4631)
         );
  NAND2_X1 U5110 ( .A1(n4811), .A2(n8035), .ZN(n4632) );
  NAND2_X1 U5111 ( .A1(n8188), .A2(n4633), .ZN(n4629) );
  INV_X1 U5112 ( .A(n8203), .ZN(n8182) );
  AND2_X1 U5113 ( .A1(n5525), .A2(n5527), .ZN(n8175) );
  INV_X1 U5114 ( .A(n8175), .ZN(n8167) );
  OR2_X1 U5115 ( .A1(n8018), .A2(n8182), .ZN(n4811) );
  AND2_X1 U5116 ( .A1(n8338), .A2(n8224), .ZN(n8034) );
  INV_X1 U5117 ( .A(n4772), .ZN(n4771) );
  OAI21_X1 U5118 ( .B1(n4774), .B2(n4258), .A(n5203), .ZN(n4772) );
  NOR2_X1 U5119 ( .A1(n5503), .A2(n4775), .ZN(n4774) );
  INV_X1 U5120 ( .A(n5506), .ZN(n4775) );
  NAND2_X1 U5121 ( .A1(n5169), .A2(n4258), .ZN(n4770) );
  NOR2_X1 U5122 ( .A1(n8274), .A2(n4622), .ZN(n4621) );
  INV_X1 U5123 ( .A(n4624), .ZN(n4622) );
  AND2_X1 U5124 ( .A1(n5501), .A2(n5500), .ZN(n8274) );
  OR2_X1 U5125 ( .A1(n7151), .A2(n8373), .ZN(n7232) );
  AND2_X1 U5126 ( .A1(n7144), .A2(n4615), .ZN(n4613) );
  OR2_X1 U5127 ( .A1(n7556), .A2(n7937), .ZN(n4615) );
  OR2_X1 U5128 ( .A1(n7140), .A2(n7139), .ZN(n4616) );
  AND2_X1 U5129 ( .A1(n5491), .A2(n5490), .ZN(n7141) );
  AND2_X1 U5130 ( .A1(n5487), .A2(n5486), .ZN(n7139) );
  AND2_X1 U5131 ( .A1(n6786), .A2(n6784), .ZN(n4597) );
  AND2_X1 U5132 ( .A1(n6567), .A2(n6566), .ZN(n6599) );
  NAND2_X1 U5133 ( .A1(n4468), .A2(n4266), .ZN(n9831) );
  INV_X1 U5134 ( .A(n9830), .ZN(n4468) );
  INV_X1 U5135 ( .A(n8266), .ZN(n8181) );
  INV_X1 U5136 ( .A(n8271), .ZN(n9842) );
  INV_X1 U5137 ( .A(n7949), .ZN(n4888) );
  OR2_X1 U5138 ( .A1(n9921), .A2(n8013), .ZN(n6752) );
  INV_X1 U5139 ( .A(n8179), .ZN(n8268) );
  NAND2_X1 U5140 ( .A1(n5333), .A2(n5332), .ZN(n8310) );
  OR2_X1 U5141 ( .A1(n5396), .A2(n7304), .ZN(n5332) );
  NOR2_X1 U5142 ( .A1(n8206), .A2(n8205), .ZN(n8343) );
  INV_X1 U5143 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5144 ( .A1(n5620), .A2(n5611), .ZN(n6250) );
  OR2_X1 U5145 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  XNOR2_X1 U5146 ( .A(n5434), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U5147 ( .A1(n4835), .A2(n4784), .ZN(n5433) );
  INV_X1 U5148 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4785) );
  INV_X1 U5149 ( .A(n5173), .ZN(n4835) );
  AND2_X1 U5150 ( .A1(n5031), .A2(n5044), .ZN(n6316) );
  INV_X1 U5151 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4987) );
  INV_X1 U5152 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4931) );
  INV_X1 U5153 ( .A(n7068), .ZN(n4707) );
  XNOR2_X1 U5154 ( .A(n5710), .B(n8448), .ZN(n5715) );
  OR2_X1 U5155 ( .A1(n8524), .A2(n7648), .ZN(n4702) );
  INV_X1 U5156 ( .A(n8552), .ZN(n4506) );
  NOR2_X1 U5157 ( .A1(n4504), .A2(n8521), .ZN(n4503) );
  NOR2_X1 U5158 ( .A1(n8436), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U5159 ( .A1(n4672), .A2(n4293), .ZN(n7624) );
  AND2_X1 U5160 ( .A1(n4503), .A2(n4500), .ZN(n4498) );
  OR2_X1 U5161 ( .A1(n4505), .A2(n4501), .ZN(n4500) );
  AND2_X1 U5162 ( .A1(n7623), .A2(n4506), .ZN(n4501) );
  AOI21_X1 U5163 ( .B1(n4701), .B2(n7648), .A(n4294), .ZN(n4699) );
  NOR2_X1 U5164 ( .A1(n8854), .A2(n9125), .ZN(n8832) );
  NAND2_X1 U5165 ( .A1(n5668), .A2(n5669), .ZN(n4521) );
  AND3_X1 U5166 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(n7656) );
  OR2_X1 U5167 ( .A1(n9217), .A2(n9011), .ZN(n9008) );
  NAND2_X1 U5168 ( .A1(n8779), .A2(n8780), .ZN(n9004) );
  INV_X1 U5169 ( .A(n8826), .ZN(n8975) );
  NOR2_X1 U5170 ( .A1(n7513), .A2(n8765), .ZN(n7528) );
  AND2_X1 U5171 ( .A1(n9036), .A2(n8520), .ZN(n9028) );
  INV_X1 U5172 ( .A(n9074), .ZN(n4643) );
  NAND2_X1 U5173 ( .A1(n4306), .A2(n8601), .ZN(n4640) );
  NAND2_X1 U5174 ( .A1(n9068), .A2(n8750), .ZN(n4645) );
  OR2_X1 U5175 ( .A1(n8803), .A2(n8802), .ZN(n9042) );
  NAND2_X1 U5176 ( .A1(n9074), .A2(n9075), .ZN(n9073) );
  AND2_X1 U5177 ( .A1(n9115), .A2(n9112), .ZN(n9107) );
  NAND2_X1 U5178 ( .A1(n9100), .A2(n4809), .ZN(n9084) );
  NAND2_X1 U5179 ( .A1(n9084), .A2(n9083), .ZN(n9082) );
  INV_X1 U5180 ( .A(n9137), .ZN(n9105) );
  AND2_X1 U5181 ( .A1(n4670), .A2(n8619), .ZN(n4669) );
  INV_X1 U5182 ( .A(n9103), .ZN(n4670) );
  OR2_X1 U5183 ( .A1(n9134), .A2(n8725), .ZN(n4671) );
  NAND2_X1 U5184 ( .A1(n9148), .A2(n9156), .ZN(n4753) );
  NOR2_X1 U5185 ( .A1(n9135), .A2(n4752), .ZN(n4751) );
  INV_X1 U5186 ( .A(n4808), .ZN(n4752) );
  NAND2_X1 U5187 ( .A1(n9531), .A2(n4275), .ZN(n7190) );
  INV_X1 U5188 ( .A(n4756), .ZN(n7351) );
  AND2_X1 U5189 ( .A1(n8678), .A2(n8677), .ZN(n8808) );
  OR2_X1 U5190 ( .A1(n6810), .A2(n8808), .ZN(n6812) );
  NAND2_X1 U5191 ( .A1(n6638), .A2(n8835), .ZN(n6639) );
  NAND2_X1 U5192 ( .A1(n6440), .A2(n6421), .ZN(n8645) );
  NAND2_X1 U5193 ( .A1(n5976), .A2(n8866), .ZN(n9687) );
  AND2_X1 U5194 ( .A1(n5913), .A2(n9574), .ZN(n6437) );
  NAND2_X1 U5195 ( .A1(n6438), .A2(n8807), .ZN(n6440) );
  INV_X1 U5196 ( .A(n9687), .ZN(n9702) );
  INV_X1 U5197 ( .A(n9208), .ZN(n4440) );
  NAND2_X1 U5198 ( .A1(n9209), .A2(n9777), .ZN(n4439) );
  NAND2_X1 U5199 ( .A1(n7449), .A2(n7448), .ZN(n9222) );
  NAND2_X1 U5200 ( .A1(n7438), .A2(n7437), .ZN(n9227) );
  NAND2_X1 U5201 ( .A1(n7387), .A2(n7386), .ZN(n9259) );
  NAND2_X1 U5202 ( .A1(n7365), .A2(n7364), .ZN(n9279) );
  NAND2_X1 U5203 ( .A1(n7355), .A2(n7354), .ZN(n9286) );
  INV_X1 U5204 ( .A(n9784), .ZN(n9777) );
  NAND2_X1 U5205 ( .A1(n5346), .A2(n5345), .ZN(n5362) );
  MUX2_X1 U5206 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4825), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5677) );
  NOR2_X1 U5207 ( .A1(n4548), .A2(n5662), .ZN(n5676) );
  XNOR2_X1 U5208 ( .A(n5362), .B(n5361), .ZN(n7464) );
  AND2_X1 U5209 ( .A1(n5630), .A2(n5639), .ZN(n4547) );
  OAI21_X1 U5210 ( .B1(n5275), .B2(n5274), .A(n5273), .ZN(n5297) );
  AND2_X1 U5211 ( .A1(n5298), .A2(n5280), .ZN(n5296) );
  XNOR2_X1 U5212 ( .A(n5255), .B(n5256), .ZN(n7404) );
  NOR2_X1 U5213 ( .A1(n5665), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5666) );
  INV_X1 U5214 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5664) );
  AOI21_X1 U5215 ( .B1(n4933), .B2(n4307), .A(n4304), .ZN(n4680) );
  INV_X1 U5216 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4748) );
  XNOR2_X1 U5217 ( .A(n4934), .B(SI_4_), .ZN(n4933) );
  INV_X1 U5218 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5628) );
  XNOR2_X1 U5219 ( .A(n4912), .B(SI_3_), .ZN(n4911) );
  INV_X1 U5220 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4517) );
  AND4_X1 U5221 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n7552)
         );
  NAND2_X1 U5222 ( .A1(n7248), .A2(n7247), .ZN(n7559) );
  NAND2_X1 U5223 ( .A1(n5159), .A2(n5158), .ZN(n8360) );
  NAND2_X1 U5224 ( .A1(n4694), .A2(n5299), .ZN(n5306) );
  NAND2_X1 U5225 ( .A1(n7313), .A2(n5427), .ZN(n4694) );
  NAND2_X1 U5226 ( .A1(n6043), .A2(n8250), .ZN(n7889) );
  AND4_X1 U5227 ( .A1(n5221), .A2(n5220), .A3(n5219), .A4(n5218), .ZN(n8033)
         );
  NAND2_X1 U5228 ( .A1(n6553), .A2(n6525), .ZN(n6735) );
  NAND2_X1 U5229 ( .A1(n7910), .A2(n7911), .ZN(n4332) );
  INV_X1 U5230 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5231 ( .A(n9850), .ZN(n6332) );
  AND2_X1 U5232 ( .A1(n6771), .A2(n8013), .ZN(n6048) );
  AND2_X1 U5233 ( .A1(n5625), .A2(n6046), .ZN(n8266) );
  INV_X1 U5234 ( .A(n8038), .ZN(n8162) );
  INV_X1 U5235 ( .A(n8030), .ZN(n8242) );
  INV_X1 U5236 ( .A(n7275), .ZN(n8243) );
  INV_X1 U5237 ( .A(n7851), .ZN(n8267) );
  INV_X1 U5238 ( .A(n7258), .ZN(n7937) );
  INV_X1 U5239 ( .A(n6896), .ZN(n7940) );
  NOR2_X1 U5240 ( .A1(n6155), .A2(n4447), .ZN(n6146) );
  AND2_X1 U5241 ( .A1(n6102), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4447) );
  NOR2_X1 U5242 ( .A1(n6133), .A2(n4316), .ZN(n6123) );
  NOR2_X1 U5243 ( .A1(n6168), .A2(n6167), .ZN(n6166) );
  NOR2_X1 U5244 ( .A1(n6215), .A2(n4452), .ZN(n6219) );
  AND2_X1 U5245 ( .A1(n6216), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4452) );
  NOR2_X1 U5246 ( .A1(n6219), .A2(n6218), .ZN(n6315) );
  NAND2_X1 U5247 ( .A1(n5178), .A2(n5177), .ZN(n8355) );
  INV_X1 U5248 ( .A(n8250), .ZN(n9834) );
  AND2_X1 U5249 ( .A1(n5845), .A2(n5797), .ZN(n5840) );
  INV_X1 U5250 ( .A(n9076), .ZN(n9106) );
  AND2_X1 U5251 ( .A1(n5789), .A2(n5765), .ZN(n9576) );
  INV_X1 U5252 ( .A(n9138), .ZN(n9171) );
  NAND2_X1 U5253 ( .A1(n7458), .A2(n7457), .ZN(n8875) );
  NAND2_X1 U5254 ( .A1(n7446), .A2(n7445), .ZN(n8876) );
  NAND2_X1 U5255 ( .A1(n7330), .A2(n7329), .ZN(n9044) );
  OR2_X1 U5256 ( .A1(n9030), .A2(n4249), .ZN(n7330) );
  INV_X1 U5257 ( .A(n7656), .ZN(n9077) );
  OR2_X1 U5258 ( .A1(n9019), .A2(n8986), .ZN(n4805) );
  NAND2_X1 U5259 ( .A1(n4441), .A2(n8990), .ZN(n9207) );
  NAND2_X1 U5260 ( .A1(n4442), .A2(n9707), .ZN(n4441) );
  NAND2_X1 U5261 ( .A1(n7315), .A2(n7314), .ZN(n9234) );
  NAND2_X1 U5262 ( .A1(n7385), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4535) );
  AND2_X1 U5263 ( .A1(n4536), .A2(n4533), .ZN(n4532) );
  AND2_X1 U5264 ( .A1(n5751), .A2(n5750), .ZN(n7223) );
  MUX2_X1 U5265 ( .A(n5439), .B(n5438), .S(n5569), .Z(n5458) );
  AND2_X1 U5266 ( .A1(n6878), .A2(n5469), .ZN(n4363) );
  INV_X1 U5267 ( .A(n5470), .ZN(n4362) );
  INV_X1 U5268 ( .A(n7096), .ZN(n4360) );
  NOR2_X1 U5269 ( .A1(n5483), .A2(n5482), .ZN(n5489) );
  NAND2_X1 U5270 ( .A1(n4357), .A2(n4356), .ZN(n5483) );
  NOR2_X1 U5271 ( .A1(n4389), .A2(n4301), .ZN(n4387) );
  INV_X1 U5272 ( .A(n4395), .ZN(n4389) );
  INV_X1 U5273 ( .A(n4396), .ZN(n4392) );
  NAND2_X1 U5274 ( .A1(n4395), .A2(n4295), .ZN(n4388) );
  NAND2_X1 U5275 ( .A1(n8714), .A2(n9184), .ZN(n4527) );
  NAND2_X1 U5276 ( .A1(n5509), .A2(n4291), .ZN(n5517) );
  OR2_X1 U5277 ( .A1(n8725), .A2(n8785), .ZN(n4558) );
  INV_X1 U5278 ( .A(n8729), .ZN(n4563) );
  NAND2_X1 U5279 ( .A1(n4355), .A2(n8201), .ZN(n4354) );
  NAND2_X1 U5280 ( .A1(n5517), .A2(n5510), .ZN(n4355) );
  OR2_X1 U5281 ( .A1(n5519), .A2(n8174), .ZN(n4352) );
  AND2_X1 U5282 ( .A1(n4554), .A2(n4552), .ZN(n8755) );
  NOR2_X1 U5283 ( .A1(n8745), .A2(n4553), .ZN(n4552) );
  OR2_X1 U5284 ( .A1(n9050), .A2(n9068), .ZN(n4553) );
  NAND2_X1 U5285 ( .A1(n5545), .A2(n5437), .ZN(n4383) );
  OAI21_X1 U5286 ( .B1(n4345), .B2(n5534), .A(n5533), .ZN(n5538) );
  AOI21_X1 U5287 ( .B1(n4349), .B2(n4346), .A(n5530), .ZN(n4345) );
  OR2_X1 U5288 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  INV_X1 U5289 ( .A(n5558), .ZN(n4708) );
  MUX2_X1 U5290 ( .A(n8765), .B(n8764), .S(n8775), .Z(n8766) );
  NAND2_X1 U5291 ( .A1(n4378), .A2(n4376), .ZN(n4710) );
  NOR2_X1 U5292 ( .A1(n4267), .A2(n4377), .ZN(n4376) );
  NOR2_X1 U5293 ( .A1(n4274), .A2(n4380), .ZN(n4379) );
  INV_X1 U5294 ( .A(n4369), .ZN(n4368) );
  INV_X1 U5295 ( .A(n4371), .ZN(n4367) );
  INV_X1 U5296 ( .A(n5243), .ZN(n4795) );
  AOI211_X1 U5297 ( .C1(n4662), .C2(n9008), .A(n8599), .B(n8983), .ZN(n8648)
         );
  NAND2_X1 U5298 ( .A1(n4434), .A2(n5311), .ZN(n4433) );
  INV_X1 U5299 ( .A(n5326), .ZN(n4434) );
  NOR2_X1 U5300 ( .A1(n4433), .A2(n4429), .ZN(n4428) );
  INV_X1 U5301 ( .A(n5296), .ZN(n4429) );
  INV_X1 U5302 ( .A(n4423), .ZN(n4422) );
  OAI21_X1 U5303 ( .B1(n4425), .B2(n4424), .A(n5244), .ZN(n4423) );
  INV_X1 U5304 ( .A(n5224), .ZN(n4424) );
  INV_X1 U5305 ( .A(n4816), .ZN(n4402) );
  INV_X1 U5306 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4343) );
  NOR2_X1 U5307 ( .A1(n8322), .A2(n4477), .ZN(n4476) );
  INV_X1 U5308 ( .A(n4478), .ZN(n4477) );
  NOR2_X1 U5309 ( .A1(n8327), .A2(n8332), .ZN(n4478) );
  OR2_X1 U5310 ( .A1(n8345), .A2(n8033), .ZN(n5520) );
  AND2_X1 U5311 ( .A1(n7139), .A2(n4615), .ZN(n4611) );
  NOR2_X1 U5312 ( .A1(n7087), .A2(n7086), .ZN(n7092) );
  NAND2_X1 U5313 ( .A1(n5047), .A2(n4277), .ZN(n5484) );
  NOR2_X1 U5314 ( .A1(n7055), .A2(n7823), .ZN(n4472) );
  NAND2_X1 U5315 ( .A1(n5469), .A2(n5478), .ZN(n6775) );
  NOR2_X1 U5316 ( .A1(n8133), .A2(n8315), .ZN(n8125) );
  INV_X1 U5317 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5609) );
  INV_X1 U5318 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U5319 ( .A1(n4511), .A2(n4510), .ZN(n7660) );
  NAND2_X1 U5320 ( .A1(n8543), .A2(n4514), .ZN(n4510) );
  NAND2_X1 U5321 ( .A1(n4513), .A2(n7657), .ZN(n4512) );
  INV_X1 U5322 ( .A(n8522), .ZN(n4505) );
  NAND2_X1 U5323 ( .A1(n4327), .A2(n4326), .ZN(n8411) );
  INV_X1 U5324 ( .A(n8531), .ZN(n4326) );
  AOI21_X1 U5325 ( .B1(n7122), .B2(n7204), .A(n4278), .ZN(n4509) );
  OAI22_X1 U5326 ( .A1(n8788), .A2(n4543), .B1(n9012), .B2(n8775), .ZN(n8783)
         );
  OR2_X1 U5327 ( .A1(n9209), .A2(n8872), .ZN(n4543) );
  NOR4_X1 U5328 ( .A1(n8829), .A2(n8828), .A3(n8984), .A4(n8827), .ZN(n8831)
         );
  OR2_X1 U5329 ( .A1(n9214), .A2(n8986), .ZN(n8780) );
  NOR2_X1 U5330 ( .A1(n9075), .A2(n9093), .ZN(n4740) );
  INV_X1 U5331 ( .A(n4810), .ZN(n4742) );
  NOR2_X1 U5332 ( .A1(n7015), .A2(n7038), .ZN(n4457) );
  OAI21_X1 U5333 ( .B1(n6638), .B2(n4540), .A(n4537), .ZN(n8674) );
  INV_X1 U5334 ( .A(n4541), .ZN(n4540) );
  NAND2_X1 U5335 ( .A1(n6422), .A2(n6584), .ZN(n4720) );
  NAND2_X1 U5336 ( .A1(n9190), .A2(n4259), .ZN(n9157) );
  NAND2_X1 U5337 ( .A1(n9542), .A2(n9557), .ZN(n9523) );
  OAI21_X1 U5338 ( .B1(n5394), .B2(n5393), .A(n5392), .ZN(n5420) );
  AND2_X1 U5339 ( .A1(n4762), .A2(n5650), .ZN(n4761) );
  NOR2_X1 U5340 ( .A1(n4646), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4549) );
  INV_X1 U5341 ( .A(n4762), .ZN(n4646) );
  AND2_X1 U5342 ( .A1(n5363), .A2(n5351), .ZN(n5361) );
  AND2_X1 U5343 ( .A1(n5345), .A2(n5331), .ZN(n5343) );
  INV_X1 U5344 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5630) );
  INV_X1 U5345 ( .A(n5256), .ZN(n4716) );
  AOI21_X1 U5346 ( .B1(n5121), .B2(n4690), .A(n4688), .ZN(n4687) );
  INV_X1 U5347 ( .A(n5143), .ZN(n4688) );
  INV_X1 U5348 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U5349 ( .A1(n6838), .A2(n7820), .ZN(n6892) );
  CLKBUF_X1 U5350 ( .A(n6888), .Z(n7820) );
  AOI21_X1 U5351 ( .B1(n4580), .B2(n4578), .A(n4285), .ZN(n4577) );
  INV_X1 U5352 ( .A(n4580), .ZN(n4579) );
  AND2_X1 U5353 ( .A1(n7726), .A2(n7721), .ZN(n4589) );
  OR2_X1 U5354 ( .A1(n5196), .A2(n5195), .ZN(n5234) );
  AND2_X1 U5355 ( .A1(n7755), .A2(n7838), .ZN(n4584) );
  NOR2_X1 U5356 ( .A1(n6047), .A2(n9850), .ZN(n6045) );
  AND3_X1 U5357 ( .A1(n5380), .A2(n5379), .A3(n5378), .ZN(n7933) );
  AND3_X1 U5358 ( .A1(n5340), .A2(n5339), .A3(n5338), .ZN(n8043) );
  AND4_X1 U5359 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n7833)
         );
  AND4_X1 U5360 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n7819)
         );
  OR2_X1 U5361 ( .A1(n4923), .A2(n4875), .ZN(n4877) );
  NAND2_X1 U5362 ( .A1(n6538), .A2(n4444), .ZN(n6540) );
  OR2_X1 U5363 ( .A1(n6539), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U5364 ( .A1(n6540), .A2(n6541), .ZN(n6669) );
  NAND2_X1 U5365 ( .A1(n6669), .A2(n4443), .ZN(n6671) );
  OR2_X1 U5366 ( .A1(n6670), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5367 ( .A1(n6671), .A2(n6672), .ZN(n6947) );
  INV_X1 U5368 ( .A(n4448), .ZN(n8001) );
  NAND2_X1 U5369 ( .A1(n5389), .A2(n5388), .ZN(n8290) );
  AND2_X1 U5370 ( .A1(n8058), .A2(n5368), .ZN(n8077) );
  AOI21_X1 U5371 ( .B1(n4779), .B2(n4781), .A(n4778), .ZN(n4777) );
  INV_X1 U5372 ( .A(n4780), .ZN(n4779) );
  OR2_X1 U5373 ( .A1(n5300), .A2(n9403), .ZN(n5320) );
  NAND2_X1 U5374 ( .A1(n8119), .A2(n8118), .ZN(n8117) );
  AND3_X1 U5375 ( .A1(n5324), .A2(n5323), .A3(n5322), .ZN(n8144) );
  NAND2_X1 U5376 ( .A1(n8189), .A2(n4474), .ZN(n8133) );
  AND2_X1 U5377 ( .A1(n4475), .A2(n4476), .ZN(n4474) );
  NAND2_X1 U5378 ( .A1(n4628), .A2(n4262), .ZN(n4625) );
  NAND2_X1 U5379 ( .A1(n8189), .A2(n4476), .ZN(n8153) );
  OR2_X1 U5380 ( .A1(n8338), .A2(n7833), .ZN(n5511) );
  NAND2_X1 U5381 ( .A1(n8200), .A2(n5243), .ZN(n4799) );
  NAND2_X1 U5382 ( .A1(n4799), .A2(n4796), .ZN(n8173) );
  NAND2_X1 U5383 ( .A1(n8189), .A2(n8018), .ZN(n8190) );
  OR2_X1 U5384 ( .A1(n8345), .A2(n8236), .ZN(n4595) );
  NAND2_X1 U5385 ( .A1(n8215), .A2(n4820), .ZN(n4596) );
  AND2_X1 U5386 ( .A1(n5511), .A2(n5513), .ZN(n8205) );
  NOR2_X1 U5387 ( .A1(n8349), .A2(n8345), .ZN(n4488) );
  AND2_X1 U5388 ( .A1(n5520), .A2(n8201), .ZN(n8223) );
  AND3_X1 U5389 ( .A1(n4491), .A2(n4489), .A3(n8233), .ZN(n8230) );
  OR3_X1 U5390 ( .A1(n5132), .A2(n5131), .A3(n7922), .ZN(n5161) );
  NOR2_X1 U5391 ( .A1(n7232), .A2(n7295), .ZN(n7277) );
  AND2_X1 U5392 ( .A1(n6874), .A2(n4268), .ZN(n7102) );
  NAND2_X1 U5393 ( .A1(n7163), .A2(n7553), .ZN(n7096) );
  AOI21_X1 U5394 ( .B1(n4767), .B2(n5473), .A(n4317), .ZN(n4766) );
  INV_X1 U5395 ( .A(n5584), .ZN(n4767) );
  OAI211_X1 U5396 ( .C1(n5047), .C2(n4618), .A(n5484), .B(n4617), .ZN(n7086)
         );
  OR2_X1 U5397 ( .A1(n5046), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5398 ( .A1(n6874), .A2(n4470), .ZN(n6937) );
  NAND2_X1 U5399 ( .A1(n4769), .A2(n5584), .ZN(n6797) );
  NAND2_X1 U5400 ( .A1(n6785), .A2(n5585), .ZN(n4769) );
  INV_X1 U5401 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U5402 ( .A1(n6874), .A2(n9907), .ZN(n6876) );
  INV_X1 U5403 ( .A(n6775), .ZN(n6571) );
  NAND2_X1 U5404 ( .A1(n6562), .A2(n6561), .ZN(n6600) );
  NAND2_X1 U5405 ( .A1(n6334), .A2(n6333), .ZN(n6575) );
  INV_X1 U5406 ( .A(n6836), .ZN(n7055) );
  OR3_X1 U5407 ( .A1(n6760), .A2(n6759), .A3(n8013), .ZN(n9880) );
  OAI211_X1 U5408 ( .C1(n4334), .C2(n6175), .A(n4974), .B(n4973), .ZN(n6763)
         );
  NAND2_X1 U5409 ( .A1(n6633), .A2(n5427), .ZN(n4974) );
  OR2_X1 U5410 ( .A1(n6621), .A2(n4885), .ZN(n4950) );
  NAND2_X1 U5411 ( .A1(n6251), .A2(n9863), .ZN(n9850) );
  NAND2_X1 U5412 ( .A1(n5431), .A2(n4801), .ZN(n4582) );
  AND2_X1 U5413 ( .A1(n4837), .A2(n4265), .ZN(n4801) );
  NAND2_X1 U5414 ( .A1(n5610), .A2(n5609), .ZN(n5620) );
  INV_X1 U5415 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5606) );
  INV_X1 U5416 ( .A(n4250), .ZN(n8643) );
  CLKBUF_X1 U5417 ( .A(n8490), .Z(n8491) );
  XNOR2_X1 U5418 ( .A(n6686), .B(n6684), .ZN(n6503) );
  NAND2_X1 U5419 ( .A1(n8504), .A2(n4675), .ZN(n4674) );
  INV_X1 U5420 ( .A(n7610), .ZN(n4675) );
  OR2_X1 U5421 ( .A1(n6713), .A2(n6712), .ZN(n6916) );
  OR2_X1 U5422 ( .A1(n8435), .A2(n8555), .ZN(n4502) );
  AND2_X1 U5423 ( .A1(n7582), .A2(n7583), .ZN(n8531) );
  CLKBUF_X1 U5424 ( .A(n8411), .Z(n8534) );
  NOR2_X1 U5425 ( .A1(n4263), .A2(n4287), .ZN(n4703) );
  XNOR2_X1 U5426 ( .A(n5729), .B(n8448), .ZN(n5732) );
  AOI21_X1 U5427 ( .B1(n4250), .B2(n7625), .A(n5730), .ZN(n5731) );
  AND2_X1 U5428 ( .A1(n8642), .A2(n5722), .ZN(n5730) );
  OR2_X1 U5429 ( .A1(n7624), .A2(n7623), .ZN(n4507) );
  CLKBUF_X1 U5430 ( .A(n8492), .Z(n8584) );
  NAND2_X1 U5431 ( .A1(n5781), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4531) );
  AND2_X1 U5432 ( .A1(n8908), .A2(n8909), .ZN(n8906) );
  NOR2_X1 U5433 ( .A1(n5928), .A2(n5929), .ZN(n5927) );
  INV_X1 U5434 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5629) );
  AOI21_X1 U5435 ( .B1(n8916), .B2(n8915), .A(n8914), .ZN(n8917) );
  AOI21_X1 U5436 ( .B1(n8951), .B2(n8950), .A(n8949), .ZN(n8953) );
  NAND2_X1 U5437 ( .A1(n5695), .A2(n7080), .ZN(n5845) );
  NOR3_X1 U5438 ( .A1(n7523), .A2(n9209), .A3(n4458), .ZN(n8991) );
  XNOR2_X1 U5439 ( .A(n8985), .B(n8980), .ZN(n4442) );
  AOI21_X1 U5440 ( .B1(n4663), .B2(n4659), .A(n8983), .ZN(n4658) );
  INV_X1 U5441 ( .A(n9004), .ZN(n9007) );
  NAND2_X1 U5442 ( .A1(n4726), .A2(n4724), .ZN(n9002) );
  INV_X1 U5443 ( .A(n4725), .ZN(n4724) );
  OAI21_X1 U5444 ( .B1(n4732), .B2(n4738), .A(n4731), .ZN(n4725) );
  INV_X1 U5445 ( .A(n4734), .ZN(n4732) );
  INV_X1 U5446 ( .A(n4735), .ZN(n4730) );
  NAND2_X1 U5447 ( .A1(n7522), .A2(n8762), .ZN(n7523) );
  NAND2_X1 U5448 ( .A1(n4635), .A2(n4636), .ZN(n7513) );
  AOI21_X1 U5449 ( .B1(n4638), .B2(n4644), .A(n4637), .ZN(n4636) );
  INV_X1 U5450 ( .A(n8602), .ZN(n4637) );
  AND2_X1 U5451 ( .A1(n9028), .A2(n8489), .ZN(n7522) );
  NOR2_X1 U5452 ( .A1(n4733), .A2(n4737), .ZN(n4722) );
  AND2_X1 U5453 ( .A1(n9107), .A2(n4269), .ZN(n9036) );
  NAND2_X1 U5454 ( .A1(n9107), .A2(n4462), .ZN(n9059) );
  AOI21_X1 U5455 ( .B1(n4669), .B2(n8725), .A(n4668), .ZN(n4667) );
  NAND2_X1 U5456 ( .A1(n9107), .A2(n9090), .ZN(n9085) );
  OR2_X1 U5457 ( .A1(n7378), .A2(n7318), .ZN(n7388) );
  AND2_X1 U5458 ( .A1(n9190), .A2(n4270), .ZN(n9115) );
  NAND2_X1 U5459 ( .A1(n9190), .A2(n4256), .ZN(n9142) );
  AOI21_X1 U5460 ( .B1(n4649), .B2(n4653), .A(n4651), .ZN(n4648) );
  INV_X1 U5461 ( .A(n8650), .ZN(n4651) );
  NOR2_X1 U5462 ( .A1(n7483), .A2(n4650), .ZN(n4649) );
  NOR2_X1 U5463 ( .A1(n9524), .A2(n9286), .ZN(n9190) );
  NAND2_X1 U5464 ( .A1(n4654), .A2(n8711), .ZN(n9168) );
  NAND2_X1 U5465 ( .A1(n4654), .A2(n4652), .ZN(n9170) );
  INV_X1 U5466 ( .A(n4647), .ZN(n4652) );
  INV_X1 U5467 ( .A(n9518), .ZN(n9172) );
  INV_X1 U5468 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7178) );
  OR2_X1 U5469 ( .A1(n7179), .A2(n7178), .ZN(n7357) );
  NAND2_X1 U5470 ( .A1(n4756), .A2(n4754), .ZN(n9510) );
  AND2_X1 U5471 ( .A1(n9511), .A2(n4755), .ZN(n4754) );
  INV_X1 U5472 ( .A(n4759), .ZN(n4755) );
  INV_X1 U5473 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U5474 ( .A1(n4457), .A2(n4456), .ZN(n9541) );
  INV_X1 U5475 ( .A(n4457), .ZN(n7042) );
  NAND2_X1 U5476 ( .A1(n4743), .A2(n4744), .ZN(n6723) );
  NAND2_X1 U5477 ( .A1(n4745), .A2(n4273), .ZN(n4744) );
  NAND2_X1 U5478 ( .A1(n8810), .A2(n4746), .ZN(n4745) );
  AND2_X1 U5479 ( .A1(n6706), .A2(n8681), .ZN(n7011) );
  NAND2_X1 U5480 ( .A1(n4655), .A2(n4656), .ZN(n6706) );
  AND2_X1 U5481 ( .A1(n4657), .A2(n8657), .ZN(n4655) );
  INV_X1 U5482 ( .A(n8810), .ZN(n4657) );
  NAND2_X1 U5483 ( .A1(n4656), .A2(n8657), .ZN(n6641) );
  NOR2_X1 U5484 ( .A1(n9673), .A2(n8567), .ZN(n6813) );
  OR2_X1 U5485 ( .A1(n9672), .A2(n9676), .ZN(n9673) );
  NAND2_X1 U5486 ( .A1(n8837), .A2(n8835), .ZN(n8804) );
  NAND2_X1 U5487 ( .A1(n9695), .A2(n9750), .ZN(n9672) );
  NOR2_X1 U5488 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  INV_X1 U5489 ( .A(n5856), .ZN(n4534) );
  NAND2_X1 U5490 ( .A1(n8645), .A2(n6422), .ZN(n9706) );
  INV_X1 U5491 ( .A(n8887), .ZN(n6586) );
  OAI22_X1 U5492 ( .A1(n8664), .A2(n8663), .B1(n8662), .B2(n8661), .ZN(n9203)
         );
  NAND2_X1 U5493 ( .A1(n7466), .A2(n7465), .ZN(n9217) );
  AND2_X1 U5494 ( .A1(n5975), .A2(n7218), .ZN(n9778) );
  INV_X1 U5495 ( .A(n9778), .ZN(n9786) );
  OR2_X1 U5496 ( .A1(n5978), .A2(n5767), .ZN(n9784) );
  INV_X1 U5497 ( .A(n8642), .ZN(n9738) );
  NOR2_X1 U5498 ( .A1(n5972), .A2(n6399), .ZN(n7224) );
  NAND2_X1 U5499 ( .A1(n5798), .A2(n9466), .ZN(n5682) );
  INV_X1 U5500 ( .A(n5749), .ZN(n5874) );
  XNOR2_X1 U5501 ( .A(n5420), .B(n5419), .ZN(n5417) );
  CLKBUF_X1 U5502 ( .A(n5777), .Z(n8866) );
  NAND2_X1 U5503 ( .A1(n4430), .A2(n5311), .ZN(n5327) );
  NAND2_X1 U5504 ( .A1(n4437), .A2(n4435), .ZN(n4430) );
  NAND2_X1 U5505 ( .A1(n4437), .A2(n5298), .ZN(n5313) );
  NAND2_X1 U5506 ( .A1(n4421), .A2(n5224), .ZN(n5245) );
  NAND2_X1 U5507 ( .A1(n4715), .A2(n4425), .ZN(n4421) );
  NAND2_X1 U5508 ( .A1(n4715), .A2(n5208), .ZN(n5223) );
  AND2_X1 U5509 ( .A1(n6412), .A2(n6580), .ZN(n8926) );
  NAND2_X1 U5510 ( .A1(n4692), .A2(n5120), .ZN(n5145) );
  NAND2_X1 U5511 ( .A1(n4693), .A2(n5117), .ZN(n4692) );
  INV_X1 U5512 ( .A(n5122), .ZN(n4693) );
  AND2_X1 U5513 ( .A1(n6211), .A2(n6309), .ZN(n8933) );
  NAND2_X1 U5514 ( .A1(n4400), .A2(n4404), .ZN(n5041) );
  OR2_X1 U5515 ( .A1(n5005), .A2(n4407), .ZN(n4400) );
  OR2_X1 U5516 ( .A1(n5005), .A2(n5004), .ZN(n4408) );
  NAND2_X1 U5517 ( .A1(n4944), .A2(n4943), .ZN(n4948) );
  NAND2_X1 U5518 ( .A1(n6735), .A2(n6734), .ZN(n6743) );
  INV_X1 U5519 ( .A(n7766), .ZN(n4587) );
  NAND2_X1 U5520 ( .A1(n5353), .A2(n5352), .ZN(n8303) );
  AND4_X1 U5521 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n8180)
         );
  OR2_X1 U5522 ( .A1(n4882), .A2(n5866), .ZN(n4350) );
  OR2_X1 U5523 ( .A1(n6497), .A2(n4885), .ZN(n4351) );
  NAND2_X1 U5524 ( .A1(n7847), .A2(n7721), .ZN(n7859) );
  AND4_X1 U5525 ( .A1(n4984), .A2(n4983), .A3(n4982), .A4(n4981), .ZN(n6896)
         );
  AND4_X1 U5526 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n7258)
         );
  NAND2_X1 U5527 ( .A1(n7559), .A2(n7252), .ZN(n7254) );
  AND4_X1 U5528 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n7890)
         );
  NAND2_X1 U5529 ( .A1(n4572), .A2(n4570), .ZN(n7248) );
  OR2_X1 U5530 ( .A1(n4882), .A2(n5857), .ZN(n4871) );
  OR2_X1 U5531 ( .A1(n7924), .A2(n8179), .ZN(n7904) );
  OR2_X1 U5532 ( .A1(n7924), .A2(n8181), .ZN(n7903) );
  NAND2_X1 U5533 ( .A1(n6523), .A2(n6522), .ZN(n6553) );
  NAND2_X1 U5534 ( .A1(n6254), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7886) );
  INV_X1 U5535 ( .A(n5600), .ZN(n5601) );
  INV_X1 U5536 ( .A(n7890), .ZN(n8195) );
  INV_X1 U5537 ( .A(n7819), .ZN(n7941) );
  CLKBUF_X1 U5538 ( .A(n6055), .Z(n7947) );
  INV_X2 U5539 ( .A(P2_U3966), .ZN(n7948) );
  OR2_X1 U5540 ( .A1(n5357), .A2(n4791), .ZN(n4788) );
  INV_X1 U5541 ( .A(n4790), .ZN(n4789) );
  NOR2_X1 U5542 ( .A1(n6157), .A2(n6156), .ZN(n6155) );
  INV_X1 U5543 ( .A(n4446), .ZN(n6144) );
  NAND2_X1 U5544 ( .A1(n6086), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4445) );
  INV_X1 U5545 ( .A(n4451), .ZN(n6121) );
  AND2_X1 U5546 ( .A1(n4451), .A2(n4450), .ZN(n6168) );
  NAND2_X1 U5547 ( .A1(n6088), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4450) );
  NOR2_X1 U5548 ( .A1(n6315), .A2(n4322), .ZN(n6317) );
  NAND2_X1 U5549 ( .A1(n6317), .A2(n6318), .ZN(n6457) );
  NOR2_X1 U5550 ( .A1(n7970), .A2(n4449), .ZN(n7973) );
  AND2_X1 U5551 ( .A1(n7976), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4449) );
  NOR2_X1 U5552 ( .A1(n7973), .A2(n7972), .ZN(n7985) );
  AND2_X1 U5553 ( .A1(n6097), .A2(n6094), .ZN(n9814) );
  NAND2_X1 U5554 ( .A1(n4481), .A2(n8288), .ZN(n4480) );
  NAND2_X1 U5555 ( .A1(n8086), .A2(n4286), .ZN(n4482) );
  OR2_X1 U5556 ( .A1(n8086), .A2(n4484), .ZN(n4483) );
  AOI21_X1 U5557 ( .B1(n4272), .B2(n4605), .A(n4603), .ZN(n4602) );
  OAI21_X1 U5558 ( .B1(n8084), .B2(n4605), .A(n4272), .ZN(n8071) );
  NAND2_X1 U5559 ( .A1(n8083), .A2(n8045), .ZN(n8073) );
  INV_X1 U5560 ( .A(n8303), .ZN(n8091) );
  NAND2_X1 U5561 ( .A1(n8138), .A2(n5536), .ZN(n8122) );
  NAND2_X1 U5562 ( .A1(n4629), .A2(n4630), .ZN(n8150) );
  OAI21_X1 U5563 ( .B1(n8188), .B2(n8035), .A(n4811), .ZN(n8168) );
  NAND2_X1 U5564 ( .A1(n4770), .A2(n4773), .ZN(n4822) );
  AND2_X1 U5565 ( .A1(n4623), .A2(n4264), .ZN(n8247) );
  NAND2_X1 U5566 ( .A1(n5169), .A2(n5501), .ZN(n8241) );
  NAND2_X1 U5567 ( .A1(n8027), .A2(n4624), .ZN(n8273) );
  AND2_X1 U5568 ( .A1(n7147), .A2(n5490), .ZN(n7229) );
  NAND2_X1 U5569 ( .A1(n5094), .A2(n5093), .ZN(n8373) );
  NAND2_X1 U5570 ( .A1(n4616), .A2(n4613), .ZN(n7228) );
  NAND2_X1 U5571 ( .A1(n4616), .A2(n4615), .ZN(n7142) );
  NAND2_X1 U5572 ( .A1(n6873), .A2(n6784), .ZN(n4600) );
  OR2_X1 U5573 ( .A1(n6575), .A2(n7798), .ZN(n8062) );
  OR2_X1 U5574 ( .A1(n4885), .A2(n5858), .ZN(n4902) );
  INV_X1 U5575 ( .A(n8262), .ZN(n8284) );
  NAND2_X1 U5576 ( .A1(n6332), .A2(n6042), .ZN(n8250) );
  AND2_X1 U5577 ( .A1(n8253), .A2(n9835), .ZN(n8255) );
  INV_X1 U5578 ( .A(n8062), .ZN(n8277) );
  NAND2_X1 U5580 ( .A1(n8253), .A2(n9845), .ZN(n8262) );
  AND2_X1 U5581 ( .A1(n6250), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9863) );
  INV_X1 U5582 ( .A(n9857), .ZN(n9860) );
  XNOR2_X1 U5583 ( .A(n5619), .B(n4802), .ZN(n7305) );
  INV_X1 U5584 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7169) );
  XNOR2_X1 U5585 ( .A(n5622), .B(n5621), .ZN(n7170) );
  INV_X1 U5586 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U5587 ( .A1(n5620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5622) );
  INV_X1 U5588 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7051) );
  INV_X1 U5589 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6929) );
  INV_X1 U5590 ( .A(n5403), .ZN(n5404) );
  CLKBUF_X1 U5591 ( .A(n5402), .Z(n5403) );
  INV_X1 U5592 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6772) );
  INV_X1 U5593 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U5594 ( .A1(n4333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U5595 ( .A1(n4835), .A2(n4276), .ZN(n4333) );
  NOR2_X1 U5596 ( .A1(n4619), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8398) );
  INV_X1 U5597 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6331) );
  INV_X1 U5598 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6214) );
  INV_X1 U5599 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6203) );
  INV_X1 U5600 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5981) );
  INV_X1 U5601 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5936) );
  INV_X1 U5602 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5878) );
  INV_X1 U5603 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5869) );
  INV_X1 U5604 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5866) );
  INV_X1 U5605 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U5606 ( .A1(n7427), .A2(n7426), .ZN(n9237) );
  NAND2_X1 U5607 ( .A1(n4704), .A2(n7067), .ZN(n7109) );
  AND2_X1 U5608 ( .A1(n7696), .A2(n7695), .ZN(n8465) );
  AND2_X1 U5609 ( .A1(n4702), .A2(n4701), .ZN(n8471) );
  NAND2_X1 U5610 ( .A1(n7406), .A2(n7405), .ZN(n9248) );
  INV_X1 U5611 ( .A(n8878), .ZN(n9189) );
  NAND2_X1 U5612 ( .A1(n7375), .A2(n7374), .ZN(n9276) );
  INV_X1 U5613 ( .A(n9234), .ZN(n8520) );
  AND2_X1 U5614 ( .A1(n4676), .A2(n4283), .ZN(n6278) );
  NAND2_X1 U5615 ( .A1(n6907), .A2(n6906), .ZN(n7069) );
  NAND2_X1 U5616 ( .A1(n4496), .A2(n4497), .ZN(n8524) );
  AOI21_X1 U5617 ( .B1(n7624), .B2(n4499), .A(n4498), .ZN(n4497) );
  AND2_X1 U5618 ( .A1(n4503), .A2(n4506), .ZN(n4499) );
  OR2_X1 U5619 ( .A1(n4700), .A2(n4514), .ZN(n8542) );
  OR2_X1 U5620 ( .A1(n7121), .A2(n7122), .ZN(n7205) );
  INV_X1 U5621 ( .A(n9094), .ZN(n9123) );
  INV_X1 U5622 ( .A(n8591), .ZN(n9575) );
  AND2_X1 U5623 ( .A1(n5787), .A2(n6010), .ZN(n8587) );
  AND2_X1 U5624 ( .A1(n8576), .A2(n8573), .ZN(n7686) );
  AND2_X1 U5625 ( .A1(n7469), .A2(n7452), .ZN(n8580) );
  INV_X1 U5626 ( .A(n9576), .ZN(n8596) );
  NAND2_X1 U5627 ( .A1(n5787), .A2(n8866), .ZN(n8590) );
  NAND2_X1 U5628 ( .A1(n5772), .A2(n6074), .ZN(n8594) );
  INV_X1 U5629 ( .A(n4565), .ZN(n4564) );
  OAI21_X1 U5630 ( .B1(n8864), .B2(n8863), .A(n8865), .ZN(n4565) );
  NAND2_X1 U5631 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5689) );
  AOI21_X1 U5632 ( .B1(n4261), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_21__SCAN_IN), .ZN(n4519) );
  AND3_X1 U5633 ( .A1(n5898), .A2(n5897), .A3(n5896), .ZN(n8966) );
  AND3_X1 U5634 ( .A1(n5894), .A2(n5893), .A3(n5892), .ZN(n8988) );
  OR2_X1 U5635 ( .A1(n7478), .A2(n4249), .ZN(n7476) );
  NAND2_X1 U5636 ( .A1(n5778), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5703) );
  OR2_X2 U5637 ( .A1(n5845), .A2(n4246), .ZN(n8888) );
  NAND2_X1 U5638 ( .A1(n5778), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5660) );
  AOI21_X1 U5639 ( .B1(n5942), .B2(n5939), .A(n9619), .ZN(n5941) );
  AOI21_X1 U5640 ( .B1(n9560), .B2(n6230), .A(n6229), .ZN(n6232) );
  AND2_X1 U5641 ( .A1(n5818), .A2(n5840), .ZN(n9661) );
  INV_X1 U5642 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4860) );
  NAND2_X1 U5643 ( .A1(n8668), .A2(n8667), .ZN(n9199) );
  NAND2_X1 U5644 ( .A1(n4665), .A2(n8598), .ZN(n7491) );
  INV_X1 U5645 ( .A(n9222), .ZN(n8762) );
  INV_X1 U5646 ( .A(n9227), .ZN(n8489) );
  NAND2_X1 U5647 ( .A1(n4641), .A2(n4640), .ZN(n9023) );
  NAND2_X1 U5648 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5649 ( .A1(n9073), .A2(n8750), .ZN(n9041) );
  NAND2_X1 U5650 ( .A1(n9069), .A2(n9068), .ZN(n9067) );
  NAND2_X1 U5651 ( .A1(n9082), .A2(n4810), .ZN(n9069) );
  NAND2_X1 U5652 ( .A1(n4671), .A2(n8619), .ZN(n9102) );
  AND2_X1 U5653 ( .A1(n9126), .A2(n4753), .ZN(n4749) );
  AND2_X1 U5654 ( .A1(n4750), .A2(n4753), .ZN(n9127) );
  NAND2_X1 U5655 ( .A1(n9151), .A2(n4808), .ZN(n9133) );
  INV_X1 U5656 ( .A(n4750), .ZN(n9132) );
  INV_X1 U5657 ( .A(n9279), .ZN(n9178) );
  NAND2_X1 U5658 ( .A1(n7350), .A2(n7349), .ZN(n9522) );
  NAND2_X1 U5659 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  NAND2_X1 U5660 ( .A1(n7116), .A2(n7115), .ZN(n9540) );
  INV_X1 U5661 ( .A(n9776), .ZN(n7010) );
  NAND2_X1 U5662 ( .A1(n9719), .A2(n9675), .ZN(n9717) );
  INV_X1 U5663 ( .A(n9118), .ZN(n9714) );
  NAND2_X1 U5664 ( .A1(n6812), .A2(n6622), .ZN(n6722) );
  NAND2_X1 U5665 ( .A1(n6639), .A2(n8837), .ZN(n9680) );
  OAI21_X1 U5666 ( .B1(n5864), .B2(n4619), .A(n4455), .ZN(n4453) );
  NAND2_X1 U5667 ( .A1(n4619), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4455) );
  OR2_X1 U5668 ( .A1(n5971), .A2(n5790), .ZN(n9118) );
  NAND2_X1 U5669 ( .A1(n6655), .A2(n9118), .ZN(n9719) );
  INV_X1 U5670 ( .A(n5973), .ZN(n9574) );
  INV_X1 U5671 ( .A(n9717), .ZN(n9539) );
  AND2_X1 U5672 ( .A1(n9144), .A2(n9778), .ZN(n9698) );
  INV_X2 U5673 ( .A(n9719), .ZN(n9715) );
  AND2_X2 U5674 ( .A1(n7224), .A2(n7223), .ZN(n9811) );
  NOR2_X1 U5675 ( .A1(n9207), .A2(n4438), .ZN(n9210) );
  NAND2_X1 U5676 ( .A1(n4440), .A2(n4439), .ZN(n4438) );
  AOI211_X1 U5677 ( .C1(n9777), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9215)
         );
  AND2_X2 U5678 ( .A1(n7224), .A2(n6400), .ZN(n9794) );
  AND2_X1 U5679 ( .A1(n5768), .A2(n5763), .ZN(n5969) );
  INV_X1 U5680 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U5681 ( .A1(n4414), .A2(n4412), .ZN(n9460) );
  NAND2_X1 U5682 ( .A1(n4415), .A2(n4413), .ZN(n4412) );
  INV_X1 U5683 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U5684 ( .A1(n4714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5647) );
  XNOR2_X1 U5685 ( .A(n5297), .B(n5296), .ZN(n7425) );
  INV_X1 U5686 ( .A(n5764), .ZN(n8798) );
  INV_X1 U5687 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6932) );
  INV_X1 U5688 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6774) );
  INV_X1 U5689 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6663) );
  INV_X1 U5690 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6413) );
  INV_X1 U5691 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6212) );
  INV_X1 U5692 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6194) );
  INV_X1 U5693 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5989) );
  INV_X1 U5694 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5919) );
  INV_X1 U5695 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5868) );
  NOR2_X1 U5696 ( .A1(n5724), .A2(n4747), .ZN(n5807) );
  NAND2_X1 U5697 ( .A1(n5628), .A2(n4748), .ZN(n4747) );
  INV_X1 U5698 ( .A(n4933), .ZN(n4466) );
  NOR2_X2 U5699 ( .A1(n5726), .A2(n5725), .ZN(n6013) );
  INV_X1 U5700 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4344) );
  AND2_X1 U5701 ( .A1(n7812), .A2(n7814), .ZN(n4335) );
  INV_X1 U5702 ( .A(n7917), .ZN(n4330) );
  NAND2_X1 U5703 ( .A1(n4332), .A2(n7919), .ZN(n4331) );
  NAND2_X1 U5704 ( .A1(n4338), .A2(n4336), .ZN(P1_U3260) );
  AOI21_X1 U5705 ( .B1(n8959), .B2(n9125), .A(n4337), .ZN(n4336) );
  NAND2_X1 U5706 ( .A1(n8960), .A2(n9679), .ZN(n4338) );
  OAI21_X1 U5707 ( .B1(n4860), .B2(n9605), .A(n8961), .ZN(n4337) );
  INV_X1 U5708 ( .A(n8355), .ZN(n4489) );
  AND2_X1 U5709 ( .A1(n4259), .A2(n9148), .ZN(n4256) );
  AND3_X1 U5710 ( .A1(n4837), .A2(n4265), .A3(n4313), .ZN(n4257) );
  INV_X2 U5711 ( .A(n4249), .ZN(n6918) );
  INV_X1 U5712 ( .A(n8233), .ZN(n8349) );
  AND2_X1 U5713 ( .A1(n5506), .A2(n5501), .ZN(n4258) );
  AND2_X1 U5714 ( .A1(n9178), .A2(n9162), .ZN(n4259) );
  OR2_X1 U5715 ( .A1(n7462), .A2(n7518), .ZN(n4260) );
  XNOR2_X1 U5716 ( .A(n5689), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5764) );
  OR2_X1 U5717 ( .A1(n5667), .A2(n4521), .ZN(n4261) );
  NAND2_X1 U5718 ( .A1(n8322), .A2(n8036), .ZN(n4262) );
  AND2_X1 U5719 ( .A1(n7108), .A2(n4705), .ZN(n4263) );
  AOI21_X1 U5720 ( .B1(n7754), .B2(n7864), .A(n4303), .ZN(n7841) );
  INV_X1 U5721 ( .A(n5473), .ZN(n4768) );
  AND2_X1 U5722 ( .A1(n4672), .A2(n4674), .ZN(n8503) );
  NAND2_X1 U5723 ( .A1(n8360), .A2(n8243), .ZN(n4264) );
  AND2_X1 U5724 ( .A1(n4838), .A2(n4802), .ZN(n4265) );
  NAND2_X1 U5725 ( .A1(n5725), .A2(n5628), .ZN(n5810) );
  AND2_X1 U5726 ( .A1(n9887), .A2(n9893), .ZN(n4266) );
  NOR2_X1 U5727 ( .A1(n4381), .A2(n5557), .ZN(n4267) );
  AND2_X1 U5728 ( .A1(n8636), .A2(n8635), .ZN(n8997) );
  INV_X1 U5729 ( .A(n8997), .ZN(n9209) );
  INV_X1 U5730 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5646) );
  AND2_X1 U5731 ( .A1(n4470), .A2(n4469), .ZN(n4268) );
  AND2_X1 U5732 ( .A1(n4462), .A2(n4461), .ZN(n4269) );
  AND2_X1 U5733 ( .A1(n4256), .A2(n4460), .ZN(n4270) );
  NOR2_X1 U5734 ( .A1(n9004), .A2(n8982), .ZN(n4663) );
  NOR2_X1 U5735 ( .A1(n8276), .A2(n8360), .ZN(n4491) );
  NAND2_X1 U5736 ( .A1(n9107), .A2(n4464), .ZN(n4465) );
  INV_X1 U5737 ( .A(n5722), .ZN(n5711) );
  INV_X1 U5738 ( .A(n8835), .ZN(n4539) );
  NAND2_X1 U5739 ( .A1(n6874), .A2(n4472), .ZN(n4473) );
  AND2_X1 U5740 ( .A1(n5381), .A2(n5361), .ZN(n4271) );
  INV_X1 U5741 ( .A(n8093), .ZN(n4713) );
  NAND2_X2 U5742 ( .A1(n4848), .A2(n4845), .ZN(n5357) );
  AND4_X1 U5743 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n7553)
         );
  INV_X1 U5744 ( .A(n7553), .ZN(n4618) );
  AND2_X1 U5745 ( .A1(n8072), .A2(n4604), .ZN(n4272) );
  INV_X1 U5746 ( .A(n7657), .ZN(n4514) );
  AND2_X1 U5747 ( .A1(n4507), .A2(n4506), .ZN(n8435) );
  OR2_X1 U5748 ( .A1(n8884), .A2(n6721), .ZN(n4273) );
  NAND2_X1 U5749 ( .A1(n4713), .A2(n4712), .ZN(n4274) );
  INV_X2 U5750 ( .A(n6283), .ZN(n8455) );
  INV_X2 U5751 ( .A(n5015), .ZN(n4953) );
  OR2_X1 U5752 ( .A1(n9561), .A2(n8700), .ZN(n4275) );
  INV_X1 U5753 ( .A(n4774), .ZN(n4773) );
  NAND2_X1 U5754 ( .A1(n4502), .A2(n8436), .ZN(n8434) );
  INV_X1 U5755 ( .A(n4714), .ZN(n5645) );
  AND2_X1 U5756 ( .A1(n4834), .A2(n4785), .ZN(n4276) );
  NAND2_X1 U5757 ( .A1(n5579), .A2(n5578), .ZN(n6344) );
  INV_X1 U5758 ( .A(n8598), .ZN(n4662) );
  AND2_X1 U5759 ( .A1(n5046), .A2(n4618), .ZN(n4277) );
  AND2_X1 U5760 ( .A1(n7565), .A2(n7563), .ZN(n4278) );
  INV_X1 U5761 ( .A(n8724), .ZN(n4668) );
  OR3_X1 U5762 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4279) );
  OR2_X1 U5763 ( .A1(n4650), .A2(n8775), .ZN(n4280) );
  OR2_X1 U5764 ( .A1(n9286), .A2(n9172), .ZN(n8711) );
  INV_X1 U5765 ( .A(n8711), .ZN(n4650) );
  AND2_X1 U5766 ( .A1(n4446), .A2(n4445), .ZN(n4281) );
  AND2_X1 U5767 ( .A1(n4664), .A2(n4663), .ZN(n4282) );
  NAND2_X1 U5768 ( .A1(n6266), .A2(n6265), .ZN(n4283) );
  AND2_X1 U5769 ( .A1(n4911), .A2(n4933), .ZN(n4284) );
  NAND2_X1 U5770 ( .A1(n5248), .A2(n5247), .ZN(n8332) );
  AND2_X1 U5771 ( .A1(n7743), .A2(n7742), .ZN(n4285) );
  NAND2_X1 U5772 ( .A1(n5366), .A2(n5365), .ZN(n8298) );
  AND2_X1 U5773 ( .A1(n4484), .A2(n4485), .ZN(n4286) );
  AND2_X1 U5774 ( .A1(n7112), .A2(n7111), .ZN(n4287) );
  INV_X1 U5775 ( .A(n4375), .ZN(n4374) );
  NAND2_X1 U5776 ( .A1(n5282), .A2(n5281), .ZN(n8322) );
  CLKBUF_X3 U5777 ( .A(n4861), .Z(n4619) );
  INV_X1 U5778 ( .A(n9893), .ZN(n9836) );
  AND3_X1 U5779 ( .A1(n4351), .A2(n4350), .A3(n4311), .ZN(n9893) );
  OR2_X1 U5780 ( .A1(n5552), .A2(n5553), .ZN(n4288) );
  AND2_X1 U5781 ( .A1(n4799), .A2(n5511), .ZN(n4289) );
  INV_X1 U5782 ( .A(n4664), .ZN(n9006) );
  AND2_X1 U5783 ( .A1(n8086), .A2(n4485), .ZN(n4290) );
  AND2_X1 U5784 ( .A1(n5508), .A2(n5510), .ZN(n4291) );
  NAND2_X1 U5785 ( .A1(n7520), .A2(n7459), .ZN(n4292) );
  INV_X1 U5786 ( .A(n4644), .ZN(n4642) );
  NAND2_X1 U5787 ( .A1(n8750), .A2(n8601), .ZN(n4644) );
  INV_X1 U5788 ( .A(n9253), .ZN(n9090) );
  NAND2_X1 U5789 ( .A1(n7396), .A2(n7395), .ZN(n9253) );
  AND2_X1 U5790 ( .A1(n5216), .A2(n5215), .ZN(n8221) );
  INV_X1 U5791 ( .A(n8221), .ZN(n8345) );
  AND2_X1 U5792 ( .A1(n4674), .A2(n7619), .ZN(n4293) );
  AND2_X1 U5793 ( .A1(n7655), .A2(n7654), .ZN(n4294) );
  INV_X1 U5794 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5669) );
  INV_X1 U5795 ( .A(n9064), .ZN(n9244) );
  AND2_X1 U5796 ( .A1(n7417), .A2(n7416), .ZN(n9064) );
  NAND2_X1 U5797 ( .A1(n5705), .A2(n4517), .ZN(n5724) );
  NAND3_X1 U5798 ( .A1(n4391), .A2(n7141), .A3(n4390), .ZN(n4295) );
  AND2_X1 U5799 ( .A1(n4629), .A2(n4627), .ZN(n4296) );
  OR2_X1 U5800 ( .A1(n5602), .A2(n5601), .ZN(n4297) );
  INV_X1 U5801 ( .A(n4459), .ZN(n9014) );
  NOR2_X1 U5802 ( .A1(n7523), .A2(n9217), .ZN(n4459) );
  AND2_X1 U5803 ( .A1(n4671), .A2(n4669), .ZN(n4298) );
  OR2_X1 U5804 ( .A1(n5916), .A2(n5667), .ZN(n4299) );
  AND2_X1 U5805 ( .A1(n4708), .A2(n5535), .ZN(n4300) );
  AND2_X1 U5806 ( .A1(n4393), .A2(n4392), .ZN(n4301) );
  NAND2_X1 U5807 ( .A1(n4700), .A2(n4514), .ZN(n4302) );
  AND2_X1 U5808 ( .A1(n5529), .A2(n8141), .ZN(n8151) );
  INV_X1 U5809 ( .A(n4797), .ZN(n4796) );
  NAND2_X1 U5810 ( .A1(n4798), .A2(n5511), .ZN(n4797) );
  AND2_X1 U5811 ( .A1(n7866), .A2(n7868), .ZN(n4303) );
  AND2_X1 U5812 ( .A1(n4935), .A2(SI_4_), .ZN(n4304) );
  NAND2_X1 U5813 ( .A1(n8976), .A2(n8975), .ZN(n4305) );
  NOR2_X1 U5814 ( .A1(n7264), .A2(n7552), .ZN(n4614) );
  MUX2_X1 U5815 ( .A(n5571), .B(n5570), .S(n5569), .Z(n5572) );
  NAND2_X1 U5816 ( .A1(n4645), .A2(n8628), .ZN(n4306) );
  INV_X1 U5817 ( .A(n6055), .ZN(n6345) );
  INV_X1 U5818 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5819 ( .A1(n4630), .A2(n8159), .ZN(n4628) );
  INV_X1 U5820 ( .A(n5306), .ZN(n4475) );
  AND2_X1 U5821 ( .A1(n4913), .A2(SI_3_), .ZN(n4307) );
  INV_X1 U5822 ( .A(n5557), .ZN(n4711) );
  AND2_X1 U5823 ( .A1(n4633), .A2(n4262), .ZN(n4308) );
  AND2_X1 U5824 ( .A1(n7268), .A2(n5497), .ZN(n4309) );
  NOR2_X1 U5825 ( .A1(n8841), .A2(n4542), .ZN(n4310) );
  OR2_X1 U5826 ( .A1(n4334), .A2(n6141), .ZN(n4311) );
  AND2_X1 U5827 ( .A1(n4273), .A2(n6622), .ZN(n4312) );
  NOR2_X1 U5828 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4313) );
  AND2_X1 U5829 ( .A1(n4761), .A2(n4760), .ZN(n4314) );
  OR2_X1 U5830 ( .A1(n4660), .A2(n8600), .ZN(n4315) );
  INV_X1 U5831 ( .A(n4608), .ZN(n4607) );
  OAI21_X1 U5832 ( .B1(n4609), .B2(n4947), .A(n4972), .ZN(n4608) );
  INV_X1 U5833 ( .A(n5778), .ZN(n5891) );
  INV_X1 U5834 ( .A(n9237), .ZN(n4461) );
  INV_X1 U5835 ( .A(n8194), .ZN(n4798) );
  INV_X1 U5836 ( .A(n5782), .ZN(n6283) );
  NAND2_X1 U5837 ( .A1(n4835), .A2(n4834), .ZN(n5175) );
  NAND2_X1 U5838 ( .A1(n7333), .A2(n7332), .ZN(n9266) );
  INV_X1 U5839 ( .A(n9266), .ZN(n4460) );
  INV_X1 U5840 ( .A(n5585), .ZN(n4765) );
  AND2_X1 U5841 ( .A1(n6100), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U5842 ( .A1(n7205), .A2(n7204), .ZN(n7564) );
  NAND2_X1 U5843 ( .A1(n7342), .A2(n7341), .ZN(n9271) );
  INV_X1 U5844 ( .A(n9271), .ZN(n9148) );
  AND2_X1 U5845 ( .A1(n6824), .A2(n6997), .ZN(n4317) );
  NOR2_X1 U5846 ( .A1(n8216), .A2(n8338), .ZN(n8189) );
  AND2_X1 U5847 ( .A1(n8711), .A2(n8710), .ZN(n4318) );
  NAND2_X1 U5848 ( .A1(n9190), .A2(n9178), .ZN(n4319) );
  NAND2_X1 U5849 ( .A1(n8493), .A2(n7610), .ZN(n8502) );
  INV_X1 U5850 ( .A(n4690), .ZN(n4689) );
  NOR2_X1 U5851 ( .A1(n5144), .A2(n4691), .ZN(n4690) );
  OR2_X1 U5852 ( .A1(n8315), .A2(n8144), .ZN(n5539) );
  INV_X1 U5853 ( .A(n5539), .ZN(n4778) );
  NAND2_X1 U5854 ( .A1(n8189), .A2(n4478), .ZN(n4479) );
  INV_X1 U5855 ( .A(n4490), .ZN(n8258) );
  NAND2_X1 U5856 ( .A1(n4491), .A2(n4489), .ZN(n4490) );
  NOR2_X1 U5857 ( .A1(n9072), .A2(n7414), .ZN(n4320) );
  INV_X1 U5858 ( .A(n4737), .ZN(n4736) );
  NOR2_X1 U5859 ( .A1(n8520), .A2(n8603), .ZN(n4737) );
  NOR2_X1 U5860 ( .A1(n7911), .A2(n4584), .ZN(n4321) );
  INV_X1 U5861 ( .A(n4738), .ZN(n4733) );
  NAND2_X1 U5862 ( .A1(n9237), .A2(n9055), .ZN(n4738) );
  AND2_X1 U5863 ( .A1(n6045), .A2(n6041), .ZN(n7919) );
  XNOR2_X1 U5864 ( .A(n5687), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U5865 ( .A1(n6892), .A2(n6843), .ZN(n6999) );
  NAND2_X1 U5866 ( .A1(n5614), .A2(n4838), .ZN(n5617) );
  INV_X1 U5867 ( .A(n4251), .ZN(n5015) );
  INV_X1 U5868 ( .A(n8836), .ZN(n4538) );
  AND2_X1 U5869 ( .A1(n5431), .A2(n4837), .ZN(n5614) );
  AND2_X1 U5870 ( .A1(n6316), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4322) );
  INV_X1 U5871 ( .A(n5363), .ZN(n4411) );
  AND2_X1 U5872 ( .A1(n5194), .A2(n5193), .ZN(n8233) );
  AND2_X1 U5873 ( .A1(n5381), .A2(n4411), .ZN(n4323) );
  NAND2_X1 U5874 ( .A1(n4551), .A2(n5638), .ZN(n4550) );
  INV_X1 U5875 ( .A(n7186), .ZN(n4456) );
  INV_X1 U5876 ( .A(n7163), .ZN(n4469) );
  OR2_X1 U5877 ( .A1(n5764), .A2(n9125), .ZN(n8785) );
  INV_X1 U5878 ( .A(n8785), .ZN(n8775) );
  INV_X1 U5879 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4802) );
  AND2_X1 U5880 ( .A1(n7986), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4324) );
  NAND2_X1 U5881 ( .A1(n5692), .A2(n5691), .ZN(n9125) );
  INV_X1 U5882 ( .A(n9125), .ZN(n9679) );
  INV_X1 U5883 ( .A(n6759), .ZN(n6771) );
  INV_X1 U5884 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n4791) );
  INV_X1 U5885 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4792) );
  AND2_X2 U5886 ( .A1(n7624), .A2(n7623), .ZN(n8555) );
  NAND2_X1 U5887 ( .A1(n6493), .A2(n6492), .ZN(n6686) );
  NAND2_X1 U5888 ( .A1(n7662), .A2(n7661), .ZN(n8425) );
  NAND2_X1 U5889 ( .A1(n8563), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U5890 ( .A1(n6859), .A2(n6858), .ZN(n4494) );
  NAND2_X1 U5891 ( .A1(n8511), .A2(n7673), .ZN(n8479) );
  NAND2_X1 U5892 ( .A1(n4325), .A2(n4703), .ZN(n7121) );
  NAND3_X1 U5893 ( .A1(n6907), .A2(n4706), .A3(n6906), .ZN(n4325) );
  NAND2_X1 U5894 ( .A1(n6003), .A2(n5698), .ZN(n6006) );
  NAND2_X1 U5895 ( .A1(n8562), .A2(n8564), .ZN(n8563) );
  INV_X1 U5896 ( .A(n8530), .ZN(n4327) );
  NAND2_X2 U5897 ( .A1(n7218), .A2(n5762), .ZN(n5693) );
  XNOR2_X2 U5898 ( .A(n5670), .B(n5669), .ZN(n7218) );
  INV_X1 U5899 ( .A(n5698), .ZN(n6004) );
  AND2_X2 U5900 ( .A1(n4342), .A2(n4340), .ZN(n4861) );
  NAND2_X1 U5901 ( .A1(n4948), .A2(n4607), .ZN(n4399) );
  NAND2_X1 U5902 ( .A1(n4665), .A2(n4661), .ZN(n4664) );
  NAND2_X1 U5903 ( .A1(n4339), .A2(n4284), .ZN(n4679) );
  OAI21_X2 U5904 ( .B1(n7791), .B2(n7786), .A(n7790), .ZN(n7877) );
  XNOR2_X1 U5905 ( .A(n6836), .B(n7749), .ZN(n6839) );
  NAND2_X1 U5906 ( .A1(n4408), .A2(n5006), .ZN(n5022) );
  NAND2_X1 U5907 ( .A1(n4573), .A2(n4576), .ZN(n4571) );
  NOR2_X1 U5908 ( .A1(n7776), .A2(n4329), .ZN(n7754) );
  NAND2_X1 U5909 ( .A1(n8235), .A2(n5516), .ZN(n8222) );
  NAND2_X2 U5910 ( .A1(n8158), .A2(n5295), .ZN(n8139) );
  NAND2_X2 U5911 ( .A1(n5104), .A2(n7141), .ZN(n7147) );
  NAND2_X1 U5912 ( .A1(n6723), .A2(n8812), .ZN(n7009) );
  NAND2_X1 U5913 ( .A1(n4750), .A2(n4749), .ZN(n9262) );
  AOI22_X2 U5914 ( .A1(n9183), .A2(n9185), .B1(n9195), .B2(n9172), .ZN(n9166)
         );
  INV_X1 U5915 ( .A(n4729), .ZN(n8977) );
  NAND2_X1 U5916 ( .A1(n4403), .A2(n4401), .ZN(n5043) );
  OAI21_X1 U5917 ( .B1(n5085), .B2(n5084), .A(n5086), .ZN(n5105) );
  NAND2_X1 U5918 ( .A1(n4427), .A2(n4431), .ZN(n5344) );
  INV_X1 U5919 ( .A(n5604), .ZN(n5602) );
  INV_X4 U5920 ( .A(n7749), .ZN(n7799) );
  OAI21_X1 U5921 ( .B1(n7908), .B2(n4331), .A(n4330), .ZN(P2_U3242) );
  NAND2_X1 U5922 ( .A1(n4784), .A2(n4783), .ZN(n4782) );
  NAND2_X2 U5923 ( .A1(n8222), .A2(n8223), .ZN(n8200) );
  NAND2_X1 U5924 ( .A1(n4763), .A2(n4766), .ZN(n6935) );
  NOR2_X2 U5925 ( .A1(n5173), .A2(n4782), .ZN(n5402) );
  NAND3_X1 U5926 ( .A1(n7815), .A2(n7813), .A3(n4335), .ZN(P2_U3222) );
  NAND2_X1 U5927 ( .A1(n4399), .A2(n4606), .ZN(n4996) );
  NAND2_X1 U5928 ( .A1(n7756), .A2(n7838), .ZN(n4586) );
  INV_X1 U5929 ( .A(n4588), .ZN(n7908) );
  AND2_X1 U5930 ( .A1(n7000), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5931 ( .A1(n8479), .A2(n8480), .ZN(n8574) );
  NAND2_X1 U5932 ( .A1(n6273), .A2(n6274), .ZN(n6275) );
  OR2_X2 U5933 ( .A1(n8530), .A2(n7581), .ZN(n7589) );
  NAND2_X1 U5934 ( .A1(n4494), .A2(n6861), .ZN(n6905) );
  INV_X1 U5935 ( .A(n7660), .ZN(n7662) );
  NAND2_X1 U5936 ( .A1(n7672), .A2(n4492), .ZN(n8511) );
  OR3_X1 U5937 ( .A1(n8454), .A2(n8466), .A3(n4495), .ZN(n8470) );
  NAND3_X1 U5938 ( .A1(n4676), .A2(n4283), .A3(n6277), .ZN(n6493) );
  NAND2_X1 U5939 ( .A1(n5674), .A2(n5673), .ZN(n5777) );
  AOI21_X1 U5940 ( .B1(n4339), .B2(n4911), .A(n4307), .ZN(n4467) );
  XNOR2_X1 U5941 ( .A(n4339), .B(n4911), .ZN(n5858) );
  NAND3_X1 U5942 ( .A1(n4341), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4340) );
  NAND3_X1 U5943 ( .A1(n4860), .A2(n4344), .A3(n4343), .ZN(n4342) );
  NAND3_X1 U5944 ( .A1(n5515), .A2(n5525), .A3(n5535), .ZN(n4349) );
  NAND2_X1 U5945 ( .A1(n7943), .A2(n9893), .ZN(n5575) );
  NAND2_X1 U5946 ( .A1(n4709), .A2(n4366), .ZN(n4364) );
  NAND2_X1 U5947 ( .A1(n4364), .A2(n4365), .ZN(n5604) );
  NOR2_X1 U5948 ( .A1(n5559), .A2(n5569), .ZN(n4375) );
  NAND2_X1 U5949 ( .A1(n5547), .A2(n4379), .ZN(n4378) );
  NAND2_X1 U5950 ( .A1(n4384), .A2(n4394), .ZN(n4385) );
  NAND2_X1 U5951 ( .A1(n4309), .A2(n4388), .ZN(n4384) );
  NAND3_X1 U5952 ( .A1(n5489), .A2(n4394), .A3(n4387), .ZN(n4386) );
  AND2_X1 U5953 ( .A1(n5487), .A2(n5569), .ZN(n4398) );
  NAND2_X1 U5954 ( .A1(n5005), .A2(n4404), .ZN(n4403) );
  AOI21_X1 U5955 ( .B1(n5362), .B2(n4271), .A(n4323), .ZN(n4414) );
  NAND2_X1 U5956 ( .A1(n4415), .A2(n5363), .ZN(n5382) );
  NOR2_X1 U5957 ( .A1(n5381), .A2(n4411), .ZN(n4413) );
  NAND2_X1 U5958 ( .A1(n4715), .A2(n4422), .ZN(n4420) );
  NAND2_X1 U5959 ( .A1(n5297), .A2(n5296), .ZN(n4437) );
  NAND2_X1 U5960 ( .A1(n5297), .A2(n4428), .ZN(n4427) );
  NAND2_X1 U5961 ( .A1(n5798), .A2(n4453), .ZN(n4454) );
  OAI21_X2 U5962 ( .B1(n5798), .B2(n5863), .A(n4454), .ZN(n6076) );
  INV_X1 U5963 ( .A(n5798), .ZN(n6269) );
  INV_X1 U5964 ( .A(n4465), .ZN(n9058) );
  INV_X1 U5965 ( .A(n4473), .ZN(n6803) );
  INV_X1 U5966 ( .A(n4479), .ZN(n8169) );
  NAND2_X1 U5967 ( .A1(n8086), .A2(n4487), .ZN(n8060) );
  NAND2_X1 U5968 ( .A1(n8086), .A2(n8079), .ZN(n8074) );
  NAND3_X1 U5969 ( .A1(n4483), .A2(n4482), .A3(n4480), .ZN(n8286) );
  NAND3_X1 U5970 ( .A1(n4491), .A2(n4489), .A3(n4488), .ZN(n8216) );
  INV_X1 U5971 ( .A(n4491), .ZN(n8275) );
  AOI21_X1 U5972 ( .B1(n8425), .B2(n4492), .A(n8512), .ZN(n8513) );
  NAND2_X1 U5973 ( .A1(n8426), .A2(n8428), .ZN(n4492) );
  INV_X1 U5974 ( .A(n4494), .ZN(n4493) );
  AND2_X2 U5975 ( .A1(n8575), .A2(n4821), .ZN(n8454) );
  NAND2_X2 U5976 ( .A1(n8574), .A2(n7686), .ZN(n8575) );
  NAND2_X1 U5977 ( .A1(n8555), .A2(n4503), .ZN(n4496) );
  INV_X1 U5978 ( .A(n4507), .ZN(n8553) );
  NAND2_X1 U5979 ( .A1(n7121), .A2(n7204), .ZN(n4508) );
  NAND2_X1 U5980 ( .A1(n4508), .A2(n4509), .ZN(n7569) );
  NAND2_X1 U5981 ( .A1(n4700), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U5982 ( .A1(n5805), .A2(n5630), .ZN(n5662) );
  INV_X1 U5983 ( .A(n5916), .ZN(n4518) );
  OAI21_X1 U5984 ( .B1(n5916), .B2(n4261), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5687) );
  OAI21_X1 U5985 ( .B1(n4518), .B2(n6206), .A(n4519), .ZN(n5688) );
  INV_X1 U5986 ( .A(n4520), .ZN(n5692) );
  NOR2_X2 U5989 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4522) );
  NOR2_X2 U5990 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4523) );
  NAND2_X1 U5991 ( .A1(n6269), .A2(n6013), .ZN(n4536) );
  NAND3_X1 U5992 ( .A1(n4534), .A2(n5852), .A3(n5798), .ZN(n4533) );
  INV_X1 U5993 ( .A(n8837), .ZN(n4542) );
  AOI21_X1 U5994 ( .B1(n4541), .B2(n4539), .A(n4538), .ZN(n4537) );
  NOR2_X1 U5995 ( .A1(n6817), .A2(n4542), .ZN(n4541) );
  INV_X1 U5996 ( .A(n8674), .ZN(n8673) );
  AND2_X1 U5997 ( .A1(n5805), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5998 ( .A1(n5638), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U5999 ( .A1(n5638), .A2(n4546), .ZN(n4714) );
  NAND3_X1 U6000 ( .A1(n4560), .A2(n4556), .A3(n4555), .ZN(n4554) );
  NAND2_X1 U6001 ( .A1(n4566), .A2(n4564), .ZN(n8871) );
  NAND2_X1 U6002 ( .A1(n4569), .A2(n4567), .ZN(n4566) );
  INV_X1 U6003 ( .A(n4568), .ZN(n4567) );
  OAI21_X1 U6004 ( .B1(n8862), .B2(n8861), .A(n8863), .ZN(n4568) );
  NAND2_X1 U6005 ( .A1(n8860), .A2(n8859), .ZN(n4569) );
  NAND2_X1 U6006 ( .A1(n6888), .A2(n4573), .ZN(n4572) );
  AOI21_X2 U6007 ( .B1(n6843), .B2(n4575), .A(n4574), .ZN(n4573) );
  OAI21_X1 U6008 ( .B1(n7877), .B2(n4579), .A(n4577), .ZN(n7747) );
  XNOR2_X1 U6009 ( .A(n7747), .B(n7745), .ZN(n7891) );
  OAI21_X1 U6010 ( .B1(n7877), .B2(n7876), .A(n7740), .ZN(n7830) );
  NAND2_X1 U6011 ( .A1(n7876), .A2(n7740), .ZN(n4581) );
  AND2_X2 U6012 ( .A1(n5402), .A2(n4836), .ZN(n5431) );
  NAND2_X1 U6013 ( .A1(n7756), .A2(n7755), .ZN(n4585) );
  NAND2_X1 U6014 ( .A1(n4588), .A2(n4587), .ZN(n7769) );
  NAND3_X1 U6015 ( .A1(n4586), .A2(n4585), .A3(n4321), .ZN(n4588) );
  NAND3_X1 U6016 ( .A1(n4586), .A2(n4585), .A3(n4583), .ZN(n7910) );
  NAND2_X1 U6017 ( .A1(n7847), .A2(n4589), .ZN(n7856) );
  OAI211_X2 U6018 ( .C1(n4885), .C2(n5864), .A(n4593), .B(n4592), .ZN(n6470)
         );
  OR2_X1 U6019 ( .A1(n6112), .A2(n9476), .ZN(n4592) );
  NAND2_X2 U6020 ( .A1(n6112), .A2(n5852), .ZN(n4882) );
  NAND2_X2 U6021 ( .A1(n6112), .A2(n4619), .ZN(n4885) );
  OR2_X1 U6022 ( .A1(n4885), .A2(n5856), .ZN(n4594) );
  INV_X2 U6023 ( .A(n4885), .ZN(n5427) );
  OAI22_X1 U6024 ( .A1(n8663), .A2(n4885), .B1(n9415), .B2(n5396), .ZN(n8023)
         );
  NAND2_X1 U6025 ( .A1(n6873), .A2(n4597), .ZN(n6795) );
  NAND2_X1 U6026 ( .A1(n6795), .A2(n4598), .ZN(n7054) );
  NAND2_X1 U6027 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  INV_X1 U6028 ( .A(n6786), .ZN(n4599) );
  NAND2_X1 U6029 ( .A1(n4601), .A2(n4602), .ZN(n8048) );
  NAND2_X1 U6030 ( .A1(n8084), .A2(n4272), .ZN(n4601) );
  NAND2_X1 U6031 ( .A1(n8084), .A2(n8093), .ZN(n8083) );
  OAI21_X1 U6032 ( .B1(n4948), .B2(n4609), .A(n4607), .ZN(n4993) );
  NAND2_X1 U6033 ( .A1(n4948), .A2(n4947), .ZN(n4969) );
  INV_X1 U6034 ( .A(n4968), .ZN(n4609) );
  NAND2_X1 U6035 ( .A1(n7140), .A2(n4613), .ZN(n4610) );
  NAND2_X1 U6036 ( .A1(n5047), .A2(n5046), .ZN(n7163) );
  INV_X8 U6037 ( .A(n4861), .ZN(n5852) );
  MUX2_X1 U6038 ( .A(n4914), .B(n5861), .S(n4619), .Z(n4934) );
  MUX2_X1 U6039 ( .A(n4901), .B(n5859), .S(n4619), .Z(n4912) );
  NAND2_X1 U6040 ( .A1(n8027), .A2(n4621), .ZN(n4623) );
  INV_X1 U6041 ( .A(n4623), .ZN(n8272) );
  OR2_X1 U6042 ( .A1(n8028), .A2(n8267), .ZN(n4624) );
  NAND2_X1 U6043 ( .A1(n8188), .A2(n4308), .ZN(n4626) );
  NAND2_X1 U6044 ( .A1(n9074), .A2(n4638), .ZN(n4635) );
  OAI21_X1 U6045 ( .B1(n9513), .B2(n4647), .A(n4648), .ZN(n9154) );
  INV_X1 U6046 ( .A(n9167), .ZN(n4653) );
  NAND2_X1 U6047 ( .A1(n6639), .A2(n4310), .ZN(n4656) );
  INV_X1 U6048 ( .A(n8807), .ZN(n6420) );
  OR2_X1 U6049 ( .A1(n7528), .A2(n8600), .ZN(n4665) );
  OAI21_X1 U6050 ( .B1(n7528), .B2(n4315), .A(n4658), .ZN(n8985) );
  NAND2_X1 U6051 ( .A1(n9134), .A2(n4669), .ZN(n4666) );
  NAND2_X1 U6052 ( .A1(n4666), .A2(n4667), .ZN(n9092) );
  NAND3_X1 U6053 ( .A1(n8490), .A2(n8492), .A3(n4673), .ZN(n4672) );
  NAND3_X1 U6054 ( .A1(n8491), .A2(n8492), .A3(n7609), .ZN(n8493) );
  NAND3_X1 U6055 ( .A1(n4678), .A2(n4677), .A3(n6267), .ZN(n4676) );
  OAI21_X1 U6056 ( .B1(n6195), .B2(n6196), .A(n5733), .ZN(n6268) );
  NAND2_X1 U6057 ( .A1(n6196), .A2(n5733), .ZN(n4677) );
  NAND2_X1 U6058 ( .A1(n6195), .A2(n5733), .ZN(n4678) );
  NAND2_X1 U6059 ( .A1(n4695), .A2(n5627), .ZN(P2_U3244) );
  NAND2_X1 U6060 ( .A1(n4696), .A2(n5612), .ZN(n4695) );
  NAND2_X1 U6061 ( .A1(n4697), .A2(n4297), .ZN(n4696) );
  NOR2_X1 U6062 ( .A1(n5605), .A2(n5613), .ZN(n4697) );
  NAND2_X1 U6063 ( .A1(n8524), .A2(n4701), .ZN(n4698) );
  INV_X1 U6064 ( .A(n4702), .ZN(n8473) );
  INV_X1 U6065 ( .A(n8472), .ZN(n4701) );
  NAND3_X1 U6066 ( .A1(n6907), .A2(n6906), .A3(n4707), .ZN(n4704) );
  NAND2_X2 U6067 ( .A1(n4996), .A2(n4995), .ZN(n5005) );
  OAI21_X2 U6068 ( .B1(n4714), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5644) );
  OAI21_X2 U6069 ( .B1(n5255), .B2(n4716), .A(n5259), .ZN(n5275) );
  OAI21_X2 U6070 ( .B1(n5059), .B2(n5058), .A(n5057), .ZN(n5085) );
  INV_X2 U6071 ( .A(n8451), .ZN(n7625) );
  NAND2_X2 U6072 ( .A1(n5694), .A2(n7649), .ZN(n8451) );
  AND2_X2 U6073 ( .A1(n5768), .A2(n5693), .ZN(n7649) );
  OR2_X2 U6074 ( .A1(n5746), .A2(n4717), .ZN(n5768) );
  INV_X1 U6075 ( .A(n6584), .ZN(n4721) );
  NAND2_X1 U6076 ( .A1(n6585), .A2(n6584), .ZN(n9692) );
  NAND2_X1 U6077 ( .A1(n6417), .A2(n8805), .ZN(n6585) );
  AND2_X1 U6078 ( .A1(n6436), .A2(n6415), .ZN(n6417) );
  NAND2_X1 U6079 ( .A1(n9035), .A2(n7435), .ZN(n4723) );
  NAND2_X1 U6080 ( .A1(n9035), .A2(n4727), .ZN(n4726) );
  NAND2_X1 U6081 ( .A1(n4723), .A2(n4722), .ZN(n7507) );
  AOI21_X2 U6082 ( .B1(n9022), .B2(n4730), .A(n4732), .ZN(n4729) );
  NAND2_X1 U6083 ( .A1(n4739), .A2(n4741), .ZN(n9049) );
  NAND2_X1 U6084 ( .A1(n9084), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U6085 ( .A1(n6810), .A2(n4312), .ZN(n4743) );
  NAND2_X1 U6086 ( .A1(n9151), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U6087 ( .A1(n7190), .A2(n4757), .ZN(n4756) );
  NOR2_X1 U6088 ( .A1(n7351), .A2(n4759), .ZN(n9512) );
  AND2_X1 U6089 ( .A1(n7352), .A2(n9517), .ZN(n4759) );
  AND2_X2 U6090 ( .A1(n5645), .A2(n4314), .ZN(n5672) );
  NAND2_X1 U6091 ( .A1(n5645), .A2(n4761), .ZN(n5675) );
  NAND2_X1 U6092 ( .A1(n6785), .A2(n4764), .ZN(n4763) );
  OAI21_X2 U6093 ( .B1(n5169), .B2(n4774), .A(n4771), .ZN(n8235) );
  NAND2_X1 U6094 ( .A1(n8139), .A2(n4779), .ZN(n4776) );
  NAND2_X1 U6095 ( .A1(n4776), .A2(n4777), .ZN(n8105) );
  NAND2_X4 U6096 ( .A1(n4848), .A2(n8401), .ZN(n5398) );
  INV_X1 U6097 ( .A(n4923), .ZN(n5409) );
  OAI21_X2 U6098 ( .B1(n8200), .B2(n4797), .A(n4793), .ZN(n8158) );
  NAND2_X2 U6099 ( .A1(n7147), .A2(n4800), .ZN(n7272) );
  OAI21_X2 U6100 ( .B1(n8092), .B2(n8093), .A(n5549), .ZN(n8067) );
  NAND2_X1 U6101 ( .A1(n5431), .A2(n4257), .ZN(n4842) );
  NAND2_X1 U6102 ( .A1(n6795), .A2(n6794), .ZN(n7095) );
  NAND2_X1 U6103 ( .A1(n8833), .A2(n8832), .ZN(n8860) );
  NAND2_X1 U6104 ( .A1(n8862), .A2(n8799), .ZN(n8833) );
  NAND2_X1 U6105 ( .A1(n8784), .A2(n8852), .ZN(n8787) );
  NAND2_X1 U6106 ( .A1(n8858), .A2(n9125), .ZN(n8859) );
  CLKBUF_X1 U6107 ( .A(n7856), .Z(n7897) );
  CLKBUF_X1 U6108 ( .A(n7536), .Z(n7538) );
  XNOR2_X1 U6109 ( .A(n6470), .B(n7749), .ZN(n6058) );
  NAND2_X1 U6110 ( .A1(n5714), .A2(n5715), .ZN(n6069) );
  AOI21_X2 U6111 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(n6515) );
  OR2_X1 U6112 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U6113 ( .A1(n8052), .A2(n8051), .ZN(n8057) );
  AOI21_X1 U6114 ( .B1(n7507), .B2(n7520), .A(n7519), .ZN(n7521) );
  OAI21_X1 U6115 ( .B1(n9839), .B2(n5462), .A(n5574), .ZN(n6603) );
  NOR2_X1 U6116 ( .A1(n9870), .A2(n7540), .ZN(n6375) );
  OR2_X1 U6117 ( .A1(n4334), .A2(n6152), .ZN(n4803) );
  AND2_X1 U6118 ( .A1(n7798), .A2(n6337), .ZN(n4804) );
  INV_X1 U6119 ( .A(n8332), .ZN(n8018) );
  OR2_X1 U6120 ( .A1(n8866), .A2(n6425), .ZN(n9685) );
  INV_X1 U6121 ( .A(n9685), .ZN(n9700) );
  INV_X1 U6122 ( .A(n9898), .ZN(n9919) );
  OR2_X1 U6123 ( .A1(n9178), .A2(n9189), .ZN(n4806) );
  NOR2_X1 U6124 ( .A1(n5141), .A2(n7268), .ZN(n4807) );
  OR2_X1 U6125 ( .A1(n9162), .A2(n9171), .ZN(n4808) );
  OR2_X1 U6126 ( .A1(n9112), .A2(n9123), .ZN(n4809) );
  OR2_X1 U6127 ( .A1(n9090), .A2(n9106), .ZN(n4810) );
  AND2_X1 U6128 ( .A1(n7811), .A2(n7919), .ZN(n4812) );
  OR2_X1 U6129 ( .A1(n6112), .A2(n5855), .ZN(n4813) );
  NOR2_X1 U6130 ( .A1(n6419), .A2(n8448), .ZN(n4814) );
  INV_X1 U6131 ( .A(n6824), .ZN(n6802) );
  INV_X2 U6132 ( .A(n9846), .ZN(n9848) );
  AND2_X1 U6133 ( .A1(n5023), .A2(n5011), .ZN(n4815) );
  AND2_X1 U6134 ( .A1(n5042), .A2(n5027), .ZN(n4816) );
  INV_X1 U6135 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5639) );
  INV_X1 U6136 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4836) );
  AND2_X1 U6137 ( .A1(n6424), .A2(n6423), .ZN(n9682) );
  AND2_X1 U6138 ( .A1(n5106), .A2(n5090), .ZN(n4817) );
  INV_X1 U6139 ( .A(n8234), .ZN(n5203) );
  AND2_X1 U6140 ( .A1(n4916), .A2(n4803), .ZN(n4818) );
  INV_X1 U6141 ( .A(n7934), .ZN(n8269) );
  AND4_X1 U6142 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n7934)
         );
  OR2_X1 U6143 ( .A1(n8291), .A2(n9921), .ZN(n4819) );
  OR2_X1 U6144 ( .A1(n8221), .A2(n8033), .ZN(n4820) );
  AND2_X1 U6145 ( .A1(n7700), .A2(n7699), .ZN(n4821) );
  OR2_X1 U6146 ( .A1(n8233), .A2(n8030), .ZN(n4823) );
  AND3_X1 U6147 ( .A1(n5457), .A2(n5460), .A3(n5456), .ZN(n4824) );
  OR2_X1 U6148 ( .A1(n6768), .A2(n6758), .ZN(n9927) );
  INV_X2 U6149 ( .A(n9940), .ZN(n9943) );
  INV_X2 U6150 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR2_X1 U6151 ( .A1(n5676), .A2(n6206), .ZN(n4825) );
  NAND2_X1 U6152 ( .A1(n5441), .A2(n5535), .ZN(n5466) );
  AND2_X1 U6153 ( .A1(n6571), .A2(n5466), .ZN(n5467) );
  NAND2_X1 U6154 ( .A1(n4778), .A2(n5535), .ZN(n5541) );
  AND2_X1 U6155 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  MUX2_X1 U6156 ( .A(n8768), .B(n8785), .S(n9222), .Z(n8769) );
  INV_X1 U6157 ( .A(n5535), .ZN(n5569) );
  NOR2_X1 U6158 ( .A1(n8828), .A2(n8775), .ZN(n8786) );
  INV_X1 U6159 ( .A(n8106), .ZN(n5341) );
  NOR3_X1 U6160 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4837) );
  NAND2_X1 U6161 ( .A1(n8790), .A2(n8775), .ZN(n8791) );
  OR4_X1 U6162 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5757) );
  INV_X1 U6163 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5650) );
  INV_X1 U6164 ( .A(n6742), .ZN(n6740) );
  INV_X1 U6165 ( .A(n6064), .ZN(n6061) );
  INV_X1 U6166 ( .A(n6878), .ZN(n6782) );
  INV_X1 U6167 ( .A(P2_B_REG_SCAN_IN), .ZN(n6024) );
  AND2_X1 U6168 ( .A1(n8425), .A2(n8512), .ZN(n7672) );
  OR2_X1 U6169 ( .A1(n7418), .A2(n8545), .ZN(n7429) );
  INV_X1 U6170 ( .A(SI_20_), .ZN(n5225) );
  INV_X1 U6171 ( .A(SI_16_), .ZN(n5148) );
  AND2_X1 U6172 ( .A1(n5983), .A2(n5982), .ZN(n6205) );
  INV_X1 U6173 ( .A(n7255), .ZN(n7253) );
  INV_X1 U6174 ( .A(n7849), .ZN(n7717) );
  OR2_X1 U6175 ( .A1(n5075), .A2(n5074), .ZN(n5097) );
  INV_X1 U6176 ( .A(n6555), .ZN(n6522) );
  OR2_X1 U6177 ( .A1(n5249), .A2(n7831), .ZN(n5286) );
  OR2_X1 U6178 ( .A1(n5016), .A2(n6894), .ZN(n5035) );
  INV_X1 U6179 ( .A(n8055), .ZN(n8056) );
  NAND2_X1 U6180 ( .A1(n5608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5610) );
  INV_X1 U6181 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5069) );
  INV_X1 U6182 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7356) );
  INV_X1 U6183 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6712) );
  OR2_X1 U6184 ( .A1(n7439), .A2(n8484), .ZN(n7451) );
  NOR2_X1 U6185 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  NAND2_X1 U6186 ( .A1(n7484), .A2(n8719), .ZN(n9134) );
  OR2_X1 U6187 ( .A1(n7186), .A2(n8881), .ZN(n7187) );
  OR2_X1 U6188 ( .A1(n6309), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6310) );
  OR2_X1 U6189 ( .A1(n6205), .A2(n6206), .ZN(n5986) );
  OR2_X1 U6190 ( .A1(n5396), .A2(n7312), .ZN(n5352) );
  INV_X1 U6191 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9346) );
  OR2_X1 U6192 ( .A1(n6091), .A2(n6048), .ZN(n6751) );
  INV_X1 U6193 ( .A(n8028), .ZN(n8366) );
  OR2_X1 U6194 ( .A1(n5398), .A2(n6081), .ZN(n4876) );
  INV_X1 U6195 ( .A(n4334), .ZN(n5886) );
  OR2_X1 U6196 ( .A1(n8349), .A2(n8242), .ZN(n8031) );
  OR2_X1 U6197 ( .A1(n7095), .A2(n7088), .ZN(n6933) );
  AND2_X1 U6198 ( .A1(n9865), .A2(n6040), .ZN(n9898) );
  OR2_X1 U6199 ( .A1(n4989), .A2(n4988), .ZN(n5012) );
  OR2_X1 U6200 ( .A1(n7357), .A2(n7356), .ZN(n7367) );
  INV_X1 U6201 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U6202 ( .A1(n7317), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7378) );
  OR2_X1 U6203 ( .A1(n7398), .A2(n7397), .ZN(n7408) );
  AND3_X1 U6204 ( .A1(n6399), .A2(n7223), .A3(n6397), .ZN(n5789) );
  NAND2_X1 U6205 ( .A1(n5840), .A2(n5839), .ZN(n9656) );
  INV_X1 U6206 ( .A(n8874), .ZN(n9011) );
  INV_X1 U6207 ( .A(n8876), .ZN(n9027) );
  NOR2_X1 U6208 ( .A1(n9244), .A2(n9077), .ZN(n7423) );
  INV_X1 U6209 ( .A(n8877), .ZN(n9156) );
  OR2_X1 U6210 ( .A1(n7030), .A2(n7029), .ZN(n7126) );
  INV_X1 U6211 ( .A(n5969), .ZN(n5790) );
  AND2_X1 U6212 ( .A1(n5775), .A2(n5774), .ZN(n6419) );
  AND2_X1 U6213 ( .A1(n8703), .A2(n8702), .ZN(n8814) );
  INV_X1 U6214 ( .A(n8881), .ZN(n9536) );
  AND2_X1 U6215 ( .A1(n6816), .A2(n8836), .ZN(n9681) );
  NAND2_X1 U6216 ( .A1(n4814), .A2(n9125), .ZN(n9726) );
  OR2_X1 U6217 ( .A1(n5874), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5751) );
  XNOR2_X1 U6218 ( .A(n5648), .B(n5639), .ZN(n7080) );
  INV_X1 U6219 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5668) );
  AND2_X1 U6220 ( .A1(n5172), .A2(n5151), .ZN(n5170) );
  OR3_X1 U6221 ( .A1(n7299), .A2(n7305), .A3(n7170), .ZN(n6251) );
  INV_X1 U6222 ( .A(n8310), .ZN(n8114) );
  AND3_X1 U6223 ( .A1(n5360), .A2(n5359), .A3(n5358), .ZN(n8108) );
  AND4_X1 U6224 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n7851)
         );
  INV_X1 U6225 ( .A(n9817), .ZN(n9812) );
  INV_X1 U6226 ( .A(n9814), .ZN(n9483) );
  INV_X1 U6227 ( .A(n8037), .ZN(n8140) );
  AND2_X1 U6228 ( .A1(n7228), .A2(n7143), .ZN(n8372) );
  INV_X1 U6229 ( .A(n7280), .ZN(n8259) );
  AND2_X1 U6230 ( .A1(n8253), .A2(n6367), .ZN(n7159) );
  NAND2_X1 U6231 ( .A1(n6338), .A2(n6337), .ZN(n8271) );
  NAND2_X1 U6232 ( .A1(n6039), .A2(n6038), .ZN(n6767) );
  INV_X1 U6233 ( .A(n9921), .ZN(n9899) );
  INV_X1 U6234 ( .A(n9925), .ZN(n9904) );
  NAND2_X1 U6235 ( .A1(n6883), .A2(n9880), .ZN(n9925) );
  AND2_X1 U6236 ( .A1(n6027), .A2(n6026), .ZN(n9849) );
  INV_X1 U6237 ( .A(n5616), .ZN(n5618) );
  AND2_X1 U6238 ( .A1(n5127), .A2(n5110), .ZN(n6948) );
  AND2_X1 U6239 ( .A1(n4619), .A2(P2_U3152), .ZN(n8405) );
  AND2_X1 U6240 ( .A1(n5970), .A2(n5969), .ZN(n6398) );
  AND2_X1 U6241 ( .A1(n7501), .A2(n7500), .ZN(n8986) );
  OR2_X1 U6242 ( .A1(n8482), .A2(n4249), .ZN(n7446) );
  INV_X1 U6243 ( .A(n9656), .ZN(n9634) );
  INV_X1 U6244 ( .A(n9605), .ZN(n9659) );
  INV_X1 U6245 ( .A(n8956), .ZN(n9665) );
  AND2_X1 U6246 ( .A1(n9719), .A2(n9125), .ZN(n9144) );
  INV_X1 U6247 ( .A(n9682), .ZN(n9707) );
  INV_X1 U6248 ( .A(n9179), .ZN(n9699) );
  NAND2_X1 U6249 ( .A1(n8798), .A2(n6931), .ZN(n5978) );
  INV_X1 U6250 ( .A(n9790), .ZN(n9288) );
  NAND2_X1 U6251 ( .A1(n9726), .A2(n9730), .ZN(n9790) );
  INV_X1 U6252 ( .A(n7223), .ZN(n6400) );
  INV_X1 U6253 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5643) );
  AND2_X1 U6254 ( .A1(n5987), .A2(n6192), .ZN(n7172) );
  OAI21_X1 U6255 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9951), .ZN(n9980) );
  INV_X1 U6256 ( .A(n9472), .ZN(n9820) );
  AOI22_X1 U6257 ( .A1(n7769), .A2(n7919), .B1(n7768), .B2(n7767), .ZN(n7775)
         );
  INV_X1 U6258 ( .A(n7919), .ZN(n7909) );
  INV_X1 U6259 ( .A(n8144), .ZN(n8041) );
  INV_X1 U6260 ( .A(n7833), .ZN(n8224) );
  INV_X1 U6261 ( .A(n8255), .ZN(n8281) );
  NAND2_X1 U6262 ( .A1(n6575), .A2(n8250), .ZN(n9846) );
  AND2_X1 U6263 ( .A1(n6360), .A2(n6359), .ZN(n9885) );
  OR2_X1 U6264 ( .A1(n6768), .A2(n6767), .ZN(n9940) );
  AND2_X1 U6265 ( .A1(n9885), .A2(n9884), .ZN(n9932) );
  NOR2_X1 U6266 ( .A1(n9850), .A2(n9849), .ZN(n9857) );
  INV_X1 U6267 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9858) );
  INV_X1 U6268 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7300) );
  INV_X1 U6269 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6452) );
  INV_X1 U6270 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5920) );
  INV_X1 U6271 ( .A(n9259), .ZN(n9112) );
  INV_X1 U6272 ( .A(n8594), .ZN(n8483) );
  AND2_X1 U6273 ( .A1(n5791), .A2(n9118), .ZN(n8591) );
  NAND2_X1 U6274 ( .A1(n7476), .A2(n7475), .ZN(n8874) );
  INV_X1 U6275 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9604) );
  INV_X1 U6276 ( .A(n9661), .ZN(n9622) );
  INV_X1 U6277 ( .A(n9698), .ZN(n8974) );
  AND2_X1 U6278 ( .A1(n6720), .A2(n6719), .ZN(n9781) );
  NAND2_X1 U6279 ( .A1(n9719), .A2(n4814), .ZN(n9198) );
  INV_X1 U6280 ( .A(n9811), .ZN(n9809) );
  AND3_X1 U6281 ( .A1(n9782), .A2(n9781), .A3(n9780), .ZN(n9808) );
  INV_X1 U6282 ( .A(n9794), .ZN(n9792) );
  NAND2_X1 U6283 ( .A1(n5874), .A2(n5969), .ZN(n9725) );
  INV_X1 U6284 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5875) );
  INV_X1 U6285 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7053) );
  INV_X1 U6286 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5923) );
  AND2_X1 U6288 ( .A1(n5800), .A2(n9863), .ZN(P2_U3966) );
  INV_X1 U6289 ( .A(n8888), .ZN(P1_U4006) );
  NOR2_X1 U6290 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4829) );
  NOR2_X1 U6291 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4831) );
  AND2_X2 U6292 ( .A1(n4869), .A2(n4831), .ZN(n4932) );
  NOR2_X2 U6293 ( .A1(n4842), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4841) );
  OR2_X2 U6294 ( .A1(n4841), .A2(n5069), .ZN(n4840) );
  INV_X1 U6295 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4839) );
  XNOR2_X2 U6296 ( .A(n4840), .B(n4839), .ZN(n4846) );
  INV_X1 U6297 ( .A(n4841), .ZN(n8396) );
  NAND2_X1 U6298 ( .A1(n4842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4843) );
  MUX2_X1 U6299 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4843), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4844) );
  NAND2_X1 U6300 ( .A1(n4919), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4852) );
  INV_X2 U6301 ( .A(n4846), .ZN(n4848) );
  INV_X2 U6302 ( .A(n4845), .ZN(n8401) );
  INV_X1 U6303 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4847) );
  OR2_X1 U6304 ( .A1(n4923), .A2(n4847), .ZN(n4850) );
  INV_X1 U6305 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9362) );
  OR2_X1 U6306 ( .A1(n5398), .A2(n9362), .ZN(n4849) );
  NAND2_X1 U6307 ( .A1(n4857), .A2(n4853), .ZN(n4856) );
  INV_X1 U6308 ( .A(n4857), .ZN(n4858) );
  NAND2_X1 U6309 ( .A1(n4858), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4859) );
  AND2_X1 U6310 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6311 ( .A1(n5852), .A2(n4862), .ZN(n5680) );
  NAND3_X1 U6312 ( .A1(n4619), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4863) );
  NAND2_X1 U6313 ( .A1(n5680), .A2(n4863), .ZN(n4865) );
  INV_X1 U6314 ( .A(SI_1_), .ZN(n4864) );
  XNOR2_X1 U6315 ( .A(n4865), .B(n4864), .ZN(n4884) );
  MUX2_X1 U6316 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5852), .Z(n4883) );
  NAND2_X1 U6317 ( .A1(n4884), .A2(n4883), .ZN(n4867) );
  NAND2_X1 U6318 ( .A1(n4865), .A2(SI_1_), .ZN(n4866) );
  NAND2_X1 U6319 ( .A1(n4867), .A2(n4866), .ZN(n4897) );
  MUX2_X1 U6320 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n4619), .Z(n4898) );
  INV_X1 U6321 ( .A(SI_2_), .ZN(n4868) );
  XNOR2_X1 U6322 ( .A(n4898), .B(n4868), .ZN(n4896) );
  XNOR2_X1 U6323 ( .A(n4897), .B(n4896), .ZN(n5856) );
  INV_X1 U6324 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5857) );
  OR2_X1 U6325 ( .A1(n4869), .A2(n5069), .ZN(n4870) );
  XNOR2_X1 U6326 ( .A(n4870), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9488) );
  INV_X1 U6327 ( .A(n9488), .ZN(n5855) );
  INV_X1 U6328 ( .A(n6373), .ZN(n4890) );
  NAND2_X1 U6329 ( .A1(n4919), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4874) );
  INV_X1 U6330 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4872) );
  INV_X1 U6331 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4875) );
  INV_X1 U6332 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6081) );
  NAND3_X2 U6333 ( .A1(n4878), .A2(n4877), .A3(n4876), .ZN(n6055) );
  NAND2_X1 U6334 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4879) );
  MUX2_X1 U6335 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4879), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4881) );
  INV_X1 U6336 ( .A(n4869), .ZN(n4880) );
  NAND2_X1 U6337 ( .A1(n4881), .A2(n4880), .ZN(n9476) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U6339 ( .A(n4884), .B(n4883), .ZN(n5864) );
  NAND2_X1 U6340 ( .A1(n4919), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4886) );
  INV_X1 U6341 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U6342 ( .A1(n4619), .A2(SI_0_), .ZN(n4887) );
  XNOR2_X1 U6343 ( .A(n4887), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8409) );
  MUX2_X1 U6344 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8409), .S(n6112), .Z(n9864) );
  NAND2_X1 U6345 ( .A1(n4888), .A2(n9864), .ZN(n6467) );
  NAND2_X1 U6346 ( .A1(n5579), .A2(n6467), .ZN(n5445) );
  INV_X1 U6347 ( .A(n6470), .ZN(n6346) );
  NAND2_X1 U6348 ( .A1(n5445), .A2(n5578), .ZN(n6372) );
  INV_X1 U6349 ( .A(n6372), .ZN(n4889) );
  NAND2_X1 U6350 ( .A1(n4890), .A2(n4889), .ZN(n6352) );
  NAND2_X1 U6351 ( .A1(n6352), .A2(n6353), .ZN(n4904) );
  NAND2_X1 U6352 ( .A1(n4251), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U6353 ( .A1(n5288), .A2(n9318), .ZN(n4893) );
  OR2_X1 U6354 ( .A1(n4924), .A2(n9886), .ZN(n4892) );
  INV_X1 U6355 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6361) );
  OR2_X1 U6356 ( .A1(n5398), .A2(n6361), .ZN(n4891) );
  AND4_X2 U6357 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n6480)
         );
  NAND2_X1 U6358 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4279), .ZN(n4895) );
  XNOR2_X1 U6359 ( .A(n4895), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6102) );
  INV_X1 U6360 ( .A(n6102), .ZN(n6163) );
  INV_X1 U6361 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5859) );
  OR2_X1 U6362 ( .A1(n4882), .A2(n5859), .ZN(n4903) );
  NAND2_X1 U6363 ( .A1(n4897), .A2(n4896), .ZN(n4900) );
  NAND2_X1 U6364 ( .A1(n4898), .A2(SI_2_), .ZN(n4899) );
  INV_X1 U6365 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4901) );
  OAI211_X1 U6366 ( .C1(n4334), .C2(n6163), .A(n4903), .B(n4902), .ZN(n6365)
         );
  NAND2_X1 U6367 ( .A1(n7945), .A2(n6257), .ZN(n5459) );
  NAND2_X1 U6368 ( .A1(n6480), .A2(n6365), .ZN(n5440) );
  NAND2_X2 U6369 ( .A1(n5459), .A2(n5440), .ZN(n6478) );
  INV_X1 U6370 ( .A(n6478), .ZN(n5448) );
  NAND2_X1 U6371 ( .A1(n4904), .A2(n5448), .ZN(n6355) );
  NAND2_X1 U6372 ( .A1(n4953), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U6373 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4921) );
  OAI21_X1 U6374 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n4921), .ZN(n6483) );
  INV_X1 U6375 ( .A(n6483), .ZN(n4905) );
  NAND2_X1 U6376 ( .A1(n4252), .A2(n4905), .ZN(n4909) );
  INV_X1 U6377 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n4906) );
  OR2_X1 U6378 ( .A1(n4924), .A2(n4906), .ZN(n4908) );
  INV_X1 U6379 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6085) );
  OR2_X1 U6380 ( .A1(n5398), .A2(n6085), .ZN(n4907) );
  AND4_X2 U6381 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n6563)
         );
  OR2_X1 U6382 ( .A1(n4882), .A2(n5861), .ZN(n4917) );
  INV_X1 U6383 ( .A(n4912), .ZN(n4913) );
  INV_X1 U6384 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4914) );
  OR2_X1 U6385 ( .A1(n4932), .A2(n5069), .ZN(n4915) );
  XNOR2_X1 U6386 ( .A(n4915), .B(n4931), .ZN(n6152) );
  INV_X1 U6387 ( .A(n5577), .ZN(n4918) );
  INV_X1 U6388 ( .A(n6563), .ZN(n7944) );
  NAND2_X1 U6389 ( .A1(n4251), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4930) );
  INV_X1 U6390 ( .A(n4921), .ZN(n4920) );
  NAND2_X1 U6391 ( .A1(n4920), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n4957) );
  INV_X1 U6392 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U6393 ( .A1(n4921), .A2(n6556), .ZN(n4922) );
  AND2_X1 U6394 ( .A1(n4957), .A2(n4922), .ZN(n9833) );
  NAND2_X1 U6395 ( .A1(n4252), .A2(n9833), .ZN(n4929) );
  INV_X1 U6396 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n4925) );
  OR2_X1 U6397 ( .A1(n4924), .A2(n4925), .ZN(n4928) );
  INV_X1 U6398 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4926) );
  OR2_X1 U6399 ( .A1(n5398), .A2(n4926), .ZN(n4927) );
  INV_X1 U6400 ( .A(n6565), .ZN(n7943) );
  NAND2_X1 U6401 ( .A1(n4932), .A2(n4931), .ZN(n4989) );
  NAND2_X1 U6402 ( .A1(n4989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4941) );
  XNOR2_X1 U6403 ( .A(n4941), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6100) );
  INV_X1 U6404 ( .A(n6100), .ZN(n6141) );
  INV_X1 U6405 ( .A(n4934), .ZN(n4935) );
  INV_X1 U6406 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4936) );
  MUX2_X1 U6407 ( .A(n5866), .B(n4936), .S(n5852), .Z(n4945) );
  XNOR2_X1 U6408 ( .A(n4945), .B(SI_5_), .ZN(n4943) );
  XNOR2_X1 U6409 ( .A(n4944), .B(n4943), .ZN(n6497) );
  INV_X1 U6410 ( .A(n5575), .ZN(n5462) );
  NAND2_X1 U6411 ( .A1(n6565), .A2(n9836), .ZN(n5574) );
  NAND2_X1 U6412 ( .A1(n5409), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U6413 ( .A1(n4953), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U6414 ( .A(n4957), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U6415 ( .A1(n4252), .A2(n6530), .ZN(n4938) );
  NAND2_X1 U6416 ( .A1(n5408), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4937) );
  NAND4_X1 U6417 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n7942)
         );
  INV_X1 U6418 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6419 ( .A1(n4941), .A2(n4986), .ZN(n4942) );
  NAND2_X1 U6420 ( .A1(n4942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4965) );
  XNOR2_X1 U6421 ( .A(n4965), .B(n4987), .ZN(n6130) );
  INV_X1 U6422 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6423 ( .A1(n4946), .A2(SI_5_), .ZN(n4947) );
  MUX2_X1 U6424 ( .A(n5869), .B(n5868), .S(n5852), .Z(n4970) );
  XNOR2_X1 U6425 ( .A(n4970), .B(SI_6_), .ZN(n4968) );
  XNOR2_X1 U6426 ( .A(n4969), .B(n4968), .ZN(n6621) );
  OR2_X1 U6427 ( .A1(n5396), .A2(n5869), .ZN(n4949) );
  OAI211_X1 U6428 ( .C1(n4334), .C2(n6130), .A(n4950), .B(n4949), .ZN(n9897)
         );
  XNOR2_X1 U6429 ( .A(n7942), .B(n9897), .ZN(n6602) );
  NAND2_X1 U6430 ( .A1(n6603), .A2(n6602), .ZN(n4952) );
  INV_X1 U6431 ( .A(n7942), .ZN(n4951) );
  NAND2_X1 U6432 ( .A1(n4951), .A2(n9897), .ZN(n5465) );
  NAND2_X1 U6433 ( .A1(n4952), .A2(n5465), .ZN(n6572) );
  NAND2_X1 U6434 ( .A1(n4953), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4964) );
  INV_X1 U6435 ( .A(n4957), .ZN(n4955) );
  AND2_X1 U6436 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n4954) );
  NAND2_X1 U6437 ( .A1(n4955), .A2(n4954), .ZN(n4977) );
  INV_X1 U6438 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4956) );
  INV_X1 U6439 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6744) );
  OAI21_X1 U6440 ( .B1(n4957), .B2(n4956), .A(n6744), .ZN(n4958) );
  AND2_X1 U6441 ( .A1(n4977), .A2(n4958), .ZN(n6746) );
  NAND2_X1 U6442 ( .A1(n4252), .A2(n6746), .ZN(n4963) );
  INV_X1 U6443 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n4959) );
  OR2_X1 U6444 ( .A1(n4924), .A2(n4959), .ZN(n4962) );
  INV_X1 U6445 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4960) );
  OR2_X1 U6446 ( .A1(n5398), .A2(n4960), .ZN(n4961) );
  NAND2_X1 U6447 ( .A1(n4965), .A2(n4987), .ZN(n4966) );
  NAND2_X1 U6448 ( .A1(n4966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4967) );
  XNOR2_X1 U6449 ( .A(n4967), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6099) );
  INV_X1 U6450 ( .A(n6099), .ZN(n6175) );
  INV_X1 U6451 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6452 ( .A1(n4971), .A2(SI_6_), .ZN(n4972) );
  MUX2_X1 U6453 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5852), .Z(n4994) );
  XNOR2_X1 U6454 ( .A(n4994), .B(SI_7_), .ZN(n4992) );
  XNOR2_X1 U6455 ( .A(n4993), .B(n4992), .ZN(n6633) );
  INV_X1 U6456 ( .A(n6633), .ZN(n5873) );
  INV_X1 U6457 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5872) );
  OR2_X1 U6458 ( .A1(n5396), .A2(n5872), .ZN(n4973) );
  INV_X1 U6459 ( .A(n6763), .ZN(n6779) );
  NAND2_X1 U6460 ( .A1(n7941), .A2(n6779), .ZN(n5469) );
  NAND2_X1 U6461 ( .A1(n6572), .A2(n5469), .ZN(n4975) );
  NAND2_X1 U6462 ( .A1(n7819), .A2(n6763), .ZN(n5478) );
  NAND2_X1 U6463 ( .A1(n4975), .A2(n5478), .ZN(n6879) );
  NAND2_X1 U6464 ( .A1(n4953), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4984) );
  INV_X1 U6465 ( .A(n4977), .ZN(n4976) );
  NAND2_X1 U6466 ( .A1(n4976), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5016) );
  INV_X1 U6467 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U6468 ( .A1(n4977), .A2(n9365), .ZN(n4978) );
  AND2_X1 U6469 ( .A1(n5016), .A2(n4978), .ZN(n7824) );
  NAND2_X1 U6470 ( .A1(n4252), .A2(n7824), .ZN(n4983) );
  INV_X1 U6471 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n4979) );
  OR2_X1 U6472 ( .A1(n4924), .A2(n4979), .ZN(n4982) );
  INV_X1 U6473 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n4980) );
  OR2_X1 U6474 ( .A1(n5398), .A2(n4980), .ZN(n4981) );
  INV_X1 U6475 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4985) );
  NAND3_X1 U6476 ( .A1(n4987), .A2(n4986), .A3(n4985), .ZN(n4988) );
  NAND2_X1 U6477 ( .A1(n5012), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4991) );
  INV_X1 U6478 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4990) );
  XNOR2_X1 U6479 ( .A(n4991), .B(n4990), .ZN(n6185) );
  NAND2_X1 U6480 ( .A1(n4994), .A2(SI_7_), .ZN(n4995) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5881) );
  MUX2_X1 U6482 ( .A(n5878), .B(n5881), .S(n5852), .Z(n4998) );
  INV_X1 U6483 ( .A(SI_8_), .ZN(n4997) );
  NAND2_X1 U6484 ( .A1(n4998), .A2(n4997), .ZN(n5006) );
  INV_X1 U6485 ( .A(n4998), .ZN(n4999) );
  NAND2_X1 U6486 ( .A1(n4999), .A2(SI_8_), .ZN(n5000) );
  NAND2_X1 U6487 ( .A1(n5006), .A2(n5000), .ZN(n5004) );
  XNOR2_X1 U6488 ( .A(n5005), .B(n5004), .ZN(n6708) );
  NAND2_X1 U6489 ( .A1(n5427), .A2(n6708), .ZN(n5002) );
  OR2_X1 U6490 ( .A1(n5396), .A2(n5878), .ZN(n5001) );
  OAI211_X1 U6491 ( .C1(n4334), .C2(n6185), .A(n5002), .B(n5001), .ZN(n7823)
         );
  NAND2_X1 U6492 ( .A1(n6896), .A2(n7823), .ZN(n5470) );
  INV_X1 U6493 ( .A(n7823), .ZN(n9907) );
  NAND2_X1 U6494 ( .A1(n9907), .A2(n7940), .ZN(n5476) );
  NAND2_X1 U6495 ( .A1(n6879), .A2(n6878), .ZN(n5003) );
  NAND2_X1 U6496 ( .A1(n5003), .A2(n5470), .ZN(n6785) );
  INV_X1 U6497 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5901) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5007) );
  MUX2_X1 U6499 ( .A(n5901), .B(n5007), .S(n5852), .Z(n5009) );
  INV_X1 U6500 ( .A(SI_9_), .ZN(n5008) );
  NAND2_X1 U6501 ( .A1(n5009), .A2(n5008), .ZN(n5023) );
  INV_X1 U6502 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6503 ( .A1(n5010), .A2(SI_9_), .ZN(n5011) );
  NAND2_X1 U6504 ( .A1(n6908), .A2(n5427), .ZN(n5014) );
  NOR2_X1 U6505 ( .A1(n5012), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6506 ( .A1(n5068), .A2(n5069), .ZN(n5028) );
  XNOR2_X1 U6507 ( .A(n5028), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U6508 ( .A1(n5426), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5886), .B2(
        n6216), .ZN(n5013) );
  AND2_X2 U6509 ( .A1(n5014), .A2(n5013), .ZN(n6836) );
  NAND2_X1 U6510 ( .A1(n5409), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6511 ( .A1(n4953), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6512 ( .A1(n5016), .A2(n6894), .ZN(n5017) );
  AND2_X1 U6513 ( .A1(n5035), .A2(n5017), .ZN(n6893) );
  NAND2_X1 U6514 ( .A1(n4252), .A2(n6893), .ZN(n5019) );
  NAND2_X1 U6515 ( .A1(n5408), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5018) );
  NAND4_X1 U6516 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n7939)
         );
  NAND2_X1 U6517 ( .A1(n6836), .A2(n7939), .ZN(n5585) );
  INV_X1 U6518 ( .A(n7939), .ZN(n6846) );
  NAND2_X1 U6519 ( .A1(n6846), .A2(n7055), .ZN(n5584) );
  MUX2_X1 U6520 ( .A(n5920), .B(n5919), .S(n5852), .Z(n5025) );
  INV_X1 U6521 ( .A(SI_10_), .ZN(n5024) );
  NAND2_X1 U6522 ( .A1(n5025), .A2(n5024), .ZN(n5042) );
  INV_X1 U6523 ( .A(n5025), .ZN(n5026) );
  NAND2_X1 U6524 ( .A1(n5026), .A2(SI_10_), .ZN(n5027) );
  NAND2_X1 U6525 ( .A1(n7025), .A2(n5427), .ZN(n5033) );
  NAND2_X1 U6526 ( .A1(n5028), .A2(n5065), .ZN(n5029) );
  NAND2_X1 U6527 ( .A1(n5029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5030) );
  OR2_X1 U6528 ( .A1(n5030), .A2(n5066), .ZN(n5031) );
  NAND2_X1 U6529 ( .A1(n5030), .A2(n5066), .ZN(n5044) );
  AOI22_X1 U6530 ( .A1(n5426), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5886), .B2(
        n6316), .ZN(n5032) );
  NAND2_X2 U6531 ( .A1(n5033), .A2(n5032), .ZN(n6824) );
  NAND2_X1 U6532 ( .A1(n5409), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6533 ( .A1(n4953), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5039) );
  INV_X1 U6534 ( .A(n5035), .ZN(n5034) );
  NAND2_X1 U6535 ( .A1(n5034), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5075) );
  INV_X1 U6536 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U6537 ( .A1(n5035), .A2(n9332), .ZN(n5036) );
  AND2_X1 U6538 ( .A1(n5075), .A2(n5036), .ZN(n6849) );
  NAND2_X1 U6539 ( .A1(n4252), .A2(n6849), .ZN(n5038) );
  NAND2_X1 U6540 ( .A1(n5408), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5037) );
  NAND4_X1 U6541 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n7938)
         );
  INV_X1 U6542 ( .A(n7938), .ZN(n6997) );
  OR2_X1 U6543 ( .A1(n6824), .A2(n6997), .ZN(n5473) );
  NAND2_X1 U6544 ( .A1(n5043), .A2(n5042), .ZN(n5059) );
  MUX2_X1 U6545 ( .A(n5936), .B(n5923), .S(n5852), .Z(n5055) );
  XNOR2_X1 U6546 ( .A(n5055), .B(SI_11_), .ZN(n5054) );
  XNOR2_X1 U6547 ( .A(n5059), .B(n5054), .ZN(n7113) );
  NAND2_X1 U6548 ( .A1(n7113), .A2(n5427), .ZN(n5047) );
  NAND2_X1 U6549 ( .A1(n5044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5045) );
  XNOR2_X1 U6550 ( .A(n5045), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6458) );
  AOI22_X1 U6551 ( .A1(n5426), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5886), .B2(
        n6458), .ZN(n5046) );
  NAND2_X1 U6552 ( .A1(n4953), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6553 ( .A(n5075), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U6554 ( .A1(n4252), .A2(n7006), .ZN(n5051) );
  INV_X1 U6555 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5048) );
  OR2_X1 U6556 ( .A1(n4924), .A2(n5048), .ZN(n5050) );
  INV_X1 U6557 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6941) );
  OR2_X1 U6558 ( .A1(n5398), .A2(n6941), .ZN(n5049) );
  INV_X1 U6559 ( .A(n7086), .ZN(n5053) );
  NAND2_X1 U6560 ( .A1(n6935), .A2(n5053), .ZN(n7097) );
  INV_X1 U6561 ( .A(n5054), .ZN(n5058) );
  INV_X1 U6562 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6563 ( .A1(n5056), .A2(SI_11_), .ZN(n5057) );
  MUX2_X1 U6564 ( .A(n5981), .B(n5989), .S(n5852), .Z(n5061) );
  INV_X1 U6565 ( .A(SI_12_), .ZN(n5060) );
  NAND2_X1 U6566 ( .A1(n5061), .A2(n5060), .ZN(n5086) );
  INV_X1 U6567 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6568 ( .A1(n5062), .A2(SI_12_), .ZN(n5063) );
  NAND2_X1 U6569 ( .A1(n5086), .A2(n5063), .ZN(n5084) );
  XNOR2_X1 U6570 ( .A(n5085), .B(n5084), .ZN(n7171) );
  NAND2_X1 U6571 ( .A1(n7171), .A2(n5427), .ZN(n5072) );
  INV_X1 U6572 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5064) );
  AND3_X1 U6573 ( .A1(n5066), .A2(n5065), .A3(n5064), .ZN(n5067) );
  AND2_X1 U6574 ( .A1(n5068), .A2(n5067), .ZN(n5092) );
  OR2_X1 U6575 ( .A1(n5092), .A2(n5069), .ZN(n5070) );
  XNOR2_X1 U6576 ( .A(n5070), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6539) );
  AOI22_X1 U6577 ( .A1(n5426), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5886), .B2(
        n6539), .ZN(n5071) );
  NAND2_X1 U6578 ( .A1(n5072), .A2(n5071), .ZN(n7556) );
  NAND2_X1 U6579 ( .A1(n4953), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5082) );
  INV_X1 U6580 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7003) );
  INV_X1 U6581 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6582 ( .B1(n5075), .B2(n7003), .A(n5073), .ZN(n5076) );
  NAND2_X1 U6583 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5074) );
  AND2_X1 U6584 ( .A1(n5076), .A2(n5097), .ZN(n7549) );
  NAND2_X1 U6585 ( .A1(n4252), .A2(n7549), .ZN(n5081) );
  INV_X1 U6586 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5077) );
  OR2_X1 U6587 ( .A1(n4923), .A2(n5077), .ZN(n5080) );
  INV_X1 U6588 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5078) );
  OR2_X1 U6589 ( .A1(n5398), .A2(n5078), .ZN(n5079) );
  OR2_X1 U6590 ( .A1(n7556), .A2(n7258), .ZN(n5487) );
  NAND2_X1 U6591 ( .A1(n7556), .A2(n7258), .ZN(n5486) );
  AND2_X1 U6592 ( .A1(n7139), .A2(n7096), .ZN(n5083) );
  NAND2_X1 U6593 ( .A1(n7097), .A2(n5083), .ZN(n7098) );
  NAND2_X1 U6594 ( .A1(n7098), .A2(n5487), .ZN(n7145) );
  INV_X1 U6595 ( .A(n7145), .ZN(n5104) );
  MUX2_X1 U6596 ( .A(n6203), .B(n6194), .S(n5852), .Z(n5088) );
  NAND2_X1 U6597 ( .A1(n5088), .A2(n5087), .ZN(n5106) );
  INV_X1 U6598 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6599 ( .A1(n5089), .A2(SI_13_), .ZN(n5090) );
  XNOR2_X1 U6600 ( .A(n5105), .B(n4817), .ZN(n7347) );
  NAND2_X1 U6601 ( .A1(n7347), .A2(n5427), .ZN(n5094) );
  NAND2_X1 U6602 ( .A1(n5092), .A2(n5091), .ZN(n5156) );
  NAND2_X1 U6603 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  XNOR2_X1 U6604 ( .A(n5107), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U6605 ( .A1(n5426), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5886), .B2(
        n6670), .ZN(n5093) );
  NAND2_X1 U6606 ( .A1(n4953), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5103) );
  INV_X1 U6607 ( .A(n5097), .ZN(n5095) );
  NAND2_X1 U6608 ( .A1(n5095), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5132) );
  INV_X1 U6609 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6610 ( .A1(n5097), .A2(n5096), .ZN(n5098) );
  AND2_X1 U6611 ( .A1(n5132), .A2(n5098), .ZN(n7261) );
  NAND2_X1 U6612 ( .A1(n4252), .A2(n7261), .ZN(n5102) );
  INV_X1 U6613 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5099) );
  OR2_X1 U6614 ( .A1(n4924), .A2(n5099), .ZN(n5101) );
  INV_X1 U6615 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7154) );
  OR2_X1 U6616 ( .A1(n5398), .A2(n7154), .ZN(n5100) );
  OR2_X1 U6617 ( .A1(n8373), .A2(n7552), .ZN(n5491) );
  NAND2_X1 U6618 ( .A1(n8373), .A2(n7552), .ZN(n5490) );
  INV_X1 U6619 ( .A(n7141), .ZN(n7144) );
  MUX2_X1 U6620 ( .A(n6214), .B(n6212), .S(n5852), .Z(n5118) );
  XNOR2_X1 U6621 ( .A(n5118), .B(SI_14_), .ZN(n5117) );
  XNOR2_X1 U6622 ( .A(n5122), .B(n5117), .ZN(n7353) );
  NAND2_X1 U6623 ( .A1(n7353), .A2(n5427), .ZN(n5112) );
  INV_X1 U6624 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6625 ( .A1(n5107), .A2(n5154), .ZN(n5108) );
  NAND2_X1 U6626 ( .A1(n5108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6627 ( .A1(n5109), .A2(n5153), .ZN(n5127) );
  OR2_X1 U6628 ( .A1(n5109), .A2(n5153), .ZN(n5110) );
  AOI22_X1 U6629 ( .A1(n5426), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5886), .B2(
        n6948), .ZN(n5111) );
  NAND2_X1 U6630 ( .A1(n5409), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6631 ( .A1(n4251), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5115) );
  XNOR2_X1 U6632 ( .A(n5132), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U6633 ( .A1(n4252), .A2(n7235), .ZN(n5114) );
  NAND2_X1 U6634 ( .A1(n5408), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5113) );
  NAND4_X1 U6635 ( .A1(n5116), .A2(n5115), .A3(n5114), .A4(n5113), .ZN(n7935)
         );
  XNOR2_X1 U6636 ( .A(n7295), .B(n7935), .ZN(n7265) );
  INV_X1 U6637 ( .A(n7265), .ZN(n5495) );
  INV_X1 U6638 ( .A(n7935), .ZN(n7257) );
  OR2_X1 U6639 ( .A1(n7295), .A2(n7257), .ZN(n7270) );
  INV_X1 U6640 ( .A(n5117), .ZN(n5121) );
  INV_X1 U6641 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6642 ( .A1(n5119), .A2(SI_14_), .ZN(n5120) );
  INV_X1 U6643 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5123) );
  MUX2_X1 U6644 ( .A(n6331), .B(n5123), .S(n5852), .Z(n5124) );
  NAND2_X1 U6645 ( .A1(n5124), .A2(n9321), .ZN(n5143) );
  INV_X1 U6646 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6647 ( .A1(n5125), .A2(SI_15_), .ZN(n5126) );
  NAND2_X1 U6648 ( .A1(n5143), .A2(n5126), .ZN(n5144) );
  XNOR2_X1 U6649 ( .A(n5145), .B(n5144), .ZN(n7363) );
  NAND2_X1 U6650 ( .A1(n7363), .A2(n5427), .ZN(n5130) );
  NAND2_X1 U6651 ( .A1(n5127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  XNOR2_X1 U6652 ( .A(n5128), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7951) );
  AOI22_X1 U6653 ( .A1(n5426), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5886), .B2(
        n7951), .ZN(n5129) );
  NAND2_X1 U6654 ( .A1(n5130), .A2(n5129), .ZN(n8028) );
  NAND2_X1 U6655 ( .A1(n4251), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5139) );
  INV_X1 U6656 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5131) );
  INV_X1 U6657 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7922) );
  OAI21_X1 U6658 ( .B1(n5132), .B2(n5131), .A(n7922), .ZN(n5133) );
  AND2_X1 U6659 ( .A1(n5133), .A2(n5161), .ZN(n7928) );
  NAND2_X1 U6660 ( .A1(n4252), .A2(n7928), .ZN(n5138) );
  INV_X1 U6661 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5134) );
  OR2_X1 U6662 ( .A1(n4923), .A2(n5134), .ZN(n5137) );
  INV_X1 U6663 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5135) );
  OR2_X1 U6664 ( .A1(n5398), .A2(n5135), .ZN(n5136) );
  NAND2_X1 U6665 ( .A1(n8366), .A2(n8267), .ZN(n5140) );
  AND2_X1 U6666 ( .A1(n7270), .A2(n5140), .ZN(n5142) );
  INV_X1 U6667 ( .A(n5140), .ZN(n5141) );
  XNOR2_X1 U6668 ( .A(n8028), .B(n7851), .ZN(n7271) );
  INV_X1 U6669 ( .A(n7271), .ZN(n7268) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5147) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5146) );
  MUX2_X1 U6672 ( .A(n5147), .B(n5146), .S(n5852), .Z(n5149) );
  NAND2_X1 U6673 ( .A1(n5149), .A2(n5148), .ZN(n5172) );
  INV_X1 U6674 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6675 ( .A1(n5150), .A2(SI_16_), .ZN(n5151) );
  XNOR2_X1 U6676 ( .A(n5171), .B(n5170), .ZN(n7373) );
  NAND2_X1 U6677 ( .A1(n7373), .A2(n5427), .ZN(n5159) );
  INV_X1 U6678 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5152) );
  NAND3_X1 U6679 ( .A1(n5154), .A2(n5153), .A3(n5152), .ZN(n5155) );
  OAI21_X1 U6680 ( .B1(n5156), .B2(n5155), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5157) );
  XNOR2_X1 U6681 ( .A(n5157), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7976) );
  AOI22_X1 U6682 ( .A1(n5426), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5886), .B2(
        n7976), .ZN(n5158) );
  NAND2_X1 U6683 ( .A1(n4251), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5168) );
  INV_X1 U6684 ( .A(n5161), .ZN(n5160) );
  NAND2_X1 U6685 ( .A1(n5160), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5180) );
  INV_X1 U6686 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U6687 ( .A1(n5161), .A2(n7956), .ZN(n5162) );
  AND2_X1 U6688 ( .A1(n5180), .A2(n5162), .ZN(n8278) );
  NAND2_X1 U6689 ( .A1(n4252), .A2(n8278), .ZN(n5167) );
  INV_X1 U6690 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5163) );
  OR2_X1 U6691 ( .A1(n4924), .A2(n5163), .ZN(n5166) );
  INV_X1 U6692 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5164) );
  OR2_X1 U6693 ( .A1(n5398), .A2(n5164), .ZN(n5165) );
  NAND2_X1 U6694 ( .A1(n8360), .A2(n7275), .ZN(n5500) );
  OR2_X1 U6695 ( .A1(n8360), .A2(n7275), .ZN(n5501) );
  MUX2_X1 U6696 ( .A(n6452), .B(n6413), .S(n5852), .Z(n5187) );
  XNOR2_X1 U6697 ( .A(n5187), .B(SI_17_), .ZN(n5186) );
  XNOR2_X1 U6698 ( .A(n5191), .B(n5186), .ZN(n7340) );
  NAND2_X1 U6699 ( .A1(n7340), .A2(n5427), .ZN(n5178) );
  NAND2_X1 U6700 ( .A1(n5173), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5174) );
  MUX2_X1 U6701 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5174), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5176) );
  AND2_X1 U6702 ( .A1(n5176), .A2(n5175), .ZN(n7986) );
  AOI22_X1 U6703 ( .A1(n5426), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5886), .B2(
        n7986), .ZN(n5177) );
  NAND2_X1 U6704 ( .A1(n4953), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5185) );
  INV_X1 U6705 ( .A(n5180), .ZN(n5179) );
  NAND2_X1 U6706 ( .A1(n5179), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5196) );
  INV_X1 U6707 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U6708 ( .A1(n5180), .A2(n7974), .ZN(n5181) );
  AND2_X1 U6709 ( .A1(n5196), .A2(n5181), .ZN(n8249) );
  NAND2_X1 U6710 ( .A1(n4252), .A2(n8249), .ZN(n5184) );
  INV_X1 U6711 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9404) );
  OR2_X1 U6712 ( .A1(n4923), .A2(n9404), .ZN(n5183) );
  INV_X1 U6713 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8252) );
  OR2_X1 U6714 ( .A1(n5398), .A2(n8252), .ZN(n5182) );
  XNOR2_X1 U6715 ( .A(n8355), .B(n7934), .ZN(n8246) );
  INV_X1 U6716 ( .A(n8246), .ZN(n5503) );
  OR2_X1 U6717 ( .A1(n8355), .A2(n7934), .ZN(n5506) );
  INV_X1 U6718 ( .A(n5186), .ZN(n5190) );
  INV_X1 U6719 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6720 ( .A1(n5188), .A2(SI_17_), .ZN(n5189) );
  OAI21_X2 U6721 ( .B1(n5191), .B2(n5190), .A(n5189), .ZN(n5206) );
  MUX2_X1 U6722 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5852), .Z(n5207) );
  XNOR2_X1 U6723 ( .A(n5207), .B(SI_18_), .ZN(n5204) );
  XNOR2_X1 U6724 ( .A(n5206), .B(n5204), .ZN(n7331) );
  NAND2_X1 U6725 ( .A1(n7331), .A2(n5427), .ZN(n5194) );
  NAND2_X1 U6726 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  XNOR2_X1 U6727 ( .A(n5192), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7993) );
  AOI22_X1 U6728 ( .A1(n5426), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5886), .B2(
        n7993), .ZN(n5193) );
  NAND2_X1 U6729 ( .A1(n4251), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5202) );
  INV_X1 U6730 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6731 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  AND2_X1 U6732 ( .A1(n5234), .A2(n5197), .ZN(n8231) );
  NAND2_X1 U6733 ( .A1(n4252), .A2(n8231), .ZN(n5201) );
  INV_X1 U6734 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6735 ( .A1(n4924), .A2(n5198), .ZN(n5200) );
  INV_X1 U6736 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9412) );
  OR2_X1 U6737 ( .A1(n5398), .A2(n9412), .ZN(n5199) );
  OR2_X1 U6738 ( .A1(n8349), .A2(n8030), .ZN(n5510) );
  NAND2_X1 U6739 ( .A1(n8349), .A2(n8030), .ZN(n5516) );
  NAND2_X1 U6740 ( .A1(n5510), .A2(n5516), .ZN(n8234) );
  INV_X1 U6741 ( .A(n5204), .ZN(n5205) );
  NAND2_X1 U6742 ( .A1(n5207), .A2(SI_18_), .ZN(n5208) );
  MUX2_X1 U6743 ( .A(n6661), .B(n6663), .S(n5852), .Z(n5210) );
  INV_X1 U6744 ( .A(SI_19_), .ZN(n5209) );
  NAND2_X1 U6745 ( .A1(n5210), .A2(n5209), .ZN(n5224) );
  INV_X1 U6746 ( .A(n5210), .ZN(n5211) );
  NAND2_X1 U6747 ( .A1(n5211), .A2(SI_19_), .ZN(n5212) );
  NAND2_X1 U6748 ( .A1(n5224), .A2(n5212), .ZN(n5222) );
  XNOR2_X1 U6749 ( .A(n5223), .B(n5222), .ZN(n7383) );
  NAND2_X1 U6750 ( .A1(n7383), .A2(n5427), .ZN(n5216) );
  XNOR2_X2 U6751 ( .A(n5214), .B(n5213), .ZN(n8013) );
  AOI22_X1 U6752 ( .A1(n5426), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9838), .B2(
        n5886), .ZN(n5215) );
  NAND2_X1 U6753 ( .A1(n4251), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6754 ( .A(n5234), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U6755 ( .A1(n4252), .A2(n8219), .ZN(n5220) );
  INV_X1 U6756 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5217) );
  OR2_X1 U6757 ( .A1(n5398), .A2(n5217), .ZN(n5219) );
  INV_X1 U6758 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9430) );
  OR2_X1 U6759 ( .A1(n4923), .A2(n9430), .ZN(n5218) );
  NAND2_X1 U6760 ( .A1(n8345), .A2(n8033), .ZN(n8201) );
  MUX2_X1 U6761 ( .A(n6772), .B(n6774), .S(n5852), .Z(n5226) );
  NAND2_X1 U6762 ( .A1(n5226), .A2(n5225), .ZN(n5246) );
  INV_X1 U6763 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6764 ( .A1(n5227), .A2(SI_20_), .ZN(n5228) );
  XNOR2_X1 U6765 ( .A(n5245), .B(n5244), .ZN(n7394) );
  NAND2_X1 U6766 ( .A1(n7394), .A2(n5427), .ZN(n5230) );
  OR2_X1 U6767 ( .A1(n5396), .A2(n6772), .ZN(n5229) );
  NAND2_X1 U6768 ( .A1(n4251), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5241) );
  INV_X1 U6769 ( .A(n5234), .ZN(n5232) );
  AND2_X1 U6770 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5231) );
  NAND2_X1 U6771 ( .A1(n5232), .A2(n5231), .ZN(n5249) );
  INV_X1 U6772 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5233) );
  INV_X1 U6773 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7878) );
  OAI21_X1 U6774 ( .B1(n5234), .B2(n5233), .A(n7878), .ZN(n5235) );
  AND2_X1 U6775 ( .A1(n5249), .A2(n5235), .ZN(n8209) );
  NAND2_X1 U6776 ( .A1(n4252), .A2(n8209), .ZN(n5240) );
  INV_X1 U6777 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5236) );
  OR2_X1 U6778 ( .A1(n4924), .A2(n5236), .ZN(n5239) );
  INV_X1 U6779 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6780 ( .A1(n5398), .A2(n5237), .ZN(n5238) );
  NAND2_X1 U6781 ( .A1(n8338), .A2(n7833), .ZN(n5513) );
  INV_X1 U6782 ( .A(n8205), .ZN(n5242) );
  INV_X1 U6783 ( .A(n8201), .ZN(n5518) );
  NOR2_X1 U6784 ( .A1(n5242), .A2(n5518), .ZN(n5243) );
  MUX2_X1 U6785 ( .A(n6929), .B(n6932), .S(n5852), .Z(n5257) );
  XNOR2_X1 U6786 ( .A(n5257), .B(SI_21_), .ZN(n5256) );
  NAND2_X1 U6787 ( .A1(n7404), .A2(n5427), .ZN(n5248) );
  OR2_X1 U6788 ( .A1(n5396), .A2(n6929), .ZN(n5247) );
  NAND2_X1 U6789 ( .A1(n4953), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6790 ( .A1(n5409), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5253) );
  INV_X1 U6791 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U6792 ( .A1(n5249), .A2(n7831), .ZN(n5250) );
  AND2_X1 U6793 ( .A1(n5286), .A2(n5250), .ZN(n8192) );
  NAND2_X1 U6794 ( .A1(n4252), .A2(n8192), .ZN(n5252) );
  NAND2_X1 U6795 ( .A1(n5408), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5251) );
  NAND4_X1 U6796 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n8203)
         );
  XNOR2_X1 U6797 ( .A(n8332), .B(n8182), .ZN(n8194) );
  INV_X1 U6798 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6799 ( .A1(n5258), .A2(SI_21_), .ZN(n5259) );
  MUX2_X1 U6800 ( .A(n7051), .B(n7053), .S(n5852), .Z(n5261) );
  INV_X1 U6801 ( .A(SI_22_), .ZN(n5260) );
  NAND2_X1 U6802 ( .A1(n5261), .A2(n5260), .ZN(n5273) );
  INV_X1 U6803 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6804 ( .A1(n5262), .A2(SI_22_), .ZN(n5263) );
  NAND2_X1 U6805 ( .A1(n5273), .A2(n5263), .ZN(n5274) );
  XNOR2_X1 U6806 ( .A(n5275), .B(n5274), .ZN(n7415) );
  NAND2_X1 U6807 ( .A1(n7415), .A2(n5427), .ZN(n5265) );
  OR2_X1 U6808 ( .A1(n5396), .A2(n7051), .ZN(n5264) );
  NAND2_X1 U6809 ( .A1(n4251), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6810 ( .A(n5286), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U6811 ( .A1(n4252), .A2(n8170), .ZN(n5270) );
  INV_X1 U6812 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6813 ( .A1(n5398), .A2(n5266), .ZN(n5269) );
  INV_X1 U6814 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6815 ( .A1(n4923), .A2(n5267), .ZN(n5268) );
  NAND2_X1 U6816 ( .A1(n8327), .A2(n7890), .ZN(n5527) );
  AND2_X1 U6817 ( .A1(n8332), .A2(n8182), .ZN(n8174) );
  NOR2_X1 U6818 ( .A1(n8167), .A2(n8174), .ZN(n5272) );
  INV_X1 U6819 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7085) );
  INV_X1 U6820 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5276) );
  MUX2_X1 U6821 ( .A(n7085), .B(n5276), .S(n5852), .Z(n5278) );
  INV_X1 U6822 ( .A(SI_23_), .ZN(n5277) );
  NAND2_X1 U6823 ( .A1(n5278), .A2(n5277), .ZN(n5298) );
  INV_X1 U6824 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6825 ( .A1(n5279), .A2(SI_23_), .ZN(n5280) );
  NAND2_X1 U6826 ( .A1(n7425), .A2(n5427), .ZN(n5282) );
  OR2_X1 U6827 ( .A1(n5396), .A2(n7085), .ZN(n5281) );
  NAND2_X1 U6828 ( .A1(n4251), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5294) );
  INV_X1 U6829 ( .A(n5286), .ZN(n5284) );
  AND2_X1 U6830 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5283) );
  NAND2_X1 U6831 ( .A1(n5284), .A2(n5283), .ZN(n5300) );
  INV_X1 U6832 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7884) );
  INV_X1 U6833 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6834 ( .B1(n5286), .B2(n7884), .A(n5285), .ZN(n5287) );
  AND2_X1 U6835 ( .A1(n5300), .A2(n5287), .ZN(n8155) );
  NAND2_X1 U6836 ( .A1(n4252), .A2(n8155), .ZN(n5293) );
  INV_X1 U6837 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5289) );
  OR2_X1 U6838 ( .A1(n4923), .A2(n5289), .ZN(n5292) );
  INV_X1 U6839 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5290) );
  OR2_X1 U6840 ( .A1(n5398), .A2(n5290), .ZN(n5291) );
  OR2_X1 U6841 ( .A1(n8322), .A2(n8180), .ZN(n5529) );
  NAND2_X1 U6842 ( .A1(n8322), .A2(n8180), .ZN(n8141) );
  INV_X1 U6843 ( .A(n8151), .ZN(n8159) );
  INV_X1 U6844 ( .A(n5525), .ZN(n8160) );
  NOR2_X1 U6845 ( .A1(n8159), .A2(n8160), .ZN(n5295) );
  INV_X1 U6846 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7199) );
  MUX2_X1 U6847 ( .A(n7169), .B(n7199), .S(n5852), .Z(n5309) );
  XNOR2_X1 U6848 ( .A(n5309), .B(SI_24_), .ZN(n5308) );
  OR2_X1 U6849 ( .A1(n5396), .A2(n7169), .ZN(n5299) );
  INV_X1 U6850 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U6851 ( .A1(n5300), .A2(n9403), .ZN(n5301) );
  NAND2_X1 U6852 ( .A1(n5320), .A2(n5301), .ZN(n8135) );
  OR2_X1 U6853 ( .A1(n5357), .A2(n8135), .ZN(n5305) );
  NAND2_X1 U6854 ( .A1(n4953), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6855 ( .A1(n5408), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6856 ( .A1(n5409), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6857 ( .A1(n5306), .A2(n8038), .ZN(n5531) );
  NAND2_X1 U6858 ( .A1(n5536), .A2(n5531), .ZN(n8037) );
  INV_X1 U6859 ( .A(n8141), .ZN(n5532) );
  NOR2_X1 U6860 ( .A1(n8037), .A2(n5532), .ZN(n5307) );
  INV_X1 U6861 ( .A(n5308), .ZN(n5312) );
  INV_X1 U6862 ( .A(n5309), .ZN(n5310) );
  NAND2_X1 U6863 ( .A1(n5310), .A2(SI_24_), .ZN(n5311) );
  INV_X1 U6864 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7303) );
  MUX2_X1 U6865 ( .A(n7300), .B(n7303), .S(n5852), .Z(n5315) );
  INV_X1 U6866 ( .A(SI_25_), .ZN(n5314) );
  NAND2_X1 U6867 ( .A1(n5315), .A2(n5314), .ZN(n5325) );
  INV_X1 U6868 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6869 ( .A1(n5316), .A2(SI_25_), .ZN(n5317) );
  NAND2_X1 U6870 ( .A1(n5325), .A2(n5317), .ZN(n5326) );
  XNOR2_X1 U6871 ( .A(n5327), .B(n5326), .ZN(n7436) );
  NAND2_X1 U6872 ( .A1(n7436), .A2(n5427), .ZN(n5319) );
  OR2_X1 U6873 ( .A1(n5396), .A2(n7300), .ZN(n5318) );
  NAND2_X1 U6874 ( .A1(n5320), .A2(n9346), .ZN(n5321) );
  AND2_X1 U6875 ( .A1(n5336), .A2(n5321), .ZN(n8126) );
  NAND2_X1 U6876 ( .A1(n8126), .A2(n4252), .ZN(n5324) );
  AOI22_X1 U6877 ( .A1(n4251), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n5409), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6878 ( .A1(n5408), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6879 ( .A1(n8315), .A2(n8144), .ZN(n5544) );
  NAND2_X1 U6880 ( .A1(n5539), .A2(n5544), .ZN(n8118) );
  INV_X1 U6881 ( .A(n8118), .ZN(n8121) );
  INV_X1 U6882 ( .A(n8105), .ZN(n5342) );
  INV_X1 U6883 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7304) );
  INV_X1 U6884 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7307) );
  MUX2_X1 U6885 ( .A(n7304), .B(n7307), .S(n5852), .Z(n5329) );
  INV_X1 U6886 ( .A(SI_26_), .ZN(n5328) );
  NAND2_X1 U6887 ( .A1(n5329), .A2(n5328), .ZN(n5345) );
  INV_X1 U6888 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U6889 ( .A1(n5330), .A2(SI_26_), .ZN(n5331) );
  XNOR2_X1 U6890 ( .A(n5344), .B(n5343), .ZN(n7447) );
  NAND2_X1 U6891 ( .A1(n7447), .A2(n5427), .ZN(n5333) );
  INV_X1 U6892 ( .A(n5336), .ZN(n5334) );
  NAND2_X1 U6893 ( .A1(n5334), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5355) );
  INV_X1 U6894 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6895 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U6896 ( .A1(n5355), .A2(n5337), .ZN(n7912) );
  OR2_X1 U6897 ( .A1(n7912), .A2(n5357), .ZN(n5340) );
  AOI22_X1 U6898 ( .A1(n4251), .A2(P2_REG1_REG_26__SCAN_IN), .B1(n5409), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6899 ( .A1(n5408), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5338) );
  OR2_X1 U6900 ( .A1(n8310), .A2(n8043), .ZN(n5540) );
  NAND2_X1 U6901 ( .A1(n8310), .A2(n8043), .ZN(n5546) );
  NAND2_X1 U6902 ( .A1(n5540), .A2(n5546), .ZN(n8106) );
  NAND2_X1 U6903 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  INV_X1 U6904 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7312) );
  INV_X1 U6905 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5347) );
  MUX2_X1 U6906 ( .A(n7312), .B(n5347), .S(n5852), .Z(n5349) );
  INV_X1 U6907 ( .A(SI_27_), .ZN(n5348) );
  NAND2_X1 U6908 ( .A1(n5349), .A2(n5348), .ZN(n5363) );
  INV_X1 U6909 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6910 ( .A1(n5350), .A2(SI_27_), .ZN(n5351) );
  NAND2_X1 U6911 ( .A1(n7464), .A2(n5427), .ZN(n5353) );
  INV_X1 U6912 ( .A(n5355), .ZN(n5354) );
  NAND2_X1 U6913 ( .A1(n5354), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5367) );
  INV_X1 U6914 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U6915 ( .A1(n5355), .A2(n7770), .ZN(n5356) );
  NAND2_X1 U6916 ( .A1(n5367), .A2(n5356), .ZN(n8088) );
  OR2_X1 U6917 ( .A1(n8088), .A2(n5357), .ZN(n5360) );
  AOI22_X1 U6918 ( .A1(n4953), .A2(P2_REG1_REG_27__SCAN_IN), .B1(n5409), .B2(
        P2_REG0_REG_27__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6919 ( .A1(n5408), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6920 ( .A(n8303), .B(n8108), .ZN(n8093) );
  OR2_X1 U6921 ( .A1(n8303), .A2(n8108), .ZN(n5549) );
  INV_X1 U6922 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5364) );
  INV_X1 U6923 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8408) );
  MUX2_X1 U6924 ( .A(n5364), .B(n8408), .S(n4619), .Z(n5384) );
  XNOR2_X1 U6925 ( .A(n5384), .B(SI_28_), .ZN(n5381) );
  NAND2_X1 U6926 ( .A1(n9460), .A2(n5427), .ZN(n5366) );
  OR2_X1 U6927 ( .A1(n5396), .A2(n8408), .ZN(n5365) );
  INV_X1 U6928 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U6929 ( .A1(n5367), .A2(n7803), .ZN(n5368) );
  NAND2_X1 U6930 ( .A1(n8077), .A2(n4252), .ZN(n5374) );
  INV_X1 U6931 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6932 ( .A1(n5408), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6933 ( .A1(n5409), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5369) );
  OAI211_X1 U6934 ( .C1(n5015), .C2(n5371), .A(n5370), .B(n5369), .ZN(n5372)
         );
  INV_X1 U6935 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6936 ( .A1(n5374), .A2(n5373), .ZN(n8095) );
  NAND2_X1 U6937 ( .A1(n8298), .A2(n8095), .ZN(n5375) );
  INV_X1 U6938 ( .A(n8072), .ZN(n5376) );
  INV_X1 U6939 ( .A(n8095), .ZN(n7771) );
  NOR2_X1 U6940 ( .A1(n8298), .A2(n7771), .ZN(n5553) );
  INV_X1 U6941 ( .A(n8058), .ZN(n5377) );
  NAND2_X1 U6942 ( .A1(n5377), .A2(n4252), .ZN(n5380) );
  AOI22_X1 U6943 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(n4953), .B1(n5409), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6944 ( .A1(n5408), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6945 ( .A1(n5382), .A2(n5381), .ZN(n5386) );
  INV_X1 U6946 ( .A(SI_28_), .ZN(n5383) );
  NAND2_X1 U6947 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  INV_X1 U6948 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7535) );
  INV_X1 U6949 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8403) );
  MUX2_X1 U6950 ( .A(n7535), .B(n8403), .S(n4619), .Z(n5390) );
  XNOR2_X1 U6951 ( .A(n5390), .B(SI_29_), .ZN(n5387) );
  XNOR2_X1 U6952 ( .A(n5394), .B(n5387), .ZN(n8634) );
  NAND2_X1 U6953 ( .A1(n8634), .A2(n5427), .ZN(n5389) );
  OR2_X1 U6954 ( .A1(n5396), .A2(n8403), .ZN(n5388) );
  OR2_X1 U6955 ( .A1(n7933), .A2(n8290), .ZN(n5558) );
  NAND2_X1 U6956 ( .A1(n8290), .A2(n7933), .ZN(n5559) );
  NAND2_X1 U6957 ( .A1(n5558), .A2(n5559), .ZN(n8047) );
  INV_X1 U6958 ( .A(n8047), .ZN(n8049) );
  NAND2_X1 U6959 ( .A1(n8050), .A2(n8049), .ZN(n8052) );
  INV_X1 U6960 ( .A(n8052), .ZN(n5415) );
  INV_X1 U6961 ( .A(n5390), .ZN(n5391) );
  NOR2_X1 U6962 ( .A1(n5391), .A2(SI_29_), .ZN(n5393) );
  NAND2_X1 U6963 ( .A1(n5391), .A2(SI_29_), .ZN(n5392) );
  MUX2_X1 U6964 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4619), .Z(n5419) );
  INV_X1 U6965 ( .A(SI_30_), .ZN(n5395) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9415) );
  INV_X1 U6967 ( .A(n8023), .ZN(n9497) );
  INV_X1 U6968 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6969 ( .A1(n4953), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5400) );
  INV_X1 U6970 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6971 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  OAI211_X1 U6972 ( .C1(n4924), .C2(n5401), .A(n5400), .B(n5399), .ZN(n8020)
         );
  INV_X1 U6973 ( .A(n8020), .ZN(n5406) );
  NAND2_X1 U6974 ( .A1(n5404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6975 ( .A1(n5406), .A2(n6053), .ZN(n5407) );
  OAI21_X1 U6976 ( .B1(n9497), .B2(n5407), .A(n5559), .ZN(n5414) );
  INV_X1 U6977 ( .A(n5407), .ZN(n5413) );
  INV_X1 U6978 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6979 ( .A1(n5408), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6980 ( .A1(n5409), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5410) );
  OAI211_X1 U6981 ( .C1(n5015), .C2(n5412), .A(n5411), .B(n5410), .ZN(n8053)
         );
  NAND2_X1 U6982 ( .A1(n9497), .A2(n8053), .ZN(n5563) );
  OAI22_X1 U6983 ( .A1(n5415), .A2(n5414), .B1(n5413), .B2(n5563), .ZN(n5428)
         );
  INV_X1 U6984 ( .A(n8053), .ZN(n5416) );
  NAND2_X1 U6985 ( .A1(n8023), .A2(n5416), .ZN(n5560) );
  INV_X1 U6986 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6987 ( .A1(n5418), .A2(SI_30_), .ZN(n5422) );
  NAND2_X1 U6988 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U6989 ( .A1(n5422), .A2(n5421), .ZN(n5425) );
  MUX2_X1 U6990 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4619), .Z(n5423) );
  XNOR2_X1 U6991 ( .A(n5423), .B(SI_31_), .ZN(n5424) );
  NAND2_X1 U6992 ( .A1(n8288), .A2(n8020), .ZN(n5568) );
  NAND2_X1 U6993 ( .A1(n5560), .A2(n5568), .ZN(n5565) );
  INV_X1 U6994 ( .A(n5565), .ZN(n5596) );
  NAND2_X1 U6995 ( .A1(n5428), .A2(n5596), .ZN(n5429) );
  OR2_X1 U6996 ( .A1(n8288), .A2(n8020), .ZN(n5564) );
  INV_X1 U6997 ( .A(n5564), .ZN(n5571) );
  NAND2_X1 U6998 ( .A1(n5429), .A2(n5564), .ZN(n5430) );
  XNOR2_X1 U6999 ( .A(n5430), .B(n8013), .ZN(n5435) );
  INV_X1 U7000 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7002 ( .A1(n7050), .A2(n6928), .ZN(n6052) );
  NAND2_X1 U7003 ( .A1(n5433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5434) );
  OR2_X2 U7004 ( .A1(n6052), .A2(n6759), .ZN(n9921) );
  NAND2_X1 U7005 ( .A1(n6053), .A2(n6759), .ZN(n6337) );
  NOR2_X1 U7006 ( .A1(n5435), .A2(n4804), .ZN(n5613) );
  NOR2_X1 U7007 ( .A1(n6928), .A2(n8013), .ZN(n5436) );
  NAND2_X1 U7008 ( .A1(n7050), .A2(n5436), .ZN(n5437) );
  INV_X1 U7009 ( .A(n5540), .ZN(n5548) );
  INV_X1 U7010 ( .A(n5437), .ZN(n5535) );
  NAND2_X1 U7011 ( .A1(n5574), .A2(n5577), .ZN(n5439) );
  NAND2_X1 U7012 ( .A1(n5575), .A2(n5576), .ZN(n5438) );
  AOI21_X1 U7013 ( .B1(n5577), .B2(n5440), .A(n5458), .ZN(n5443) );
  INV_X1 U7014 ( .A(n5574), .ZN(n5442) );
  INV_X1 U7015 ( .A(n5465), .ZN(n5441) );
  NOR3_X1 U7016 ( .A1(n5443), .A2(n5442), .A3(n5441), .ZN(n5451) );
  INV_X1 U7017 ( .A(n9864), .ZN(n5444) );
  NAND2_X1 U7018 ( .A1(n5444), .A2(n7949), .ZN(n6051) );
  AOI21_X1 U7019 ( .B1(n6053), .B2(n6051), .A(n5445), .ZN(n5447) );
  NAND2_X1 U7020 ( .A1(n5578), .A2(n5454), .ZN(n5446) );
  OAI211_X1 U7021 ( .C1(n5447), .C2(n5446), .A(n6353), .B(n5437), .ZN(n5449)
         );
  NAND2_X1 U7022 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  OAI22_X1 U7023 ( .A1(n5451), .A2(n5535), .B1(n5450), .B2(n5458), .ZN(n5457)
         );
  INV_X1 U7024 ( .A(n9897), .ZN(n6609) );
  NAND2_X1 U7025 ( .A1(n6609), .A2(n7942), .ZN(n5460) );
  INV_X1 U7026 ( .A(n5578), .ZN(n5453) );
  INV_X1 U7027 ( .A(n6051), .ZN(n5452) );
  OAI211_X1 U7028 ( .C1(n5453), .C2(n5452), .A(n6353), .B(n5579), .ZN(n5455)
         );
  NAND3_X1 U7029 ( .A1(n5455), .A2(n5535), .A3(n5454), .ZN(n5456) );
  AOI21_X1 U7030 ( .B1(n5576), .B2(n5459), .A(n5458), .ZN(n5463) );
  INV_X1 U7031 ( .A(n5460), .ZN(n5461) );
  NOR3_X1 U7032 ( .A1(n5463), .A2(n5462), .A3(n5461), .ZN(n5464) );
  NAND2_X1 U7033 ( .A1(n6824), .A2(n7938), .ZN(n7090) );
  OR2_X1 U7034 ( .A1(n6824), .A2(n7938), .ZN(n5471) );
  NAND2_X1 U7035 ( .A1(n7090), .A2(n5471), .ZN(n7088) );
  MUX2_X1 U7036 ( .A(n5584), .B(n5585), .S(n5535), .Z(n5472) );
  NAND2_X1 U7037 ( .A1(n7088), .A2(n5472), .ZN(n5480) );
  INV_X1 U7038 ( .A(n5484), .ZN(n5474) );
  AOI211_X1 U7039 ( .C1(n4765), .C2(n7088), .A(n4768), .B(n5474), .ZN(n5475)
         );
  OAI21_X1 U7040 ( .B1(n5476), .B2(n5480), .A(n5475), .ZN(n5477) );
  NAND4_X1 U7041 ( .A1(n5479), .A2(n6878), .A3(n5437), .A4(n5478), .ZN(n5481)
         );
  AOI21_X1 U7042 ( .B1(n5481), .B2(n5584), .A(n5480), .ZN(n5482) );
  NAND2_X1 U7043 ( .A1(n5487), .A2(n5484), .ZN(n5485) );
  NAND2_X1 U7044 ( .A1(n5486), .A2(n7096), .ZN(n5488) );
  INV_X1 U7045 ( .A(n5490), .ZN(n5493) );
  INV_X1 U7046 ( .A(n5491), .ZN(n5492) );
  MUX2_X1 U7047 ( .A(n5493), .B(n5492), .S(n5569), .Z(n5494) );
  NAND2_X1 U7048 ( .A1(n7295), .A2(n7257), .ZN(n5496) );
  MUX2_X1 U7049 ( .A(n7270), .B(n5496), .S(n5569), .Z(n5497) );
  MUX2_X1 U7050 ( .A(n8028), .B(n8267), .S(n5569), .Z(n5498) );
  OAI21_X1 U7051 ( .B1(n8366), .B2(n7851), .A(n5498), .ZN(n5499) );
  MUX2_X1 U7052 ( .A(n5501), .B(n5500), .S(n5569), .Z(n5502) );
  NAND3_X1 U7053 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(n5509) );
  INV_X1 U7054 ( .A(n5516), .ZN(n5505) );
  AOI21_X1 U7055 ( .B1(n7934), .B2(n8355), .A(n5505), .ZN(n5507) );
  MUX2_X1 U7056 ( .A(n5507), .B(n5506), .S(n5569), .Z(n5508) );
  INV_X1 U7057 ( .A(n5511), .ZN(n5523) );
  INV_X1 U7058 ( .A(n5520), .ZN(n5512) );
  INV_X1 U7059 ( .A(n5513), .ZN(n5519) );
  NOR2_X1 U7060 ( .A1(n8332), .A2(n8182), .ZN(n5522) );
  OAI21_X1 U7061 ( .B1(n5514), .B2(n5522), .A(n5527), .ZN(n5515) );
  NAND2_X1 U7062 ( .A1(n5517), .A2(n5516), .ZN(n5521) );
  AOI211_X1 U7063 ( .C1(n5521), .C2(n5520), .A(n5519), .B(n5518), .ZN(n5524)
         );
  NOR3_X1 U7064 ( .A1(n5524), .A2(n5523), .A3(n5522), .ZN(n5526) );
  OAI21_X1 U7065 ( .B1(n5526), .B2(n8174), .A(n5525), .ZN(n5528) );
  AOI21_X1 U7066 ( .B1(n8140), .B2(n5529), .A(n5437), .ZN(n5530) );
  INV_X1 U7067 ( .A(n5531), .ZN(n5534) );
  OAI21_X1 U7068 ( .B1(n5534), .B2(n5532), .A(n5437), .ZN(n5533) );
  NAND3_X1 U7069 ( .A1(n5538), .A2(n8121), .A3(n5537), .ZN(n5543) );
  NAND2_X1 U7070 ( .A1(n5543), .A2(n5542), .ZN(n5547) );
  NAND2_X1 U7071 ( .A1(n5546), .A2(n5544), .ZN(n5545) );
  INV_X1 U7072 ( .A(n5549), .ZN(n5551) );
  INV_X1 U7073 ( .A(n8108), .ZN(n8068) );
  NAND2_X1 U7074 ( .A1(n8298), .A2(n7771), .ZN(n5554) );
  OAI21_X1 U7075 ( .B1(n8091), .B2(n8068), .A(n5554), .ZN(n5550) );
  MUX2_X1 U7076 ( .A(n5551), .B(n5550), .S(n5569), .Z(n5552) );
  INV_X1 U7077 ( .A(n8298), .ZN(n8079) );
  INV_X1 U7078 ( .A(n5554), .ZN(n5555) );
  AOI21_X1 U7079 ( .B1(n8079), .B2(n5437), .A(n5555), .ZN(n5556) );
  AOI21_X1 U7080 ( .B1(n7771), .B2(n5437), .A(n5556), .ZN(n5557) );
  INV_X1 U7081 ( .A(n5563), .ZN(n5562) );
  INV_X1 U7082 ( .A(n5560), .ZN(n5561) );
  NOR2_X1 U7083 ( .A1(n5562), .A2(n5561), .ZN(n5567) );
  NAND2_X1 U7084 ( .A1(n5564), .A2(n5563), .ZN(n5573) );
  MUX2_X1 U7085 ( .A(n5565), .B(n5573), .S(n5569), .Z(n5566) );
  INV_X1 U7086 ( .A(n5568), .ZN(n5570) );
  INV_X1 U7087 ( .A(n5573), .ZN(n5597) );
  NAND2_X1 U7088 ( .A1(n5575), .A2(n5574), .ZN(n9840) );
  NOR2_X1 U7089 ( .A1(n9840), .A2(n9825), .ZN(n5582) );
  NOR2_X1 U7090 ( .A1(n4328), .A2(n6344), .ZN(n5581) );
  AND2_X1 U7091 ( .A1(n6467), .A2(n6051), .ZN(n6343) );
  NOR2_X1 U7092 ( .A1(n6478), .A2(n6771), .ZN(n5580) );
  AND4_X1 U7093 ( .A1(n5582), .A2(n5581), .A3(n6343), .A4(n5580), .ZN(n5583)
         );
  NAND4_X1 U7094 ( .A1(n5583), .A2(n6571), .A3(n6878), .A4(n6602), .ZN(n5587)
         );
  INV_X1 U7095 ( .A(n7088), .ZN(n5586) );
  NAND2_X1 U7096 ( .A1(n5585), .A2(n5584), .ZN(n6786) );
  NOR4_X1 U7097 ( .A1(n5587), .A2(n7086), .A3(n5586), .A4(n6786), .ZN(n5588)
         );
  AND4_X1 U7098 ( .A1(n7265), .A2(n7141), .A3(n7139), .A4(n5588), .ZN(n5589)
         );
  NAND3_X1 U7099 ( .A1(n8274), .A2(n5589), .A3(n7268), .ZN(n5590) );
  NOR3_X1 U7100 ( .A1(n8234), .A2(n8246), .A3(n5590), .ZN(n5591) );
  NAND4_X1 U7101 ( .A1(n8175), .A2(n8205), .A3(n8223), .A4(n5591), .ZN(n5592)
         );
  NOR4_X1 U7102 ( .A1(n8037), .A2(n8159), .A3(n8194), .A4(n5592), .ZN(n5593)
         );
  NAND2_X1 U7103 ( .A1(n8121), .A2(n5593), .ZN(n5594) );
  NOR4_X1 U7104 ( .A1(n8072), .A2(n8093), .A3(n8106), .A4(n5594), .ZN(n5595)
         );
  NAND4_X1 U7105 ( .A1(n5597), .A2(n8049), .A3(n5596), .A4(n5595), .ZN(n5598)
         );
  XNOR2_X1 U7106 ( .A(n5598), .B(n8013), .ZN(n5599) );
  NAND2_X1 U7107 ( .A1(n6760), .A2(n9838), .ZN(n6338) );
  OAI22_X1 U7108 ( .A1(n5599), .A2(n6053), .B1(n6759), .B2(n6338), .ZN(n5600)
         );
  INV_X1 U7109 ( .A(n6338), .ZN(n5603) );
  INV_X1 U7110 ( .A(n6052), .ZN(n9865) );
  NOR3_X1 U7111 ( .A1(n5604), .A2(n5603), .A3(n9865), .ZN(n5605) );
  NAND2_X1 U7112 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  OR2_X1 U7113 ( .A1(n6250), .A2(P2_U3152), .ZN(n7083) );
  INV_X1 U7114 ( .A(n7083), .ZN(n5612) );
  NOR2_X1 U7115 ( .A1(n5614), .A2(n5069), .ZN(n5615) );
  MUX2_X1 U7116 ( .A(n5069), .B(n5615), .S(P2_IR_REG_25__SCAN_IN), .Z(n5616)
         );
  NAND2_X1 U7117 ( .A1(n5618), .A2(n5617), .ZN(n7299) );
  NAND2_X1 U7118 ( .A1(n5617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5619) );
  INV_X1 U7119 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7120 ( .A1(n6760), .A2(n6053), .ZN(n6091) );
  INV_X1 U7121 ( .A(n6091), .ZN(n6046) );
  INV_X1 U7122 ( .A(n7310), .ZN(n8019) );
  NAND4_X1 U7123 ( .A1(n6332), .A2(n8266), .A3(n8019), .A4(n6048), .ZN(n5626)
         );
  OAI211_X1 U7124 ( .C1(n6760), .C2(n7083), .A(n5626), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5627) );
  NOR2_X2 U7125 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6204) );
  NOR2_X1 U7126 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5636) );
  NOR2_X1 U7127 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5635) );
  NOR2_X1 U7128 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5634) );
  NAND4_X1 U7129 ( .A1(n5636), .A2(n5635), .A3(n5634), .A4(n5669), .ZN(n5637)
         );
  NAND2_X1 U7130 ( .A1(n5644), .A2(n5643), .ZN(n5640) );
  INV_X1 U7131 ( .A(n5768), .ZN(n5695) );
  NAND2_X1 U7132 ( .A1(n4550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7133 ( .A1(n5672), .A2(n5651), .ZN(n5654) );
  INV_X1 U7134 ( .A(n5657), .ZN(n7560) );
  AND2_X2 U7135 ( .A1(n7560), .A2(n7534), .ZN(n5781) );
  NAND2_X1 U7136 ( .A1(n5781), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5661) );
  AND2_X2 U7137 ( .A1(n7560), .A2(n5656), .ZN(n5778) );
  AND2_X2 U7138 ( .A1(n5656), .A2(n5657), .ZN(n6644) );
  NAND2_X1 U7139 ( .A1(n6644), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5659) );
  AND2_X2 U7140 ( .A1(n5657), .A2(n7534), .ZN(n5782) );
  NAND2_X1 U7141 ( .A1(n5782), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7142 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  INV_X1 U7143 ( .A(n5693), .ZN(n5774) );
  NAND2_X1 U7144 ( .A1(n5913), .A2(n5722), .ZN(n5686) );
  NAND2_X1 U7145 ( .A1(n5675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5671) );
  MUX2_X1 U7146 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5671), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5674) );
  INV_X1 U7147 ( .A(n5672), .ZN(n5673) );
  INV_X1 U7148 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9587) );
  INV_X1 U7149 ( .A(SI_0_), .ZN(n5679) );
  INV_X1 U7150 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5678) );
  OAI21_X1 U7151 ( .B1(n4619), .B2(n5679), .A(n5678), .ZN(n5681) );
  NAND2_X1 U7152 ( .A1(n5681), .A2(n5680), .ZN(n9466) );
  OAI21_X2 U7153 ( .B1(n5798), .B2(P1_IR_REG_0__SCAN_IN), .A(n5682), .ZN(n5973) );
  INV_X1 U7154 ( .A(n7649), .ZN(n5683) );
  INV_X1 U7155 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9327) );
  OAI22_X1 U7156 ( .A1(n5973), .A2(n5683), .B1(n5768), .B2(n9327), .ZN(n5684)
         );
  INV_X1 U7157 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U7158 ( .A1(n5686), .A2(n5685), .ZN(n5698) );
  NAND2_X1 U7159 ( .A1(n4299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5690) );
  MUX2_X1 U7160 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5690), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5691) );
  NAND2_X1 U7161 ( .A1(n5764), .A2(n9125), .ZN(n5773) );
  NAND2_X4 U7162 ( .A1(n5773), .A2(n5693), .ZN(n7680) );
  NAND2_X1 U7163 ( .A1(n6004), .A2(n7680), .ZN(n5699) );
  NAND2_X1 U7164 ( .A1(n8798), .A2(n5767), .ZN(n5694) );
  NAND2_X1 U7165 ( .A1(n5913), .A2(n7614), .ZN(n5697) );
  AOI22_X1 U7166 ( .A1(n9574), .A2(n5722), .B1(n5695), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5696) );
  AND2_X1 U7167 ( .A1(n5697), .A2(n5696), .ZN(n6003) );
  NAND2_X1 U7168 ( .A1(n5699), .A2(n6006), .ZN(n5714) );
  NAND2_X1 U7169 ( .A1(n6644), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7170 ( .A1(n5782), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7171 ( .A1(n6414), .A2(n5722), .ZN(n5709) );
  NAND2_X1 U7172 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5704) );
  MUX2_X1 U7173 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5704), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5707) );
  INV_X1 U7174 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7175 ( .A1(n5707), .A2(n5706), .ZN(n5863) );
  INV_X1 U7176 ( .A(n5863), .ZN(n8889) );
  NAND2_X1 U7177 ( .A1(n6076), .A2(n7674), .ZN(n5708) );
  NAND2_X1 U7178 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  NAND2_X1 U7179 ( .A1(n6414), .A2(n7614), .ZN(n5713) );
  NAND2_X1 U7180 ( .A1(n6076), .A2(n5722), .ZN(n5712) );
  NAND2_X1 U7181 ( .A1(n5713), .A2(n5712), .ZN(n6072) );
  NAND2_X1 U7182 ( .A1(n6069), .A2(n6072), .ZN(n5718) );
  INV_X1 U7183 ( .A(n5714), .ZN(n5717) );
  INV_X1 U7184 ( .A(n5715), .ZN(n5716) );
  NAND2_X1 U7185 ( .A1(n5717), .A2(n5716), .ZN(n6070) );
  NAND2_X1 U7186 ( .A1(n5718), .A2(n6070), .ZN(n6195) );
  NAND2_X1 U7187 ( .A1(n5778), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7188 ( .A1(n6644), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7189 ( .A1(n5782), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7190 ( .A1(n6075), .A2(n5722), .ZN(n5728) );
  NOR2_X1 U7191 ( .A1(n5705), .A2(n6206), .ZN(n5723) );
  MUX2_X1 U7192 ( .A(n6206), .B(n5723), .S(P1_IR_REG_2__SCAN_IN), .Z(n5726) );
  INV_X1 U7193 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U7194 ( .A1(n8642), .A2(n7649), .ZN(n5727) );
  NAND2_X1 U7195 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  XNOR2_X1 U7196 ( .A(n5732), .B(n5731), .ZN(n6196) );
  NAND2_X1 U7197 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  NAND2_X1 U7198 ( .A1(n7385), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7199 ( .A1(n5724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X1 U7200 ( .A(n5734), .B(P1_IR_REG_3__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U7201 ( .A1(n6269), .A2(n8902), .ZN(n5735) );
  NAND2_X1 U7202 ( .A1(n9693), .A2(n7674), .ZN(n5742) );
  NAND2_X1 U7203 ( .A1(n5778), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5740) );
  INV_X1 U7204 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U7205 ( .A1(n6644), .A2(n9713), .ZN(n5739) );
  NAND2_X1 U7206 ( .A1(n5781), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7207 ( .A1(n5782), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5737) );
  NAND4_X1 U7208 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n8887)
         );
  NAND2_X1 U7209 ( .A1(n8887), .A2(n5722), .ZN(n5741) );
  NAND2_X1 U7210 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  XNOR2_X1 U7211 ( .A(n5743), .B(n7680), .ZN(n6264) );
  AND2_X1 U7212 ( .A1(n9693), .A2(n5722), .ZN(n5744) );
  AOI21_X1 U7213 ( .B1(n8887), .B2(n7625), .A(n5744), .ZN(n6265) );
  XNOR2_X1 U7214 ( .A(n6264), .B(n6265), .ZN(n6267) );
  XOR2_X1 U7215 ( .A(n6267), .B(n6268), .Z(n5766) );
  NAND2_X1 U7216 ( .A1(n7301), .A2(P1_B_REG_SCAN_IN), .ZN(n5745) );
  MUX2_X1 U7217 ( .A(P1_B_REG_SCAN_IN), .B(n5745), .S(n7198), .Z(n5748) );
  INV_X1 U7218 ( .A(n5746), .ZN(n5747) );
  AND2_X1 U7219 ( .A1(n5746), .A2(n7301), .ZN(n5876) );
  NAND2_X1 U7220 ( .A1(n5746), .A2(n7198), .ZN(n5750) );
  NOR4_X1 U7221 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5760) );
  NOR4_X1 U7222 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5759) );
  NOR4_X1 U7223 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5755) );
  NOR4_X1 U7224 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5754) );
  NOR4_X1 U7225 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5753) );
  NOR4_X1 U7226 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5752) );
  NAND4_X1 U7227 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n5756)
         );
  NOR4_X1 U7228 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5757), .A4(n5756), .ZN(n5758) );
  AND3_X1 U7229 ( .A1(n5760), .A2(n5759), .A3(n5758), .ZN(n5761) );
  OR2_X1 U7230 ( .A1(n5874), .A2(n5761), .ZN(n6397) );
  INV_X1 U7231 ( .A(n5762), .ZN(n6931) );
  AND2_X1 U7232 ( .A1(n7080), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7233 ( .A1(n5764), .A2(n5762), .ZN(n6425) );
  AND3_X1 U7234 ( .A1(n9784), .A2(n5969), .A3(n6425), .ZN(n5765) );
  NOR2_X1 U7235 ( .A1(n5766), .A2(n8596), .ZN(n5795) );
  OR2_X1 U7236 ( .A1(n6425), .A2(n5767), .ZN(n5970) );
  AND3_X1 U7237 ( .A1(n5970), .A2(n5768), .A3(n7080), .ZN(n5769) );
  INV_X1 U7238 ( .A(n5789), .ZN(n5776) );
  NAND2_X1 U7239 ( .A1(n5776), .A2(n9784), .ZN(n6073) );
  NAND2_X1 U7240 ( .A1(n5769), .A2(n6073), .ZN(n5770) );
  NAND2_X1 U7241 ( .A1(n5770), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5772) );
  OR2_X1 U7242 ( .A1(n5978), .A2(n7218), .ZN(n6403) );
  NOR2_X1 U7243 ( .A1(n6403), .A2(n5790), .ZN(n5771) );
  NAND2_X1 U7244 ( .A1(n5776), .A2(n5771), .ZN(n6074) );
  MUX2_X1 U7245 ( .A(n4246), .B(n8594), .S(n9713), .Z(n5794) );
  INV_X1 U7246 ( .A(n5773), .ZN(n5775) );
  NAND2_X1 U7247 ( .A1(n6419), .A2(n5969), .ZN(n8867) );
  NOR2_X1 U7248 ( .A1(n5776), .A2(n8867), .ZN(n5787) );
  INV_X1 U7249 ( .A(n8866), .ZN(n6010) );
  AND2_X1 U7250 ( .A1(n8587), .A2(n4250), .ZN(n5793) );
  NAND2_X1 U7251 ( .A1(n5778), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5786) );
  INV_X1 U7252 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7253 ( .A1(n5779), .A2(n9713), .ZN(n5780) );
  NAND2_X1 U7254 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6281) );
  AND2_X1 U7255 ( .A1(n5780), .A2(n6281), .ZN(n6590) );
  NAND2_X1 U7256 ( .A1(n6644), .A2(n6590), .ZN(n5785) );
  NAND2_X1 U7257 ( .A1(n5781), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7258 ( .A1(n5782), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5783) );
  NAND4_X1 U7259 ( .A1(n5786), .A2(n5785), .A3(n5784), .A4(n5783), .ZN(n9701)
         );
  INV_X1 U7260 ( .A(n9701), .ZN(n9684) );
  NOR2_X1 U7261 ( .A1(n6403), .A2(n5790), .ZN(n5788) );
  NAND2_X1 U7262 ( .A1(n5789), .A2(n5788), .ZN(n5791) );
  INV_X1 U7263 ( .A(n5978), .ZN(n5975) );
  NAND2_X1 U7264 ( .A1(n9778), .A2(n9679), .ZN(n5971) );
  INV_X1 U7265 ( .A(n9693), .ZN(n9744) );
  OAI22_X1 U7266 ( .A1(n9684), .A2(n8590), .B1(n8591), .B2(n9744), .ZN(n5792)
         );
  OR4_X1 U7267 ( .A1(n5795), .A2(n5794), .A3(n5793), .A4(n5792), .ZN(P1_U3216)
         );
  INV_X1 U7268 ( .A(n7080), .ZN(n5796) );
  OR2_X1 U7269 ( .A1(n6425), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U7270 ( .A1(n5840), .A2(n5798), .ZN(n5799) );
  NAND2_X1 U7271 ( .A1(n5799), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7272 ( .A(n6251), .ZN(n5800) );
  INV_X1 U7273 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9357) );
  NOR2_X1 U7274 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9357), .ZN(n6863) );
  OR2_X1 U7275 ( .A1(n5662), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7276 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  INV_X1 U7277 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U7278 ( .A1(n5802), .A2(n9320), .ZN(n5882) );
  OR2_X1 U7279 ( .A1(n5802), .A2(n9320), .ZN(n5803) );
  NAND2_X1 U7280 ( .A1(n5882), .A2(n5803), .ZN(n5879) );
  INV_X1 U7281 ( .A(n5879), .ZN(n6707) );
  NOR2_X1 U7282 ( .A1(n6707), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7283 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U7284 ( .A(n5804), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6634) );
  INV_X1 U7285 ( .A(n6634), .ZN(n5960) );
  INV_X1 U7286 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U7287 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6634), .B1(n5960), .B2(
        n9805), .ZN(n5965) );
  OR2_X1 U7288 ( .A1(n5805), .A2(n6206), .ZN(n5806) );
  XNOR2_X1 U7289 ( .A(n5806), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6618) );
  OR2_X1 U7290 ( .A1(n5807), .A2(n6206), .ZN(n5808) );
  XNOR2_X1 U7291 ( .A(n5808), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7292 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6494), .ZN(n5809) );
  OAI21_X1 U7293 ( .B1(n6494), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5809), .ZN(
        n5928) );
  NAND2_X1 U7294 ( .A1(n5810), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5811) );
  XNOR2_X1 U7295 ( .A(n5811), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9595) );
  INV_X1 U7296 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9797) );
  XNOR2_X1 U7297 ( .A(n6013), .B(n9797), .ZN(n6019) );
  XNOR2_X1 U7298 ( .A(n5863), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n8893) );
  AND2_X1 U7299 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5812) );
  NAND2_X1 U7300 ( .A1(n8893), .A2(n5812), .ZN(n8897) );
  NAND2_X1 U7301 ( .A1(n8889), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7302 ( .A1(n8897), .A2(n5813), .ZN(n6018) );
  NAND2_X1 U7303 ( .A1(n6019), .A2(n6018), .ZN(n6017) );
  NAND2_X1 U7304 ( .A1(n6013), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7305 ( .A1(n6017), .A2(n5814), .ZN(n8908) );
  INV_X1 U7306 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U7307 ( .A(n8902), .B(n5815), .ZN(n8909) );
  AOI21_X1 U7308 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n8902), .A(n8906), .ZN(
        n9593) );
  INV_X1 U7309 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5816) );
  MUX2_X1 U7310 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5816), .S(n9595), .Z(n9592)
         );
  NAND2_X1 U7311 ( .A1(n9593), .A2(n9592), .ZN(n9591) );
  OAI21_X1 U7312 ( .B1(n9595), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9591), .ZN(
        n5929) );
  AOI21_X1 U7313 ( .B1(n6494), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5927), .ZN(
        n5904) );
  INV_X1 U7314 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9803) );
  INV_X1 U7315 ( .A(n6618), .ZN(n5867) );
  AOI22_X1 U7316 ( .A1(n6618), .A2(P1_REG1_REG_6__SCAN_IN), .B1(n9803), .B2(
        n5867), .ZN(n5903) );
  NAND2_X1 U7317 ( .A1(n5904), .A2(n5903), .ZN(n5902) );
  OAI21_X1 U7318 ( .B1(n6618), .B2(P1_REG1_REG_6__SCAN_IN), .A(n5902), .ZN(
        n5964) );
  NAND2_X1 U7319 ( .A1(n5965), .A2(n5964), .ZN(n5963) );
  OR2_X1 U7320 ( .A1(n6634), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7321 ( .A1(n5963), .A2(n5817), .ZN(n5843) );
  NOR2_X1 U7322 ( .A1(n8866), .A2(n4246), .ZN(n9461) );
  AND2_X1 U7323 ( .A1(n9461), .A2(n8964), .ZN(n5818) );
  INV_X1 U7324 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9807) );
  AOI211_X1 U7325 ( .C1(n5819), .C2(n5843), .A(n9622), .B(n9609), .ZN(n5850)
         );
  INV_X1 U7326 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7327 ( .A1(n5879), .A2(n5820), .ZN(n5833) );
  INV_X1 U7328 ( .A(n5833), .ZN(n5835) );
  NOR2_X1 U7329 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6634), .ZN(n5821) );
  AOI21_X1 U7330 ( .B1(n6634), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5821), .ZN(
        n5958) );
  NOR2_X1 U7331 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6494), .ZN(n5822) );
  AOI21_X1 U7332 ( .B1(n6494), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5822), .ZN(
        n5926) );
  INV_X1 U7333 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U7334 ( .A(n6013), .B(n6429), .ZN(n6016) );
  XNOR2_X1 U7335 ( .A(n5863), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U7336 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6008) );
  INV_X1 U7337 ( .A(n6008), .ZN(n8891) );
  NAND2_X1 U7338 ( .A1(n8892), .A2(n8891), .ZN(n8890) );
  NAND2_X1 U7339 ( .A1(n8889), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7340 ( .A1(n8890), .A2(n5823), .ZN(n6015) );
  NAND2_X1 U7341 ( .A1(n6016), .A2(n6015), .ZN(n6014) );
  NAND2_X1 U7342 ( .A1(n6013), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7343 ( .A1(n6014), .A2(n5824), .ZN(n8904) );
  NAND2_X1 U7344 ( .A1(n8902), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5826) );
  OR2_X1 U7345 ( .A1(n8902), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5825) );
  AND2_X1 U7346 ( .A1(n5826), .A2(n5825), .ZN(n8905) );
  NAND2_X1 U7347 ( .A1(n8904), .A2(n8905), .ZN(n8903) );
  NAND2_X1 U7348 ( .A1(n8903), .A2(n5826), .ZN(n9597) );
  INV_X1 U7349 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5827) );
  MUX2_X1 U7350 ( .A(n5827), .B(P1_REG2_REG_4__SCAN_IN), .S(n9595), .Z(n9596)
         );
  OR2_X1 U7351 ( .A1(n9597), .A2(n9596), .ZN(n5828) );
  OAI21_X1 U7352 ( .B1(n9595), .B2(P1_REG2_REG_4__SCAN_IN), .A(n5828), .ZN(
        n5925) );
  NAND2_X1 U7353 ( .A1(n5926), .A2(n5925), .ZN(n5924) );
  OAI21_X1 U7354 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6494), .A(n5924), .ZN(
        n5907) );
  INV_X1 U7355 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5829) );
  MUX2_X1 U7356 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n5829), .S(n6618), .Z(n5830)
         );
  INV_X1 U7357 ( .A(n5830), .ZN(n5906) );
  NOR2_X1 U7358 ( .A1(n5907), .A2(n5906), .ZN(n5905) );
  AOI21_X1 U7359 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6618), .A(n5905), .ZN(
        n5957) );
  NAND2_X1 U7360 ( .A1(n5958), .A2(n5957), .ZN(n5956) );
  OR2_X1 U7361 ( .A1(n6634), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7362 ( .A1(n5956), .A2(n5831), .ZN(n5836) );
  INV_X1 U7363 ( .A(n8964), .ZN(n9582) );
  AND2_X1 U7364 ( .A1(n9461), .A2(n9582), .ZN(n5832) );
  NAND2_X1 U7365 ( .A1(n5832), .A2(n5840), .ZN(n8956) );
  OAI21_X1 U7366 ( .B1(n5820), .B2(n5879), .A(n5836), .ZN(n5834) );
  AND2_X1 U7367 ( .A1(n5834), .A2(n5833), .ZN(n9613) );
  AOI211_X1 U7368 ( .C1(n5835), .C2(n5836), .A(n8956), .B(n9613), .ZN(n5849)
         );
  NAND2_X1 U7369 ( .A1(n9661), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5842) );
  INV_X1 U7370 ( .A(n5836), .ZN(n5838) );
  NOR2_X1 U7371 ( .A1(n8956), .A2(n5820), .ZN(n5837) );
  NAND2_X1 U7372 ( .A1(n5838), .A2(n5837), .ZN(n5841) );
  NOR2_X1 U7373 ( .A1(n8964), .A2(P1_U3084), .ZN(n7308) );
  AND2_X1 U7374 ( .A1(n7308), .A2(n8866), .ZN(n5839) );
  OAI211_X1 U7375 ( .C1(n5843), .C2(n5842), .A(n5841), .B(n9656), .ZN(n5844)
         );
  INV_X1 U7376 ( .A(n5844), .ZN(n5847) );
  INV_X1 U7377 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6980) );
  INV_X1 U7378 ( .A(n5845), .ZN(n5846) );
  OR2_X1 U7379 ( .A1(P1_U3083), .A2(n5846), .ZN(n9605) );
  OAI22_X1 U7380 ( .A1(n5847), .A2(n5879), .B1(n6980), .B2(n9605), .ZN(n5848)
         );
  OR4_X1 U7381 ( .A1(n6863), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(P1_U3249)
         );
  INV_X2 U7382 ( .A(n8398), .ZN(n8404) );
  INV_X2 U7383 ( .A(n8405), .ZN(n8400) );
  OAI222_X1 U7384 ( .A1(n8404), .A2(n5851), .B1(n8400), .B2(n5864), .C1(
        P2_U3152), .C2(n9476), .ZN(P2_U3357) );
  AOI22_X1 U7385 ( .A1(n4244), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n8902), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n5853) );
  OAI21_X1 U7386 ( .B1(n5858), .B2(n9464), .A(n5853), .ZN(P1_U3350) );
  AOI22_X1 U7387 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6013), .B1(n4244), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n5854) );
  OAI21_X1 U7388 ( .B1(n5856), .B2(n9464), .A(n5854), .ZN(P1_U3351) );
  OAI222_X1 U7389 ( .A1(n8404), .A2(n5857), .B1(n8400), .B2(n5856), .C1(
        P2_U3152), .C2(n5855), .ZN(P2_U3356) );
  OAI222_X1 U7390 ( .A1(n8404), .A2(n5859), .B1(n8400), .B2(n5858), .C1(
        P2_U3152), .C2(n6163), .ZN(P2_U3355) );
  AOI22_X1 U7391 ( .A1(n9595), .A2(P1_STATE_REG_SCAN_IN), .B1(n4244), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U7392 ( .B1(n6272), .B2(n9464), .A(n5860), .ZN(P1_U3349) );
  OAI222_X1 U7393 ( .A1(n8404), .A2(n5861), .B1(n8400), .B2(n6272), .C1(
        P2_U3152), .C2(n6152), .ZN(P2_U3354) );
  AOI22_X1 U7394 ( .A1(n6494), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n4244), .ZN(n5862) );
  OAI21_X1 U7395 ( .B1(n6497), .B2(n9464), .A(n5862), .ZN(P1_U3348) );
  INV_X1 U7396 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5865) );
  OAI222_X1 U7397 ( .A1(n9462), .A2(n5865), .B1(n9464), .B2(n5864), .C1(n4246), 
        .C2(n5863), .ZN(P1_U3352) );
  OAI222_X1 U7398 ( .A1(n8404), .A2(n5866), .B1(n8400), .B2(n6497), .C1(
        P2_U3152), .C2(n6141), .ZN(P2_U3353) );
  OAI222_X1 U7399 ( .A1(n9462), .A2(n5868), .B1(n9464), .B2(n6621), .C1(n4246), 
        .C2(n5867), .ZN(P1_U3347) );
  OAI222_X1 U7400 ( .A1(n8404), .A2(n5869), .B1(n8400), .B2(n6621), .C1(
        P2_U3152), .C2(n6130), .ZN(P2_U3352) );
  INV_X1 U7401 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7402 ( .A1(n7223), .A2(n5969), .ZN(n5870) );
  OAI21_X1 U7403 ( .B1(n5969), .B2(n5871), .A(n5870), .ZN(P1_U3440) );
  OAI222_X1 U7404 ( .A1(n8404), .A2(n5872), .B1(n8400), .B2(n5873), .C1(
        P2_U3152), .C2(n6175), .ZN(P2_U3351) );
  INV_X1 U7405 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6637) );
  OAI222_X1 U7406 ( .A1(n9462), .A2(n6637), .B1(n9464), .B2(n5873), .C1(
        P1_U3084), .C2(n5960), .ZN(P1_U3346) );
  AND2_X1 U7407 ( .A1(n9725), .A2(n5875), .ZN(n5877) );
  OAI22_X1 U7408 ( .A1(n5877), .A2(n5876), .B1(n5969), .B2(n5875), .ZN(
        P1_U3441) );
  INV_X1 U7409 ( .A(n6708), .ZN(n5880) );
  OAI222_X1 U7410 ( .A1(n8404), .A2(n5878), .B1(n8400), .B2(n5880), .C1(
        P2_U3152), .C2(n6185), .ZN(P2_U3350) );
  OAI222_X1 U7411 ( .A1(n9462), .A2(n5881), .B1(n9464), .B2(n5880), .C1(
        P1_U3084), .C2(n5879), .ZN(P1_U3345) );
  INV_X1 U7412 ( .A(n6908), .ZN(n5900) );
  NAND2_X1 U7413 ( .A1(n5882), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7414 ( .A(n5883), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9606) );
  AOI22_X1 U7415 ( .A1(n9606), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n4244), .ZN(n5884) );
  OAI21_X1 U7416 ( .B1(n5900), .B2(n9464), .A(n5884), .ZN(P1_U3344) );
  NAND2_X1 U7417 ( .A1(n9850), .A2(n7083), .ZN(n5885) );
  NAND2_X1 U7418 ( .A1(n5886), .A2(n5885), .ZN(n5888) );
  NAND2_X1 U7419 ( .A1(n6332), .A2(n6046), .ZN(n5887) );
  AND2_X1 U7420 ( .A1(n5888), .A2(n5887), .ZN(n9472) );
  NOR2_X1 U7421 ( .A1(n9820), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7422 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7423 ( .A1(n8020), .A2(P2_U3966), .ZN(n5889) );
  OAI21_X1 U7424 ( .B1(n5890), .B2(P2_U3966), .A(n5889), .ZN(P2_U3583) );
  INV_X2 U7425 ( .A(n5891), .ZN(n7471) );
  NAND2_X1 U7426 ( .A1(n7471), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7427 ( .A1(n8455), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7428 ( .A1(n8456), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7429 ( .A1(n8888), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U7430 ( .B1(n8988), .B2(n8888), .A(n5895), .ZN(P1_U3585) );
  NAND2_X1 U7431 ( .A1(n7471), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7432 ( .A1(n8455), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7433 ( .A1(n8456), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7434 ( .A1(n8888), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5899) );
  OAI21_X1 U7435 ( .B1(n8966), .B2(n8888), .A(n5899), .ZN(P1_U3586) );
  INV_X1 U7436 ( .A(n6216), .ZN(n6221) );
  OAI222_X1 U7437 ( .A1(n8404), .A2(n5901), .B1(n8400), .B2(n5900), .C1(n6221), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7438 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U7439 ( .B1(n5904), .B2(n5903), .A(n5902), .ZN(n5909) );
  AOI211_X1 U7440 ( .C1(n5907), .C2(n5906), .A(n5905), .B(n8956), .ZN(n5908)
         );
  AOI21_X1 U7441 ( .B1(n9661), .B2(n5909), .A(n5908), .ZN(n5911) );
  AND2_X1 U7442 ( .A1(n4246), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8566) );
  AOI21_X1 U7443 ( .B1(n9634), .B2(n6618), .A(n8566), .ZN(n5910) );
  OAI211_X1 U7444 ( .C1(n9605), .C2(n5912), .A(n5911), .B(n5910), .ZN(P1_U3247) );
  INV_X1 U7445 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U7446 ( .A1(n5913), .A2(P1_U4006), .ZN(n5914) );
  OAI21_X1 U7447 ( .B1(P1_U4006), .B2(n9348), .A(n5914), .ZN(P1_U3555) );
  INV_X1 U7448 ( .A(n7025), .ZN(n5921) );
  NAND2_X1 U7449 ( .A1(n5916), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5915) );
  MUX2_X1 U7450 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5915), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5918) );
  NOR2_X1 U7451 ( .A1(n5916), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5983) );
  INV_X1 U7452 ( .A(n5983), .ZN(n5917) );
  NAND2_X1 U7453 ( .A1(n5918), .A2(n5917), .ZN(n5942) );
  OAI222_X1 U7454 ( .A1(n9464), .A2(n5921), .B1(n5942), .B2(P1_U3084), .C1(
        n5919), .C2(n9462), .ZN(P1_U3343) );
  INV_X1 U7455 ( .A(n6316), .ZN(n6321) );
  OAI222_X1 U7456 ( .A1(P2_U3152), .A2(n6321), .B1(n8400), .B2(n5921), .C1(
        n5920), .C2(n8404), .ZN(P2_U3348) );
  INV_X1 U7457 ( .A(n7113), .ZN(n5935) );
  OR2_X1 U7458 ( .A1(n5983), .A2(n6206), .ZN(n5922) );
  XNOR2_X1 U7459 ( .A(n5922), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7114) );
  INV_X1 U7460 ( .A(n7114), .ZN(n5991) );
  OAI222_X1 U7461 ( .A1(n9464), .A2(n5935), .B1(n5991), .B2(n4246), .C1(n5923), 
        .C2(n9462), .ZN(P1_U3342) );
  INV_X1 U7462 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5934) );
  OAI21_X1 U7463 ( .B1(n5926), .B2(n5925), .A(n5924), .ZN(n5931) );
  AOI211_X1 U7464 ( .C1(n5929), .C2(n5928), .A(n5927), .B(n9622), .ZN(n5930)
         );
  AOI21_X1 U7465 ( .B1(n9665), .B2(n5931), .A(n5930), .ZN(n5933) );
  AND2_X1 U7466 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6510) );
  AOI21_X1 U7467 ( .B1(n9634), .B2(n6494), .A(n6510), .ZN(n5932) );
  OAI211_X1 U7468 ( .C1(n9605), .C2(n5934), .A(n5933), .B(n5932), .ZN(P1_U3246) );
  INV_X1 U7469 ( .A(n6458), .ZN(n6454) );
  OAI222_X1 U7470 ( .A1(n8404), .A2(n5936), .B1(n8400), .B2(n5935), .C1(n6454), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7471 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5939) );
  NOR2_X1 U7472 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9606), .ZN(n5938) );
  INV_X1 U7473 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5937) );
  MUX2_X1 U7474 ( .A(n5937), .B(P1_REG1_REG_9__SCAN_IN), .S(n9606), .Z(n9608)
         );
  NOR2_X1 U7475 ( .A1(n9609), .A2(n9608), .ZN(n9607) );
  NOR2_X1 U7476 ( .A1(n5938), .A2(n9607), .ZN(n9621) );
  MUX2_X1 U7477 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n5939), .S(n5942), .Z(n9620)
         );
  NOR2_X1 U7478 ( .A1(n9621), .A2(n9620), .ZN(n9619) );
  INV_X1 U7479 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U7480 ( .A1(n7114), .A2(n9566), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n5991), .ZN(n5940) );
  NOR2_X1 U7481 ( .A1(n5941), .A2(n5940), .ZN(n5990) );
  AOI21_X1 U7482 ( .B1(n5941), .B2(n5940), .A(n5990), .ZN(n5955) );
  INV_X1 U7483 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9431) );
  AOI22_X1 U7484 ( .A1(n7114), .A2(n9431), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n5991), .ZN(n5948) );
  INV_X1 U7485 ( .A(n5942), .ZN(n9618) );
  NAND2_X1 U7486 ( .A1(n9618), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5946) );
  INV_X1 U7487 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5943) );
  MUX2_X1 U7488 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n5943), .S(n5942), .Z(n5944)
         );
  INV_X1 U7489 ( .A(n5944), .ZN(n9625) );
  INV_X1 U7490 ( .A(n9606), .ZN(n5945) );
  INV_X1 U7491 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9307) );
  MUX2_X1 U7492 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9307), .S(n9606), .Z(n9612)
         );
  NAND2_X1 U7493 ( .A1(n9612), .A2(n9613), .ZN(n9611) );
  OAI21_X1 U7494 ( .B1(n5945), .B2(n9307), .A(n9611), .ZN(n9626) );
  NAND2_X1 U7495 ( .A1(n9625), .A2(n9626), .ZN(n9624) );
  NAND2_X1 U7496 ( .A1(n5946), .A2(n9624), .ZN(n5947) );
  NOR2_X1 U7497 ( .A1(n5948), .A2(n5947), .ZN(n5996) );
  AOI21_X1 U7498 ( .B1(n5948), .B2(n5947), .A(n5996), .ZN(n5949) );
  INV_X1 U7499 ( .A(n5949), .ZN(n5953) );
  INV_X1 U7500 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n5951) );
  AND2_X1 U7501 ( .A1(n4246), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7132) );
  AOI21_X1 U7502 ( .B1(n9634), .B2(n7114), .A(n7132), .ZN(n5950) );
  OAI21_X1 U7503 ( .B1(n9605), .B2(n5951), .A(n5950), .ZN(n5952) );
  AOI21_X1 U7504 ( .B1(n5953), .B2(n9665), .A(n5952), .ZN(n5954) );
  OAI21_X1 U7505 ( .B1(n5955), .B2(n9622), .A(n5954), .ZN(P1_U3252) );
  OAI21_X1 U7506 ( .B1(n5958), .B2(n5957), .A(n5956), .ZN(n5962) );
  NAND2_X1 U7507 ( .A1(n9659), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7508 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6700) );
  OAI211_X1 U7509 ( .C1(n9656), .C2(n5960), .A(n5959), .B(n6700), .ZN(n5961)
         );
  AOI21_X1 U7510 ( .B1(n9665), .B2(n5962), .A(n5961), .ZN(n5968) );
  OAI21_X1 U7511 ( .B1(n5965), .B2(n5964), .A(n5963), .ZN(n5966) );
  NAND2_X1 U7512 ( .A1(n5966), .A2(n9661), .ZN(n5967) );
  NAND2_X1 U7513 ( .A1(n5968), .A2(n5967), .ZN(P1_U3248) );
  NAND3_X1 U7514 ( .A1(n5971), .A2(n6398), .A3(n6397), .ZN(n5972) );
  INV_X1 U7515 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5980) );
  INV_X1 U7516 ( .A(n5913), .ZN(n5974) );
  AOI21_X1 U7517 ( .B1(n5974), .B2(n5973), .A(n6437), .ZN(n8806) );
  NOR2_X1 U7518 ( .A1(n6419), .A2(n5975), .ZN(n5977) );
  INV_X1 U7519 ( .A(n6425), .ZN(n5976) );
  AOI22_X1 U7520 ( .A1(n8806), .A2(n5977), .B1(n9702), .B2(n6414), .ZN(n6406)
         );
  OAI21_X1 U7521 ( .B1(n5973), .B2(n5978), .A(n6406), .ZN(n9290) );
  NAND2_X1 U7522 ( .A1(n9290), .A2(n9794), .ZN(n5979) );
  OAI21_X1 U7523 ( .B1(n9794), .B2(n5980), .A(n5979), .ZN(P1_U3454) );
  INV_X1 U7524 ( .A(n7171), .ZN(n5988) );
  INV_X1 U7525 ( .A(n6539), .ZN(n6544) );
  OAI222_X1 U7526 ( .A1(n8404), .A2(n5981), .B1(n8400), .B2(n5988), .C1(
        P2_U3152), .C2(n6544), .ZN(P2_U3346) );
  INV_X1 U7527 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5982) );
  INV_X1 U7528 ( .A(n5986), .ZN(n5984) );
  NAND2_X1 U7529 ( .A1(n5984), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5987) );
  INV_X1 U7530 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7531 ( .A1(n5986), .A2(n5985), .ZN(n6192) );
  INV_X1 U7532 ( .A(n7172), .ZN(n6230) );
  OAI222_X1 U7533 ( .A1(n9462), .A2(n5989), .B1(n9464), .B2(n5988), .C1(n4246), 
        .C2(n6230), .ZN(P1_U3341) );
  AOI21_X1 U7534 ( .B1(n5991), .B2(n9566), .A(n5990), .ZN(n5993) );
  INV_X1 U7535 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U7536 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6230), .B1(n7172), .B2(
        n9560), .ZN(n5992) );
  NOR2_X1 U7537 ( .A1(n5993), .A2(n5992), .ZN(n6229) );
  AOI21_X1 U7538 ( .B1(n5993), .B2(n5992), .A(n6229), .ZN(n6002) );
  INV_X1 U7539 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7125) );
  NOR2_X1 U7540 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7125), .ZN(n7211) );
  NOR2_X1 U7541 ( .A1(n9656), .A2(n6230), .ZN(n5994) );
  AOI211_X1 U7542 ( .C1(n9659), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7211), .B(
        n5994), .ZN(n6001) );
  NOR2_X1 U7543 ( .A1(n7114), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5995) );
  NOR2_X1 U7544 ( .A1(n5996), .A2(n5995), .ZN(n5999) );
  INV_X1 U7545 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5997) );
  MUX2_X1 U7546 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n5997), .S(n7172), .Z(n5998)
         );
  NAND2_X1 U7547 ( .A1(n5998), .A2(n5999), .ZN(n6234) );
  OAI211_X1 U7548 ( .C1(n5999), .C2(n5998), .A(n9665), .B(n6234), .ZN(n6000)
         );
  OAI211_X1 U7549 ( .C1(n6002), .C2(n9622), .A(n6001), .B(n6000), .ZN(P1_U3253) );
  INV_X1 U7550 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6964) );
  INV_X1 U7551 ( .A(n6003), .ZN(n6005) );
  NAND2_X1 U7552 ( .A1(n6005), .A2(n6004), .ZN(n6007) );
  NAND2_X1 U7553 ( .A1(n6007), .A2(n6006), .ZN(n9577) );
  MUX2_X1 U7554 ( .A(n9577), .B(n6008), .S(n9582), .Z(n6012) );
  INV_X1 U7555 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U7556 ( .A1(n9582), .A2(n6401), .ZN(n6009) );
  NAND2_X1 U7557 ( .A1(n6010), .A2(n6009), .ZN(n9581) );
  AND2_X1 U7558 ( .A1(n9581), .A2(n9587), .ZN(n9583) );
  NOR2_X1 U7559 ( .A1(n9583), .A2(n8888), .ZN(n6011) );
  OAI21_X1 U7560 ( .B1(n6012), .B2(n8866), .A(n6011), .ZN(n9601) );
  AOI22_X1 U7561 ( .A1(n9634), .A2(n6013), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6022) );
  OAI211_X1 U7562 ( .C1(n6016), .C2(n6015), .A(n9665), .B(n6014), .ZN(n6021)
         );
  OAI211_X1 U7563 ( .C1(n6019), .C2(n6018), .A(n9661), .B(n6017), .ZN(n6020)
         );
  AND3_X1 U7564 ( .A1(n6022), .A2(n6021), .A3(n6020), .ZN(n6023) );
  OAI211_X1 U7565 ( .C1(n6964), .C2(n9605), .A(n9601), .B(n6023), .ZN(P1_U3243) );
  INV_X1 U7566 ( .A(n7305), .ZN(n6027) );
  XOR2_X1 U7567 ( .A(n7170), .B(n6024), .Z(n6025) );
  NAND2_X1 U7568 ( .A1(n7299), .A2(n6025), .ZN(n6026) );
  INV_X1 U7569 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9861) );
  AND2_X1 U7570 ( .A1(n7299), .A2(n7305), .ZN(n9862) );
  AOI21_X1 U7571 ( .B1(n9849), .B2(n9861), .A(n9862), .ZN(n6757) );
  NOR4_X1 U7572 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6031) );
  NOR4_X1 U7573 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6030) );
  NOR4_X1 U7574 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6029) );
  NOR4_X1 U7575 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6028) );
  NAND4_X1 U7576 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n6037)
         );
  NOR2_X1 U7577 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n6035) );
  NOR4_X1 U7578 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6034) );
  NOR4_X1 U7579 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6033) );
  NOR4_X1 U7580 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7581 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6036)
         );
  OAI21_X1 U7582 ( .B1(n6037), .B2(n6036), .A(n9849), .ZN(n6755) );
  AND2_X1 U7583 ( .A1(n6757), .A2(n6755), .ZN(n6334) );
  AND2_X1 U7584 ( .A1(n7170), .A2(n7305), .ZN(n9859) );
  INV_X1 U7585 ( .A(n9859), .ZN(n6039) );
  NAND2_X1 U7586 ( .A1(n9849), .A2(n9858), .ZN(n6038) );
  INV_X1 U7587 ( .A(n6767), .ZN(n6758) );
  NAND2_X1 U7588 ( .A1(n6334), .A2(n6758), .ZN(n6047) );
  INV_X1 U7589 ( .A(n6048), .ZN(n6040) );
  NOR2_X1 U7590 ( .A1(n9898), .A2(n6046), .ZN(n6041) );
  NAND2_X1 U7591 ( .A1(n7919), .A2(n7798), .ZN(n7898) );
  AOI21_X1 U7592 ( .B1(n7949), .B2(n7798), .A(n7909), .ZN(n6044) );
  NOR2_X1 U7593 ( .A1(n6052), .A2(n6771), .ZN(n9835) );
  NAND2_X1 U7594 ( .A1(n6045), .A2(n9835), .ZN(n6043) );
  INV_X1 U7595 ( .A(n6752), .ZN(n6042) );
  OAI21_X1 U7596 ( .B1(n6044), .B2(n7889), .A(n9864), .ZN(n6050) );
  NAND2_X1 U7597 ( .A1(n6045), .A2(n6048), .ZN(n7924) );
  NAND2_X1 U7598 ( .A1(n5624), .A2(n6046), .ZN(n8179) );
  INV_X1 U7599 ( .A(n7904), .ZN(n7913) );
  NAND2_X1 U7600 ( .A1(n6047), .A2(n6752), .ZN(n6253) );
  NAND3_X1 U7601 ( .A1(n6253), .A2(n6332), .A3(n6751), .ZN(n7539) );
  AOI22_X1 U7602 ( .A1(n7913), .A2(n7947), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7539), .ZN(n6049) );
  OAI211_X1 U7603 ( .C1(n6051), .C2(n7898), .A(n6050), .B(n6049), .ZN(P2_U3234) );
  NAND3_X1 U7604 ( .A1(n6338), .A2(n6052), .A3(n6928), .ZN(n6054) );
  NAND2_X1 U7605 ( .A1(n6053), .A2(n6771), .ZN(n6336) );
  AND2_X2 U7606 ( .A1(n6054), .A2(n6336), .ZN(n7749) );
  INV_X1 U7607 ( .A(n6058), .ZN(n6057) );
  NAND2_X1 U7608 ( .A1(n6055), .A2(n7798), .ZN(n6059) );
  INV_X1 U7609 ( .A(n6059), .ZN(n6056) );
  NAND2_X1 U7610 ( .A1(n6057), .A2(n6056), .ZN(n6060) );
  NAND2_X1 U7611 ( .A1(n6059), .A2(n6058), .ZN(n6243) );
  NAND2_X1 U7612 ( .A1(n6060), .A2(n6243), .ZN(n6065) );
  NAND2_X1 U7613 ( .A1(n7949), .A2(n9864), .ZN(n6469) );
  INV_X1 U7614 ( .A(n6065), .ZN(n6062) );
  NAND2_X1 U7615 ( .A1(n6062), .A2(n6061), .ZN(n6244) );
  INV_X1 U7616 ( .A(n6244), .ZN(n6063) );
  AOI21_X1 U7617 ( .B1(n6065), .B2(n6064), .A(n6063), .ZN(n6068) );
  INV_X1 U7618 ( .A(n7903), .ZN(n7914) );
  AOI22_X1 U7619 ( .A1(n7914), .A2(n7949), .B1(n7913), .B2(n7946), .ZN(n6067)
         );
  AOI22_X1 U7620 ( .A1(n7889), .A2(n6470), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7539), .ZN(n6066) );
  OAI211_X1 U7621 ( .C1(n6068), .C2(n7909), .A(n6067), .B(n6066), .ZN(P2_U3224) );
  NAND2_X1 U7622 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  XOR2_X1 U7623 ( .A(n6072), .B(n6071), .Z(n6080) );
  AND3_X1 U7624 ( .A1(n6074), .A2(n6073), .A3(n6398), .ZN(n9580) );
  INV_X1 U7625 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6447) );
  NOR2_X1 U7626 ( .A1(n9580), .A2(n6447), .ZN(n6078) );
  OAI22_X1 U7627 ( .A1(n8643), .A2(n8590), .B1(n8591), .B2(n9732), .ZN(n6077)
         );
  AOI211_X1 U7628 ( .C1(n8587), .C2(n5913), .A(n6078), .B(n6077), .ZN(n6079)
         );
  OAI21_X1 U7629 ( .B1(n6080), .B2(n8596), .A(n6079), .ZN(P1_U3220) );
  INV_X1 U7630 ( .A(n6130), .ZN(n6088) );
  INV_X1 U7631 ( .A(n6152), .ZN(n6086) );
  INV_X1 U7632 ( .A(n9476), .ZN(n6105) );
  INV_X1 U7633 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U7634 ( .A1(n9476), .A2(n6081), .ZN(n6083) );
  NAND2_X1 U7635 ( .A1(n6105), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7636 ( .A1(n6083), .A2(n6082), .ZN(n9470) );
  NOR3_X1 U7637 ( .A1(n9823), .A2(n9813), .A3(n9470), .ZN(n9468) );
  AOI21_X1 U7638 ( .B1(n6105), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9468), .ZN(
        n9486) );
  XNOR2_X1 U7639 ( .A(n9488), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9485) );
  NOR2_X1 U7640 ( .A1(n9486), .A2(n9485), .ZN(n9484) );
  AOI21_X1 U7641 ( .B1(n9488), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9484), .ZN(
        n6157) );
  NAND2_X1 U7642 ( .A1(n6102), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7643 ( .B1(n6102), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6084), .ZN(
        n6156) );
  MUX2_X1 U7644 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6085), .S(n6152), .Z(n6145)
         );
  NAND2_X1 U7645 ( .A1(n6100), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7646 ( .B1(n6100), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6087), .ZN(
        n6134) );
  NOR2_X1 U7647 ( .A1(n4281), .A2(n6134), .ZN(n6133) );
  INV_X1 U7648 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6605) );
  MUX2_X1 U7649 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6605), .S(n6130), .Z(n6122)
         );
  NAND2_X1 U7650 ( .A1(n6099), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7651 ( .B1(n6099), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6089), .ZN(
        n6167) );
  AOI21_X1 U7652 ( .B1(n6099), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6166), .ZN(
        n6096) );
  MUX2_X1 U7653 ( .A(n4980), .B(P2_REG2_REG_8__SCAN_IN), .S(n6185), .Z(n6090)
         );
  INV_X1 U7654 ( .A(n6090), .ZN(n6095) );
  NOR2_X1 U7655 ( .A1(n6096), .A2(n6095), .ZN(n6178) );
  OR2_X1 U7656 ( .A1(n5624), .A2(P2_U3152), .ZN(n8406) );
  NAND2_X1 U7657 ( .A1(n6332), .A2(n6091), .ZN(n6092) );
  OAI211_X1 U7658 ( .C1(n6251), .C2(n8406), .A(n6092), .B(n7083), .ZN(n6114)
         );
  NAND2_X1 U7659 ( .A1(n6114), .A2(n4334), .ZN(n6093) );
  NAND2_X1 U7660 ( .A1(n6093), .A2(n7948), .ZN(n6097) );
  NOR2_X1 U7661 ( .A1(n5624), .A2(n7310), .ZN(n6094) );
  AOI211_X1 U7662 ( .C1(n6096), .C2(n6095), .A(n6178), .B(n9483), .ZN(n6120)
         );
  NAND2_X1 U7663 ( .A1(n6097), .A2(n5624), .ZN(n9815) );
  NOR2_X1 U7664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9365), .ZN(n6098) );
  AOI21_X1 U7665 ( .B1(n9820), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6098), .ZN(
        n6118) );
  INV_X1 U7666 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9351) );
  MUX2_X1 U7667 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9351), .S(n6099), .Z(n6171)
         );
  INV_X1 U7668 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9936) );
  MUX2_X1 U7669 ( .A(n9936), .B(P2_REG1_REG_6__SCAN_IN), .S(n6130), .Z(n6126)
         );
  NAND2_X1 U7670 ( .A1(n6100), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6110) );
  INV_X1 U7671 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6101) );
  MUX2_X1 U7672 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6101), .S(n6100), .Z(n6137)
         );
  INV_X1 U7673 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U7674 ( .A(n9933), .B(P2_REG1_REG_4__SCAN_IN), .S(n6152), .Z(n6148)
         );
  NAND2_X1 U7675 ( .A1(n6102), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6109) );
  INV_X1 U7676 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U7677 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6103), .S(n6102), .Z(n6159)
         );
  NAND2_X1 U7678 ( .A1(n9488), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6108) );
  INV_X1 U7679 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6104) );
  MUX2_X1 U7680 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6104), .S(n9488), .Z(n9491)
         );
  NAND2_X1 U7681 ( .A1(n6105), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6107) );
  INV_X1 U7682 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6106) );
  MUX2_X1 U7683 ( .A(n6106), .B(P2_REG1_REG_1__SCAN_IN), .S(n9476), .Z(n9479)
         );
  NAND3_X1 U7684 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9479), .ZN(n9478) );
  NAND2_X1 U7685 ( .A1(n6107), .A2(n9478), .ZN(n9492) );
  NAND2_X1 U7686 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  NAND2_X1 U7687 ( .A1(n6108), .A2(n9490), .ZN(n6160) );
  NAND2_X1 U7688 ( .A1(n6159), .A2(n6160), .ZN(n6158) );
  NAND2_X1 U7689 ( .A1(n6109), .A2(n6158), .ZN(n6149) );
  NAND2_X1 U7690 ( .A1(n6148), .A2(n6149), .ZN(n6147) );
  OAI21_X1 U7691 ( .B1(n6152), .B2(n9933), .A(n6147), .ZN(n6138) );
  NAND2_X1 U7692 ( .A1(n6137), .A2(n6138), .ZN(n6136) );
  NAND2_X1 U7693 ( .A1(n6110), .A2(n6136), .ZN(n6127) );
  NAND2_X1 U7694 ( .A1(n6126), .A2(n6127), .ZN(n6125) );
  OAI21_X1 U7695 ( .B1(n6130), .B2(n9936), .A(n6125), .ZN(n6172) );
  NAND2_X1 U7696 ( .A1(n6171), .A2(n6172), .ZN(n6170) );
  OAI21_X1 U7697 ( .B1(n6175), .B2(n9351), .A(n6170), .ZN(n6116) );
  INV_X1 U7698 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6111) );
  MUX2_X1 U7699 ( .A(n6111), .B(P2_REG1_REG_8__SCAN_IN), .S(n6185), .Z(n6115)
         );
  AND2_X1 U7700 ( .A1(n4334), .A2(n7310), .ZN(n6113) );
  NAND2_X1 U7701 ( .A1(n6114), .A2(n6113), .ZN(n9817) );
  NAND2_X1 U7702 ( .A1(n6115), .A2(n6116), .ZN(n6184) );
  OAI211_X1 U7703 ( .C1(n6116), .C2(n6115), .A(n9812), .B(n6184), .ZN(n6117)
         );
  OAI211_X1 U7704 ( .C1(n9815), .C2(n6185), .A(n6118), .B(n6117), .ZN(n6119)
         );
  OR2_X1 U7705 ( .A1(n6120), .A2(n6119), .ZN(P2_U3253) );
  AOI211_X1 U7706 ( .C1(n6123), .C2(n6122), .A(n6121), .B(n9483), .ZN(n6132)
         );
  NAND2_X1 U7707 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6531) );
  INV_X1 U7708 ( .A(n6531), .ZN(n6124) );
  AOI21_X1 U7709 ( .B1(n9820), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6124), .ZN(
        n6129) );
  OAI211_X1 U7710 ( .C1(n6127), .C2(n6126), .A(n9812), .B(n6125), .ZN(n6128)
         );
  OAI211_X1 U7711 ( .C1(n9815), .C2(n6130), .A(n6129), .B(n6128), .ZN(n6131)
         );
  OR2_X1 U7712 ( .A1(n6132), .A2(n6131), .ZN(P2_U3251) );
  AOI211_X1 U7713 ( .C1(n4281), .C2(n6134), .A(n6133), .B(n9483), .ZN(n6143)
         );
  AND2_X1 U7714 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6135) );
  AOI21_X1 U7715 ( .B1(n9820), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6135), .ZN(
        n6140) );
  OAI211_X1 U7716 ( .C1(n6138), .C2(n6137), .A(n9812), .B(n6136), .ZN(n6139)
         );
  OAI211_X1 U7717 ( .C1(n9815), .C2(n6141), .A(n6140), .B(n6139), .ZN(n6142)
         );
  OR2_X1 U7718 ( .A1(n6143), .A2(n6142), .ZN(P2_U3250) );
  AOI211_X1 U7719 ( .C1(n6146), .C2(n6145), .A(n6144), .B(n9483), .ZN(n6154)
         );
  INV_X1 U7720 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9302) );
  NOR2_X1 U7721 ( .A1(n9302), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6303) );
  AOI21_X1 U7722 ( .B1(n9820), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6303), .ZN(
        n6151) );
  OAI211_X1 U7723 ( .C1(n6149), .C2(n6148), .A(n9812), .B(n6147), .ZN(n6150)
         );
  OAI211_X1 U7724 ( .C1(n9815), .C2(n6152), .A(n6151), .B(n6150), .ZN(n6153)
         );
  OR2_X1 U7725 ( .A1(n6154), .A2(n6153), .ZN(P2_U3249) );
  AOI211_X1 U7726 ( .C1(n6157), .C2(n6156), .A(n6155), .B(n9483), .ZN(n6165)
         );
  INV_X1 U7727 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9318) );
  NOR2_X1 U7728 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9318), .ZN(n6255) );
  AOI21_X1 U7729 ( .B1(n9820), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6255), .ZN(
        n6162) );
  OAI211_X1 U7730 ( .C1(n6160), .C2(n6159), .A(n9812), .B(n6158), .ZN(n6161)
         );
  OAI211_X1 U7731 ( .C1(n9815), .C2(n6163), .A(n6162), .B(n6161), .ZN(n6164)
         );
  OR2_X1 U7732 ( .A1(n6165), .A2(n6164), .ZN(P2_U3248) );
  AOI211_X1 U7733 ( .C1(n6168), .C2(n6167), .A(n6166), .B(n9483), .ZN(n6177)
         );
  AND2_X1 U7734 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6169) );
  AOI21_X1 U7735 ( .B1(n9820), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6169), .ZN(
        n6174) );
  OAI211_X1 U7736 ( .C1(n6172), .C2(n6171), .A(n9812), .B(n6170), .ZN(n6173)
         );
  OAI211_X1 U7737 ( .C1(n9815), .C2(n6175), .A(n6174), .B(n6173), .ZN(n6176)
         );
  OR2_X1 U7738 ( .A1(n6177), .A2(n6176), .ZN(P2_U3252) );
  INV_X1 U7739 ( .A(n6185), .ZN(n6179) );
  AOI21_X1 U7740 ( .B1(n6179), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6178), .ZN(
        n6182) );
  NAND2_X1 U7741 ( .A1(n6216), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7742 ( .B1(n6216), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6180), .ZN(
        n6181) );
  NOR2_X1 U7743 ( .A1(n6182), .A2(n6181), .ZN(n6215) );
  AOI211_X1 U7744 ( .C1(n6182), .C2(n6181), .A(n6215), .B(n9483), .ZN(n6191)
         );
  AND2_X1 U7745 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6183) );
  AOI21_X1 U7746 ( .B1(n9820), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6183), .ZN(
        n6189) );
  OAI21_X1 U7747 ( .B1(n6185), .B2(n6111), .A(n6184), .ZN(n6187) );
  MUX2_X1 U7748 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7064), .S(n6216), .Z(n6186)
         );
  NAND2_X1 U7749 ( .A1(n6186), .A2(n6187), .ZN(n6220) );
  OAI211_X1 U7750 ( .C1(n6187), .C2(n6186), .A(n9812), .B(n6220), .ZN(n6188)
         );
  OAI211_X1 U7751 ( .C1(n9815), .C2(n6221), .A(n6189), .B(n6188), .ZN(n6190)
         );
  OR2_X1 U7752 ( .A1(n6191), .A2(n6190), .ZN(P2_U3254) );
  INV_X1 U7753 ( .A(n7347), .ZN(n6202) );
  NAND2_X1 U7754 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7755 ( .A(n6193), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7348) );
  INV_X1 U7756 ( .A(n7348), .ZN(n6385) );
  OAI222_X1 U7757 ( .A1(n9464), .A2(n6202), .B1(n6385), .B2(P1_U3084), .C1(
        n6194), .C2(n9462), .ZN(P1_U3340) );
  XOR2_X1 U7758 ( .A(n6195), .B(n6196), .Z(n6201) );
  INV_X1 U7759 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6197) );
  NOR2_X1 U7760 ( .A1(n9580), .A2(n6197), .ZN(n6199) );
  OAI22_X1 U7761 ( .A1(n6586), .A2(n8590), .B1(n8591), .B2(n9738), .ZN(n6198)
         );
  AOI211_X1 U7762 ( .C1(n8587), .C2(n6414), .A(n6199), .B(n6198), .ZN(n6200)
         );
  OAI21_X1 U7763 ( .B1(n6201), .B2(n8596), .A(n6200), .ZN(P1_U3235) );
  INV_X1 U7764 ( .A(n6670), .ZN(n6666) );
  OAI222_X1 U7765 ( .A1(n8404), .A2(n6203), .B1(n8400), .B2(n6202), .C1(n6666), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7766 ( .A(n7353), .ZN(n6213) );
  NOR2_X1 U7767 ( .A1(n6210), .A2(n6206), .ZN(n6207) );
  MUX2_X1 U7768 ( .A(n6206), .B(n6207), .S(P1_IR_REG_14__SCAN_IN), .Z(n6208)
         );
  INV_X1 U7769 ( .A(n6208), .ZN(n6211) );
  INV_X1 U7770 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7771 ( .A1(n6210), .A2(n6209), .ZN(n6309) );
  INV_X1 U7772 ( .A(n8933), .ZN(n8916) );
  OAI222_X1 U7773 ( .A1(n9464), .A2(n6213), .B1(n8916), .B2(n4246), .C1(n6212), 
        .C2(n9462), .ZN(P1_U3339) );
  INV_X1 U7774 ( .A(n6948), .ZN(n6951) );
  OAI222_X1 U7775 ( .A1(n8404), .A2(n6214), .B1(n8400), .B2(n6213), .C1(n6951), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U7776 ( .A1(n6316), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7777 ( .B1(n6316), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6217), .ZN(
        n6218) );
  AOI211_X1 U7778 ( .C1(n6219), .C2(n6218), .A(n6315), .B(n9483), .ZN(n6228)
         );
  NOR2_X1 U7779 ( .A1(n9332), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6848) );
  AOI21_X1 U7780 ( .B1(n9820), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6848), .ZN(
        n6226) );
  INV_X1 U7781 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7064) );
  OAI21_X1 U7782 ( .B1(n6221), .B2(n7064), .A(n6220), .ZN(n6224) );
  INV_X1 U7783 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6222) );
  MUX2_X1 U7784 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6222), .S(n6316), .Z(n6223)
         );
  NAND2_X1 U7785 ( .A1(n6223), .A2(n6224), .ZN(n6320) );
  OAI211_X1 U7786 ( .C1(n6224), .C2(n6223), .A(n9812), .B(n6320), .ZN(n6225)
         );
  OAI211_X1 U7787 ( .C1(n9815), .C2(n6321), .A(n6226), .B(n6225), .ZN(n6227)
         );
  OR2_X1 U7788 ( .A1(n6228), .A2(n6227), .ZN(P2_U3255) );
  INV_X1 U7789 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9554) );
  AOI22_X1 U7790 ( .A1(n7348), .A2(n9554), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n6385), .ZN(n6231) );
  NOR2_X1 U7791 ( .A1(n6232), .A2(n6231), .ZN(n6384) );
  AOI21_X1 U7792 ( .B1(n6232), .B2(n6231), .A(n6384), .ZN(n6242) );
  AND2_X1 U7793 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8536) );
  NOR2_X1 U7794 ( .A1(n9656), .A2(n6385), .ZN(n6233) );
  AOI211_X1 U7795 ( .C1(n9659), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n8536), .B(
        n6233), .ZN(n6241) );
  NAND2_X1 U7796 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7172), .ZN(n6235) );
  NAND2_X1 U7797 ( .A1(n6235), .A2(n6234), .ZN(n6239) );
  INV_X1 U7798 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6236) );
  MUX2_X1 U7799 ( .A(n6236), .B(P1_REG2_REG_13__SCAN_IN), .S(n7348), .Z(n6237)
         );
  INV_X1 U7800 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7801 ( .A1(n6238), .A2(n6239), .ZN(n6389) );
  OAI211_X1 U7802 ( .C1(n6239), .C2(n6238), .A(n9665), .B(n6389), .ZN(n6240)
         );
  OAI211_X1 U7803 ( .C1(n6242), .C2(n9622), .A(n6241), .B(n6240), .ZN(P1_U3254) );
  NAND2_X1 U7804 ( .A1(n6244), .A2(n6243), .ZN(n7536) );
  NAND2_X1 U7805 ( .A1(n7946), .A2(n7798), .ZN(n6245) );
  XNOR2_X1 U7806 ( .A(n7540), .B(n7749), .ZN(n6246) );
  XNOR2_X1 U7807 ( .A(n6245), .B(n6246), .ZN(n7537) );
  INV_X1 U7808 ( .A(n6245), .ZN(n6248) );
  INV_X1 U7809 ( .A(n6246), .ZN(n6247) );
  NAND2_X1 U7810 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  NAND2_X1 U7811 ( .A1(n7945), .A2(n7798), .ZN(n6292) );
  XNOR2_X1 U7812 ( .A(n6365), .B(n7799), .ZN(n6293) );
  XNOR2_X1 U7813 ( .A(n6292), .B(n6293), .ZN(n6296) );
  XNOR2_X1 U7814 ( .A(n6297), .B(n6296), .ZN(n6261) );
  AND3_X1 U7815 ( .A1(n6251), .A2(n6250), .A3(n6751), .ZN(n6252) );
  NAND2_X1 U7816 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  INV_X1 U7817 ( .A(n6255), .ZN(n6256) );
  OAI21_X1 U7818 ( .B1(n7886), .B2(P2_REG3_REG_3__SCAN_IN), .A(n6256), .ZN(
        n6259) );
  INV_X1 U7819 ( .A(n7889), .ZN(n7925) );
  OAI22_X1 U7820 ( .A1(n7925), .A2(n6257), .B1(n7904), .B2(n6563), .ZN(n6258)
         );
  AOI211_X1 U7821 ( .C1(n7914), .C2(n7946), .A(n6259), .B(n6258), .ZN(n6260)
         );
  OAI21_X1 U7822 ( .B1(n7909), .B2(n6261), .A(n6260), .ZN(P2_U3220) );
  INV_X1 U7823 ( .A(n7363), .ZN(n6330) );
  NAND2_X1 U7824 ( .A1(n6309), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U7825 ( .A(n6262), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9633) );
  AOI22_X1 U7826 ( .A1(n9633), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n4244), .ZN(n6263) );
  OAI21_X1 U7827 ( .B1(n6330), .B2(n9464), .A(n6263), .ZN(P1_U3338) );
  INV_X1 U7828 ( .A(n6590), .ZN(n6291) );
  INV_X1 U7829 ( .A(n6264), .ZN(n6266) );
  NAND2_X1 U7830 ( .A1(n9701), .A2(n5722), .ZN(n6274) );
  NAND2_X1 U7831 ( .A1(n7385), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7832 ( .A1(n7384), .A2(n9595), .ZN(n6270) );
  NAND2_X1 U7833 ( .A1(n6591), .A2(n7674), .ZN(n6273) );
  XNOR2_X1 U7834 ( .A(n6275), .B(n7680), .ZN(n6491) );
  AND2_X1 U7835 ( .A1(n6591), .A2(n5722), .ZN(n6276) );
  AOI21_X1 U7836 ( .B1(n9701), .B2(n7625), .A(n6276), .ZN(n6489) );
  XNOR2_X1 U7837 ( .A(n6491), .B(n6489), .ZN(n6277) );
  OAI211_X1 U7838 ( .C1(n6278), .C2(n6277), .A(n6493), .B(n9576), .ZN(n6290)
         );
  AND2_X1 U7839 ( .A1(n4246), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9598) );
  INV_X1 U7840 ( .A(n8587), .ZN(n8538) );
  NAND2_X1 U7841 ( .A1(n7471), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6287) );
  INV_X1 U7842 ( .A(n6281), .ZN(n6279) );
  NAND2_X1 U7843 ( .A1(n6279), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6627) );
  INV_X1 U7844 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7845 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  AND2_X1 U7846 ( .A1(n6627), .A2(n6282), .ZN(n9677) );
  NAND2_X1 U7847 ( .A1(n6918), .A2(n9677), .ZN(n6286) );
  NAND2_X1 U7848 ( .A1(n5781), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7849 ( .A1(n5782), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6284) );
  NAND4_X1 U7850 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n8886)
         );
  INV_X1 U7851 ( .A(n8886), .ZN(n6616) );
  OAI22_X1 U7852 ( .A1(n8538), .A2(n6586), .B1(n6616), .B2(n8590), .ZN(n6288)
         );
  AOI211_X1 U7853 ( .C1(n6591), .C2(n9575), .A(n9598), .B(n6288), .ZN(n6289)
         );
  OAI211_X1 U7854 ( .C1(n8483), .C2(n6291), .A(n6290), .B(n6289), .ZN(P1_U3228) );
  INV_X1 U7855 ( .A(n6292), .ZN(n6294) );
  AND2_X1 U7856 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  NOR2_X1 U7857 ( .A1(n6563), .A2(n7759), .ZN(n6298) );
  XNOR2_X1 U7858 ( .A(n9829), .B(n7799), .ZN(n6299) );
  NAND2_X1 U7859 ( .A1(n6298), .A2(n6299), .ZN(n6514) );
  INV_X1 U7860 ( .A(n6298), .ZN(n6301) );
  INV_X1 U7861 ( .A(n6299), .ZN(n6300) );
  NAND2_X1 U7862 ( .A1(n6301), .A2(n6300), .ZN(n6516) );
  NAND2_X1 U7863 ( .A1(n6514), .A2(n6516), .ZN(n6302) );
  XNOR2_X1 U7864 ( .A(n6515), .B(n6302), .ZN(n6308) );
  INV_X1 U7865 ( .A(n6303), .ZN(n6304) );
  OAI21_X1 U7866 ( .B1(n7886), .B2(n6483), .A(n6304), .ZN(n6306) );
  OAI22_X1 U7867 ( .A1(n7925), .A2(n9887), .B1(n7904), .B2(n6565), .ZN(n6305)
         );
  AOI211_X1 U7868 ( .C1(n7914), .C2(n7945), .A(n6306), .B(n6305), .ZN(n6307)
         );
  OAI21_X1 U7869 ( .B1(n6308), .B2(n7909), .A(n6307), .ZN(P2_U3232) );
  INV_X1 U7870 ( .A(n7373), .ZN(n6313) );
  NAND2_X1 U7871 ( .A1(n6310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U7872 ( .A(n6408), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8929) );
  AOI22_X1 U7873 ( .A1(n8929), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n4244), .ZN(n6311) );
  OAI21_X1 U7874 ( .B1(n6313), .B2(n9464), .A(n6311), .ZN(P1_U3337) );
  AOI22_X1 U7875 ( .A1(n7976), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8398), .ZN(n6312) );
  OAI21_X1 U7876 ( .B1(n6313), .B2(n8400), .A(n6312), .ZN(P2_U3342) );
  MUX2_X1 U7877 ( .A(n6941), .B(P2_REG2_REG_11__SCAN_IN), .S(n6458), .Z(n6314)
         );
  INV_X1 U7878 ( .A(n6314), .ZN(n6318) );
  OAI21_X1 U7879 ( .B1(n6318), .B2(n6317), .A(n6457), .ZN(n6328) );
  NOR2_X1 U7880 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7003), .ZN(n6319) );
  AOI21_X1 U7881 ( .B1(n9820), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6319), .ZN(
        n6326) );
  OAI21_X1 U7882 ( .B1(n6321), .B2(n6222), .A(n6320), .ZN(n6324) );
  INV_X1 U7883 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U7884 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6322), .S(n6458), .Z(n6323)
         );
  NAND2_X1 U7885 ( .A1(n6323), .A2(n6324), .ZN(n6453) );
  OAI211_X1 U7886 ( .C1(n6324), .C2(n6323), .A(n9812), .B(n6453), .ZN(n6325)
         );
  OAI211_X1 U7887 ( .C1(n9815), .C2(n6454), .A(n6326), .B(n6325), .ZN(n6327)
         );
  AOI21_X1 U7888 ( .B1(n9814), .B2(n6328), .A(n6327), .ZN(n6329) );
  INV_X1 U7889 ( .A(n6329), .ZN(P2_U3256) );
  INV_X1 U7890 ( .A(n7951), .ZN(n7960) );
  OAI222_X1 U7891 ( .A1(n8404), .A2(n6331), .B1(n8400), .B2(n6330), .C1(
        P2_U3152), .C2(n7960), .ZN(P2_U3343) );
  AND3_X1 U7892 ( .A1(n6767), .A2(n6332), .A3(n6751), .ZN(n6333) );
  XNOR2_X1 U7893 ( .A(n6760), .B(n6336), .ZN(n6335) );
  NAND2_X1 U7894 ( .A1(n6335), .A2(n8013), .ZN(n6883) );
  OR2_X1 U7895 ( .A1(n6336), .A2(n8013), .ZN(n6366) );
  NAND2_X1 U7896 ( .A1(n6883), .A2(n6366), .ZN(n9845) );
  INV_X1 U7897 ( .A(n6343), .ZN(n9866) );
  AOI22_X1 U7898 ( .A1(n9866), .A2(n8271), .B1(n8268), .B2(n7947), .ZN(n9868)
         );
  OAI21_X1 U7899 ( .B1(n4791), .B2(n8250), .A(n9868), .ZN(n6340) );
  NOR2_X1 U7900 ( .A1(n8253), .A2(n9813), .ZN(n6339) );
  AOI21_X1 U7901 ( .B1(n6340), .B2(n8253), .A(n6339), .ZN(n6342) );
  OAI21_X1 U7902 ( .B1(n8255), .B2(n8277), .A(n9864), .ZN(n6341) );
  OAI211_X1 U7903 ( .C1(n6343), .C2(n8262), .A(n6342), .B(n6341), .ZN(P2_U3296) );
  NAND2_X1 U7904 ( .A1(n6344), .A2(n6469), .ZN(n6348) );
  NAND2_X1 U7905 ( .A1(n6345), .A2(n6346), .ZN(n6347) );
  NAND2_X1 U7906 ( .A1(n6348), .A2(n6347), .ZN(n6370) );
  NAND2_X1 U7907 ( .A1(n6370), .A2(n4328), .ZN(n6351) );
  NAND2_X1 U7908 ( .A1(n6356), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U7909 ( .A1(n6351), .A2(n6350), .ZN(n6479) );
  XNOR2_X1 U7910 ( .A(n6478), .B(n6479), .ZN(n9883) );
  INV_X1 U7911 ( .A(n6883), .ZN(n7150) );
  NAND2_X1 U7912 ( .A1(n9883), .A2(n7150), .ZN(n6360) );
  NAND3_X1 U7913 ( .A1(n6352), .A2(n6478), .A3(n6353), .ZN(n6354) );
  NAND2_X1 U7914 ( .A1(n6355), .A2(n6354), .ZN(n6358) );
  OAI22_X1 U7915 ( .A1(n6356), .A2(n8181), .B1(n6563), .B2(n8179), .ZN(n6357)
         );
  AOI21_X1 U7916 ( .B1(n6358), .B2(n8271), .A(n6357), .ZN(n6359) );
  OAI22_X1 U7917 ( .A1(n8253), .A2(n6361), .B1(n8250), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6364) );
  OR2_X1 U7918 ( .A1(n6470), .A2(n9864), .ZN(n9870) );
  NAND2_X1 U7919 ( .A1(n6375), .A2(n6257), .ZN(n9830) );
  OR2_X1 U7920 ( .A1(n6375), .A2(n6257), .ZN(n6362) );
  NAND2_X1 U7921 ( .A1(n9830), .A2(n6362), .ZN(n9881) );
  NOR2_X1 U7922 ( .A1(n9881), .A2(n8062), .ZN(n6363) );
  AOI211_X1 U7923 ( .C1(n8255), .C2(n6365), .A(n6364), .B(n6363), .ZN(n6369)
         );
  INV_X1 U7924 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U7925 ( .A1(n9883), .A2(n7159), .ZN(n6368) );
  OAI211_X1 U7926 ( .C1(n9885), .C2(n9848), .A(n6369), .B(n6368), .ZN(P2_U3293) );
  XNOR2_X1 U7927 ( .A(n4328), .B(n6370), .ZN(n9879) );
  INV_X1 U7928 ( .A(n9879), .ZN(n6383) );
  INV_X1 U7929 ( .A(n6352), .ZN(n6371) );
  AOI21_X1 U7930 ( .B1(n4328), .B2(n6372), .A(n6371), .ZN(n6374) );
  OAI222_X1 U7931 ( .A1(n8179), .A2(n6480), .B1(n8181), .B2(n6345), .C1(n9842), 
        .C2(n6374), .ZN(n9877) );
  AND2_X1 U7932 ( .A1(n9870), .A2(n7540), .ZN(n6376) );
  OR2_X1 U7933 ( .A1(n6376), .A2(n6375), .ZN(n9876) );
  INV_X1 U7934 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6377) );
  OAI22_X1 U7935 ( .A1(n8062), .A2(n9876), .B1(n6377), .B2(n8250), .ZN(n6378)
         );
  INV_X1 U7936 ( .A(n6378), .ZN(n6380) );
  NAND2_X1 U7937 ( .A1(n8255), .A2(n7540), .ZN(n6379) );
  OAI211_X1 U7938 ( .C1(n8253), .C2(n9362), .A(n6380), .B(n6379), .ZN(n6381)
         );
  AOI21_X1 U7939 ( .B1(n9877), .B2(n9846), .A(n6381), .ZN(n6382) );
  OAI21_X1 U7940 ( .B1(n6383), .B2(n8262), .A(n6382), .ZN(P2_U3294) );
  AOI21_X1 U7941 ( .B1(n6385), .B2(n9554), .A(n6384), .ZN(n6387) );
  INV_X1 U7942 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8915) );
  AOI22_X1 U7943 ( .A1(n8933), .A2(n8915), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8916), .ZN(n6386) );
  NOR2_X1 U7944 ( .A1(n6387), .A2(n6386), .ZN(n8914) );
  AOI21_X1 U7945 ( .B1(n6387), .B2(n6386), .A(n8914), .ZN(n6396) );
  NOR2_X1 U7946 ( .A1(n7356), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8420) );
  INV_X1 U7947 ( .A(n8420), .ZN(n6388) );
  OAI21_X1 U7948 ( .B1(n9656), .B2(n8916), .A(n6388), .ZN(n6394) );
  NAND2_X1 U7949 ( .A1(n7348), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7950 ( .A1(n6390), .A2(n6389), .ZN(n8932) );
  XNOR2_X1 U7951 ( .A(n8933), .B(n8932), .ZN(n6391) );
  NOR2_X1 U7952 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n6391), .ZN(n8934) );
  AOI21_X1 U7953 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n6391), .A(n8934), .ZN(
        n6392) );
  NOR2_X1 U7954 ( .A1(n6392), .A2(n8956), .ZN(n6393) );
  AOI211_X1 U7955 ( .C1(n9659), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n6394), .B(
        n6393), .ZN(n6395) );
  OAI21_X1 U7956 ( .B1(n6396), .B2(n9622), .A(n6395), .ZN(P1_U3255) );
  NAND4_X1 U7957 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6655)
         );
  INV_X1 U7958 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9579) );
  OAI22_X1 U7959 ( .A1(n9719), .A2(n6401), .B1(n9579), .B2(n9118), .ZN(n6402)
         );
  INV_X1 U7960 ( .A(n6402), .ZN(n6405) );
  INV_X1 U7961 ( .A(n6403), .ZN(n9675) );
  OAI21_X1 U7962 ( .B1(n9698), .B2(n9539), .A(n9574), .ZN(n6404) );
  OAI211_X1 U7963 ( .C1(n6406), .C2(n9715), .A(n6405), .B(n6404), .ZN(P1_U3291) );
  INV_X1 U7964 ( .A(n7340), .ZN(n6451) );
  INV_X1 U7965 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7966 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U7967 ( .A1(n6409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6411) );
  INV_X1 U7968 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6410) );
  OR2_X1 U7969 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  NAND2_X1 U7970 ( .A1(n6411), .A2(n6410), .ZN(n6580) );
  INV_X1 U7971 ( .A(n8926), .ZN(n9655) );
  OAI222_X1 U7972 ( .A1(n9464), .A2(n6451), .B1(n9655), .B2(P1_U3084), .C1(
        n6413), .C2(n9462), .ZN(P1_U3336) );
  NAND2_X1 U7973 ( .A1(n6420), .A2(n6437), .ZN(n6436) );
  NAND2_X1 U7974 ( .A1(n6414), .A2(n6076), .ZN(n6415) );
  NAND2_X1 U7975 ( .A1(n4250), .A2(n8642), .ZN(n6416) );
  AND2_X2 U7976 ( .A1(n6584), .A2(n6416), .ZN(n8805) );
  OAI21_X1 U7977 ( .B1(n6417), .B2(n8805), .A(n6585), .ZN(n9742) );
  INV_X1 U7978 ( .A(n9742), .ZN(n6435) );
  NOR2_X1 U7979 ( .A1(n5693), .A2(n9125), .ZN(n6418) );
  NAND2_X1 U7980 ( .A1(n9719), .A2(n6418), .ZN(n9179) );
  INV_X1 U7981 ( .A(n8805), .ZN(n6422) );
  NOR2_X1 U7982 ( .A1(n5913), .A2(n5973), .ZN(n6438) );
  INV_X1 U7983 ( .A(n6414), .ZN(n8640) );
  NAND2_X1 U7984 ( .A1(n8640), .A2(n6076), .ZN(n6421) );
  OAI21_X1 U7985 ( .B1(n6422), .B2(n8645), .A(n9706), .ZN(n6427) );
  NAND2_X1 U7986 ( .A1(n5764), .A2(n9679), .ZN(n6424) );
  INV_X1 U7987 ( .A(n7218), .ZN(n8863) );
  NAND2_X1 U7988 ( .A1(n5762), .A2(n8863), .ZN(n6423) );
  OAI22_X1 U7989 ( .A1(n8640), .A2(n9685), .B1(n6586), .B2(n9687), .ZN(n6426)
         );
  AOI21_X1 U7990 ( .B1(n6427), .B2(n9707), .A(n6426), .ZN(n6428) );
  OAI21_X1 U7991 ( .B1(n6435), .B2(n9726), .A(n6428), .ZN(n9740) );
  NAND2_X1 U7992 ( .A1(n9740), .A2(n9719), .ZN(n6434) );
  OAI22_X1 U7993 ( .A1(n9719), .A2(n6429), .B1(n6197), .B2(n9118), .ZN(n6432)
         );
  NAND2_X1 U7994 ( .A1(n9732), .A2(n5973), .ZN(n6445) );
  NAND2_X1 U7995 ( .A1(n6445), .A2(n8642), .ZN(n6430) );
  NAND2_X1 U7996 ( .A1(n9694), .A2(n6430), .ZN(n9739) );
  NOR2_X1 U7997 ( .A1(n8974), .A2(n9739), .ZN(n6431) );
  AOI211_X1 U7998 ( .C1(n9539), .C2(n8642), .A(n6432), .B(n6431), .ZN(n6433)
         );
  OAI211_X1 U7999 ( .C1(n6435), .C2(n9179), .A(n6434), .B(n6433), .ZN(P1_U3289) );
  OAI21_X1 U8000 ( .B1(n6420), .B2(n6437), .A(n6436), .ZN(n9729) );
  INV_X1 U8001 ( .A(n6438), .ZN(n6439) );
  NAND2_X1 U8002 ( .A1(n6439), .A2(n6420), .ZN(n6441) );
  NAND2_X1 U8003 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  NAND2_X1 U8004 ( .A1(n6442), .A2(n9707), .ZN(n6444) );
  AOI22_X1 U8005 ( .A1(n9702), .A2(n4250), .B1(n5913), .B2(n9700), .ZN(n6443)
         );
  NAND2_X1 U8006 ( .A1(n6444), .A2(n6443), .ZN(n9727) );
  AOI21_X1 U8007 ( .B1(n9574), .B2(n6076), .A(n9786), .ZN(n6446) );
  NAND2_X1 U8008 ( .A1(n6446), .A2(n6445), .ZN(n9731) );
  OAI22_X1 U8009 ( .A1(n9731), .A2(n9679), .B1(n6447), .B2(n9118), .ZN(n6448)
         );
  OAI21_X1 U8010 ( .B1(n9727), .B2(n6448), .A(n9719), .ZN(n6450) );
  AOI22_X1 U8011 ( .A1(n9539), .A2(n6076), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9715), .ZN(n6449) );
  OAI211_X1 U8012 ( .C1(n9198), .C2(n9729), .A(n6450), .B(n6449), .ZN(P1_U3290) );
  INV_X1 U8013 ( .A(n7986), .ZN(n7991) );
  OAI222_X1 U8014 ( .A1(n8404), .A2(n6452), .B1(n8400), .B2(n6451), .C1(n7991), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U8015 ( .B1(n6322), .B2(n6454), .A(n6453), .ZN(n6456) );
  INV_X1 U8016 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U8017 ( .A1(n6539), .A2(n9941), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n6544), .ZN(n6455) );
  NOR2_X1 U8018 ( .A1(n6456), .A2(n6455), .ZN(n6543) );
  AOI21_X1 U8019 ( .B1(n6456), .B2(n6455), .A(n6543), .ZN(n6466) );
  AOI22_X1 U8020 ( .A1(n6539), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n5078), .B2(
        n6544), .ZN(n6460) );
  OAI21_X1 U8021 ( .B1(n6458), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6457), .ZN(
        n6459) );
  NAND2_X1 U8022 ( .A1(n6460), .A2(n6459), .ZN(n6538) );
  OAI21_X1 U8023 ( .B1(n6460), .B2(n6459), .A(n6538), .ZN(n6461) );
  NAND2_X1 U8024 ( .A1(n6461), .A2(n9814), .ZN(n6465) );
  INV_X1 U8025 ( .A(n9815), .ZN(n9489) );
  INV_X1 U8026 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8027 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7550) );
  OAI21_X1 U8028 ( .B1(n9472), .B2(n6462), .A(n7550), .ZN(n6463) );
  AOI21_X1 U8029 ( .B1(n9489), .B2(n6539), .A(n6463), .ZN(n6464) );
  OAI211_X1 U8030 ( .C1(n6466), .C2(n9817), .A(n6465), .B(n6464), .ZN(P2_U3257) );
  XNOR2_X1 U8031 ( .A(n6344), .B(n6467), .ZN(n6468) );
  AOI222_X1 U8032 ( .A1(n8271), .A2(n6468), .B1(n7946), .B2(n8268), .C1(n7949), 
        .C2(n8266), .ZN(n9872) );
  XNOR2_X1 U8033 ( .A(n6344), .B(n6469), .ZN(n9875) );
  NAND2_X1 U8034 ( .A1(n6470), .A2(n9864), .ZN(n9869) );
  NAND3_X1 U8035 ( .A1(n8277), .A2(n9870), .A3(n9869), .ZN(n6471) );
  OAI21_X1 U8036 ( .B1(n8250), .B2(n4872), .A(n6471), .ZN(n6472) );
  AOI21_X1 U8037 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n9848), .A(n6472), .ZN(
        n6473) );
  OAI21_X1 U8038 ( .B1(n6346), .B2(n8281), .A(n6473), .ZN(n6474) );
  AOI21_X1 U8039 ( .B1(n8284), .B2(n9875), .A(n6474), .ZN(n6475) );
  OAI21_X1 U8040 ( .B1(n9848), .B2(n9872), .A(n6475), .ZN(P2_U3295) );
  XNOR2_X1 U8041 ( .A(n6476), .B(n9825), .ZN(n6477) );
  OAI222_X1 U8042 ( .A1(n8179), .A2(n6565), .B1(n8181), .B2(n6480), .C1(n6477), 
        .C2(n9842), .ZN(n9889) );
  INV_X1 U8043 ( .A(n9889), .ZN(n6488) );
  NAND2_X1 U8044 ( .A1(n6479), .A2(n6478), .ZN(n6482) );
  NAND2_X1 U8045 ( .A1(n6480), .A2(n6257), .ZN(n6481) );
  NAND2_X1 U8046 ( .A1(n6482), .A2(n6481), .ZN(n6562) );
  XNOR2_X1 U8047 ( .A(n6562), .B(n9825), .ZN(n9891) );
  XNOR2_X1 U8048 ( .A(n9830), .B(n9829), .ZN(n9888) );
  OAI22_X1 U8049 ( .A1(n8253), .A2(n6085), .B1(n6483), .B2(n8250), .ZN(n6484)
         );
  AOI21_X1 U8050 ( .B1(n8255), .B2(n9829), .A(n6484), .ZN(n6485) );
  OAI21_X1 U8051 ( .B1(n8062), .B2(n9888), .A(n6485), .ZN(n6486) );
  AOI21_X1 U8052 ( .B1(n9891), .B2(n8284), .A(n6486), .ZN(n6487) );
  OAI21_X1 U8053 ( .B1(n6488), .B2(n9848), .A(n6487), .ZN(P2_U3292) );
  INV_X1 U8054 ( .A(n9677), .ZN(n6513) );
  INV_X1 U8055 ( .A(n6489), .ZN(n6490) );
  NAND2_X1 U8056 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  NAND2_X1 U8057 ( .A1(n8886), .A2(n7641), .ZN(n6499) );
  NAND2_X1 U8058 ( .A1(n7385), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U8059 ( .A1(n7384), .A2(n6494), .ZN(n6495) );
  OAI211_X1 U8060 ( .C1(n8664), .C2(n6497), .A(n6496), .B(n6495), .ZN(n9676)
         );
  NAND2_X1 U8061 ( .A1(n9676), .A2(n7674), .ZN(n6498) );
  NAND2_X1 U8062 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  XNOR2_X1 U8063 ( .A(n6500), .B(n8448), .ZN(n6684) );
  AND2_X1 U8064 ( .A1(n9676), .A2(n7641), .ZN(n6501) );
  AOI21_X1 U8065 ( .B1(n8886), .B2(n7625), .A(n6501), .ZN(n6502) );
  NAND2_X1 U8066 ( .A1(n6503), .A2(n6502), .ZN(n6688) );
  OAI21_X1 U8067 ( .B1(n6503), .B2(n6502), .A(n6688), .ZN(n6504) );
  NAND2_X1 U8068 ( .A1(n6504), .A2(n9576), .ZN(n6512) );
  NAND2_X1 U8069 ( .A1(n7471), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6508) );
  XNOR2_X1 U8070 ( .A(n6627), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U8071 ( .A1(n6918), .A2(n8568), .ZN(n6507) );
  NAND2_X1 U8072 ( .A1(n5781), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8073 ( .A1(n8455), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6505) );
  NAND4_X1 U8074 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n8885)
         );
  INV_X1 U8075 ( .A(n8885), .ZN(n9686) );
  OAI22_X1 U8076 ( .A1(n8538), .A2(n9684), .B1(n9686), .B2(n8590), .ZN(n6509)
         );
  AOI211_X1 U8077 ( .C1(n9676), .C2(n9575), .A(n6510), .B(n6509), .ZN(n6511)
         );
  OAI211_X1 U8078 ( .C1(n8483), .C2(n6513), .A(n6512), .B(n6511), .ZN(P1_U3225) );
  XNOR2_X1 U8079 ( .A(n9897), .B(n7799), .ZN(n6731) );
  NAND2_X1 U8080 ( .A1(n7942), .A2(n7798), .ZN(n6732) );
  XNOR2_X1 U8081 ( .A(n6731), .B(n6732), .ZN(n6526) );
  NAND2_X1 U8082 ( .A1(n6515), .A2(n6514), .ZN(n6517) );
  NAND2_X1 U8083 ( .A1(n6517), .A2(n6516), .ZN(n6552) );
  INV_X1 U8084 ( .A(n6552), .ZN(n6523) );
  NOR2_X1 U8085 ( .A1(n6565), .A2(n7759), .ZN(n6518) );
  XNOR2_X1 U8086 ( .A(n9836), .B(n7799), .ZN(n6527) );
  NAND2_X1 U8087 ( .A1(n6518), .A2(n6527), .ZN(n6524) );
  INV_X1 U8088 ( .A(n6518), .ZN(n6520) );
  INV_X1 U8089 ( .A(n6527), .ZN(n6519) );
  NAND2_X1 U8090 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  NAND2_X1 U8091 ( .A1(n6524), .A2(n6521), .ZN(n6555) );
  AND2_X1 U8092 ( .A1(n6526), .A2(n6524), .ZN(n6525) );
  OAI21_X1 U8093 ( .B1(n6526), .B2(n6553), .A(n6735), .ZN(n6535) );
  INV_X1 U8094 ( .A(n7898), .ZN(n7918) );
  INV_X1 U8095 ( .A(n6526), .ZN(n6528) );
  NAND3_X1 U8096 ( .A1(n7918), .A2(n6528), .A3(n6527), .ZN(n6529) );
  AOI21_X1 U8097 ( .B1(n6529), .B2(n7903), .A(n6565), .ZN(n6534) );
  INV_X1 U8098 ( .A(n6530), .ZN(n6608) );
  AOI22_X1 U8099 ( .A1(n7913), .A2(n7941), .B1(n9897), .B2(n7889), .ZN(n6532)
         );
  OAI211_X1 U8100 ( .C1(n6608), .C2(n7886), .A(n6532), .B(n6531), .ZN(n6533)
         );
  AOI211_X1 U8101 ( .C1(n6535), .C2(n7919), .A(n6534), .B(n6533), .ZN(n6536)
         );
  INV_X1 U8102 ( .A(n6536), .ZN(P2_U3241) );
  NOR2_X1 U8103 ( .A1(n6670), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6537) );
  AOI21_X1 U8104 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6670), .A(n6537), .ZN(
        n6541) );
  OAI21_X1 U8105 ( .B1(n6541), .B2(n6540), .A(n6669), .ZN(n6550) );
  AND2_X1 U8106 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7260) );
  AOI21_X1 U8107 ( .B1(n9820), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7260), .ZN(
        n6542) );
  OAI21_X1 U8108 ( .B1(n9815), .B2(n6666), .A(n6542), .ZN(n6549) );
  AOI21_X1 U8109 ( .B1(n6544), .B2(n9941), .A(n6543), .ZN(n6546) );
  INV_X1 U8110 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U8111 ( .A1(n6670), .A2(n6665), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n6666), .ZN(n6545) );
  NOR2_X1 U8112 ( .A1(n6546), .A2(n6545), .ZN(n6664) );
  AOI21_X1 U8113 ( .B1(n6546), .B2(n6545), .A(n6664), .ZN(n6547) );
  NOR2_X1 U8114 ( .A1(n6547), .A2(n9817), .ZN(n6548) );
  AOI211_X1 U8115 ( .C1(n6550), .C2(n9814), .A(n6549), .B(n6548), .ZN(n6551)
         );
  INV_X1 U8116 ( .A(n6551), .ZN(P2_U3258) );
  INV_X1 U8117 ( .A(n6553), .ZN(n6554) );
  AOI211_X1 U8118 ( .C1(n6555), .C2(n6552), .A(n7909), .B(n6554), .ZN(n6560)
         );
  AOI22_X1 U8119 ( .A1(n7944), .A2(n8266), .B1(n8268), .B2(n7942), .ZN(n9841)
         );
  OAI22_X1 U8120 ( .A1(n7924), .A2(n9841), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6556), .ZN(n6559) );
  INV_X1 U8121 ( .A(n9833), .ZN(n6557) );
  OAI22_X1 U8122 ( .A1(n7925), .A2(n9893), .B1(n7886), .B2(n6557), .ZN(n6558)
         );
  OR3_X1 U8123 ( .A1(n6560), .A2(n6559), .A3(n6558), .ZN(P2_U3229) );
  AND2_X1 U8124 ( .A1(n9825), .A2(n9840), .ZN(n6561) );
  OR2_X1 U8125 ( .A1(n7942), .A2(n9897), .ZN(n6568) );
  NAND2_X1 U8126 ( .A1(n6563), .A2(n9887), .ZN(n9826) );
  INV_X1 U8127 ( .A(n9826), .ZN(n6564) );
  NAND2_X1 U8128 ( .A1(n9840), .A2(n6564), .ZN(n6567) );
  NAND2_X1 U8129 ( .A1(n6565), .A2(n9893), .ZN(n6566) );
  NAND2_X1 U8130 ( .A1(n6600), .A2(n6569), .ZN(n6778) );
  NAND2_X1 U8131 ( .A1(n7942), .A2(n9897), .ZN(n6776) );
  NAND2_X1 U8132 ( .A1(n6778), .A2(n6776), .ZN(n6570) );
  XOR2_X1 U8133 ( .A(n6571), .B(n6570), .Z(n6765) );
  XOR2_X1 U8134 ( .A(n6572), .B(n6571), .Z(n6573) );
  AOI22_X1 U8135 ( .A1(n7940), .A2(n8268), .B1(n8266), .B2(n7942), .ZN(n6745)
         );
  OAI21_X1 U8136 ( .B1(n6573), .B2(n9842), .A(n6745), .ZN(n6761) );
  NAND2_X1 U8137 ( .A1(n6761), .A2(n8253), .ZN(n6579) );
  INV_X1 U8138 ( .A(n6607), .ZN(n6574) );
  AND2_X1 U8139 ( .A1(n6607), .A2(n6779), .ZN(n6874) );
  AOI211_X1 U8140 ( .C1(n6763), .C2(n6574), .A(n9921), .B(n6874), .ZN(n6762)
         );
  OR2_X1 U8141 ( .A1(n6575), .A2(n9838), .ZN(n7280) );
  AOI22_X1 U8142 ( .A1(n9848), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n6746), .B2(
        n9834), .ZN(n6576) );
  OAI21_X1 U8143 ( .B1(n8281), .B2(n6779), .A(n6576), .ZN(n6577) );
  AOI21_X1 U8144 ( .B1(n6762), .B2(n8259), .A(n6577), .ZN(n6578) );
  OAI211_X1 U8145 ( .C1(n6765), .C2(n8262), .A(n6579), .B(n6578), .ZN(P2_U3289) );
  INV_X1 U8146 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9411) );
  INV_X1 U8147 ( .A(n7331), .ZN(n6582) );
  INV_X1 U8148 ( .A(n7993), .ZN(n8007) );
  OAI222_X1 U8149 ( .A1(n8404), .A2(n9411), .B1(n8400), .B2(n6582), .C1(
        P2_U3152), .C2(n8007), .ZN(P2_U3340) );
  INV_X1 U8150 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8151 ( .A1(n6580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6581) );
  XNOR2_X1 U8152 ( .A(n6581), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8940) );
  INV_X1 U8153 ( .A(n8940), .ZN(n8951) );
  OAI222_X1 U8154 ( .A1(n9462), .A2(n6583), .B1(n9464), .B2(n6582), .C1(
        P1_U3084), .C2(n8951), .ZN(P1_U3335) );
  NAND2_X1 U8155 ( .A1(n6586), .A2(n9693), .ZN(n8838) );
  NAND2_X1 U8156 ( .A1(n8887), .A2(n9744), .ZN(n8647) );
  NAND2_X1 U8157 ( .A1(n8838), .A2(n8647), .ZN(n9704) );
  NAND2_X1 U8158 ( .A1(n6586), .A2(n9744), .ZN(n6587) );
  NAND2_X1 U8159 ( .A1(n6588), .A2(n6587), .ZN(n6613) );
  NAND2_X1 U8160 ( .A1(n9684), .A2(n6591), .ZN(n8837) );
  INV_X1 U8161 ( .A(n6591), .ZN(n9750) );
  NAND2_X1 U8162 ( .A1(n9701), .A2(n9750), .ZN(n8835) );
  XNOR2_X1 U8163 ( .A(n6613), .B(n8804), .ZN(n9754) );
  OR2_X1 U8164 ( .A1(n9695), .A2(n9750), .ZN(n6589) );
  NAND2_X1 U8165 ( .A1(n9672), .A2(n6589), .ZN(n9751) );
  AOI22_X1 U8166 ( .A1(n9539), .A2(n6591), .B1(n9714), .B2(n6590), .ZN(n6592)
         );
  OAI21_X1 U8167 ( .B1(n9751), .B2(n8974), .A(n6592), .ZN(n6597) );
  NAND2_X1 U8168 ( .A1(n8643), .A2(n8642), .ZN(n9705) );
  NAND2_X1 U8169 ( .A1(n9706), .A2(n9705), .ZN(n8834) );
  INV_X1 U8170 ( .A(n9704), .ZN(n9691) );
  NAND2_X1 U8171 ( .A1(n8834), .A2(n9691), .ZN(n9703) );
  NAND2_X1 U8172 ( .A1(n9703), .A2(n8838), .ZN(n6638) );
  XNOR2_X1 U8173 ( .A(n6638), .B(n8804), .ZN(n6595) );
  INV_X1 U8174 ( .A(n9726), .ZN(n9537) );
  NAND2_X1 U8175 ( .A1(n9754), .A2(n9537), .ZN(n6594) );
  AOI22_X1 U8176 ( .A1(n9702), .A2(n8886), .B1(n8887), .B2(n9700), .ZN(n6593)
         );
  OAI211_X1 U8177 ( .C1(n9682), .C2(n6595), .A(n6594), .B(n6593), .ZN(n9752)
         );
  MUX2_X1 U8178 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9752), .S(n9719), .Z(n6596)
         );
  AOI211_X1 U8179 ( .C1(n9699), .C2(n9754), .A(n6597), .B(n6596), .ZN(n6598)
         );
  INV_X1 U8180 ( .A(n6598), .ZN(P1_U3287) );
  NAND2_X1 U8181 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  XNOR2_X1 U8182 ( .A(n6601), .B(n6602), .ZN(n9903) );
  XNOR2_X1 U8183 ( .A(n6603), .B(n6602), .ZN(n6604) );
  AOI222_X1 U8184 ( .A1(n8271), .A2(n6604), .B1(n7941), .B2(n8268), .C1(n7943), 
        .C2(n8266), .ZN(n9902) );
  MUX2_X1 U8185 ( .A(n6605), .B(n9902), .S(n8253), .Z(n6612) );
  AND2_X1 U8186 ( .A1(n9831), .A2(n9897), .ZN(n6606) );
  NOR2_X1 U8187 ( .A1(n6607), .A2(n6606), .ZN(n9900) );
  OAI22_X1 U8188 ( .A1(n8281), .A2(n6609), .B1(n8250), .B2(n6608), .ZN(n6610)
         );
  AOI21_X1 U8189 ( .B1(n9900), .B2(n8277), .A(n6610), .ZN(n6611) );
  OAI211_X1 U8190 ( .C1(n8262), .C2(n9903), .A(n6612), .B(n6611), .ZN(P2_U3290) );
  NAND2_X1 U8191 ( .A1(n6613), .A2(n8804), .ZN(n6615) );
  NAND2_X1 U8192 ( .A1(n9684), .A2(n9750), .ZN(n6614) );
  NAND2_X1 U8193 ( .A1(n6615), .A2(n6614), .ZN(n9671) );
  NAND2_X1 U8194 ( .A1(n6616), .A2(n9676), .ZN(n6816) );
  INV_X1 U8195 ( .A(n9676), .ZN(n9757) );
  NAND2_X1 U8196 ( .A1(n8886), .A2(n9757), .ZN(n8836) );
  NAND2_X1 U8197 ( .A1(n8886), .A2(n9676), .ZN(n6617) );
  OAI21_X2 U8198 ( .B1(n9671), .B2(n9681), .A(n6617), .ZN(n6810) );
  NAND2_X1 U8199 ( .A1(n8666), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8200 ( .A1(n7384), .A2(n6618), .ZN(n6619) );
  OAI211_X1 U8201 ( .C1(n8664), .C2(n6621), .A(n6620), .B(n6619), .ZN(n8567)
         );
  NAND2_X1 U8202 ( .A1(n9686), .A2(n8567), .ZN(n8678) );
  INV_X1 U8203 ( .A(n8567), .ZN(n9762) );
  NAND2_X1 U8204 ( .A1(n8885), .A2(n9762), .ZN(n8677) );
  NAND2_X1 U8205 ( .A1(n9686), .A2(n9762), .ZN(n6622) );
  INV_X1 U8206 ( .A(n6627), .ZN(n6624) );
  AND2_X1 U8207 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6623) );
  NAND2_X1 U8208 ( .A1(n6624), .A2(n6623), .ZN(n6646) );
  INV_X1 U8209 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6626) );
  INV_X1 U8210 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6625) );
  OAI21_X1 U8211 ( .B1(n6627), .B2(n6626), .A(n6625), .ZN(n6628) );
  AND2_X1 U8212 ( .A1(n6646), .A2(n6628), .ZN(n6679) );
  NAND2_X1 U8213 ( .A1(n6918), .A2(n6679), .ZN(n6632) );
  NAND2_X1 U8214 ( .A1(n7471), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8215 ( .A1(n8456), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U8216 ( .A1(n5782), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6629) );
  NAND4_X1 U8217 ( .A1(n6632), .A2(n6631), .A3(n6630), .A4(n6629), .ZN(n8884)
         );
  INV_X1 U8218 ( .A(n8884), .ZN(n6867) );
  INV_X1 U8219 ( .A(n8666), .ZN(n8662) );
  NAND2_X1 U8220 ( .A1(n7463), .A2(n6633), .ZN(n6636) );
  NAND2_X1 U8221 ( .A1(n7384), .A2(n6634), .ZN(n6635) );
  OAI211_X1 U8222 ( .C1(n8662), .C2(n6637), .A(n6636), .B(n6635), .ZN(n6721)
         );
  NAND2_X1 U8223 ( .A1(n6867), .A2(n6721), .ZN(n8681) );
  NAND2_X1 U8224 ( .A1(n8884), .A2(n9770), .ZN(n8680) );
  NAND2_X1 U8225 ( .A1(n8681), .A2(n8680), .ZN(n8810) );
  XNOR2_X1 U8226 ( .A(n6722), .B(n8810), .ZN(n9773) );
  INV_X1 U8227 ( .A(n9773), .ZN(n6660) );
  NAND2_X1 U8228 ( .A1(n8678), .A2(n6816), .ZN(n8841) );
  NAND2_X1 U8229 ( .A1(n8836), .A2(n8677), .ZN(n6640) );
  NAND2_X1 U8230 ( .A1(n8678), .A2(n6640), .ZN(n8657) );
  NAND2_X1 U8231 ( .A1(n6641), .A2(n8810), .ZN(n6642) );
  NAND2_X1 U8232 ( .A1(n6706), .A2(n6642), .ZN(n6643) );
  NAND2_X1 U8233 ( .A1(n6643), .A2(n9707), .ZN(n6653) );
  NAND2_X1 U8234 ( .A1(n7471), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6651) );
  INV_X1 U8235 ( .A(n6646), .ZN(n6645) );
  NAND2_X1 U8236 ( .A1(n6645), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8237 ( .A1(n6646), .A2(n9357), .ZN(n6647) );
  AND2_X1 U8238 ( .A1(n6713), .A2(n6647), .ZN(n6864) );
  NAND2_X1 U8239 ( .A1(n6918), .A2(n6864), .ZN(n6650) );
  NAND2_X1 U8240 ( .A1(n8456), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8241 ( .A1(n8455), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6648) );
  NAND4_X1 U8242 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n8883)
         );
  AOI22_X1 U8243 ( .A1(n9700), .A2(n8885), .B1(n8883), .B2(n9702), .ZN(n6652)
         );
  NAND2_X1 U8244 ( .A1(n6653), .A2(n6652), .ZN(n9771) );
  AND2_X1 U8245 ( .A1(n6813), .A2(n9770), .ZN(n6725) );
  INV_X1 U8246 ( .A(n6725), .ZN(n6654) );
  OAI211_X1 U8247 ( .C1(n9770), .C2(n6813), .A(n6654), .B(n9778), .ZN(n9769)
         );
  NOR2_X1 U8248 ( .A1(n6655), .A2(n9679), .ZN(n9191) );
  INV_X1 U8249 ( .A(n9191), .ZN(n7047) );
  AOI22_X1 U8250 ( .A1(n9715), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6679), .B2(
        n9714), .ZN(n6657) );
  NAND2_X1 U8251 ( .A1(n9539), .A2(n6721), .ZN(n6656) );
  OAI211_X1 U8252 ( .C1(n9769), .C2(n7047), .A(n6657), .B(n6656), .ZN(n6658)
         );
  AOI21_X1 U8253 ( .B1(n9771), .B2(n9719), .A(n6658), .ZN(n6659) );
  OAI21_X1 U8254 ( .B1(n6660), .B2(n9198), .A(n6659), .ZN(P1_U3284) );
  INV_X1 U8255 ( .A(n7383), .ZN(n6662) );
  OAI222_X1 U8256 ( .A1(n8404), .A2(n6661), .B1(n8400), .B2(n6662), .C1(
        P2_U3152), .C2(n8013), .ZN(P2_U3339) );
  OAI222_X1 U8257 ( .A1(n9462), .A2(n6663), .B1(n9464), .B2(n6662), .C1(n9125), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  AOI21_X1 U8258 ( .B1(n6666), .B2(n6665), .A(n6664), .ZN(n6668) );
  INV_X1 U8259 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9505) );
  AOI22_X1 U8260 ( .A1(n6948), .A2(n9505), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n6951), .ZN(n6667) );
  NOR2_X1 U8261 ( .A1(n6668), .A2(n6667), .ZN(n6950) );
  AOI21_X1 U8262 ( .B1(n6668), .B2(n6667), .A(n6950), .ZN(n6678) );
  INV_X1 U8263 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7236) );
  AOI22_X1 U8264 ( .A1(n6948), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7236), .B2(
        n6951), .ZN(n6672) );
  OAI21_X1 U8265 ( .B1(n6672), .B2(n6671), .A(n6947), .ZN(n6676) );
  NOR2_X1 U8266 ( .A1(n9815), .A2(n6951), .ZN(n6675) );
  INV_X1 U8267 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8268 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7287) );
  OAI21_X1 U8269 ( .B1(n9472), .B2(n6673), .A(n7287), .ZN(n6674) );
  AOI211_X1 U8270 ( .C1(n6676), .C2(n9814), .A(n6675), .B(n6674), .ZN(n6677)
         );
  OAI21_X1 U8271 ( .B1(n6678), .B2(n9817), .A(n6677), .ZN(P2_U3259) );
  INV_X1 U8272 ( .A(n6679), .ZN(n6705) );
  NAND2_X1 U8273 ( .A1(n8884), .A2(n7641), .ZN(n6681) );
  NAND2_X1 U8274 ( .A1(n6721), .A2(n7674), .ZN(n6680) );
  NAND2_X1 U8275 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  XNOR2_X1 U8276 ( .A(n6682), .B(n7680), .ZN(n6855) );
  AND2_X1 U8277 ( .A1(n6721), .A2(n4253), .ZN(n6683) );
  AOI21_X1 U8278 ( .B1(n8884), .B2(n7625), .A(n6683), .ZN(n6856) );
  XNOR2_X1 U8279 ( .A(n6855), .B(n6856), .ZN(n6698) );
  INV_X1 U8280 ( .A(n6684), .ZN(n6685) );
  OR2_X1 U8281 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  NAND2_X1 U8282 ( .A1(n6688), .A2(n6687), .ZN(n8562) );
  NAND2_X1 U8283 ( .A1(n8885), .A2(n4253), .ZN(n6690) );
  NAND2_X1 U8284 ( .A1(n8567), .A2(n7674), .ZN(n6689) );
  NAND2_X1 U8285 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  XNOR2_X1 U8286 ( .A(n6691), .B(n7680), .ZN(n6693) );
  AND2_X1 U8287 ( .A1(n8567), .A2(n4253), .ZN(n6692) );
  AOI21_X1 U8288 ( .B1(n8885), .B2(n7625), .A(n6692), .ZN(n6694) );
  XNOR2_X1 U8289 ( .A(n6693), .B(n6694), .ZN(n8564) );
  INV_X1 U8290 ( .A(n6693), .ZN(n6695) );
  NAND2_X1 U8291 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  NAND2_X1 U8292 ( .A1(n6697), .A2(n6698), .ZN(n6859) );
  OAI21_X1 U8293 ( .B1(n6698), .B2(n6697), .A(n6859), .ZN(n6699) );
  NAND2_X1 U8294 ( .A1(n6699), .A2(n9576), .ZN(n6704) );
  INV_X1 U8295 ( .A(n8883), .ZN(n7014) );
  NAND2_X1 U8296 ( .A1(n8587), .A2(n8885), .ZN(n6701) );
  OAI211_X1 U8297 ( .C1(n7014), .C2(n8590), .A(n6701), .B(n6700), .ZN(n6702)
         );
  AOI21_X1 U8298 ( .B1(n6721), .B2(n9575), .A(n6702), .ZN(n6703) );
  OAI211_X1 U8299 ( .C1(n8483), .C2(n6705), .A(n6704), .B(n6703), .ZN(P1_U3211) );
  AOI22_X1 U8300 ( .A1(n8666), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7384), .B2(
        n6707), .ZN(n6710) );
  NAND2_X1 U8301 ( .A1(n6708), .A2(n7463), .ZN(n6709) );
  NAND2_X1 U8302 ( .A1(n6710), .A2(n6709), .ZN(n9776) );
  NAND2_X1 U8303 ( .A1(n7014), .A2(n9776), .ZN(n8692) );
  NAND2_X1 U8304 ( .A1(n8883), .A2(n7010), .ZN(n7023) );
  NAND2_X1 U8305 ( .A1(n8692), .A2(n7023), .ZN(n8812) );
  XNOR2_X1 U8306 ( .A(n7011), .B(n8812), .ZN(n6711) );
  NAND2_X1 U8307 ( .A1(n6711), .A2(n9707), .ZN(n6720) );
  NAND2_X1 U8308 ( .A1(n7471), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U8309 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  AND2_X1 U8310 ( .A1(n6916), .A2(n6714), .ZN(n7017) );
  NAND2_X1 U8311 ( .A1(n6918), .A2(n7017), .ZN(n6717) );
  NAND2_X1 U8312 ( .A1(n8456), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8313 ( .A1(n8455), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6715) );
  NAND4_X1 U8314 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n8882)
         );
  AOI22_X1 U8315 ( .A1(n9700), .A2(n8884), .B1(n8882), .B2(n9702), .ZN(n6719)
         );
  OR2_X1 U8316 ( .A1(n6723), .A2(n8812), .ZN(n6724) );
  AND2_X1 U8317 ( .A1(n7009), .A2(n6724), .ZN(n9775) );
  INV_X1 U8318 ( .A(n9198), .ZN(n9128) );
  NAND2_X1 U8319 ( .A1(n6725), .A2(n7010), .ZN(n7015) );
  OR2_X1 U8320 ( .A1(n6725), .A2(n7010), .ZN(n6726) );
  AND2_X1 U8321 ( .A1(n7015), .A2(n6726), .ZN(n9779) );
  NAND2_X1 U8322 ( .A1(n9779), .A2(n9698), .ZN(n6728) );
  AOI22_X1 U8323 ( .A1(n9715), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6864), .B2(
        n9714), .ZN(n6727) );
  OAI211_X1 U8324 ( .C1(n7010), .C2(n9717), .A(n6728), .B(n6727), .ZN(n6729)
         );
  AOI21_X1 U8325 ( .B1(n9775), .B2(n9128), .A(n6729), .ZN(n6730) );
  OAI21_X1 U8326 ( .B1(n9715), .B2(n9781), .A(n6730), .ZN(P1_U3283) );
  INV_X1 U8327 ( .A(n6731), .ZN(n6733) );
  NAND2_X1 U8328 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NOR2_X1 U8329 ( .A1(n7819), .A2(n7759), .ZN(n6736) );
  XNOR2_X1 U8330 ( .A(n6763), .B(n7799), .ZN(n6737) );
  NAND2_X1 U8331 ( .A1(n6736), .A2(n6737), .ZN(n6829) );
  INV_X1 U8332 ( .A(n6736), .ZN(n6738) );
  INV_X1 U8333 ( .A(n6737), .ZN(n7818) );
  NAND2_X1 U8334 ( .A1(n6738), .A2(n7818), .ZN(n6739) );
  NAND2_X1 U8335 ( .A1(n6829), .A2(n6739), .ZN(n6742) );
  INV_X1 U8336 ( .A(n6830), .ZN(n6741) );
  AOI211_X1 U8337 ( .C1(n6743), .C2(n6742), .A(n7909), .B(n6741), .ZN(n6750)
         );
  OAI22_X1 U8338 ( .A1(n7924), .A2(n6745), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6744), .ZN(n6749) );
  INV_X1 U8339 ( .A(n6746), .ZN(n6747) );
  OAI22_X1 U8340 ( .A1(n7925), .A2(n6779), .B1(n7886), .B2(n6747), .ZN(n6748)
         );
  OR3_X1 U8341 ( .A1(n6750), .A2(n6749), .A3(n6748), .ZN(P2_U3215) );
  NAND2_X1 U8342 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  NOR2_X1 U8343 ( .A1(n9850), .A2(n6753), .ZN(n6754) );
  NAND2_X1 U8344 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  OR2_X1 U8345 ( .A1(n6757), .A2(n6756), .ZN(n6768) );
  INV_X2 U8346 ( .A(n9927), .ZN(n9912) );
  AOI211_X1 U8347 ( .C1(n9898), .C2(n6763), .A(n6762), .B(n6761), .ZN(n6764)
         );
  OAI21_X1 U8348 ( .B1(n9904), .B2(n6765), .A(n6764), .ZN(n6769) );
  NAND2_X1 U8349 ( .A1(n6769), .A2(n9912), .ZN(n6766) );
  OAI21_X1 U8350 ( .B1(n9912), .B2(n4959), .A(n6766), .ZN(P2_U3472) );
  NAND2_X1 U8351 ( .A1(n6769), .A2(n9943), .ZN(n6770) );
  OAI21_X1 U8352 ( .B1(n9943), .B2(n9351), .A(n6770), .ZN(P2_U3527) );
  INV_X1 U8353 ( .A(n7394), .ZN(n6773) );
  OAI222_X1 U8354 ( .A1(n8404), .A2(n6772), .B1(n8400), .B2(n6773), .C1(n6771), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U8355 ( .A1(n9462), .A2(n6774), .B1(P1_U3084), .B2(n7218), .C1(
        n9464), .C2(n6773), .ZN(P1_U3333) );
  AND2_X1 U8356 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  NAND2_X1 U8357 ( .A1(n6778), .A2(n6777), .ZN(n6781) );
  NAND2_X1 U8358 ( .A1(n7819), .A2(n6779), .ZN(n6780) );
  NAND2_X1 U8359 ( .A1(n6781), .A2(n6780), .ZN(n6871) );
  INV_X1 U8360 ( .A(n6871), .ZN(n6783) );
  NAND2_X1 U8361 ( .A1(n6783), .A2(n6782), .ZN(n6873) );
  NAND2_X1 U8362 ( .A1(n7940), .A2(n7823), .ZN(n6784) );
  OAI22_X1 U8363 ( .A1(n6997), .A2(n8179), .B1(n6896), .B2(n8181), .ZN(n6789)
         );
  XNOR2_X1 U8364 ( .A(n6785), .B(n6786), .ZN(n6787) );
  NOR2_X1 U8365 ( .A1(n6787), .A2(n9842), .ZN(n6788) );
  AOI211_X1 U8366 ( .C1(n7150), .C2(n7054), .A(n6789), .B(n6788), .ZN(n7058)
         );
  AOI21_X1 U8367 ( .B1(n7055), .B2(n6876), .A(n6803), .ZN(n7056) );
  NAND2_X1 U8368 ( .A1(n7056), .A2(n8277), .ZN(n6791) );
  AOI22_X1 U8369 ( .A1(n9848), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n6893), .B2(
        n9834), .ZN(n6790) );
  OAI211_X1 U8370 ( .C1(n6836), .C2(n8281), .A(n6791), .B(n6790), .ZN(n6792)
         );
  AOI21_X1 U8371 ( .B1(n7054), .B2(n7159), .A(n6792), .ZN(n6793) );
  OAI21_X1 U8372 ( .B1(n7058), .B2(n9848), .A(n6793), .ZN(P2_U3287) );
  NAND2_X1 U8373 ( .A1(n6836), .A2(n6846), .ZN(n6794) );
  NAND2_X1 U8374 ( .A1(n7095), .A2(n7088), .ZN(n6796) );
  NAND2_X1 U8375 ( .A1(n6933), .A2(n6796), .ZN(n6801) );
  AOI22_X1 U8376 ( .A1(n4618), .A2(n8268), .B1(n8266), .B2(n7939), .ZN(n6800)
         );
  XNOR2_X1 U8377 ( .A(n6797), .B(n7088), .ZN(n6798) );
  NAND2_X1 U8378 ( .A1(n6798), .A2(n8271), .ZN(n6799) );
  OAI211_X1 U8379 ( .C1(n6801), .C2(n6883), .A(n6800), .B(n6799), .ZN(n9914)
         );
  INV_X1 U8380 ( .A(n9914), .ZN(n6809) );
  INV_X1 U8381 ( .A(n6801), .ZN(n9916) );
  NAND2_X1 U8382 ( .A1(n4473), .A2(n6824), .ZN(n6804) );
  NAND2_X1 U8383 ( .A1(n6937), .A2(n6804), .ZN(n9913) );
  AOI22_X1 U8384 ( .A1(n9848), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n6849), .B2(
        n9834), .ZN(n6806) );
  NAND2_X1 U8385 ( .A1(n8255), .A2(n6824), .ZN(n6805) );
  OAI211_X1 U8386 ( .C1(n9913), .C2(n8062), .A(n6806), .B(n6805), .ZN(n6807)
         );
  AOI21_X1 U8387 ( .B1(n9916), .B2(n7159), .A(n6807), .ZN(n6808) );
  OAI21_X1 U8388 ( .B1(n6809), .B2(n9848), .A(n6808), .ZN(P2_U3286) );
  NAND2_X1 U8389 ( .A1(n6810), .A2(n8808), .ZN(n6811) );
  NAND2_X1 U8390 ( .A1(n6812), .A2(n6811), .ZN(n9766) );
  AND2_X1 U8391 ( .A1(n9673), .A2(n8567), .ZN(n6814) );
  OR2_X1 U8392 ( .A1(n6814), .A2(n6813), .ZN(n9763) );
  AOI22_X1 U8393 ( .A1(n9539), .A2(n8567), .B1(n8568), .B2(n9714), .ZN(n6815)
         );
  OAI21_X1 U8394 ( .B1(n9763), .B2(n8974), .A(n6815), .ZN(n6822) );
  INV_X1 U8395 ( .A(n6816), .ZN(n6817) );
  INV_X1 U8396 ( .A(n8808), .ZN(n8675) );
  XNOR2_X1 U8397 ( .A(n8673), .B(n8675), .ZN(n6820) );
  NAND2_X1 U8398 ( .A1(n9766), .A2(n9537), .ZN(n6819) );
  AOI22_X1 U8399 ( .A1(n9700), .A2(n8886), .B1(n8884), .B2(n9702), .ZN(n6818)
         );
  OAI211_X1 U8400 ( .C1(n9682), .C2(n6820), .A(n6819), .B(n6818), .ZN(n9764)
         );
  MUX2_X1 U8401 ( .A(n9764), .B(P1_REG2_REG_6__SCAN_IN), .S(n9715), .Z(n6821)
         );
  AOI211_X1 U8402 ( .C1(n9699), .C2(n9766), .A(n6822), .B(n6821), .ZN(n6823)
         );
  INV_X1 U8403 ( .A(n6823), .ZN(P1_U3285) );
  XNOR2_X1 U8404 ( .A(n6824), .B(n7799), .ZN(n6825) );
  AND2_X1 U8405 ( .A1(n7938), .A2(n7798), .ZN(n6826) );
  NAND2_X1 U8406 ( .A1(n6825), .A2(n6826), .ZN(n6998) );
  INV_X1 U8407 ( .A(n6825), .ZN(n6996) );
  INV_X1 U8408 ( .A(n6826), .ZN(n6827) );
  NAND2_X1 U8409 ( .A1(n6996), .A2(n6827), .ZN(n6828) );
  AND2_X1 U8410 ( .A1(n6998), .A2(n6828), .ZN(n6845) );
  NAND2_X1 U8411 ( .A1(n6830), .A2(n6829), .ZN(n6835) );
  NOR2_X1 U8412 ( .A1(n6896), .A2(n7759), .ZN(n6831) );
  XNOR2_X1 U8413 ( .A(n7823), .B(n7799), .ZN(n6832) );
  NAND2_X1 U8414 ( .A1(n6831), .A2(n6832), .ZN(n6837) );
  INV_X1 U8415 ( .A(n6831), .ZN(n6833) );
  INV_X1 U8416 ( .A(n6832), .ZN(n6889) );
  NAND2_X1 U8417 ( .A1(n6833), .A2(n6889), .ZN(n6834) );
  AND2_X1 U8418 ( .A1(n6837), .A2(n6834), .ZN(n7816) );
  NAND2_X1 U8419 ( .A1(n6835), .A2(n7816), .ZN(n6888) );
  NAND2_X1 U8420 ( .A1(n7939), .A2(n7798), .ZN(n6840) );
  XNOR2_X1 U8421 ( .A(n6839), .B(n6840), .ZN(n6902) );
  AND2_X1 U8422 ( .A1(n6902), .A2(n6837), .ZN(n6838) );
  INV_X1 U8423 ( .A(n6839), .ZN(n6841) );
  NAND2_X1 U8424 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  AND2_X1 U8425 ( .A1(n6892), .A2(n6842), .ZN(n6844) );
  AND2_X1 U8426 ( .A1(n6845), .A2(n6842), .ZN(n6843) );
  OAI211_X1 U8427 ( .C1(n6845), .C2(n6844), .A(n6999), .B(n7919), .ZN(n6851)
         );
  INV_X1 U8428 ( .A(n7886), .ZN(n7929) );
  OAI22_X1 U8429 ( .A1(n6846), .A2(n7903), .B1(n7904), .B2(n7553), .ZN(n6847)
         );
  AOI211_X1 U8430 ( .C1(n7929), .C2(n6849), .A(n6848), .B(n6847), .ZN(n6850)
         );
  OAI211_X1 U8431 ( .C1(n6802), .C2(n7925), .A(n6851), .B(n6850), .ZN(P2_U3219) );
  NAND2_X1 U8432 ( .A1(n8883), .A2(n4253), .ZN(n6853) );
  NAND2_X1 U8433 ( .A1(n9776), .A2(n8445), .ZN(n6852) );
  NAND2_X1 U8434 ( .A1(n6853), .A2(n6852), .ZN(n6854) );
  XNOR2_X1 U8435 ( .A(n6854), .B(n7680), .ZN(n6904) );
  INV_X1 U8436 ( .A(n6855), .ZN(n6857) );
  NAND2_X1 U8437 ( .A1(n6857), .A2(n6856), .ZN(n6858) );
  AOI22_X1 U8438 ( .A1(n8883), .A2(n7625), .B1(n4253), .B2(n9776), .ZN(n6861)
         );
  INV_X1 U8439 ( .A(n6861), .ZN(n6860) );
  NAND2_X1 U8440 ( .A1(n6906), .A2(n6905), .ZN(n6862) );
  XOR2_X1 U8441 ( .A(n6904), .B(n6862), .Z(n6870) );
  INV_X1 U8442 ( .A(n8590), .ZN(n9573) );
  AOI21_X1 U8443 ( .B1(n9573), .B2(n8882), .A(n6863), .ZN(n6866) );
  NAND2_X1 U8444 ( .A1(n8594), .A2(n6864), .ZN(n6865) );
  OAI211_X1 U8445 ( .C1(n6867), .C2(n8538), .A(n6866), .B(n6865), .ZN(n6868)
         );
  AOI21_X1 U8446 ( .B1(n9776), .B2(n9575), .A(n6868), .ZN(n6869) );
  OAI21_X1 U8447 ( .B1(n6870), .B2(n8596), .A(n6869), .ZN(P1_U3219) );
  NAND2_X1 U8448 ( .A1(n6871), .A2(n6878), .ZN(n6872) );
  NAND2_X1 U8449 ( .A1(n6873), .A2(n6872), .ZN(n6884) );
  INV_X1 U8450 ( .A(n6884), .ZN(n9911) );
  OR2_X1 U8451 ( .A1(n6874), .A2(n9907), .ZN(n6875) );
  NAND2_X1 U8452 ( .A1(n6876), .A2(n6875), .ZN(n9908) );
  AOI22_X1 U8453 ( .A1(n8255), .A2(n7823), .B1(n9834), .B2(n7824), .ZN(n6877)
         );
  OAI21_X1 U8454 ( .B1(n9908), .B2(n8062), .A(n6877), .ZN(n6886) );
  AOI22_X1 U8455 ( .A1(n7941), .A2(n8266), .B1(n8268), .B2(n7939), .ZN(n6882)
         );
  XNOR2_X1 U8456 ( .A(n6879), .B(n6878), .ZN(n6880) );
  NAND2_X1 U8457 ( .A1(n6880), .A2(n8271), .ZN(n6881) );
  OAI211_X1 U8458 ( .C1(n6884), .C2(n6883), .A(n6882), .B(n6881), .ZN(n9909)
         );
  MUX2_X1 U8459 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9909), .S(n8253), .Z(n6885)
         );
  AOI211_X1 U8460 ( .C1(n9911), .C2(n7159), .A(n6886), .B(n6885), .ZN(n6887)
         );
  INV_X1 U8461 ( .A(n6887), .ZN(P2_U3288) );
  INV_X1 U8462 ( .A(n7820), .ZN(n6891) );
  NOR3_X1 U8463 ( .A1(n7898), .A2(n6896), .A3(n6889), .ZN(n6890) );
  AOI21_X1 U8464 ( .B1(n6891), .B2(n7919), .A(n6890), .ZN(n6903) );
  NOR2_X1 U8465 ( .A1(n6892), .A2(n7909), .ZN(n6900) );
  AND2_X1 U8466 ( .A1(n7889), .A2(n7055), .ZN(n6899) );
  INV_X1 U8467 ( .A(n6893), .ZN(n6895) );
  OAI22_X1 U8468 ( .A1(n7886), .A2(n6895), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6894), .ZN(n6898) );
  OAI22_X1 U8469 ( .A1(n6896), .A2(n7903), .B1(n7904), .B2(n6997), .ZN(n6897)
         );
  NOR4_X1 U8470 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6901)
         );
  OAI21_X1 U8471 ( .B1(n6903), .B2(n6902), .A(n6901), .ZN(P2_U3233) );
  NAND2_X1 U8472 ( .A1(n6908), .A2(n7463), .ZN(n6910) );
  AOI22_X1 U8473 ( .A1(n8666), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7384), .B2(
        n9606), .ZN(n6909) );
  NAND2_X1 U8474 ( .A1(n6910), .A2(n6909), .ZN(n7038) );
  NAND2_X1 U8475 ( .A1(n7038), .A2(n8445), .ZN(n6912) );
  NAND2_X1 U8476 ( .A1(n8882), .A2(n4253), .ZN(n6911) );
  NAND2_X1 U8477 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  XNOR2_X1 U8478 ( .A(n6913), .B(n8448), .ZN(n7066) );
  AOI22_X1 U8479 ( .A1(n7038), .A2(n4253), .B1(n8882), .B2(n7625), .ZN(n7065)
         );
  XNOR2_X1 U8480 ( .A(n7066), .B(n7065), .ZN(n7068) );
  XOR2_X1 U8481 ( .A(n7069), .B(n7068), .Z(n6927) );
  INV_X1 U8482 ( .A(n7038), .ZN(n9785) );
  NOR2_X1 U8483 ( .A1(n9785), .A2(n8591), .ZN(n6925) );
  NAND2_X1 U8484 ( .A1(n7471), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6922) );
  INV_X1 U8485 ( .A(n6916), .ZN(n6914) );
  NAND2_X1 U8486 ( .A1(n6914), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7030) );
  INV_X1 U8487 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8488 ( .A1(n6916), .A2(n6915), .ZN(n6917) );
  AND2_X1 U8489 ( .A1(n7030), .A2(n6917), .ZN(n7077) );
  NAND2_X1 U8490 ( .A1(n6918), .A2(n7077), .ZN(n6921) );
  NAND2_X1 U8491 ( .A1(n8456), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U8492 ( .A1(n8455), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6919) );
  NAND4_X1 U8493 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n8881)
         );
  NAND2_X1 U8494 ( .A1(n8587), .A2(n8883), .ZN(n6923) );
  NAND2_X1 U8495 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9616) );
  OAI211_X1 U8496 ( .C1(n9536), .C2(n8590), .A(n6923), .B(n9616), .ZN(n6924)
         );
  AOI211_X1 U8497 ( .C1(n7017), .C2(n8594), .A(n6925), .B(n6924), .ZN(n6926)
         );
  OAI21_X1 U8498 ( .B1(n6927), .B2(n8596), .A(n6926), .ZN(P1_U3229) );
  INV_X1 U8499 ( .A(n7404), .ZN(n6930) );
  OAI222_X1 U8500 ( .A1(n8404), .A2(n6929), .B1(n8400), .B2(n6930), .C1(n6928), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U8501 ( .A1(n9462), .A2(n6932), .B1(n4246), .B2(n6931), .C1(n9464), 
        .C2(n6930), .ZN(P1_U3332) );
  NAND2_X1 U8502 ( .A1(n6933), .A2(n7090), .ZN(n6934) );
  XNOR2_X1 U8503 ( .A(n6934), .B(n7086), .ZN(n7165) );
  XNOR2_X1 U8504 ( .A(n6935), .B(n7086), .ZN(n6936) );
  AOI22_X1 U8505 ( .A1(n7937), .A2(n8268), .B1(n8266), .B2(n7938), .ZN(n7004)
         );
  OAI21_X1 U8506 ( .B1(n6936), .B2(n9842), .A(n7004), .ZN(n7161) );
  NAND2_X1 U8507 ( .A1(n6937), .A2(n7163), .ZN(n6938) );
  NAND2_X1 U8508 ( .A1(n6938), .A2(n9899), .ZN(n6939) );
  NOR2_X1 U8509 ( .A1(n7102), .A2(n6939), .ZN(n7162) );
  NAND2_X1 U8510 ( .A1(n7162), .A2(n8259), .ZN(n6944) );
  INV_X1 U8511 ( .A(n7006), .ZN(n6940) );
  OAI22_X1 U8512 ( .A1(n8253), .A2(n6941), .B1(n6940), .B2(n8250), .ZN(n6942)
         );
  AOI21_X1 U8513 ( .B1(n8255), .B2(n7163), .A(n6942), .ZN(n6943) );
  NAND2_X1 U8514 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  AOI21_X1 U8515 ( .B1(n7161), .B2(n8253), .A(n6945), .ZN(n6946) );
  OAI21_X1 U8516 ( .B1(n8262), .B2(n7165), .A(n6946), .ZN(P2_U3285) );
  OAI21_X1 U8517 ( .B1(n6948), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6947), .ZN(
        n7959) );
  XNOR2_X1 U8518 ( .A(n7959), .B(n7951), .ZN(n6949) );
  NAND2_X1 U8519 ( .A1(n6949), .A2(n5135), .ZN(n7961) );
  OAI21_X1 U8520 ( .B1(n6949), .B2(n5135), .A(n7961), .ZN(n6957) );
  AOI21_X1 U8521 ( .B1(n6951), .B2(n9505), .A(n6950), .ZN(n7950) );
  XNOR2_X1 U8522 ( .A(n7950), .B(n7960), .ZN(n6952) );
  NAND2_X1 U8523 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6952), .ZN(n7952) );
  OAI211_X1 U8524 ( .C1(n6952), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9812), .B(
        n7952), .ZN(n6955) );
  AND2_X1 U8525 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6953) );
  AOI21_X1 U8526 ( .B1(n9820), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n6953), .ZN(
        n6954) );
  OAI211_X1 U8527 ( .C1(n9815), .C2(n7960), .A(n6955), .B(n6954), .ZN(n6956)
         );
  AOI21_X1 U8528 ( .B1(n9814), .B2(n6957), .A(n6956), .ZN(n6958) );
  INV_X1 U8529 ( .A(n6958), .ZN(P2_U3260) );
  INV_X1 U8530 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U8531 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6959) );
  AOI21_X1 U8532 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6959), .ZN(n9953) );
  NOR2_X1 U8533 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6960) );
  AOI21_X1 U8534 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6960), .ZN(n9956) );
  NOR2_X1 U8535 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6961) );
  AOI21_X1 U8536 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6961), .ZN(n9959) );
  NOR2_X1 U8537 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6962) );
  AOI21_X1 U8538 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6962), .ZN(n9962) );
  NOR2_X1 U8539 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6963) );
  AOI21_X1 U8540 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6963), .ZN(n9965) );
  NOR2_X1 U8541 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6970) );
  XOR2_X1 U8542 ( .A(n9604), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n9993) );
  NAND2_X1 U8543 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6968) );
  XOR2_X1 U8544 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9991) );
  NAND2_X1 U8545 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6966) );
  XNOR2_X1 U8546 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n6964), .ZN(n9989) );
  AOI21_X1 U8547 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9944) );
  INV_X1 U8548 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9948) );
  NAND3_X1 U8549 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9946) );
  OAI21_X1 U8550 ( .B1(n9944), .B2(n9948), .A(n9946), .ZN(n9988) );
  NAND2_X1 U8551 ( .A1(n9989), .A2(n9988), .ZN(n6965) );
  NAND2_X1 U8552 ( .A1(n6966), .A2(n6965), .ZN(n9990) );
  NAND2_X1 U8553 ( .A1(n9991), .A2(n9990), .ZN(n6967) );
  NAND2_X1 U8554 ( .A1(n6968), .A2(n6967), .ZN(n9992) );
  NOR2_X1 U8555 ( .A1(n9993), .A2(n9992), .ZN(n6969) );
  NOR2_X1 U8556 ( .A1(n6970), .A2(n6969), .ZN(n6971) );
  NOR2_X1 U8557 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6971), .ZN(n9977) );
  AND2_X1 U8558 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6971), .ZN(n9976) );
  NOR2_X1 U8559 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9976), .ZN(n6972) );
  NOR2_X1 U8560 ( .A1(n9977), .A2(n6972), .ZN(n6973) );
  NAND2_X1 U8561 ( .A1(n6973), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6975) );
  XOR2_X1 U8562 ( .A(n6973), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9975) );
  NAND2_X1 U8563 ( .A1(n9975), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8564 ( .A1(n6975), .A2(n6974), .ZN(n6976) );
  NAND2_X1 U8565 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n6976), .ZN(n6978) );
  XOR2_X1 U8566 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n6976), .Z(n9987) );
  NAND2_X1 U8567 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9987), .ZN(n6977) );
  NAND2_X1 U8568 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  NAND2_X1 U8569 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n6979), .ZN(n6982) );
  XNOR2_X1 U8570 ( .A(n6980), .B(n6979), .ZN(n9986) );
  NAND2_X1 U8571 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9986), .ZN(n6981) );
  NAND2_X1 U8572 ( .A1(n6982), .A2(n6981), .ZN(n6983) );
  AND2_X1 U8573 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6983), .ZN(n6984) );
  INV_X1 U8574 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9985) );
  XNOR2_X1 U8575 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n6983), .ZN(n9984) );
  NOR2_X1 U8576 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NOR2_X1 U8577 ( .A1(n6984), .A2(n9983), .ZN(n9974) );
  NAND2_X1 U8578 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n6985) );
  OAI21_X1 U8579 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6985), .ZN(n9973) );
  NOR2_X1 U8580 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  AOI21_X1 U8581 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9972), .ZN(n9971) );
  NAND2_X1 U8582 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n6986) );
  OAI21_X1 U8583 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6986), .ZN(n9970) );
  NOR2_X1 U8584 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  AOI21_X1 U8585 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9969), .ZN(n9968) );
  NOR2_X1 U8586 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6987) );
  AOI21_X1 U8587 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6987), .ZN(n9967) );
  NAND2_X1 U8588 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  OAI21_X1 U8589 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9966), .ZN(n9964) );
  NAND2_X1 U8590 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  OAI21_X1 U8591 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9963), .ZN(n9961) );
  NAND2_X1 U8592 ( .A1(n9962), .A2(n9961), .ZN(n9960) );
  OAI21_X1 U8593 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9960), .ZN(n9958) );
  NAND2_X1 U8594 ( .A1(n9959), .A2(n9958), .ZN(n9957) );
  OAI21_X1 U8595 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9957), .ZN(n9955) );
  NAND2_X1 U8596 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  OAI21_X1 U8597 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9954), .ZN(n9952) );
  NAND2_X1 U8598 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  NOR2_X1 U8599 ( .A1(n9981), .A2(n9980), .ZN(n6988) );
  NAND2_X1 U8600 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  OAI21_X1 U8601 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6988), .A(n9979), .ZN(
        n6990) );
  XNOR2_X1 U8602 ( .A(n4344), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6989) );
  XNOR2_X1 U8603 ( .A(n6990), .B(n6989), .ZN(ADD_1071_U4) );
  XNOR2_X1 U8604 ( .A(n7163), .B(n7799), .ZN(n7544) );
  NOR2_X1 U8605 ( .A1(n7553), .A2(n7759), .ZN(n6991) );
  NAND2_X1 U8606 ( .A1(n7544), .A2(n6991), .ZN(n7246) );
  INV_X1 U8607 ( .A(n7544), .ZN(n6993) );
  INV_X1 U8608 ( .A(n6991), .ZN(n6992) );
  NAND2_X1 U8609 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  AND2_X1 U8610 ( .A1(n7246), .A2(n6994), .ZN(n7000) );
  INV_X1 U8611 ( .A(n7000), .ZN(n6995) );
  AOI21_X1 U8612 ( .B1(n6999), .B2(n6995), .A(n7909), .ZN(n7002) );
  NOR3_X1 U8613 ( .A1(n7898), .A2(n6997), .A3(n6996), .ZN(n7001) );
  OAI21_X1 U8614 ( .B1(n7002), .B2(n7001), .A(n7248), .ZN(n7008) );
  OAI22_X1 U8615 ( .A1(n7924), .A2(n7004), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7003), .ZN(n7005) );
  AOI21_X1 U8616 ( .B1(n7006), .B2(n7929), .A(n7005), .ZN(n7007) );
  OAI211_X1 U8617 ( .C1(n4469), .C2(n7925), .A(n7008), .B(n7007), .ZN(P2_U3238) );
  OAI21_X1 U8618 ( .B1(n7010), .B2(n7014), .A(n7009), .ZN(n7040) );
  NAND2_X1 U8619 ( .A1(n9785), .A2(n8882), .ZN(n8694) );
  INV_X1 U8620 ( .A(n8882), .ZN(n7037) );
  NAND2_X1 U8621 ( .A1(n7037), .A2(n7038), .ZN(n8693) );
  NAND2_X1 U8622 ( .A1(n8694), .A2(n8693), .ZN(n8811) );
  XOR2_X1 U8623 ( .A(n7040), .B(n8811), .Z(n9791) );
  INV_X1 U8624 ( .A(n9791), .ZN(n7022) );
  NAND2_X1 U8625 ( .A1(n7011), .A2(n8692), .ZN(n7024) );
  NAND2_X1 U8626 ( .A1(n7024), .A2(n7023), .ZN(n7012) );
  XOR2_X1 U8627 ( .A(n8811), .B(n7012), .Z(n7013) );
  OAI222_X1 U8628 ( .A1(n9687), .A2(n9536), .B1(n9685), .B2(n7014), .C1(n9682), 
        .C2(n7013), .ZN(n9788) );
  INV_X1 U8629 ( .A(n7015), .ZN(n7016) );
  OAI21_X1 U8630 ( .B1(n7016), .B2(n9785), .A(n7042), .ZN(n9787) );
  AOI22_X1 U8631 ( .A1(n9715), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7017), .B2(
        n9714), .ZN(n7019) );
  NAND2_X1 U8632 ( .A1(n9539), .A2(n7038), .ZN(n7018) );
  OAI211_X1 U8633 ( .C1(n9787), .C2(n8974), .A(n7019), .B(n7018), .ZN(n7020)
         );
  AOI21_X1 U8634 ( .B1(n9788), .B2(n9719), .A(n7020), .ZN(n7021) );
  OAI21_X1 U8635 ( .B1(n9198), .B2(n7022), .A(n7021), .ZN(P1_U3282) );
  AND2_X1 U8636 ( .A1(n8694), .A2(n7023), .ZN(n8687) );
  NAND2_X1 U8637 ( .A1(n7024), .A2(n8687), .ZN(n7175) );
  NAND2_X1 U8638 ( .A1(n7175), .A2(n8693), .ZN(n7028) );
  NAND2_X1 U8639 ( .A1(n7025), .A2(n7463), .ZN(n7027) );
  AOI22_X1 U8640 ( .A1(n8666), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7384), .B2(
        n9618), .ZN(n7026) );
  NAND2_X1 U8641 ( .A1(n7027), .A2(n7026), .ZN(n7186) );
  OR2_X1 U8642 ( .A1(n7186), .A2(n9536), .ZN(n8609) );
  NAND2_X1 U8643 ( .A1(n7186), .A2(n9536), .ZN(n8688) );
  NAND2_X1 U8644 ( .A1(n8609), .A2(n8688), .ZN(n8689) );
  INV_X1 U8645 ( .A(n8689), .ZN(n8815) );
  XNOR2_X1 U8646 ( .A(n7028), .B(n8815), .ZN(n7036) );
  NAND2_X1 U8647 ( .A1(n7471), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7035) );
  NAND2_X1 U8648 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  AND2_X1 U8649 ( .A1(n7126), .A2(n7031), .ZN(n9538) );
  NAND2_X1 U8650 ( .A1(n6918), .A2(n9538), .ZN(n7034) );
  NAND2_X1 U8651 ( .A1(n8456), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8652 ( .A1(n8455), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7032) );
  NAND4_X1 U8653 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n8880)
         );
  AOI222_X1 U8654 ( .A1(n9707), .A2(n7036), .B1(n8882), .B2(n9700), .C1(n8880), 
        .C2(n9702), .ZN(n7220) );
  NAND2_X1 U8655 ( .A1(n9785), .A2(n7037), .ZN(n7039) );
  AOI22_X1 U8656 ( .A1(n7040), .A2(n7039), .B1(n7038), .B2(n8882), .ZN(n7041)
         );
  NAND2_X1 U8657 ( .A1(n7041), .A2(n8689), .ZN(n7188) );
  OAI21_X1 U8658 ( .B1(n7041), .B2(n8689), .A(n7188), .ZN(n7222) );
  AOI21_X1 U8659 ( .B1(n7042), .B2(n7186), .A(n9786), .ZN(n7043) );
  NAND2_X1 U8660 ( .A1(n7043), .A2(n9541), .ZN(n7219) );
  INV_X1 U8661 ( .A(n7077), .ZN(n7044) );
  OAI22_X1 U8662 ( .A1(n9719), .A2(n5943), .B1(n7044), .B2(n9118), .ZN(n7045)
         );
  AOI21_X1 U8663 ( .B1(n7186), .B2(n9539), .A(n7045), .ZN(n7046) );
  OAI21_X1 U8664 ( .B1(n7219), .B2(n7047), .A(n7046), .ZN(n7048) );
  AOI21_X1 U8665 ( .B1(n7222), .B2(n9128), .A(n7048), .ZN(n7049) );
  OAI21_X1 U8666 ( .B1(n7220), .B2(n9715), .A(n7049), .ZN(P1_U3281) );
  INV_X1 U8667 ( .A(n7415), .ZN(n7052) );
  OAI222_X1 U8668 ( .A1(n8404), .A2(n7051), .B1(n8400), .B2(n7052), .C1(
        P2_U3152), .C2(n7050), .ZN(P2_U3336) );
  OAI222_X1 U8669 ( .A1(n9462), .A2(n7053), .B1(n9464), .B2(n7052), .C1(n8798), 
        .C2(n4246), .ZN(P1_U3331) );
  INV_X1 U8670 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7061) );
  INV_X1 U8671 ( .A(n7054), .ZN(n7059) );
  AOI22_X1 U8672 ( .A1(n7056), .A2(n9899), .B1(n9898), .B2(n7055), .ZN(n7057)
         );
  OAI211_X1 U8673 ( .C1(n7059), .C2(n9880), .A(n7058), .B(n7057), .ZN(n7062)
         );
  NAND2_X1 U8674 ( .A1(n7062), .A2(n9912), .ZN(n7060) );
  OAI21_X1 U8675 ( .B1(n9912), .B2(n7061), .A(n7060), .ZN(P2_U3478) );
  NAND2_X1 U8676 ( .A1(n7062), .A2(n9943), .ZN(n7063) );
  OAI21_X1 U8677 ( .B1(n9943), .B2(n7064), .A(n7063), .ZN(P2_U3529) );
  NAND2_X1 U8678 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  NAND2_X1 U8679 ( .A1(n7186), .A2(n7674), .ZN(n7071) );
  NAND2_X1 U8680 ( .A1(n8881), .A2(n4253), .ZN(n7070) );
  NAND2_X1 U8681 ( .A1(n7071), .A2(n7070), .ZN(n7072) );
  XNOR2_X1 U8682 ( .A(n7072), .B(n7680), .ZN(n7110) );
  AND2_X1 U8683 ( .A1(n8881), .A2(n7625), .ZN(n7073) );
  AOI21_X1 U8684 ( .B1(n7186), .B2(n4253), .A(n7073), .ZN(n7111) );
  XNOR2_X1 U8685 ( .A(n7110), .B(n7111), .ZN(n7108) );
  XOR2_X1 U8686 ( .A(n7109), .B(n7108), .Z(n7079) );
  INV_X1 U8687 ( .A(n8880), .ZN(n8700) );
  NAND2_X1 U8688 ( .A1(n8587), .A2(n8882), .ZN(n7074) );
  NAND2_X1 U8689 ( .A1(n4246), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9629) );
  OAI211_X1 U8690 ( .C1(n8700), .C2(n8590), .A(n7074), .B(n9629), .ZN(n7076)
         );
  NOR2_X1 U8691 ( .A1(n4456), .A2(n8591), .ZN(n7075) );
  AOI211_X1 U8692 ( .C1(n7077), .C2(n8594), .A(n7076), .B(n7075), .ZN(n7078)
         );
  OAI21_X1 U8693 ( .B1(n7079), .B2(n8596), .A(n7078), .ZN(P1_U3215) );
  INV_X1 U8694 ( .A(n7425), .ZN(n7082) );
  NOR2_X1 U8695 ( .A1(n7080), .A2(n4246), .ZN(n8865) );
  AOI21_X1 U8696 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n4244), .A(n8865), .ZN(
        n7081) );
  OAI21_X1 U8697 ( .B1(n7082), .B2(n9464), .A(n7081), .ZN(P1_U3330) );
  NAND2_X1 U8698 ( .A1(n7425), .A2(n8405), .ZN(n7084) );
  OAI211_X1 U8699 ( .C1(n7085), .C2(n8404), .A(n7084), .B(n7083), .ZN(P2_U3335) );
  NAND2_X1 U8700 ( .A1(n7163), .A2(n4618), .ZN(n7089) );
  INV_X1 U8701 ( .A(n7089), .ZN(n7087) );
  OR2_X1 U8702 ( .A1(n7088), .A2(n7092), .ZN(n7094) );
  AND2_X1 U8703 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  OR2_X1 U8704 ( .A1(n7092), .A2(n7091), .ZN(n7093) );
  OAI21_X1 U8705 ( .B1(n7095), .B2(n7094), .A(n7093), .ZN(n7140) );
  XNOR2_X1 U8706 ( .A(n7140), .B(n7139), .ZN(n9926) );
  INV_X1 U8707 ( .A(n9926), .ZN(n7107) );
  AND2_X1 U8708 ( .A1(n7097), .A2(n7096), .ZN(n7099) );
  OAI211_X1 U8709 ( .C1(n7099), .C2(n7139), .A(n7098), .B(n8271), .ZN(n7101)
         );
  NAND2_X1 U8710 ( .A1(n4618), .A2(n8266), .ZN(n7100) );
  OAI211_X1 U8711 ( .C1(n7552), .C2(n8179), .A(n7101), .B(n7100), .ZN(n9923)
         );
  INV_X1 U8712 ( .A(n7556), .ZN(n9920) );
  NAND2_X1 U8713 ( .A1(n7102), .A2(n9920), .ZN(n7151) );
  OAI21_X1 U8714 ( .B1(n7102), .B2(n9920), .A(n7151), .ZN(n9922) );
  AOI22_X1 U8715 ( .A1(n9848), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7549), .B2(
        n9834), .ZN(n7104) );
  NAND2_X1 U8716 ( .A1(n8255), .A2(n7556), .ZN(n7103) );
  OAI211_X1 U8717 ( .C1(n9922), .C2(n8062), .A(n7104), .B(n7103), .ZN(n7105)
         );
  AOI21_X1 U8718 ( .B1(n9923), .B2(n8253), .A(n7105), .ZN(n7106) );
  OAI21_X1 U8719 ( .B1(n8262), .B2(n7107), .A(n7106), .ZN(P2_U3284) );
  INV_X1 U8720 ( .A(n7110), .ZN(n7112) );
  NAND2_X1 U8721 ( .A1(n7113), .A2(n7463), .ZN(n7116) );
  AOI22_X1 U8722 ( .A1(n8666), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7384), .B2(
        n7114), .ZN(n7115) );
  NAND2_X1 U8723 ( .A1(n9540), .A2(n8445), .ZN(n7118) );
  NAND2_X1 U8724 ( .A1(n8880), .A2(n4253), .ZN(n7117) );
  NAND2_X1 U8725 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  XNOR2_X1 U8726 ( .A(n7119), .B(n8448), .ZN(n7200) );
  AND2_X1 U8727 ( .A1(n8880), .A2(n7625), .ZN(n7120) );
  AOI21_X1 U8728 ( .B1(n9540), .B2(n4253), .A(n7120), .ZN(n7201) );
  XNOR2_X1 U8729 ( .A(n7200), .B(n7201), .ZN(n7122) );
  AOI21_X1 U8730 ( .B1(n7121), .B2(n7122), .A(n8596), .ZN(n7123) );
  NAND2_X1 U8731 ( .A1(n7123), .A2(n7205), .ZN(n7138) );
  INV_X1 U8732 ( .A(n7126), .ZN(n7124) );
  NAND2_X1 U8733 ( .A1(n7124), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8734 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  AND2_X1 U8735 ( .A1(n7179), .A2(n7127), .ZN(n7212) );
  NAND2_X1 U8736 ( .A1(n6644), .A2(n7212), .ZN(n7131) );
  NAND2_X1 U8737 ( .A1(n7471), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U8738 ( .A1(n8456), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U8739 ( .A1(n8455), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7128) );
  NAND4_X1 U8740 ( .A1(n7131), .A2(n7130), .A3(n7129), .A4(n7128), .ZN(n9517)
         );
  INV_X1 U8741 ( .A(n9517), .ZN(n9535) );
  NAND2_X1 U8742 ( .A1(n8587), .A2(n8881), .ZN(n7134) );
  INV_X1 U8743 ( .A(n7132), .ZN(n7133) );
  OAI211_X1 U8744 ( .C1(n9535), .C2(n8590), .A(n7134), .B(n7133), .ZN(n7136)
         );
  INV_X1 U8745 ( .A(n9540), .ZN(n9561) );
  NOR2_X1 U8746 ( .A1(n9561), .A2(n8591), .ZN(n7135) );
  AOI211_X1 U8747 ( .C1(n9538), .C2(n8594), .A(n7136), .B(n7135), .ZN(n7137)
         );
  NAND2_X1 U8748 ( .A1(n7138), .A2(n7137), .ZN(P1_U3234) );
  NAND2_X1 U8749 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  OAI22_X1 U8750 ( .A1(n7257), .A2(n8179), .B1(n7258), .B2(n8181), .ZN(n7149)
         );
  NAND2_X1 U8751 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  AOI21_X1 U8752 ( .B1(n7147), .B2(n7146), .A(n9842), .ZN(n7148) );
  AOI211_X1 U8753 ( .C1(n8372), .C2(n7150), .A(n7149), .B(n7148), .ZN(n8376)
         );
  NAND2_X1 U8754 ( .A1(n7151), .A2(n8373), .ZN(n7152) );
  AND2_X1 U8755 ( .A1(n7232), .A2(n7152), .ZN(n8374) );
  NAND2_X1 U8756 ( .A1(n8374), .A2(n8277), .ZN(n7157) );
  INV_X1 U8757 ( .A(n7261), .ZN(n7153) );
  OAI22_X1 U8758 ( .A1(n8253), .A2(n7154), .B1(n7153), .B2(n8250), .ZN(n7155)
         );
  AOI21_X1 U8759 ( .B1(n8373), .B2(n8255), .A(n7155), .ZN(n7156) );
  NAND2_X1 U8760 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  AOI21_X1 U8761 ( .B1(n8372), .B2(n7159), .A(n7158), .ZN(n7160) );
  OAI21_X1 U8762 ( .B1(n8376), .B2(n9848), .A(n7160), .ZN(P2_U3283) );
  AOI211_X1 U8763 ( .C1(n9898), .C2(n7163), .A(n7162), .B(n7161), .ZN(n7164)
         );
  OAI21_X1 U8764 ( .B1(n9904), .B2(n7165), .A(n7164), .ZN(n7167) );
  NAND2_X1 U8765 ( .A1(n7167), .A2(n9943), .ZN(n7166) );
  OAI21_X1 U8766 ( .B1(n9943), .B2(n6322), .A(n7166), .ZN(P2_U3531) );
  NAND2_X1 U8767 ( .A1(n7167), .A2(n9912), .ZN(n7168) );
  OAI21_X1 U8768 ( .B1(n9912), .B2(n5048), .A(n7168), .ZN(P2_U3484) );
  INV_X1 U8769 ( .A(n7313), .ZN(n7197) );
  OAI222_X1 U8770 ( .A1(P2_U3152), .A2(n7170), .B1(n8400), .B2(n7197), .C1(
        n7169), .C2(n8404), .ZN(P2_U3334) );
  NAND2_X1 U8771 ( .A1(n7171), .A2(n7463), .ZN(n7174) );
  AOI22_X1 U8772 ( .A1(n8666), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7384), .B2(
        n7172), .ZN(n7173) );
  NAND2_X1 U8773 ( .A1(n7174), .A2(n7173), .ZN(n7352) );
  OR2_X1 U8774 ( .A1(n7352), .A2(n9535), .ZN(n8703) );
  NAND2_X1 U8775 ( .A1(n7352), .A2(n9535), .ZN(n8702) );
  AND2_X1 U8776 ( .A1(n8688), .A2(n8693), .ZN(n8610) );
  NAND2_X1 U8777 ( .A1(n7175), .A2(n8610), .ZN(n7176) );
  NAND2_X1 U8778 ( .A1(n7176), .A2(n8609), .ZN(n9533) );
  NAND2_X1 U8779 ( .A1(n9540), .A2(n8700), .ZN(n8607) );
  NAND2_X1 U8780 ( .A1(n9533), .A2(n8607), .ZN(n7481) );
  OR2_X1 U8781 ( .A1(n9540), .A2(n8700), .ZN(n7480) );
  NAND2_X1 U8782 ( .A1(n7481), .A2(n7480), .ZN(n7177) );
  XOR2_X1 U8783 ( .A(n8814), .B(n7177), .Z(n7185) );
  NAND2_X1 U8784 ( .A1(n7471), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7184) );
  NAND2_X1 U8785 ( .A1(n7179), .A2(n7178), .ZN(n7180) );
  AND2_X1 U8786 ( .A1(n7357), .A2(n7180), .ZN(n9521) );
  NAND2_X1 U8787 ( .A1(n6644), .A2(n9521), .ZN(n7183) );
  NAND2_X1 U8788 ( .A1(n8456), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U8789 ( .A1(n8455), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7181) );
  NAND4_X1 U8790 ( .A1(n7184), .A2(n7183), .A3(n7182), .A4(n7181), .ZN(n8879)
         );
  AOI222_X1 U8791 ( .A1(n9707), .A2(n7185), .B1(n8879), .B2(n9702), .C1(n8880), 
        .C2(n9700), .ZN(n9556) );
  NAND2_X1 U8792 ( .A1(n7188), .A2(n7187), .ZN(n9531) );
  NAND2_X1 U8793 ( .A1(n9561), .A2(n8700), .ZN(n7189) );
  AOI21_X1 U8794 ( .B1(n8814), .B2(n7191), .A(n7351), .ZN(n9559) );
  NAND2_X1 U8795 ( .A1(n9559), .A2(n9128), .ZN(n7196) );
  INV_X1 U8796 ( .A(n7352), .ZN(n9557) );
  OAI211_X1 U8797 ( .C1(n9542), .C2(n9557), .A(n9523), .B(n9778), .ZN(n9555)
         );
  INV_X1 U8798 ( .A(n9555), .ZN(n7194) );
  AOI22_X1 U8799 ( .A1(n9715), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7212), .B2(
        n9714), .ZN(n7192) );
  OAI21_X1 U8800 ( .B1(n9557), .B2(n9717), .A(n7192), .ZN(n7193) );
  AOI21_X1 U8801 ( .B1(n7194), .B2(n9191), .A(n7193), .ZN(n7195) );
  OAI211_X1 U8802 ( .C1(n9715), .C2(n9556), .A(n7196), .B(n7195), .ZN(P1_U3279) );
  OAI222_X1 U8803 ( .A1(n9462), .A2(n7199), .B1(P1_U3084), .B2(n7198), .C1(
        n9464), .C2(n7197), .ZN(P1_U3329) );
  INV_X1 U8804 ( .A(n7200), .ZN(n7203) );
  INV_X1 U8805 ( .A(n7201), .ZN(n7202) );
  NAND2_X1 U8806 ( .A1(n7203), .A2(n7202), .ZN(n7204) );
  NAND2_X1 U8807 ( .A1(n7352), .A2(n8445), .ZN(n7207) );
  NAND2_X1 U8808 ( .A1(n9517), .A2(n4253), .ZN(n7206) );
  NAND2_X1 U8809 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  XNOR2_X1 U8810 ( .A(n7208), .B(n8448), .ZN(n7565) );
  AND2_X1 U8811 ( .A1(n9517), .A2(n7625), .ZN(n7209) );
  AOI21_X1 U8812 ( .B1(n7352), .B2(n4253), .A(n7209), .ZN(n7563) );
  INV_X1 U8813 ( .A(n7563), .ZN(n7566) );
  XNOR2_X1 U8814 ( .A(n7565), .B(n7566), .ZN(n7210) );
  XNOR2_X1 U8815 ( .A(n7564), .B(n7210), .ZN(n7217) );
  AOI21_X1 U8816 ( .B1(n9573), .B2(n8879), .A(n7211), .ZN(n7214) );
  NAND2_X1 U8817 ( .A1(n8594), .A2(n7212), .ZN(n7213) );
  OAI211_X1 U8818 ( .C1(n8700), .C2(n8538), .A(n7214), .B(n7213), .ZN(n7215)
         );
  AOI21_X1 U8819 ( .B1(n7352), .B2(n9575), .A(n7215), .ZN(n7216) );
  OAI21_X1 U8820 ( .B1(n7217), .B2(n8596), .A(n7216), .ZN(P1_U3222) );
  NAND2_X1 U8821 ( .A1(n8775), .A2(n7218), .ZN(n9730) );
  OAI211_X1 U8822 ( .C1(n4456), .C2(n9784), .A(n7220), .B(n7219), .ZN(n7221)
         );
  AOI21_X1 U8823 ( .B1(n9790), .B2(n7222), .A(n7221), .ZN(n7227) );
  NAND2_X1 U8824 ( .A1(n9809), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7225) );
  OAI21_X1 U8825 ( .B1(n7227), .B2(n9809), .A(n7225), .ZN(P1_U3533) );
  NAND2_X1 U8826 ( .A1(n9792), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7226) );
  OAI21_X1 U8827 ( .B1(n7227), .B2(n9792), .A(n7226), .ZN(P1_U3484) );
  INV_X1 U8828 ( .A(n8373), .ZN(n7264) );
  XNOR2_X1 U8829 ( .A(n7266), .B(n7265), .ZN(n9504) );
  INV_X1 U8830 ( .A(n9504), .ZN(n7241) );
  OAI211_X1 U8831 ( .C1(n7229), .C2(n7265), .A(n8271), .B(n7272), .ZN(n7231)
         );
  NAND2_X1 U8832 ( .A1(n8267), .A2(n8268), .ZN(n7230) );
  OAI211_X1 U8833 ( .C1(n7552), .C2(n8181), .A(n7231), .B(n7230), .ZN(n9502)
         );
  INV_X1 U8834 ( .A(n7295), .ZN(n9500) );
  INV_X1 U8835 ( .A(n7232), .ZN(n7234) );
  INV_X1 U8836 ( .A(n7277), .ZN(n7233) );
  OAI21_X1 U8837 ( .B1(n9500), .B2(n7234), .A(n7233), .ZN(n9501) );
  INV_X1 U8838 ( .A(n7235), .ZN(n7289) );
  OAI22_X1 U8839 ( .A1(n8253), .A2(n7236), .B1(n7289), .B2(n8250), .ZN(n7237)
         );
  AOI21_X1 U8840 ( .B1(n7295), .B2(n8255), .A(n7237), .ZN(n7238) );
  OAI21_X1 U8841 ( .B1(n9501), .B2(n8062), .A(n7238), .ZN(n7239) );
  AOI21_X1 U8842 ( .B1(n9502), .B2(n8253), .A(n7239), .ZN(n7240) );
  OAI21_X1 U8843 ( .B1(n7241), .B2(n8262), .A(n7240), .ZN(P2_U3282) );
  XNOR2_X1 U8844 ( .A(n8373), .B(n7799), .ZN(n7242) );
  NOR2_X1 U8845 ( .A1(n7552), .A2(n7759), .ZN(n7243) );
  NAND2_X1 U8846 ( .A1(n7242), .A2(n7243), .ZN(n7290) );
  INV_X1 U8847 ( .A(n7242), .ZN(n7284) );
  INV_X1 U8848 ( .A(n7243), .ZN(n7244) );
  NAND2_X1 U8849 ( .A1(n7284), .A2(n7244), .ZN(n7245) );
  NAND2_X1 U8850 ( .A1(n7290), .A2(n7245), .ZN(n7255) );
  XNOR2_X1 U8851 ( .A(n7556), .B(n7799), .ZN(n7249) );
  NAND2_X1 U8852 ( .A1(n7937), .A2(n7798), .ZN(n7250) );
  XNOR2_X1 U8853 ( .A(n7249), .B(n7250), .ZN(n7546) );
  AND2_X1 U8854 ( .A1(n7546), .A2(n7246), .ZN(n7247) );
  INV_X1 U8855 ( .A(n7249), .ZN(n7251) );
  NAND2_X1 U8856 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  INV_X1 U8857 ( .A(n7292), .ZN(n7286) );
  AOI211_X1 U8858 ( .C1(n7255), .C2(n7254), .A(n7909), .B(n7286), .ZN(n7256)
         );
  INV_X1 U8859 ( .A(n7256), .ZN(n7263) );
  OAI22_X1 U8860 ( .A1(n7258), .A2(n7903), .B1(n7904), .B2(n7257), .ZN(n7259)
         );
  AOI211_X1 U8861 ( .C1(n7929), .C2(n7261), .A(n7260), .B(n7259), .ZN(n7262)
         );
  OAI211_X1 U8862 ( .C1(n7264), .C2(n7925), .A(n7263), .B(n7262), .ZN(P2_U3236) );
  OAI22_X1 U8863 ( .A1(n7266), .A2(n7265), .B1(n7295), .B2(n7935), .ZN(n7267)
         );
  NAND2_X1 U8864 ( .A1(n7267), .A2(n7271), .ZN(n8027) );
  OAI21_X1 U8865 ( .B1(n7267), .B2(n7271), .A(n8027), .ZN(n8369) );
  INV_X1 U8866 ( .A(n8369), .ZN(n7283) );
  NAND2_X1 U8867 ( .A1(n7272), .A2(n7270), .ZN(n7269) );
  NAND2_X1 U8868 ( .A1(n7269), .A2(n7268), .ZN(n7274) );
  NAND3_X1 U8869 ( .A1(n7272), .A2(n7271), .A3(n7270), .ZN(n7273) );
  NAND3_X1 U8870 ( .A1(n7274), .A2(n8271), .A3(n7273), .ZN(n7276) );
  AOI22_X1 U8871 ( .A1(n8243), .A2(n8268), .B1(n8266), .B2(n7935), .ZN(n7923)
         );
  NAND2_X1 U8872 ( .A1(n7276), .A2(n7923), .ZN(n8367) );
  NAND2_X1 U8873 ( .A1(n7277), .A2(n8366), .ZN(n8276) );
  OAI211_X1 U8874 ( .C1(n7277), .C2(n8366), .A(n8276), .B(n9899), .ZN(n8365)
         );
  AOI22_X1 U8875 ( .A1(n9848), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7928), .B2(
        n9834), .ZN(n7279) );
  NAND2_X1 U8876 ( .A1(n8028), .A2(n8255), .ZN(n7278) );
  OAI211_X1 U8877 ( .C1(n8365), .C2(n7280), .A(n7279), .B(n7278), .ZN(n7281)
         );
  AOI21_X1 U8878 ( .B1(n8367), .B2(n8253), .A(n7281), .ZN(n7282) );
  OAI21_X1 U8879 ( .B1(n7283), .B2(n8262), .A(n7282), .ZN(P2_U3281) );
  NOR3_X1 U8880 ( .A1(n7284), .A2(n7552), .A3(n7898), .ZN(n7285) );
  AOI21_X1 U8881 ( .B1(n7286), .B2(n7919), .A(n7285), .ZN(n7298) );
  XNOR2_X1 U8882 ( .A(n7295), .B(n7799), .ZN(n7707) );
  NAND2_X1 U8883 ( .A1(n7935), .A2(n7798), .ZN(n7708) );
  XNOR2_X1 U8884 ( .A(n7707), .B(n7708), .ZN(n7297) );
  INV_X1 U8885 ( .A(n7552), .ZN(n7936) );
  AOI22_X1 U8886 ( .A1(n7914), .A2(n7936), .B1(n7913), .B2(n8267), .ZN(n7288)
         );
  OAI211_X1 U8887 ( .C1(n7886), .C2(n7289), .A(n7288), .B(n7287), .ZN(n7294)
         );
  AND2_X1 U8888 ( .A1(n7297), .A2(n7290), .ZN(n7291) );
  NOR2_X1 U8889 ( .A1(n7711), .A2(n7909), .ZN(n7293) );
  AOI211_X1 U8890 ( .C1(n7295), .C2(n7889), .A(n7294), .B(n7293), .ZN(n7296)
         );
  OAI21_X1 U8891 ( .B1(n7298), .B2(n7297), .A(n7296), .ZN(P2_U3217) );
  INV_X1 U8892 ( .A(n7436), .ZN(n7302) );
  OAI222_X1 U8893 ( .A1(n8404), .A2(n7300), .B1(n8400), .B2(n7302), .C1(
        P2_U3152), .C2(n7299), .ZN(P2_U3333) );
  OAI222_X1 U8894 ( .A1(n9462), .A2(n7303), .B1(n9464), .B2(n7302), .C1(n7301), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U8895 ( .A(n7447), .ZN(n7306) );
  OAI222_X1 U8896 ( .A1(P2_U3152), .A2(n7305), .B1(n8400), .B2(n7306), .C1(
        n7304), .C2(n8404), .ZN(P2_U3332) );
  OAI222_X1 U8897 ( .A1(n9462), .A2(n7307), .B1(n4246), .B2(n5746), .C1(n9464), 
        .C2(n7306), .ZN(P1_U3327) );
  INV_X1 U8898 ( .A(n7464), .ZN(n7311) );
  AOI21_X1 U8899 ( .B1(n4244), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7308), .ZN(
        n7309) );
  OAI21_X1 U8900 ( .B1(n7311), .B2(n9464), .A(n7309), .ZN(P1_U3326) );
  OAI222_X1 U8901 ( .A1(n8404), .A2(n7312), .B1(n8400), .B2(n7311), .C1(n7310), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U8902 ( .A1(n7313), .A2(n7463), .ZN(n7315) );
  NAND2_X1 U8903 ( .A1(n8666), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7314) );
  INV_X1 U8904 ( .A(n7367), .ZN(n7316) );
  NAND2_X1 U8905 ( .A1(n7316), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7376) );
  INV_X1 U8906 ( .A(n7376), .ZN(n7317) );
  NAND2_X1 U8907 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n7318) );
  INV_X1 U8908 ( .A(n7388), .ZN(n7319) );
  NAND2_X1 U8909 ( .A1(n7319), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7398) );
  INV_X1 U8910 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7397) );
  INV_X1 U8911 ( .A(n7408), .ZN(n7320) );
  NAND2_X1 U8912 ( .A1(n7320), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7418) );
  INV_X1 U8913 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8545) );
  INV_X1 U8914 ( .A(n7429), .ZN(n7321) );
  NAND2_X1 U8915 ( .A1(n7321), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7431) );
  INV_X1 U8916 ( .A(n7431), .ZN(n7322) );
  NAND2_X1 U8917 ( .A1(n7322), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7439) );
  INV_X1 U8918 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U8919 ( .A1(n7431), .A2(n7323), .ZN(n7324) );
  NAND2_X1 U8920 ( .A1(n7439), .A2(n7324), .ZN(n9030) );
  INV_X1 U8921 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U8922 ( .A1(n8455), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7326) );
  NAND2_X1 U8923 ( .A1(n8456), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7325) );
  OAI211_X1 U8924 ( .C1(n5891), .C2(n7327), .A(n7326), .B(n7325), .ZN(n7328)
         );
  INV_X1 U8925 ( .A(n7328), .ZN(n7329) );
  NAND2_X1 U8926 ( .A1(n7331), .A2(n7463), .ZN(n7333) );
  AOI22_X1 U8927 ( .A1(n8940), .A2(n7384), .B1(n8666), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U8928 ( .A1(n7471), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7339) );
  INV_X1 U8929 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8506) );
  INV_X1 U8930 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7334) );
  OAI21_X1 U8931 ( .B1(n7378), .B2(n8506), .A(n7334), .ZN(n7335) );
  AND2_X1 U8932 ( .A1(n7335), .A2(n7388), .ZN(n9116) );
  NAND2_X1 U8933 ( .A1(n6918), .A2(n9116), .ZN(n7338) );
  NAND2_X1 U8934 ( .A1(n8456), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U8935 ( .A1(n8455), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7336) );
  NAND4_X1 U8936 ( .A1(n7339), .A2(n7338), .A3(n7337), .A4(n7336), .ZN(n9137)
         );
  NAND2_X1 U8937 ( .A1(n7340), .A2(n7463), .ZN(n7342) );
  AOI22_X1 U8938 ( .A1(n7384), .A2(n8926), .B1(n8666), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U8939 ( .A1(n7471), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7346) );
  XNOR2_X1 U8940 ( .A(n7378), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U8941 ( .A1(n6918), .A2(n9145), .ZN(n7345) );
  NAND2_X1 U8942 ( .A1(n8456), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7344) );
  NAND2_X1 U8943 ( .A1(n8455), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7343) );
  NAND4_X1 U8944 ( .A1(n7346), .A2(n7345), .A3(n7344), .A4(n7343), .ZN(n8877)
         );
  NAND2_X1 U8945 ( .A1(n7347), .A2(n7463), .ZN(n7350) );
  AOI22_X1 U8946 ( .A1(n8666), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7384), .B2(
        n7348), .ZN(n7349) );
  INV_X1 U8947 ( .A(n8879), .ZN(n9188) );
  OR2_X1 U8948 ( .A1(n9522), .A2(n9188), .ZN(n8710) );
  NAND2_X1 U8949 ( .A1(n9522), .A2(n9188), .ZN(n9184) );
  NAND2_X1 U8950 ( .A1(n8710), .A2(n9184), .ZN(n9511) );
  OAI21_X1 U8951 ( .B1(n8879), .B2(n9522), .A(n9510), .ZN(n9183) );
  NAND2_X1 U8952 ( .A1(n7353), .A2(n7463), .ZN(n7355) );
  AOI22_X1 U8953 ( .A1(n8666), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7384), .B2(
        n8933), .ZN(n7354) );
  NAND2_X1 U8954 ( .A1(n7471), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U8955 ( .A1(n7357), .A2(n7356), .ZN(n7358) );
  AND2_X1 U8956 ( .A1(n7367), .A2(n7358), .ZN(n9192) );
  NAND2_X1 U8957 ( .A1(n6918), .A2(n9192), .ZN(n7361) );
  NAND2_X1 U8958 ( .A1(n8456), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U8959 ( .A1(n8455), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7359) );
  NAND4_X1 U8960 ( .A1(n7362), .A2(n7361), .A3(n7360), .A4(n7359), .ZN(n9518)
         );
  NAND2_X1 U8961 ( .A1(n9286), .A2(n9172), .ZN(n8708) );
  NAND2_X1 U8962 ( .A1(n8711), .A2(n8708), .ZN(n9185) );
  INV_X1 U8963 ( .A(n9286), .ZN(n9195) );
  NAND2_X1 U8964 ( .A1(n7363), .A2(n7463), .ZN(n7365) );
  AOI22_X1 U8965 ( .A1(n8666), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7384), .B2(
        n9633), .ZN(n7364) );
  NAND2_X1 U8966 ( .A1(n7471), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7372) );
  INV_X1 U8967 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U8968 ( .A1(n7367), .A2(n7366), .ZN(n7368) );
  AND2_X1 U8969 ( .A1(n7376), .A2(n7368), .ZN(n9176) );
  NAND2_X1 U8970 ( .A1(n6918), .A2(n9176), .ZN(n7371) );
  NAND2_X1 U8971 ( .A1(n8456), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U8972 ( .A1(n8455), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7369) );
  NAND4_X1 U8973 ( .A1(n7372), .A2(n7371), .A3(n7370), .A4(n7369), .ZN(n8878)
         );
  OR2_X1 U8974 ( .A1(n9279), .A2(n9189), .ZN(n8606) );
  NAND2_X1 U8975 ( .A1(n9279), .A2(n9189), .ZN(n8650) );
  NAND2_X1 U8976 ( .A1(n8606), .A2(n8650), .ZN(n9167) );
  NAND2_X1 U8977 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  NAND2_X1 U8978 ( .A1(n9165), .A2(n4806), .ZN(n9152) );
  NAND2_X1 U8979 ( .A1(n7373), .A2(n7463), .ZN(n7375) );
  AOI22_X1 U8980 ( .A1(n8666), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7384), .B2(
        n8929), .ZN(n7374) );
  NAND2_X1 U8981 ( .A1(n7471), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7382) );
  INV_X1 U8982 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U8983 ( .A1(n7376), .A2(n9433), .ZN(n7377) );
  AND2_X1 U8984 ( .A1(n7378), .A2(n7377), .ZN(n9159) );
  NAND2_X1 U8985 ( .A1(n6918), .A2(n9159), .ZN(n7381) );
  NAND2_X1 U8986 ( .A1(n8456), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U8987 ( .A1(n8455), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7379) );
  NAND4_X1 U8988 ( .A1(n7382), .A2(n7381), .A3(n7380), .A4(n7379), .ZN(n9138)
         );
  OR2_X1 U8989 ( .A1(n9276), .A2(n9171), .ZN(n8721) );
  NAND2_X1 U8990 ( .A1(n9276), .A2(n9171), .ZN(n8719) );
  NAND2_X1 U8991 ( .A1(n8721), .A2(n8719), .ZN(n9153) );
  NAND2_X1 U8992 ( .A1(n9152), .A2(n9153), .ZN(n9151) );
  INV_X1 U8993 ( .A(n9276), .ZN(n9162) );
  NOR2_X1 U8994 ( .A1(n9271), .A2(n9156), .ZN(n9120) );
  AND2_X1 U8995 ( .A1(n9271), .A2(n9156), .ZN(n7485) );
  OR2_X1 U8996 ( .A1(n9266), .A2(n9105), .ZN(n7488) );
  NAND2_X1 U8997 ( .A1(n9266), .A2(n9105), .ZN(n7489) );
  NAND2_X1 U8998 ( .A1(n7488), .A2(n7489), .ZN(n9126) );
  OAI21_X1 U8999 ( .B1(n4460), .B2(n9105), .A(n9262), .ZN(n9101) );
  NAND2_X1 U9000 ( .A1(n7383), .A2(n7463), .ZN(n7387) );
  AOI22_X1 U9001 ( .A1(n8666), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9679), .B2(
        n7384), .ZN(n7386) );
  NAND2_X1 U9002 ( .A1(n7471), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7393) );
  INV_X1 U9003 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U9004 ( .A1(n7388), .A2(n9366), .ZN(n7389) );
  AND2_X1 U9005 ( .A1(n7398), .A2(n7389), .ZN(n9109) );
  NAND2_X1 U9006 ( .A1(n6918), .A2(n9109), .ZN(n7392) );
  NAND2_X1 U9007 ( .A1(n8456), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U9008 ( .A1(n8455), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7390) );
  NAND4_X1 U9009 ( .A1(n7393), .A2(n7392), .A3(n7391), .A4(n7390), .ZN(n9094)
         );
  OR2_X1 U9010 ( .A1(n9259), .A2(n9123), .ZN(n8728) );
  NAND2_X1 U9011 ( .A1(n9259), .A2(n9123), .ZN(n8724) );
  NAND2_X1 U9012 ( .A1(n8728), .A2(n8724), .ZN(n9103) );
  NAND2_X1 U9013 ( .A1(n9101), .A2(n9103), .ZN(n9100) );
  NAND2_X1 U9014 ( .A1(n7394), .A2(n7463), .ZN(n7396) );
  NAND2_X1 U9015 ( .A1(n8666), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U9016 ( .A1(n7471), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9017 ( .A1(n7398), .A2(n7397), .ZN(n7399) );
  AND2_X1 U9018 ( .A1(n7408), .A2(n7399), .ZN(n9088) );
  NAND2_X1 U9019 ( .A1(n6918), .A2(n9088), .ZN(n7402) );
  NAND2_X1 U9020 ( .A1(n8456), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U9021 ( .A1(n8455), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7400) );
  NAND4_X1 U9022 ( .A1(n7403), .A2(n7402), .A3(n7401), .A4(n7400), .ZN(n9076)
         );
  OR2_X1 U9023 ( .A1(n9253), .A2(n9106), .ZN(n8744) );
  NAND2_X1 U9024 ( .A1(n9253), .A2(n9106), .ZN(n8731) );
  NAND2_X1 U9025 ( .A1(n8744), .A2(n8731), .ZN(n9083) );
  NAND2_X1 U9026 ( .A1(n7404), .A2(n7463), .ZN(n7406) );
  NAND2_X1 U9027 ( .A1(n8666), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7405) );
  INV_X1 U9028 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U9029 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  AND2_X1 U9030 ( .A1(n7418), .A2(n7409), .ZN(n9070) );
  NAND2_X1 U9031 ( .A1(n9070), .A2(n6918), .ZN(n7413) );
  NAND2_X1 U9032 ( .A1(n8456), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U9033 ( .A1(n8455), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U9034 ( .A1(n7471), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7410) );
  NAND4_X1 U9035 ( .A1(n7413), .A2(n7412), .A3(n7411), .A4(n7410), .ZN(n9095)
         );
  INV_X1 U9036 ( .A(n9095), .ZN(n7414) );
  OR2_X1 U9037 ( .A1(n9248), .A2(n7414), .ZN(n8624) );
  NAND2_X1 U9038 ( .A1(n9248), .A2(n7414), .ZN(n9051) );
  NAND2_X1 U9039 ( .A1(n8624), .A2(n9051), .ZN(n9068) );
  INV_X1 U9040 ( .A(n9248), .ZN(n9072) );
  INV_X1 U9041 ( .A(n9049), .ZN(n7424) );
  NAND2_X1 U9042 ( .A1(n7415), .A2(n7463), .ZN(n7417) );
  NAND2_X1 U9043 ( .A1(n8666), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U9044 ( .A1(n7418), .A2(n8545), .ZN(n7419) );
  AND2_X1 U9045 ( .A1(n7429), .A2(n7419), .ZN(n9061) );
  NAND2_X1 U9046 ( .A1(n9061), .A2(n6918), .ZN(n7422) );
  AOI22_X1 U9047 ( .A1(n8455), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n8456), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U9048 ( .A1(n7471), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7420) );
  OAI22_X2 U9049 ( .A1(n7424), .A2(n7423), .B1(n7656), .B2(n9064), .ZN(n9035)
         );
  NAND2_X1 U9050 ( .A1(n7425), .A2(n7463), .ZN(n7427) );
  NAND2_X1 U9051 ( .A1(n8666), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7426) );
  INV_X1 U9052 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7434) );
  INV_X1 U9053 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7428) );
  NAND2_X1 U9054 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  NAND2_X1 U9055 ( .A1(n7431), .A2(n7430), .ZN(n9037) );
  OR2_X1 U9056 ( .A1(n9037), .A2(n4249), .ZN(n7433) );
  AOI22_X1 U9057 ( .A1(n7471), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n8456), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n7432) );
  OAI211_X1 U9058 ( .C1(n6283), .C2(n7434), .A(n7433), .B(n7432), .ZN(n9055)
         );
  INV_X1 U9059 ( .A(n9055), .ZN(n9026) );
  NAND2_X1 U9060 ( .A1(n4461), .A2(n9026), .ZN(n7435) );
  NAND2_X1 U9061 ( .A1(n8520), .A2(n8603), .ZN(n7508) );
  NAND2_X1 U9062 ( .A1(n7436), .A2(n7463), .ZN(n7438) );
  NAND2_X1 U9063 ( .A1(n8666), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9064 ( .A1(n7439), .A2(n8484), .ZN(n7440) );
  NAND2_X1 U9065 ( .A1(n7451), .A2(n7440), .ZN(n8482) );
  INV_X1 U9066 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U9067 ( .A1(n8456), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9068 ( .A1(n8455), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7441) );
  OAI211_X1 U9069 ( .C1(n5891), .C2(n7443), .A(n7442), .B(n7441), .ZN(n7444)
         );
  INV_X1 U9070 ( .A(n7444), .ZN(n7445) );
  NAND2_X1 U9071 ( .A1(n8489), .A2(n9027), .ZN(n7460) );
  AND2_X1 U9072 ( .A1(n7508), .A2(n7460), .ZN(n7520) );
  NAND2_X1 U9073 ( .A1(n7447), .A2(n7463), .ZN(n7449) );
  NAND2_X1 U9074 ( .A1(n8666), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7448) );
  INV_X1 U9075 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9076 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  NAND2_X1 U9077 ( .A1(n8580), .A2(n6918), .ZN(n7458) );
  INV_X1 U9078 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U9079 ( .A1(n8456), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U9080 ( .A1(n8455), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7453) );
  OAI211_X1 U9081 ( .C1(n5891), .C2(n7455), .A(n7454), .B(n7453), .ZN(n7456)
         );
  INV_X1 U9082 ( .A(n7456), .ZN(n7457) );
  NOR2_X1 U9083 ( .A1(n9222), .A2(n8875), .ZN(n7462) );
  INV_X1 U9084 ( .A(n7462), .ZN(n7459) );
  INV_X1 U9085 ( .A(n7460), .ZN(n7461) );
  NAND2_X1 U9086 ( .A1(n9227), .A2(n9027), .ZN(n8605) );
  NAND2_X1 U9087 ( .A1(n7527), .A2(n8605), .ZN(n8823) );
  OR2_X1 U9088 ( .A1(n7461), .A2(n8823), .ZN(n7518) );
  NAND2_X1 U9089 ( .A1(n9222), .A2(n8875), .ZN(n8976) );
  NAND2_X1 U9090 ( .A1(n8977), .A2(n8976), .ZN(n7477) );
  NAND2_X1 U9091 ( .A1(n7464), .A2(n7463), .ZN(n7466) );
  NAND2_X1 U9092 ( .A1(n8666), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7465) );
  INV_X1 U9093 ( .A(n7469), .ZN(n7467) );
  NAND2_X1 U9094 ( .A1(n7467), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7494) );
  INV_X1 U9095 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9096 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  NAND2_X1 U9097 ( .A1(n7494), .A2(n7470), .ZN(n7478) );
  INV_X1 U9098 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U9099 ( .A1(n7471), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U9100 ( .A1(n8456), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7472) );
  OAI211_X1 U9101 ( .C1(n9330), .C2(n6283), .A(n7473), .B(n7472), .ZN(n7474)
         );
  INV_X1 U9102 ( .A(n7474), .ZN(n7475) );
  NAND2_X1 U9103 ( .A1(n9217), .A2(n9011), .ZN(n8776) );
  XNOR2_X1 U9104 ( .A(n7477), .B(n8975), .ZN(n9221) );
  OR2_X1 U9105 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  AOI21_X1 U9106 ( .B1(n9217), .B2(n7523), .A(n4459), .ZN(n9218) );
  INV_X1 U9107 ( .A(n9217), .ZN(n8978) );
  INV_X1 U9108 ( .A(n7478), .ZN(n7704) );
  AOI22_X1 U9109 ( .A1(n7704), .A2(n9714), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9715), .ZN(n7479) );
  OAI21_X1 U9110 ( .B1(n8978), .B2(n9717), .A(n7479), .ZN(n7505) );
  AND2_X1 U9111 ( .A1(n8703), .A2(n7480), .ZN(n8612) );
  NAND2_X1 U9112 ( .A1(n7481), .A2(n8612), .ZN(n7482) );
  NAND2_X1 U9113 ( .A1(n7482), .A2(n8702), .ZN(n9514) );
  INV_X1 U9114 ( .A(n9511), .ZN(n9515) );
  NAND2_X1 U9115 ( .A1(n9514), .A2(n9515), .ZN(n9513) );
  INV_X1 U9116 ( .A(n9184), .ZN(n8709) );
  NOR2_X1 U9117 ( .A1(n9185), .A2(n8709), .ZN(n7483) );
  NAND2_X1 U9118 ( .A1(n9154), .A2(n8721), .ZN(n7484) );
  INV_X1 U9119 ( .A(n7485), .ZN(n7486) );
  NAND2_X1 U9120 ( .A1(n7489), .A2(n7486), .ZN(n8725) );
  INV_X1 U9121 ( .A(n9120), .ZN(n7487) );
  NAND2_X1 U9122 ( .A1(n7488), .A2(n7487), .ZN(n8729) );
  NAND2_X1 U9123 ( .A1(n8729), .A2(n7489), .ZN(n8619) );
  INV_X1 U9124 ( .A(n9083), .ZN(n9093) );
  NAND2_X1 U9125 ( .A1(n9092), .A2(n9093), .ZN(n9091) );
  NAND2_X1 U9126 ( .A1(n9091), .A2(n8731), .ZN(n9074) );
  INV_X1 U9127 ( .A(n9068), .ZN(n9075) );
  OR2_X1 U9128 ( .A1(n9064), .A2(n9077), .ZN(n8747) );
  AND2_X1 U9129 ( .A1(n8747), .A2(n9051), .ZN(n8750) );
  OR2_X1 U9130 ( .A1(n9237), .A2(n9026), .ZN(n8801) );
  NAND2_X1 U9131 ( .A1(n9064), .A2(n9077), .ZN(n9040) );
  AND2_X1 U9132 ( .A1(n8801), .A2(n9040), .ZN(n8628) );
  AND2_X1 U9133 ( .A1(n9237), .A2(n9026), .ZN(n8802) );
  XNOR2_X1 U9134 ( .A(n9234), .B(n8603), .ZN(n9024) );
  NAND2_X1 U9135 ( .A1(n9234), .A2(n8603), .ZN(n8602) );
  INV_X1 U9136 ( .A(n8605), .ZN(n8765) );
  INV_X1 U9137 ( .A(n8875), .ZN(n8763) );
  OR2_X1 U9138 ( .A1(n9222), .A2(n8763), .ZN(n7490) );
  NAND2_X1 U9139 ( .A1(n7490), .A2(n7527), .ZN(n8600) );
  NAND2_X1 U9140 ( .A1(n9222), .A2(n8763), .ZN(n8598) );
  AOI211_X1 U9141 ( .C1(n8975), .C2(n7491), .A(n9682), .B(n9006), .ZN(n7503)
         );
  INV_X1 U9142 ( .A(n7494), .ZN(n7492) );
  NAND2_X1 U9143 ( .A1(n7492), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8993) );
  INV_X1 U9144 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U9145 ( .A1(n7494), .A2(n7493), .ZN(n7495) );
  NAND2_X1 U9146 ( .A1(n8993), .A2(n7495), .ZN(n9015) );
  OR2_X1 U9147 ( .A1(n9015), .A2(n4249), .ZN(n7501) );
  INV_X1 U9148 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U9149 ( .A1(n8455), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U9150 ( .A1(n8456), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7496) );
  OAI211_X1 U9151 ( .C1(n5891), .C2(n7498), .A(n7497), .B(n7496), .ZN(n7499)
         );
  INV_X1 U9152 ( .A(n7499), .ZN(n7500) );
  OAI22_X1 U9153 ( .A1(n8986), .A2(n9687), .B1(n8763), .B2(n9685), .ZN(n7502)
         );
  NOR2_X1 U9154 ( .A1(n7503), .A2(n7502), .ZN(n9220) );
  NOR2_X1 U9155 ( .A1(n9220), .A2(n9715), .ZN(n7504) );
  AOI211_X1 U9156 ( .C1(n9218), .C2(n9698), .A(n7505), .B(n7504), .ZN(n7506)
         );
  OAI21_X1 U9157 ( .B1(n9221), .B2(n9198), .A(n7506), .ZN(P1_U3264) );
  OAI222_X1 U9158 ( .A1(P2_U3152), .A2(n4846), .B1(n8400), .B2(n8663), .C1(
        n9415), .C2(n8404), .ZN(P2_U3328) );
  NAND2_X1 U9159 ( .A1(n7507), .A2(n7508), .ZN(n7509) );
  XOR2_X1 U9160 ( .A(n8823), .B(n7509), .Z(n9231) );
  INV_X1 U9161 ( .A(n9028), .ZN(n7510) );
  AOI21_X1 U9162 ( .B1(n9227), .B2(n7510), .A(n7522), .ZN(n9228) );
  INV_X1 U9163 ( .A(n8482), .ZN(n7511) );
  AOI22_X1 U9164 ( .A1(n7511), .A2(n9714), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9715), .ZN(n7512) );
  OAI21_X1 U9165 ( .B1(n8489), .B2(n9717), .A(n7512), .ZN(n7516) );
  XOR2_X1 U9166 ( .A(n8823), .B(n7513), .Z(n7514) );
  AOI222_X1 U9167 ( .A1(n9707), .A2(n7514), .B1(n8875), .B2(n9702), .C1(n9044), 
        .C2(n9700), .ZN(n9230) );
  NOR2_X1 U9168 ( .A1(n9230), .A2(n9715), .ZN(n7515) );
  AOI211_X1 U9169 ( .C1(n9698), .C2(n9228), .A(n7516), .B(n7515), .ZN(n7517)
         );
  OAI21_X1 U9170 ( .B1(n9231), .B2(n9198), .A(n7517), .ZN(P1_U3266) );
  INV_X1 U9171 ( .A(n7518), .ZN(n7519) );
  XNOR2_X1 U9172 ( .A(n9222), .B(n8875), .ZN(n8824) );
  XNOR2_X1 U9173 ( .A(n7521), .B(n8824), .ZN(n9226) );
  INV_X1 U9174 ( .A(n7522), .ZN(n7525) );
  INV_X1 U9175 ( .A(n7523), .ZN(n7524) );
  AOI21_X1 U9176 ( .B1(n9222), .B2(n7525), .A(n7524), .ZN(n9223) );
  AOI22_X1 U9177 ( .A1(n8580), .A2(n9714), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9715), .ZN(n7526) );
  OAI21_X1 U9178 ( .B1(n8762), .B2(n9717), .A(n7526), .ZN(n7532) );
  INV_X1 U9179 ( .A(n7527), .ZN(n8764) );
  NOR2_X1 U9180 ( .A1(n7528), .A2(n8764), .ZN(n7529) );
  XNOR2_X1 U9181 ( .A(n7529), .B(n8824), .ZN(n7530) );
  AOI222_X1 U9182 ( .A1(n9707), .A2(n7530), .B1(n8874), .B2(n9702), .C1(n8876), 
        .C2(n9700), .ZN(n9225) );
  NOR2_X1 U9183 ( .A1(n9225), .A2(n9715), .ZN(n7531) );
  AOI211_X1 U9184 ( .C1(n9698), .C2(n9223), .A(n7532), .B(n7531), .ZN(n7533)
         );
  OAI21_X1 U9185 ( .B1(n9226), .B2(n9198), .A(n7533), .ZN(P1_U3265) );
  INV_X1 U9186 ( .A(n8634), .ZN(n8402) );
  OAI222_X1 U9187 ( .A1(n9462), .A2(n7535), .B1(n7534), .B2(n4246), .C1(n9464), 
        .C2(n8402), .ZN(P1_U3324) );
  XNOR2_X1 U9188 ( .A(n7538), .B(n7537), .ZN(n7543) );
  AOI22_X1 U9189 ( .A1(n7914), .A2(n7947), .B1(n7913), .B2(n7945), .ZN(n7542)
         );
  AOI22_X1 U9190 ( .A1(n7889), .A2(n7540), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7539), .ZN(n7541) );
  OAI211_X1 U9191 ( .C1(n7543), .C2(n7909), .A(n7542), .B(n7541), .ZN(P2_U3239) );
  NAND3_X1 U9192 ( .A1(n7918), .A2(n4618), .A3(n7544), .ZN(n7545) );
  OAI21_X1 U9193 ( .B1(n7248), .B2(n7909), .A(n7545), .ZN(n7548) );
  INV_X1 U9194 ( .A(n7546), .ZN(n7547) );
  NAND2_X1 U9195 ( .A1(n7548), .A2(n7547), .ZN(n7558) );
  INV_X1 U9196 ( .A(n7549), .ZN(n7551) );
  OAI21_X1 U9197 ( .B1(n7886), .B2(n7551), .A(n7550), .ZN(n7555) );
  OAI22_X1 U9198 ( .A1(n7553), .A2(n7903), .B1(n7904), .B2(n7552), .ZN(n7554)
         );
  AOI211_X1 U9199 ( .C1(n7556), .C2(n7889), .A(n7555), .B(n7554), .ZN(n7557)
         );
  OAI211_X1 U9200 ( .C1(n7909), .C2(n7559), .A(n7558), .B(n7557), .ZN(P2_U3226) );
  INV_X1 U9201 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8661) );
  OAI222_X1 U9202 ( .A1(n9462), .A2(n8661), .B1(n9464), .B2(n8663), .C1(n4246), 
        .C2(n7560), .ZN(P1_U3323) );
  AOI22_X1 U9203 ( .A1(n9244), .A2(n8445), .B1(n7641), .B2(n9077), .ZN(n7562)
         );
  XNOR2_X1 U9204 ( .A(n7562), .B(n7680), .ZN(n8543) );
  INV_X1 U9205 ( .A(n7565), .ZN(n7567) );
  NAND2_X1 U9206 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  NAND2_X1 U9207 ( .A1(n7569), .A2(n7568), .ZN(n8530) );
  NAND2_X1 U9208 ( .A1(n9522), .A2(n7674), .ZN(n7571) );
  NAND2_X1 U9209 ( .A1(n8879), .A2(n7641), .ZN(n7570) );
  NAND2_X1 U9210 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  XNOR2_X1 U9211 ( .A(n7572), .B(n7680), .ZN(n7582) );
  NAND2_X1 U9212 ( .A1(n9522), .A2(n4253), .ZN(n7574) );
  NAND2_X1 U9213 ( .A1(n8879), .A2(n7625), .ZN(n7573) );
  NAND2_X1 U9214 ( .A1(n7574), .A2(n7573), .ZN(n7583) );
  NAND2_X1 U9215 ( .A1(n9286), .A2(n4253), .ZN(n7576) );
  NAND2_X1 U9216 ( .A1(n9518), .A2(n7625), .ZN(n7575) );
  NAND2_X1 U9217 ( .A1(n7576), .A2(n7575), .ZN(n8414) );
  INV_X1 U9218 ( .A(n8414), .ZN(n7580) );
  NAND2_X1 U9219 ( .A1(n9286), .A2(n7674), .ZN(n7578) );
  NAND2_X1 U9220 ( .A1(n9518), .A2(n4253), .ZN(n7577) );
  NAND2_X1 U9221 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  XNOR2_X1 U9222 ( .A(n7579), .B(n8448), .ZN(n8412) );
  NOR2_X1 U9223 ( .A1(n7580), .A2(n8412), .ZN(n7587) );
  OR2_X1 U9224 ( .A1(n8531), .A2(n7587), .ZN(n7581) );
  INV_X1 U9225 ( .A(n7582), .ZN(n7585) );
  INV_X1 U9226 ( .A(n7583), .ZN(n7584) );
  NAND2_X1 U9227 ( .A1(n7585), .A2(n7584), .ZN(n8529) );
  AND2_X1 U9228 ( .A1(n8529), .A2(n8414), .ZN(n7586) );
  OR2_X1 U9229 ( .A1(n7587), .A2(n7586), .ZN(n7588) );
  NAND2_X2 U9230 ( .A1(n7589), .A2(n7588), .ZN(n8418) );
  INV_X1 U9231 ( .A(n8412), .ZN(n7590) );
  AND2_X1 U9232 ( .A1(n7590), .A2(n8529), .ZN(n7591) );
  NAND2_X1 U9233 ( .A1(n9279), .A2(n8445), .ZN(n7593) );
  NAND2_X1 U9234 ( .A1(n8878), .A2(n7641), .ZN(n7592) );
  NAND2_X1 U9235 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  XNOR2_X1 U9236 ( .A(n7594), .B(n8448), .ZN(n7606) );
  NAND3_X1 U9237 ( .A1(n8418), .A2(n8410), .A3(n7606), .ZN(n8583) );
  NAND2_X1 U9238 ( .A1(n9279), .A2(n7641), .ZN(n7596) );
  NAND2_X1 U9239 ( .A1(n8878), .A2(n7625), .ZN(n7595) );
  NAND2_X1 U9240 ( .A1(n7596), .A2(n7595), .ZN(n8586) );
  NAND2_X1 U9241 ( .A1(n8583), .A2(n8586), .ZN(n8490) );
  NAND2_X1 U9242 ( .A1(n9276), .A2(n8445), .ZN(n7598) );
  NAND2_X1 U9243 ( .A1(n9138), .A2(n4253), .ZN(n7597) );
  NAND2_X1 U9244 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  XNOR2_X1 U9245 ( .A(n7599), .B(n8448), .ZN(n7601) );
  AND2_X1 U9246 ( .A1(n9138), .A2(n7625), .ZN(n7600) );
  AOI21_X1 U9247 ( .B1(n9276), .B2(n4253), .A(n7600), .ZN(n7602) );
  NAND2_X1 U9248 ( .A1(n7601), .A2(n7602), .ZN(n7610) );
  INV_X1 U9249 ( .A(n7601), .ZN(n7604) );
  INV_X1 U9250 ( .A(n7602), .ZN(n7603) );
  NAND2_X1 U9251 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  NAND2_X1 U9252 ( .A1(n7610), .A2(n7605), .ZN(n8495) );
  INV_X1 U9253 ( .A(n8495), .ZN(n7609) );
  NAND2_X1 U9254 ( .A1(n8410), .A2(n8418), .ZN(n7608) );
  INV_X1 U9255 ( .A(n7606), .ZN(n7607) );
  NAND2_X1 U9256 ( .A1(n7608), .A2(n7607), .ZN(n8492) );
  NAND2_X1 U9257 ( .A1(n9271), .A2(n7674), .ZN(n7612) );
  NAND2_X1 U9258 ( .A1(n8877), .A2(n4253), .ZN(n7611) );
  NAND2_X1 U9259 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  XNOR2_X1 U9260 ( .A(n7613), .B(n7680), .ZN(n7616) );
  AND2_X1 U9261 ( .A1(n8877), .A2(n7614), .ZN(n7615) );
  AOI21_X1 U9262 ( .B1(n9271), .B2(n4253), .A(n7615), .ZN(n7617) );
  XNOR2_X1 U9263 ( .A(n7616), .B(n7617), .ZN(n8504) );
  INV_X1 U9264 ( .A(n7616), .ZN(n7618) );
  NAND2_X1 U9265 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U9266 ( .A1(n9266), .A2(n8445), .ZN(n7621) );
  NAND2_X1 U9267 ( .A1(n9137), .A2(n4253), .ZN(n7620) );
  NAND2_X1 U9268 ( .A1(n7621), .A2(n7620), .ZN(n7622) );
  XNOR2_X1 U9269 ( .A(n7622), .B(n8448), .ZN(n7623) );
  NAND2_X1 U9270 ( .A1(n9266), .A2(n7641), .ZN(n7627) );
  NAND2_X1 U9271 ( .A1(n9137), .A2(n7625), .ZN(n7626) );
  NAND2_X1 U9272 ( .A1(n7627), .A2(n7626), .ZN(n8552) );
  NAND2_X1 U9273 ( .A1(n9259), .A2(n8445), .ZN(n7629) );
  NAND2_X1 U9274 ( .A1(n9094), .A2(n7641), .ZN(n7628) );
  NAND2_X1 U9275 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  XNOR2_X1 U9276 ( .A(n7630), .B(n8448), .ZN(n7632) );
  AND2_X1 U9277 ( .A1(n9094), .A2(n7625), .ZN(n7631) );
  AOI21_X1 U9278 ( .B1(n9259), .B2(n7641), .A(n7631), .ZN(n7633) );
  NAND2_X1 U9279 ( .A1(n7632), .A2(n7633), .ZN(n8522) );
  INV_X1 U9280 ( .A(n7632), .ZN(n7635) );
  INV_X1 U9281 ( .A(n7633), .ZN(n7634) );
  NAND2_X1 U9282 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  AND2_X1 U9283 ( .A1(n8522), .A2(n7636), .ZN(n8436) );
  NAND2_X1 U9284 ( .A1(n9253), .A2(n7674), .ZN(n7638) );
  NAND2_X1 U9285 ( .A1(n9076), .A2(n4253), .ZN(n7637) );
  NAND2_X1 U9286 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  XNOR2_X1 U9287 ( .A(n7639), .B(n8448), .ZN(n7642) );
  AND2_X1 U9288 ( .A1(n9076), .A2(n7625), .ZN(n7640) );
  AOI21_X1 U9289 ( .B1(n9253), .B2(n4253), .A(n7640), .ZN(n7643) );
  NAND2_X1 U9290 ( .A1(n7642), .A2(n7643), .ZN(n7647) );
  INV_X1 U9291 ( .A(n7642), .ZN(n7645) );
  INV_X1 U9292 ( .A(n7643), .ZN(n7644) );
  NAND2_X1 U9293 ( .A1(n7645), .A2(n7644), .ZN(n7646) );
  NAND2_X1 U9294 ( .A1(n7647), .A2(n7646), .ZN(n8521) );
  INV_X1 U9295 ( .A(n7647), .ZN(n7648) );
  AOI22_X1 U9296 ( .A1(n9248), .A2(n4253), .B1(n7625), .B2(n9095), .ZN(n7654)
         );
  NAND2_X1 U9297 ( .A1(n9248), .A2(n7649), .ZN(n7651) );
  NAND2_X1 U9298 ( .A1(n9095), .A2(n7641), .ZN(n7650) );
  NAND2_X1 U9299 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  XNOR2_X1 U9300 ( .A(n7652), .B(n7680), .ZN(n7653) );
  XOR2_X1 U9301 ( .A(n7654), .B(n7653), .Z(n8472) );
  INV_X1 U9302 ( .A(n7653), .ZN(n7655) );
  OAI22_X1 U9303 ( .A1(n9064), .A2(n5711), .B1(n7656), .B2(n8451), .ZN(n7657)
         );
  AOI22_X1 U9304 ( .A1(n9237), .A2(n8445), .B1(n4253), .B2(n9055), .ZN(n7658)
         );
  XOR2_X1 U9305 ( .A(n7680), .B(n7658), .Z(n7661) );
  INV_X1 U9306 ( .A(n7661), .ZN(n7659) );
  NAND2_X1 U9307 ( .A1(n7660), .A2(n7659), .ZN(n8426) );
  OAI22_X1 U9308 ( .A1(n4461), .A2(n5711), .B1(n9026), .B2(n8451), .ZN(n8428)
         );
  NAND2_X1 U9309 ( .A1(n9234), .A2(n8445), .ZN(n7664) );
  NAND2_X1 U9310 ( .A1(n9044), .A2(n7641), .ZN(n7663) );
  NAND2_X1 U9311 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  XNOR2_X1 U9312 ( .A(n7665), .B(n8448), .ZN(n7667) );
  AND2_X1 U9313 ( .A1(n9044), .A2(n7614), .ZN(n7666) );
  AOI21_X1 U9314 ( .B1(n9234), .B2(n4253), .A(n7666), .ZN(n7668) );
  NAND2_X1 U9315 ( .A1(n7667), .A2(n7668), .ZN(n7673) );
  INV_X1 U9316 ( .A(n7667), .ZN(n7670) );
  INV_X1 U9317 ( .A(n7668), .ZN(n7669) );
  NAND2_X1 U9318 ( .A1(n7670), .A2(n7669), .ZN(n7671) );
  AND2_X1 U9319 ( .A1(n7673), .A2(n7671), .ZN(n8512) );
  NAND2_X1 U9320 ( .A1(n9227), .A2(n7674), .ZN(n7676) );
  NAND2_X1 U9321 ( .A1(n8876), .A2(n4253), .ZN(n7675) );
  NAND2_X1 U9322 ( .A1(n7676), .A2(n7675), .ZN(n7677) );
  XNOR2_X1 U9323 ( .A(n7677), .B(n7680), .ZN(n7683) );
  AOI22_X1 U9324 ( .A1(n9227), .A2(n4253), .B1(n7625), .B2(n8876), .ZN(n7684)
         );
  XNOR2_X1 U9325 ( .A(n7683), .B(n7684), .ZN(n8480) );
  NAND2_X1 U9326 ( .A1(n9222), .A2(n8445), .ZN(n7679) );
  NAND2_X1 U9327 ( .A1(n8875), .A2(n7641), .ZN(n7678) );
  NAND2_X1 U9328 ( .A1(n7679), .A2(n7678), .ZN(n7681) );
  XNOR2_X1 U9329 ( .A(n7681), .B(n7680), .ZN(n7689) );
  AND2_X1 U9330 ( .A1(n8875), .A2(n7614), .ZN(n7682) );
  AOI21_X1 U9331 ( .B1(n9222), .B2(n4253), .A(n7682), .ZN(n7687) );
  XNOR2_X1 U9332 ( .A(n7689), .B(n7687), .ZN(n8576) );
  INV_X1 U9333 ( .A(n7683), .ZN(n7685) );
  NAND2_X1 U9334 ( .A1(n7685), .A2(n7684), .ZN(n8573) );
  INV_X1 U9335 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U9336 ( .A1(n7689), .A2(n7688), .ZN(n7699) );
  NAND2_X1 U9337 ( .A1(n9217), .A2(n8445), .ZN(n7691) );
  NAND2_X1 U9338 ( .A1(n8874), .A2(n7641), .ZN(n7690) );
  NAND2_X1 U9339 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  XNOR2_X1 U9340 ( .A(n7692), .B(n8448), .ZN(n7696) );
  INV_X1 U9341 ( .A(n7696), .ZN(n7698) );
  AND2_X1 U9342 ( .A1(n8874), .A2(n7625), .ZN(n7693) );
  AOI21_X1 U9343 ( .B1(n9217), .B2(n7641), .A(n7693), .ZN(n7695) );
  INV_X1 U9344 ( .A(n7695), .ZN(n7697) );
  AOI21_X1 U9345 ( .B1(n7698), .B2(n7697), .A(n8465), .ZN(n7700) );
  AOI21_X1 U9346 ( .B1(n8575), .B2(n7699), .A(n7700), .ZN(n7701) );
  OAI21_X1 U9347 ( .B1(n7701), .B2(n8454), .A(n9576), .ZN(n7706) );
  AOI22_X1 U9348 ( .A1(n8875), .A2(n8587), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        n4246), .ZN(n7702) );
  OAI21_X1 U9349 ( .B1(n8986), .B2(n8590), .A(n7702), .ZN(n7703) );
  AOI21_X1 U9350 ( .B1(n7704), .B2(n8594), .A(n7703), .ZN(n7705) );
  OAI211_X1 U9351 ( .C1(n8978), .C2(n8591), .A(n7706), .B(n7705), .ZN(P1_U3212) );
  NOR2_X1 U9352 ( .A1(n8038), .A2(n7759), .ZN(n7753) );
  XNOR2_X1 U9353 ( .A(n5306), .B(n7799), .ZN(n7752) );
  INV_X1 U9354 ( .A(n7707), .ZN(n7709) );
  NAND2_X1 U9355 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  XNOR2_X1 U9356 ( .A(n8028), .B(n7799), .ZN(n7713) );
  NOR2_X1 U9357 ( .A1(n7851), .A2(n7759), .ZN(n7712) );
  NAND2_X1 U9358 ( .A1(n7920), .A2(n7712), .ZN(n7921) );
  INV_X1 U9359 ( .A(n7713), .ZN(n7714) );
  OR2_X1 U9360 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  NAND2_X1 U9361 ( .A1(n7921), .A2(n7716), .ZN(n7846) );
  INV_X1 U9362 ( .A(n7846), .ZN(n7718) );
  XNOR2_X1 U9363 ( .A(n8360), .B(n7749), .ZN(n7720) );
  NAND2_X1 U9364 ( .A1(n8243), .A2(n7798), .ZN(n7719) );
  XNOR2_X1 U9365 ( .A(n7720), .B(n7719), .ZN(n7849) );
  NAND2_X1 U9366 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  XNOR2_X1 U9367 ( .A(n8355), .B(n7799), .ZN(n7722) );
  NOR2_X1 U9368 ( .A1(n7934), .A2(n7759), .ZN(n7723) );
  NAND2_X1 U9369 ( .A1(n7722), .A2(n7723), .ZN(n7727) );
  INV_X1 U9370 ( .A(n7722), .ZN(n7899) );
  INV_X1 U9371 ( .A(n7723), .ZN(n7724) );
  NAND2_X1 U9372 ( .A1(n7899), .A2(n7724), .ZN(n7725) );
  NAND2_X1 U9373 ( .A1(n7727), .A2(n7725), .ZN(n7858) );
  INV_X1 U9374 ( .A(n7858), .ZN(n7726) );
  NAND2_X1 U9375 ( .A1(n7856), .A2(n7727), .ZN(n7728) );
  XNOR2_X1 U9376 ( .A(n8233), .B(n7749), .ZN(n7731) );
  NAND2_X1 U9377 ( .A1(n8242), .A2(n7798), .ZN(n7729) );
  XNOR2_X1 U9378 ( .A(n7731), .B(n7729), .ZN(n7895) );
  NAND2_X1 U9379 ( .A1(n7728), .A2(n7895), .ZN(n7900) );
  INV_X1 U9380 ( .A(n7729), .ZN(n7730) );
  NAND2_X1 U9381 ( .A1(n7731), .A2(n7730), .ZN(n7732) );
  NAND2_X1 U9382 ( .A1(n7900), .A2(n7732), .ZN(n7791) );
  XNOR2_X1 U9383 ( .A(n8221), .B(n7749), .ZN(n7788) );
  NOR2_X1 U9384 ( .A1(n8033), .A2(n7759), .ZN(n7733) );
  AND2_X1 U9385 ( .A1(n7788), .A2(n7733), .ZN(n7786) );
  INV_X1 U9386 ( .A(n7788), .ZN(n7735) );
  INV_X1 U9387 ( .A(n7733), .ZN(n7734) );
  NAND2_X1 U9388 ( .A1(n7735), .A2(n7734), .ZN(n7790) );
  XNOR2_X1 U9389 ( .A(n8338), .B(n7749), .ZN(n7736) );
  NAND2_X1 U9390 ( .A1(n8224), .A2(n7798), .ZN(n7737) );
  XNOR2_X1 U9391 ( .A(n7736), .B(n7737), .ZN(n7876) );
  INV_X1 U9392 ( .A(n7736), .ZN(n7739) );
  INV_X1 U9393 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U9394 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  XNOR2_X1 U9395 ( .A(n8332), .B(n7799), .ZN(n7743) );
  NAND2_X1 U9396 ( .A1(n8203), .A2(n7798), .ZN(n7741) );
  XNOR2_X1 U9397 ( .A(n7743), .B(n7741), .ZN(n7829) );
  INV_X1 U9398 ( .A(n7741), .ZN(n7742) );
  XNOR2_X1 U9399 ( .A(n8327), .B(n7749), .ZN(n7745) );
  NAND2_X1 U9400 ( .A1(n8195), .A2(n7798), .ZN(n7744) );
  NAND2_X1 U9401 ( .A1(n7891), .A2(n7744), .ZN(n7894) );
  INV_X1 U9402 ( .A(n7745), .ZN(n7746) );
  OR2_X1 U9403 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  NAND2_X1 U9404 ( .A1(n7894), .A2(n7748), .ZN(n7751) );
  XNOR2_X1 U9405 ( .A(n8322), .B(n7749), .ZN(n7750) );
  NOR2_X1 U9406 ( .A1(n7751), .A2(n7750), .ZN(n7776) );
  NAND2_X1 U9407 ( .A1(n7751), .A2(n7750), .ZN(n7777) );
  NOR2_X1 U9408 ( .A1(n8180), .A2(n7759), .ZN(n7779) );
  NAND2_X1 U9409 ( .A1(n7777), .A2(n7779), .ZN(n7864) );
  INV_X1 U9410 ( .A(n7752), .ZN(n7866) );
  INV_X1 U9411 ( .A(n7753), .ZN(n7868) );
  XOR2_X1 U9412 ( .A(n7799), .B(n8315), .Z(n7755) );
  INV_X1 U9413 ( .A(n7755), .ZN(n7839) );
  INV_X1 U9414 ( .A(n7841), .ZN(n7756) );
  NAND2_X1 U9415 ( .A1(n8041), .A2(n7798), .ZN(n7838) );
  XNOR2_X1 U9416 ( .A(n8310), .B(n7799), .ZN(n7767) );
  NOR2_X1 U9417 ( .A1(n8043), .A2(n7759), .ZN(n7757) );
  NAND2_X1 U9418 ( .A1(n7767), .A2(n7757), .ZN(n7758) );
  OAI21_X1 U9419 ( .B1(n7767), .B2(n7757), .A(n7758), .ZN(n7911) );
  INV_X1 U9420 ( .A(n7758), .ZN(n7765) );
  XNOR2_X1 U9421 ( .A(n8303), .B(n7799), .ZN(n7760) );
  NOR2_X1 U9422 ( .A1(n8108), .A2(n7759), .ZN(n7761) );
  NAND2_X1 U9423 ( .A1(n7760), .A2(n7761), .ZN(n7809) );
  INV_X1 U9424 ( .A(n7760), .ZN(n7763) );
  INV_X1 U9425 ( .A(n7761), .ZN(n7762) );
  NAND2_X1 U9426 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  AND2_X1 U9427 ( .A1(n7809), .A2(n7764), .ZN(n7766) );
  INV_X1 U9428 ( .A(n7808), .ZN(n7802) );
  NOR2_X1 U9429 ( .A1(n7898), .A2(n8043), .ZN(n7768) );
  OAI22_X1 U9430 ( .A1(n7886), .A2(n8088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7770), .ZN(n7773) );
  OAI22_X1 U9431 ( .A1(n8043), .A2(n7903), .B1(n7904), .B2(n7771), .ZN(n7772)
         );
  AOI211_X1 U9432 ( .C1(n8303), .C2(n7889), .A(n7773), .B(n7772), .ZN(n7774)
         );
  OAI21_X1 U9433 ( .B1(n7802), .B2(n7775), .A(n7774), .ZN(P2_U3216) );
  INV_X1 U9434 ( .A(n7776), .ZN(n7865) );
  AND2_X1 U9435 ( .A1(n7865), .A2(n7777), .ZN(n7778) );
  NOR3_X1 U9436 ( .A1(n7778), .A2(n8180), .A3(n7898), .ZN(n7785) );
  INV_X1 U9437 ( .A(n7778), .ZN(n7780) );
  NOR3_X1 U9438 ( .A1(n7780), .A2(n7779), .A3(n7909), .ZN(n7784) );
  INV_X1 U9439 ( .A(n8322), .ZN(n8157) );
  AOI22_X1 U9440 ( .A1(n7929), .A2(n8155), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7782) );
  AOI22_X1 U9441 ( .A1(n7914), .A2(n8195), .B1(n7913), .B2(n8162), .ZN(n7781)
         );
  OAI211_X1 U9442 ( .C1(n8157), .C2(n7925), .A(n7782), .B(n7781), .ZN(n7783)
         );
  OR3_X1 U9443 ( .A1(n7785), .A2(n7784), .A3(n7783), .ZN(P2_U3218) );
  INV_X1 U9444 ( .A(n7790), .ZN(n7787) );
  NOR3_X1 U9445 ( .A1(n7787), .A2(n7786), .A3(n7909), .ZN(n7793) );
  INV_X1 U9446 ( .A(n8033), .ZN(n8236) );
  NAND3_X1 U9447 ( .A1(n7788), .A2(n7918), .A3(n8236), .ZN(n7789) );
  OAI21_X1 U9448 ( .B1(n7790), .B2(n7909), .A(n7789), .ZN(n7792) );
  MUX2_X1 U9449 ( .A(n7793), .B(n7792), .S(n7791), .Z(n7797) );
  AOI22_X1 U9450 ( .A1(n7929), .A2(n8219), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n7795) );
  AOI22_X1 U9451 ( .A1(n7914), .A2(n8242), .B1(n7913), .B2(n8224), .ZN(n7794)
         );
  OAI211_X1 U9452 ( .C1(n8221), .C2(n7925), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OR2_X1 U9453 ( .A1(n7797), .A2(n7796), .ZN(P2_U3221) );
  NAND2_X1 U9454 ( .A1(n8095), .A2(n7798), .ZN(n7800) );
  XNOR2_X1 U9455 ( .A(n7800), .B(n7799), .ZN(n7801) );
  XNOR2_X1 U9456 ( .A(n8298), .B(n7801), .ZN(n7807) );
  INV_X1 U9457 ( .A(n7807), .ZN(n7811) );
  NAND2_X1 U9458 ( .A1(n7802), .A2(n4812), .ZN(n7815) );
  INV_X1 U9459 ( .A(n8077), .ZN(n7804) );
  OAI22_X1 U9460 ( .A1(n7886), .A2(n7804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7803), .ZN(n7806) );
  OAI22_X1 U9461 ( .A1(n8108), .A2(n7903), .B1(n7904), .B2(n7933), .ZN(n7805)
         );
  AOI211_X1 U9462 ( .C1(n8298), .C2(n7889), .A(n7806), .B(n7805), .ZN(n7814)
         );
  NAND4_X1 U9463 ( .A1(n7808), .A2(n7919), .A3(n7809), .A4(n7807), .ZN(n7813)
         );
  INV_X1 U9464 ( .A(n7809), .ZN(n7810) );
  NAND3_X1 U9465 ( .A1(n7811), .A2(n7810), .A3(n7919), .ZN(n7812) );
  INV_X1 U9466 ( .A(n7816), .ZN(n7817) );
  AOI21_X1 U9467 ( .B1(n6830), .B2(n7817), .A(n7909), .ZN(n7822) );
  NOR3_X1 U9468 ( .A1(n7898), .A2(n7819), .A3(n7818), .ZN(n7821) );
  OAI21_X1 U9469 ( .B1(n7822), .B2(n7821), .A(n7820), .ZN(n7828) );
  AOI22_X1 U9470 ( .A1(n7913), .A2(n7939), .B1(n7823), .B2(n7889), .ZN(n7827)
         );
  AOI22_X1 U9471 ( .A1(n7929), .A2(n7824), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7826) );
  NAND2_X1 U9472 ( .A1(n7914), .A2(n7941), .ZN(n7825) );
  NAND4_X1 U9473 ( .A1(n7828), .A2(n7827), .A3(n7826), .A4(n7825), .ZN(
        P2_U3223) );
  XNOR2_X1 U9474 ( .A(n7830), .B(n7829), .ZN(n7837) );
  INV_X1 U9475 ( .A(n8192), .ZN(n7832) );
  OAI22_X1 U9476 ( .A1(n7886), .A2(n7832), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7831), .ZN(n7835) );
  OAI22_X1 U9477 ( .A1(n7833), .A2(n7903), .B1(n7904), .B2(n7890), .ZN(n7834)
         );
  AOI211_X1 U9478 ( .C1(n8332), .C2(n7889), .A(n7835), .B(n7834), .ZN(n7836)
         );
  OAI21_X1 U9479 ( .B1(n7837), .B2(n7909), .A(n7836), .ZN(P2_U3225) );
  XNOR2_X1 U9480 ( .A(n7839), .B(n7838), .ZN(n7840) );
  XNOR2_X1 U9481 ( .A(n7841), .B(n7840), .ZN(n7845) );
  INV_X1 U9482 ( .A(n8043), .ZN(n8094) );
  AOI22_X1 U9483 ( .A1(n8094), .A2(n8268), .B1(n8266), .B2(n8162), .ZN(n8123)
         );
  OAI22_X1 U9484 ( .A1(n8123), .A2(n7924), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9346), .ZN(n7842) );
  AOI21_X1 U9485 ( .B1(n8126), .B2(n7929), .A(n7842), .ZN(n7844) );
  NAND2_X1 U9486 ( .A1(n8315), .A2(n7889), .ZN(n7843) );
  OAI211_X1 U9487 ( .C1(n7845), .C2(n7909), .A(n7844), .B(n7843), .ZN(P2_U3227) );
  INV_X1 U9488 ( .A(n7847), .ZN(n7848) );
  AOI21_X1 U9489 ( .B1(n7849), .B2(n7846), .A(n7848), .ZN(n7855) );
  INV_X1 U9490 ( .A(n8278), .ZN(n7850) );
  OAI22_X1 U9491 ( .A1(n7886), .A2(n7850), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7956), .ZN(n7853) );
  OAI22_X1 U9492 ( .A1(n7851), .A2(n7903), .B1(n7904), .B2(n7934), .ZN(n7852)
         );
  AOI211_X1 U9493 ( .C1(n8360), .C2(n7889), .A(n7853), .B(n7852), .ZN(n7854)
         );
  OAI21_X1 U9494 ( .B1(n7855), .B2(n7909), .A(n7854), .ZN(P2_U3228) );
  INV_X1 U9495 ( .A(n7897), .ZN(n7857) );
  AOI211_X1 U9496 ( .C1(n7859), .C2(n7858), .A(n7909), .B(n7857), .ZN(n7863)
         );
  AOI22_X1 U9497 ( .A1(n7929), .A2(n8249), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7861) );
  AOI22_X1 U9498 ( .A1(n7913), .A2(n8242), .B1(n7914), .B2(n8243), .ZN(n7860)
         );
  OAI211_X1 U9499 ( .C1(n4489), .C2(n7925), .A(n7861), .B(n7860), .ZN(n7862)
         );
  OR2_X1 U9500 ( .A1(n7863), .A2(n7862), .ZN(P2_U3230) );
  NAND2_X1 U9501 ( .A1(n7865), .A2(n7864), .ZN(n7867) );
  XNOR2_X1 U9502 ( .A(n7867), .B(n7866), .ZN(n7869) );
  NAND3_X1 U9503 ( .A1(n7869), .A2(n7919), .A3(n7868), .ZN(n7875) );
  INV_X1 U9504 ( .A(n7869), .ZN(n7870) );
  NAND3_X1 U9505 ( .A1(n7870), .A2(n7918), .A3(n8162), .ZN(n7874) );
  OAI22_X1 U9506 ( .A1(n7886), .A2(n8135), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9403), .ZN(n7872) );
  OAI22_X1 U9507 ( .A1(n8180), .A2(n7903), .B1(n7904), .B2(n8144), .ZN(n7871)
         );
  AOI211_X1 U9508 ( .C1(n5306), .C2(n7889), .A(n7872), .B(n7871), .ZN(n7873)
         );
  NAND3_X1 U9509 ( .A1(n7875), .A2(n7874), .A3(n7873), .ZN(P2_U3231) );
  XNOR2_X1 U9510 ( .A(n7877), .B(n7876), .ZN(n7883) );
  INV_X1 U9511 ( .A(n8209), .ZN(n7879) );
  OAI22_X1 U9512 ( .A1(n7886), .A2(n7879), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7878), .ZN(n7881) );
  OAI22_X1 U9513 ( .A1(n8182), .A2(n7904), .B1(n7903), .B2(n8033), .ZN(n7880)
         );
  AOI211_X1 U9514 ( .C1(n8338), .C2(n7889), .A(n7881), .B(n7880), .ZN(n7882)
         );
  OAI21_X1 U9515 ( .B1(n7883), .B2(n7909), .A(n7882), .ZN(P2_U3235) );
  INV_X1 U9516 ( .A(n8170), .ZN(n7885) );
  OAI22_X1 U9517 ( .A1(n7886), .A2(n7885), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7884), .ZN(n7888) );
  OAI22_X1 U9518 ( .A1(n8182), .A2(n7903), .B1(n7904), .B2(n8180), .ZN(n7887)
         );
  AOI211_X1 U9519 ( .C1(n8327), .C2(n7889), .A(n7888), .B(n7887), .ZN(n7893)
         );
  OR3_X1 U9520 ( .A1(n7891), .A2(n7890), .A3(n7898), .ZN(n7892) );
  OAI211_X1 U9521 ( .C1(n7894), .C2(n7909), .A(n7893), .B(n7892), .ZN(P2_U3237) );
  INV_X1 U9522 ( .A(n7895), .ZN(n7896) );
  AOI21_X1 U9523 ( .B1(n7897), .B2(n7896), .A(n7909), .ZN(n7902) );
  NOR3_X1 U9524 ( .A1(n7899), .A2(n7934), .A3(n7898), .ZN(n7901) );
  OAI21_X1 U9525 ( .B1(n7902), .B2(n7901), .A(n7900), .ZN(n7907) );
  AND2_X1 U9526 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7988) );
  OAI22_X1 U9527 ( .A1(n8033), .A2(n7904), .B1(n7903), .B2(n7934), .ZN(n7905)
         );
  AOI211_X1 U9528 ( .C1(n7929), .C2(n8231), .A(n7988), .B(n7905), .ZN(n7906)
         );
  OAI211_X1 U9529 ( .C1(n8233), .C2(n7925), .A(n7907), .B(n7906), .ZN(P2_U3240) );
  INV_X1 U9530 ( .A(n7912), .ZN(n8111) );
  AOI22_X1 U9531 ( .A1(n7929), .A2(n8111), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n7916) );
  AOI22_X1 U9532 ( .A1(n7914), .A2(n8041), .B1(n7913), .B2(n8068), .ZN(n7915)
         );
  OAI211_X1 U9533 ( .C1(n8114), .C2(n7925), .A(n7916), .B(n7915), .ZN(n7917)
         );
  AOI22_X1 U9534 ( .A1(n7920), .A2(n7919), .B1(n7918), .B2(n8267), .ZN(n7932)
         );
  INV_X1 U9535 ( .A(n7921), .ZN(n7931) );
  OAI22_X1 U9536 ( .A1(n7924), .A2(n7923), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7922), .ZN(n7927) );
  NOR2_X1 U9537 ( .A1(n8366), .A2(n7925), .ZN(n7926) );
  AOI211_X1 U9538 ( .C1(n7929), .C2(n7928), .A(n7927), .B(n7926), .ZN(n7930)
         );
  OAI21_X1 U9539 ( .B1(n7932), .B2(n7931), .A(n7930), .ZN(P2_U3243) );
  MUX2_X1 U9540 ( .A(n8053), .B(P2_DATAO_REG_30__SCAN_IN), .S(n7948), .Z(
        P2_U3582) );
  INV_X1 U9541 ( .A(n7933), .ZN(n8069) );
  MUX2_X1 U9542 ( .A(n8069), .B(P2_DATAO_REG_29__SCAN_IN), .S(n7948), .Z(
        P2_U3581) );
  MUX2_X1 U9543 ( .A(n8095), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7948), .Z(
        P2_U3580) );
  MUX2_X1 U9544 ( .A(n8068), .B(P2_DATAO_REG_27__SCAN_IN), .S(n7948), .Z(
        P2_U3579) );
  MUX2_X1 U9545 ( .A(n8094), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7948), .Z(
        P2_U3578) );
  MUX2_X1 U9546 ( .A(n8041), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7948), .Z(
        P2_U3577) );
  MUX2_X1 U9547 ( .A(n8162), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7948), .Z(
        P2_U3576) );
  INV_X1 U9548 ( .A(n8180), .ZN(n8036) );
  MUX2_X1 U9549 ( .A(n8036), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7948), .Z(
        P2_U3575) );
  MUX2_X1 U9550 ( .A(n8195), .B(P2_DATAO_REG_22__SCAN_IN), .S(n7948), .Z(
        P2_U3574) );
  MUX2_X1 U9551 ( .A(n8203), .B(P2_DATAO_REG_21__SCAN_IN), .S(n7948), .Z(
        P2_U3573) );
  MUX2_X1 U9552 ( .A(n8224), .B(P2_DATAO_REG_20__SCAN_IN), .S(n7948), .Z(
        P2_U3572) );
  MUX2_X1 U9553 ( .A(n8236), .B(P2_DATAO_REG_19__SCAN_IN), .S(n7948), .Z(
        P2_U3571) );
  MUX2_X1 U9554 ( .A(n8242), .B(P2_DATAO_REG_18__SCAN_IN), .S(n7948), .Z(
        P2_U3570) );
  MUX2_X1 U9555 ( .A(n8269), .B(P2_DATAO_REG_17__SCAN_IN), .S(n7948), .Z(
        P2_U3569) );
  MUX2_X1 U9556 ( .A(n8243), .B(P2_DATAO_REG_16__SCAN_IN), .S(n7948), .Z(
        P2_U3568) );
  MUX2_X1 U9557 ( .A(n8267), .B(P2_DATAO_REG_15__SCAN_IN), .S(n7948), .Z(
        P2_U3567) );
  MUX2_X1 U9558 ( .A(n7935), .B(P2_DATAO_REG_14__SCAN_IN), .S(n7948), .Z(
        P2_U3566) );
  MUX2_X1 U9559 ( .A(n7936), .B(P2_DATAO_REG_13__SCAN_IN), .S(n7948), .Z(
        P2_U3565) );
  MUX2_X1 U9560 ( .A(n7937), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7948), .Z(
        P2_U3564) );
  MUX2_X1 U9561 ( .A(n4618), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7948), .Z(
        P2_U3563) );
  MUX2_X1 U9562 ( .A(n7938), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7948), .Z(
        P2_U3562) );
  MUX2_X1 U9563 ( .A(n7939), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7948), .Z(
        P2_U3561) );
  MUX2_X1 U9564 ( .A(n7940), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7948), .Z(
        P2_U3560) );
  MUX2_X1 U9565 ( .A(n7941), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7948), .Z(
        P2_U3559) );
  MUX2_X1 U9566 ( .A(n7942), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7948), .Z(
        P2_U3558) );
  MUX2_X1 U9567 ( .A(n7943), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7948), .Z(
        P2_U3557) );
  MUX2_X1 U9568 ( .A(n7944), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7948), .Z(
        P2_U3556) );
  MUX2_X1 U9569 ( .A(n7945), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7948), .Z(
        P2_U3555) );
  MUX2_X1 U9570 ( .A(n7946), .B(P2_DATAO_REG_2__SCAN_IN), .S(n7948), .Z(
        P2_U3554) );
  MUX2_X1 U9571 ( .A(n7947), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7948), .Z(
        P2_U3553) );
  MUX2_X1 U9572 ( .A(n7949), .B(P2_DATAO_REG_0__SCAN_IN), .S(n7948), .Z(
        P2_U3552) );
  NAND2_X1 U9573 ( .A1(n7951), .A2(n7950), .ZN(n7953) );
  NAND2_X1 U9574 ( .A1(n7953), .A2(n7952), .ZN(n7955) );
  XNOR2_X1 U9575 ( .A(n7976), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7954) );
  NOR2_X1 U9576 ( .A1(n7954), .A2(n7955), .ZN(n7977) );
  AOI21_X1 U9577 ( .B1(n7955), .B2(n7954), .A(n7977), .ZN(n7969) );
  NOR2_X1 U9578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7956), .ZN(n7957) );
  AOI21_X1 U9579 ( .B1(n9820), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7957), .ZN(
        n7958) );
  INV_X1 U9580 ( .A(n7958), .ZN(n7967) );
  NAND2_X1 U9581 ( .A1(n7960), .A2(n7959), .ZN(n7962) );
  NAND2_X1 U9582 ( .A1(n7962), .A2(n7961), .ZN(n7965) );
  NAND2_X1 U9583 ( .A1(n7976), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7963) );
  OAI21_X1 U9584 ( .B1(n7976), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7963), .ZN(
        n7964) );
  NOR2_X1 U9585 ( .A1(n7964), .A2(n7965), .ZN(n7970) );
  AOI211_X1 U9586 ( .C1(n7965), .C2(n7964), .A(n7970), .B(n9483), .ZN(n7966)
         );
  AOI211_X1 U9587 ( .C1(n9489), .C2(n7976), .A(n7967), .B(n7966), .ZN(n7968)
         );
  OAI21_X1 U9588 ( .B1(n7969), .B2(n9817), .A(n7968), .ZN(P2_U3261) );
  NAND2_X1 U9589 ( .A1(n7986), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7971) );
  OAI21_X1 U9590 ( .B1(n7986), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7971), .ZN(
        n7972) );
  AOI211_X1 U9591 ( .C1(n7973), .C2(n7972), .A(n7985), .B(n9483), .ZN(n7984)
         );
  NOR2_X1 U9592 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7974), .ZN(n7975) );
  AOI21_X1 U9593 ( .B1(n9820), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7975), .ZN(
        n7982) );
  INV_X1 U9594 ( .A(n7976), .ZN(n7978) );
  INV_X1 U9595 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9409) );
  AOI21_X1 U9596 ( .B1(n7978), .B2(n9409), .A(n7977), .ZN(n7980) );
  XNOR2_X1 U9597 ( .A(n7991), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U9598 ( .A1(n7979), .A2(n7980), .ZN(n7990) );
  OAI211_X1 U9599 ( .C1(n7980), .C2(n7979), .A(n9812), .B(n7990), .ZN(n7981)
         );
  OAI211_X1 U9600 ( .C1(n9815), .C2(n7991), .A(n7982), .B(n7981), .ZN(n7983)
         );
  OR2_X1 U9601 ( .A1(n7984), .A2(n7983), .ZN(P2_U3262) );
  NAND2_X1 U9602 ( .A1(n7987), .A2(n9412), .ZN(n8003) );
  OAI21_X1 U9603 ( .B1(n7987), .B2(n9412), .A(n8003), .ZN(n7999) );
  AOI21_X1 U9604 ( .B1(n9820), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7988), .ZN(
        n7989) );
  OAI21_X1 U9605 ( .B1(n9815), .B2(n8007), .A(n7989), .ZN(n7998) );
  INV_X1 U9606 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7992) );
  OAI21_X1 U9607 ( .B1(n7992), .B2(n7991), .A(n7990), .ZN(n7995) );
  INV_X1 U9608 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8006) );
  AOI22_X1 U9609 ( .A1(n7993), .A2(n8006), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8007), .ZN(n7994) );
  NOR2_X1 U9610 ( .A1(n7995), .A2(n7994), .ZN(n8005) );
  AOI21_X1 U9611 ( .B1(n7995), .B2(n7994), .A(n8005), .ZN(n7996) );
  NOR2_X1 U9612 ( .A1(n7996), .A2(n9817), .ZN(n7997) );
  AOI211_X1 U9613 ( .C1(n7999), .C2(n9814), .A(n7998), .B(n7997), .ZN(n8000)
         );
  INV_X1 U9614 ( .A(n8000), .ZN(P2_U3263) );
  NAND2_X1 U9615 ( .A1(n8001), .A2(n8007), .ZN(n8002) );
  NAND2_X1 U9616 ( .A1(n8003), .A2(n8002), .ZN(n8004) );
  XNOR2_X1 U9617 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8004), .ZN(n8012) );
  INV_X1 U9618 ( .A(n8012), .ZN(n8010) );
  AOI21_X1 U9619 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8008) );
  XOR2_X1 U9620 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8008), .Z(n8011) );
  OAI21_X1 U9621 ( .B1(n8011), .B2(n9817), .A(n9815), .ZN(n8009) );
  AOI21_X1 U9622 ( .B1(n8010), .B2(n9814), .A(n8009), .ZN(n8015) );
  AOI22_X1 U9623 ( .A1(n8012), .A2(n9814), .B1(n9812), .B2(n8011), .ZN(n8014)
         );
  MUX2_X1 U9624 ( .A(n8015), .B(n8014), .S(n8013), .Z(n8017) );
  NAND2_X1 U9625 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8016) );
  OAI211_X1 U9626 ( .C1(n9472), .C2(n4344), .A(n8017), .B(n8016), .ZN(P2_U3264) );
  NAND2_X1 U9627 ( .A1(n8286), .A2(n8277), .ZN(n8022) );
  AOI21_X1 U9628 ( .B1(n8019), .B2(P2_B_REG_SCAN_IN), .A(n8179), .ZN(n8054) );
  NAND2_X1 U9629 ( .A1(n8020), .A2(n8054), .ZN(n9496) );
  NOR2_X1 U9630 ( .A1(n9848), .A2(n9496), .ZN(n8024) );
  AOI21_X1 U9631 ( .B1(n9848), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8024), .ZN(
        n8021) );
  OAI211_X1 U9632 ( .C1(n8288), .C2(n8281), .A(n8022), .B(n8021), .ZN(P2_U3265) );
  AOI21_X1 U9633 ( .B1(n8060), .B2(n8023), .A(n4290), .ZN(n9499) );
  NAND2_X1 U9634 ( .A1(n9499), .A2(n8277), .ZN(n8026) );
  AOI21_X1 U9635 ( .B1(n9848), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8024), .ZN(
        n8025) );
  OAI211_X1 U9636 ( .C1(n9497), .C2(n8281), .A(n8026), .B(n8025), .ZN(P2_U3266) );
  NAND2_X1 U9637 ( .A1(n4489), .A2(n7934), .ZN(n8029) );
  NAND2_X1 U9638 ( .A1(n8245), .A2(n8029), .ZN(n8229) );
  NAND2_X1 U9639 ( .A1(n8229), .A2(n4823), .ZN(n8032) );
  NOR2_X1 U9640 ( .A1(n8332), .A2(n8203), .ZN(n8035) );
  NAND2_X1 U9641 ( .A1(n8132), .A2(n8037), .ZN(n8040) );
  NAND2_X1 U9642 ( .A1(n4475), .A2(n8038), .ZN(n8039) );
  NAND2_X1 U9643 ( .A1(n8040), .A2(n8039), .ZN(n8119) );
  NAND2_X1 U9644 ( .A1(n8117), .A2(n8042), .ZN(n8101) );
  NAND2_X1 U9645 ( .A1(n8101), .A2(n8106), .ZN(n8100) );
  NAND2_X1 U9646 ( .A1(n8114), .A2(n8043), .ZN(n8044) );
  NAND2_X1 U9647 ( .A1(n8100), .A2(n8044), .ZN(n8084) );
  NAND2_X1 U9648 ( .A1(n8091), .A2(n8108), .ZN(n8045) );
  XNOR2_X1 U9649 ( .A(n8048), .B(n8047), .ZN(n8289) );
  INV_X1 U9650 ( .A(n8289), .ZN(n8066) );
  AOI22_X1 U9651 ( .A1(n8095), .A2(n8266), .B1(n8054), .B2(n8053), .ZN(n8055)
         );
  OAI21_X1 U9652 ( .B1(n8058), .B2(n8250), .A(n8292), .ZN(n8064) );
  NAND2_X1 U9653 ( .A1(n8074), .A2(n8290), .ZN(n8059) );
  NAND2_X1 U9654 ( .A1(n8060), .A2(n8059), .ZN(n8291) );
  AOI22_X1 U9655 ( .A1(n8290), .A2(n8255), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9848), .ZN(n8061) );
  OAI21_X1 U9656 ( .B1(n8291), .B2(n8062), .A(n8061), .ZN(n8063) );
  AOI21_X1 U9657 ( .B1(n8064), .B2(n9846), .A(n8063), .ZN(n8065) );
  OAI21_X1 U9658 ( .B1(n8066), .B2(n8262), .A(n8065), .ZN(P2_U3267) );
  XNOR2_X1 U9659 ( .A(n8067), .B(n8072), .ZN(n8070) );
  AOI222_X1 U9660 ( .A1(n8271), .A2(n8070), .B1(n8069), .B2(n8268), .C1(n8068), 
        .C2(n8266), .ZN(n8301) );
  OAI21_X1 U9661 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8297) );
  NAND2_X1 U9662 ( .A1(n8297), .A2(n8284), .ZN(n8082) );
  INV_X1 U9663 ( .A(n8086), .ZN(n8076) );
  INV_X1 U9664 ( .A(n8074), .ZN(n8075) );
  AOI21_X1 U9665 ( .B1(n8298), .B2(n8076), .A(n8075), .ZN(n8299) );
  AOI22_X1 U9666 ( .A1(n9848), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8077), .B2(
        n9834), .ZN(n8078) );
  OAI21_X1 U9667 ( .B1(n8079), .B2(n8281), .A(n8078), .ZN(n8080) );
  AOI21_X1 U9668 ( .B1(n8299), .B2(n8277), .A(n8080), .ZN(n8081) );
  OAI211_X1 U9669 ( .C1(n9848), .C2(n8301), .A(n8082), .B(n8081), .ZN(P2_U3268) );
  OAI21_X1 U9670 ( .B1(n8084), .B2(n8093), .A(n8083), .ZN(n8085) );
  INV_X1 U9671 ( .A(n8085), .ZN(n8307) );
  INV_X1 U9672 ( .A(n8109), .ZN(n8087) );
  AOI21_X1 U9673 ( .B1(n8303), .B2(n8087), .A(n8086), .ZN(n8304) );
  INV_X1 U9674 ( .A(n8088), .ZN(n8089) );
  AOI22_X1 U9675 ( .A1(n9848), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8089), .B2(
        n9834), .ZN(n8090) );
  OAI21_X1 U9676 ( .B1(n8091), .B2(n8281), .A(n8090), .ZN(n8098) );
  XOR2_X1 U9677 ( .A(n8093), .B(n8092), .Z(n8096) );
  AOI222_X1 U9678 ( .A1(n8271), .A2(n8096), .B1(n8095), .B2(n8268), .C1(n8094), 
        .C2(n8266), .ZN(n8306) );
  NOR2_X1 U9679 ( .A1(n8306), .A2(n9848), .ZN(n8097) );
  AOI211_X1 U9680 ( .C1(n8304), .C2(n8277), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI21_X1 U9681 ( .B1(n8307), .B2(n8262), .A(n8099), .ZN(P2_U3269) );
  OAI21_X1 U9682 ( .B1(n8101), .B2(n8106), .A(n8100), .ZN(n8102) );
  INV_X1 U9683 ( .A(n8102), .ZN(n8312) );
  INV_X1 U9684 ( .A(n8103), .ZN(n8104) );
  AOI21_X1 U9685 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8107) );
  OAI222_X1 U9686 ( .A1(n8179), .A2(n8108), .B1(n8181), .B2(n8144), .C1(n9842), 
        .C2(n8107), .ZN(n8308) );
  INV_X1 U9687 ( .A(n8125), .ZN(n8110) );
  AOI211_X1 U9688 ( .C1(n8310), .C2(n8110), .A(n9921), .B(n8109), .ZN(n8309)
         );
  NAND2_X1 U9689 ( .A1(n8309), .A2(n8259), .ZN(n8113) );
  AOI22_X1 U9690 ( .A1(n9848), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8111), .B2(
        n9834), .ZN(n8112) );
  OAI211_X1 U9691 ( .C1(n8114), .C2(n8281), .A(n8113), .B(n8112), .ZN(n8115)
         );
  AOI21_X1 U9692 ( .B1(n8308), .B2(n9846), .A(n8115), .ZN(n8116) );
  OAI21_X1 U9693 ( .B1(n8312), .B2(n8262), .A(n8116), .ZN(P2_U3270) );
  OAI21_X1 U9694 ( .B1(n8119), .B2(n8118), .A(n8117), .ZN(n8120) );
  INV_X1 U9695 ( .A(n8120), .ZN(n8317) );
  XNOR2_X1 U9696 ( .A(n8122), .B(n8121), .ZN(n8124) );
  OAI21_X1 U9697 ( .B1(n8124), .B2(n9842), .A(n8123), .ZN(n8313) );
  INV_X1 U9698 ( .A(n8315), .ZN(n8129) );
  AOI211_X1 U9699 ( .C1(n8315), .C2(n8133), .A(n9921), .B(n8125), .ZN(n8314)
         );
  NAND2_X1 U9700 ( .A1(n8314), .A2(n8259), .ZN(n8128) );
  AOI22_X1 U9701 ( .A1(n9848), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8126), .B2(
        n9834), .ZN(n8127) );
  OAI211_X1 U9702 ( .C1(n8129), .C2(n8281), .A(n8128), .B(n8127), .ZN(n8130)
         );
  AOI21_X1 U9703 ( .B1(n8313), .B2(n9846), .A(n8130), .ZN(n8131) );
  OAI21_X1 U9704 ( .B1(n8317), .B2(n8262), .A(n8131), .ZN(P2_U3271) );
  XNOR2_X1 U9705 ( .A(n8132), .B(n8140), .ZN(n8321) );
  INV_X1 U9706 ( .A(n8133), .ZN(n8134) );
  AOI21_X1 U9707 ( .B1(n5306), .B2(n8153), .A(n8134), .ZN(n8318) );
  INV_X1 U9708 ( .A(n8135), .ZN(n8136) );
  AOI22_X1 U9709 ( .A1(n9848), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8136), .B2(
        n9834), .ZN(n8137) );
  OAI21_X1 U9710 ( .B1(n4475), .B2(n8281), .A(n8137), .ZN(n8148) );
  INV_X1 U9711 ( .A(n8138), .ZN(n8143) );
  AOI21_X1 U9712 ( .B1(n8139), .B2(n8141), .A(n8140), .ZN(n8142) );
  NOR3_X1 U9713 ( .A1(n8143), .A2(n8142), .A3(n9842), .ZN(n8146) );
  OAI22_X1 U9714 ( .A1(n8144), .A2(n8179), .B1(n8180), .B2(n8181), .ZN(n8145)
         );
  NOR2_X1 U9715 ( .A1(n8146), .A2(n8145), .ZN(n8320) );
  NOR2_X1 U9716 ( .A1(n8320), .A2(n9848), .ZN(n8147) );
  AOI211_X1 U9717 ( .C1(n8318), .C2(n8277), .A(n8148), .B(n8147), .ZN(n8149)
         );
  OAI21_X1 U9718 ( .B1(n8321), .B2(n8262), .A(n8149), .ZN(P2_U3272) );
  AOI21_X1 U9719 ( .B1(n8151), .B2(n8150), .A(n4296), .ZN(n8152) );
  INV_X1 U9720 ( .A(n8152), .ZN(n8326) );
  INV_X1 U9721 ( .A(n8153), .ZN(n8154) );
  AOI21_X1 U9722 ( .B1(n8322), .B2(n4479), .A(n8154), .ZN(n8323) );
  AOI22_X1 U9723 ( .A1(n9848), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8155), .B2(
        n9834), .ZN(n8156) );
  OAI21_X1 U9724 ( .B1(n8157), .B2(n8281), .A(n8156), .ZN(n8165) );
  INV_X1 U9725 ( .A(n8158), .ZN(n8178) );
  OAI21_X1 U9726 ( .B1(n8178), .B2(n8160), .A(n8159), .ZN(n8161) );
  NAND2_X1 U9727 ( .A1(n8161), .A2(n8139), .ZN(n8163) );
  AOI222_X1 U9728 ( .A1(n8271), .A2(n8163), .B1(n8162), .B2(n8268), .C1(n8195), 
        .C2(n8266), .ZN(n8325) );
  NOR2_X1 U9729 ( .A1(n8325), .A2(n9848), .ZN(n8164) );
  AOI211_X1 U9730 ( .C1(n8323), .C2(n8277), .A(n8165), .B(n8164), .ZN(n8166)
         );
  OAI21_X1 U9731 ( .B1(n8326), .B2(n8262), .A(n8166), .ZN(P2_U3273) );
  XNOR2_X1 U9732 ( .A(n8168), .B(n8167), .ZN(n8331) );
  AOI21_X1 U9733 ( .B1(n8327), .B2(n8190), .A(n8169), .ZN(n8328) );
  INV_X1 U9734 ( .A(n8327), .ZN(n8172) );
  AOI22_X1 U9735 ( .A1(n9848), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8170), .B2(
        n9834), .ZN(n8171) );
  OAI21_X1 U9736 ( .B1(n8172), .B2(n8281), .A(n8171), .ZN(n8186) );
  INV_X1 U9737 ( .A(n8174), .ZN(n8176) );
  AOI21_X1 U9738 ( .B1(n8173), .B2(n8176), .A(n8175), .ZN(n8177) );
  NOR3_X1 U9739 ( .A1(n8178), .A2(n8177), .A3(n9842), .ZN(n8184) );
  OAI22_X1 U9740 ( .A1(n8182), .A2(n8181), .B1(n8180), .B2(n8179), .ZN(n8183)
         );
  NOR2_X1 U9741 ( .A1(n8184), .A2(n8183), .ZN(n8330) );
  NOR2_X1 U9742 ( .A1(n8330), .A2(n9848), .ZN(n8185) );
  AOI211_X1 U9743 ( .C1(n8328), .C2(n8277), .A(n8186), .B(n8185), .ZN(n8187)
         );
  OAI21_X1 U9744 ( .B1(n8331), .B2(n8262), .A(n8187), .ZN(P2_U3274) );
  XOR2_X1 U9745 ( .A(n8194), .B(n8188), .Z(n8336) );
  INV_X1 U9746 ( .A(n8189), .ZN(n8208) );
  INV_X1 U9747 ( .A(n8190), .ZN(n8191) );
  AOI21_X1 U9748 ( .B1(n8332), .B2(n8208), .A(n8191), .ZN(n8333) );
  AOI22_X1 U9749 ( .A1(n9848), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8192), .B2(
        n9834), .ZN(n8193) );
  OAI21_X1 U9750 ( .B1(n8018), .B2(n8281), .A(n8193), .ZN(n8198) );
  OAI21_X1 U9751 ( .B1(n4289), .B2(n4798), .A(n8173), .ZN(n8196) );
  AOI222_X1 U9752 ( .A1(n8271), .A2(n8196), .B1(n8195), .B2(n8268), .C1(n8224), 
        .C2(n8266), .ZN(n8335) );
  NOR2_X1 U9753 ( .A1(n8335), .A2(n9848), .ZN(n8197) );
  AOI211_X1 U9754 ( .C1(n8333), .C2(n8277), .A(n8198), .B(n8197), .ZN(n8199)
         );
  OAI21_X1 U9755 ( .B1(n8336), .B2(n8262), .A(n8199), .ZN(P2_U3275) );
  NAND2_X1 U9756 ( .A1(n8200), .A2(n8201), .ZN(n8202) );
  XNOR2_X1 U9757 ( .A(n8202), .B(n8205), .ZN(n8204) );
  AOI222_X1 U9758 ( .A1(n8271), .A2(n8204), .B1(n8236), .B2(n8266), .C1(n8203), 
        .C2(n8268), .ZN(n8341) );
  INV_X1 U9759 ( .A(n8343), .ZN(n8207) );
  NAND2_X1 U9760 ( .A1(n8206), .A2(n8205), .ZN(n8337) );
  NAND3_X1 U9761 ( .A1(n8207), .A2(n8284), .A3(n8337), .ZN(n8214) );
  AOI21_X1 U9762 ( .B1(n8338), .B2(n8216), .A(n8189), .ZN(n8339) );
  INV_X1 U9763 ( .A(n8338), .ZN(n8211) );
  AOI22_X1 U9764 ( .A1(n9848), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8209), .B2(
        n9834), .ZN(n8210) );
  OAI21_X1 U9765 ( .B1(n8211), .B2(n8281), .A(n8210), .ZN(n8212) );
  AOI21_X1 U9766 ( .B1(n8339), .B2(n8277), .A(n8212), .ZN(n8213) );
  OAI211_X1 U9767 ( .C1(n9848), .C2(n8341), .A(n8214), .B(n8213), .ZN(P2_U3276) );
  XNOR2_X1 U9768 ( .A(n8215), .B(n8223), .ZN(n8348) );
  INV_X1 U9769 ( .A(n8230), .ZN(n8218) );
  INV_X1 U9770 ( .A(n8216), .ZN(n8217) );
  AOI211_X1 U9771 ( .C1(n8345), .C2(n8218), .A(n9921), .B(n8217), .ZN(n8344)
         );
  AOI22_X1 U9772 ( .A1(n9848), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8219), .B2(
        n9834), .ZN(n8220) );
  OAI21_X1 U9773 ( .B1(n8221), .B2(n8281), .A(n8220), .ZN(n8227) );
  OAI21_X1 U9774 ( .B1(n8223), .B2(n8222), .A(n8200), .ZN(n8225) );
  AOI222_X1 U9775 ( .A1(n8271), .A2(n8225), .B1(n8224), .B2(n8268), .C1(n8242), 
        .C2(n8266), .ZN(n8347) );
  NOR2_X1 U9776 ( .A1(n8347), .A2(n9848), .ZN(n8226) );
  AOI211_X1 U9777 ( .C1(n8344), .C2(n8259), .A(n8227), .B(n8226), .ZN(n8228)
         );
  OAI21_X1 U9778 ( .B1(n8348), .B2(n8262), .A(n8228), .ZN(P2_U3277) );
  XOR2_X1 U9779 ( .A(n8234), .B(n8229), .Z(n8353) );
  AOI21_X1 U9780 ( .B1(n8349), .B2(n4490), .A(n8230), .ZN(n8350) );
  AOI22_X1 U9781 ( .A1(n9848), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8231), .B2(
        n9834), .ZN(n8232) );
  OAI21_X1 U9782 ( .B1(n8233), .B2(n8281), .A(n8232), .ZN(n8239) );
  OAI21_X1 U9783 ( .B1(n4822), .B2(n5203), .A(n8235), .ZN(n8237) );
  AOI222_X1 U9784 ( .A1(n8271), .A2(n8237), .B1(n8269), .B2(n8266), .C1(n8236), 
        .C2(n8268), .ZN(n8352) );
  NOR2_X1 U9785 ( .A1(n8352), .A2(n9848), .ZN(n8238) );
  AOI211_X1 U9786 ( .C1(n8350), .C2(n8277), .A(n8239), .B(n8238), .ZN(n8240)
         );
  OAI21_X1 U9787 ( .B1(n8353), .B2(n8262), .A(n8240), .ZN(P2_U3278) );
  XNOR2_X1 U9788 ( .A(n8241), .B(n8246), .ZN(n8244) );
  AOI222_X1 U9789 ( .A1(n8271), .A2(n8244), .B1(n8243), .B2(n8266), .C1(n8242), 
        .C2(n8268), .ZN(n8357) );
  OAI21_X1 U9790 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8248) );
  INV_X1 U9791 ( .A(n8248), .ZN(n8358) );
  INV_X1 U9792 ( .A(n8249), .ZN(n8251) );
  OAI22_X1 U9793 ( .A1(n8253), .A2(n8252), .B1(n8251), .B2(n8250), .ZN(n8254)
         );
  AOI21_X1 U9794 ( .B1(n8355), .B2(n8255), .A(n8254), .ZN(n8261) );
  NAND2_X1 U9795 ( .A1(n8275), .A2(n8355), .ZN(n8256) );
  NAND2_X1 U9796 ( .A1(n8256), .A2(n9899), .ZN(n8257) );
  NOR2_X1 U9797 ( .A1(n8258), .A2(n8257), .ZN(n8354) );
  NAND2_X1 U9798 ( .A1(n8354), .A2(n8259), .ZN(n8260) );
  OAI211_X1 U9799 ( .C1(n8358), .C2(n8262), .A(n8261), .B(n8260), .ZN(n8263)
         );
  INV_X1 U9800 ( .A(n8263), .ZN(n8264) );
  OAI21_X1 U9801 ( .B1(n9848), .B2(n8357), .A(n8264), .ZN(P2_U3279) );
  XOR2_X1 U9802 ( .A(n8265), .B(n8274), .Z(n8270) );
  AOI222_X1 U9803 ( .A1(n8271), .A2(n8270), .B1(n8269), .B2(n8268), .C1(n8267), 
        .C2(n8266), .ZN(n8363) );
  AOI21_X1 U9804 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8359) );
  INV_X1 U9805 ( .A(n8360), .ZN(n8282) );
  AOI21_X1 U9806 ( .B1(n8360), .B2(n8276), .A(n4491), .ZN(n8361) );
  NAND2_X1 U9807 ( .A1(n8361), .A2(n8277), .ZN(n8280) );
  AOI22_X1 U9808 ( .A1(n9848), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8278), .B2(
        n9834), .ZN(n8279) );
  OAI211_X1 U9809 ( .C1(n8282), .C2(n8281), .A(n8280), .B(n8279), .ZN(n8283)
         );
  AOI21_X1 U9810 ( .B1(n8359), .B2(n8284), .A(n8283), .ZN(n8285) );
  OAI21_X1 U9811 ( .B1(n9848), .B2(n8363), .A(n8285), .ZN(P2_U3280) );
  NAND2_X1 U9812 ( .A1(n8286), .A2(n9899), .ZN(n8287) );
  OAI211_X1 U9813 ( .C1(n8288), .C2(n9919), .A(n8287), .B(n9496), .ZN(n8378)
         );
  MUX2_X1 U9814 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8378), .S(n9943), .Z(
        P2_U3551) );
  NAND2_X1 U9815 ( .A1(n8289), .A2(n9925), .ZN(n8296) );
  INV_X1 U9816 ( .A(n8290), .ZN(n8293) );
  OAI211_X1 U9817 ( .C1(n9919), .C2(n8293), .A(n4819), .B(n8292), .ZN(n8294)
         );
  INV_X1 U9818 ( .A(n8294), .ZN(n8295) );
  NAND2_X1 U9819 ( .A1(n8296), .A2(n8295), .ZN(n8379) );
  MUX2_X1 U9820 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8379), .S(n9943), .Z(
        P2_U3549) );
  NAND2_X1 U9821 ( .A1(n8297), .A2(n9925), .ZN(n8302) );
  AOI22_X1 U9822 ( .A1(n8299), .A2(n9899), .B1(n9898), .B2(n8298), .ZN(n8300)
         );
  NAND3_X1 U9823 ( .A1(n8302), .A2(n8301), .A3(n8300), .ZN(n8380) );
  MUX2_X1 U9824 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8380), .S(n9943), .Z(
        P2_U3548) );
  AOI22_X1 U9825 ( .A1(n8304), .A2(n9899), .B1(n9898), .B2(n8303), .ZN(n8305)
         );
  OAI211_X1 U9826 ( .C1(n8307), .C2(n9904), .A(n8306), .B(n8305), .ZN(n8381)
         );
  MUX2_X1 U9827 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8381), .S(n9943), .Z(
        P2_U3547) );
  AOI211_X1 U9828 ( .C1(n9898), .C2(n8310), .A(n8309), .B(n8308), .ZN(n8311)
         );
  OAI21_X1 U9829 ( .B1(n8312), .B2(n9904), .A(n8311), .ZN(n8382) );
  MUX2_X1 U9830 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8382), .S(n9943), .Z(
        P2_U3546) );
  AOI211_X1 U9831 ( .C1(n9898), .C2(n8315), .A(n8314), .B(n8313), .ZN(n8316)
         );
  OAI21_X1 U9832 ( .B1(n8317), .B2(n9904), .A(n8316), .ZN(n8383) );
  MUX2_X1 U9833 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8383), .S(n9943), .Z(
        P2_U3545) );
  AOI22_X1 U9834 ( .A1(n8318), .A2(n9899), .B1(n9898), .B2(n5306), .ZN(n8319)
         );
  OAI211_X1 U9835 ( .C1(n8321), .C2(n9904), .A(n8320), .B(n8319), .ZN(n8384)
         );
  MUX2_X1 U9836 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8384), .S(n9943), .Z(
        P2_U3544) );
  AOI22_X1 U9837 ( .A1(n8323), .A2(n9899), .B1(n9898), .B2(n8322), .ZN(n8324)
         );
  OAI211_X1 U9838 ( .C1(n8326), .C2(n9904), .A(n8325), .B(n8324), .ZN(n8385)
         );
  MUX2_X1 U9839 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8385), .S(n9943), .Z(
        P2_U3543) );
  AOI22_X1 U9840 ( .A1(n8328), .A2(n9899), .B1(n9898), .B2(n8327), .ZN(n8329)
         );
  OAI211_X1 U9841 ( .C1(n8331), .C2(n9904), .A(n8330), .B(n8329), .ZN(n8386)
         );
  MUX2_X1 U9842 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8386), .S(n9943), .Z(
        P2_U3542) );
  AOI22_X1 U9843 ( .A1(n8333), .A2(n9899), .B1(n9898), .B2(n8332), .ZN(n8334)
         );
  OAI211_X1 U9844 ( .C1(n8336), .C2(n9904), .A(n8335), .B(n8334), .ZN(n8387)
         );
  MUX2_X1 U9845 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8387), .S(n9943), .Z(
        P2_U3541) );
  NAND2_X1 U9846 ( .A1(n8337), .A2(n9925), .ZN(n8342) );
  AOI22_X1 U9847 ( .A1(n8339), .A2(n9899), .B1(n9898), .B2(n8338), .ZN(n8340)
         );
  OAI211_X1 U9848 ( .C1(n8343), .C2(n8342), .A(n8341), .B(n8340), .ZN(n8388)
         );
  MUX2_X1 U9849 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8388), .S(n9943), .Z(
        P2_U3540) );
  AOI21_X1 U9850 ( .B1(n9898), .B2(n8345), .A(n8344), .ZN(n8346) );
  OAI211_X1 U9851 ( .C1(n8348), .C2(n9904), .A(n8347), .B(n8346), .ZN(n8389)
         );
  MUX2_X1 U9852 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8389), .S(n9943), .Z(
        P2_U3539) );
  AOI22_X1 U9853 ( .A1(n8350), .A2(n9899), .B1(n9898), .B2(n8349), .ZN(n8351)
         );
  OAI211_X1 U9854 ( .C1(n8353), .C2(n9904), .A(n8352), .B(n8351), .ZN(n8390)
         );
  MUX2_X1 U9855 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8390), .S(n9943), .Z(
        P2_U3538) );
  AOI21_X1 U9856 ( .B1(n9898), .B2(n8355), .A(n8354), .ZN(n8356) );
  OAI211_X1 U9857 ( .C1(n8358), .C2(n9904), .A(n8357), .B(n8356), .ZN(n8391)
         );
  MUX2_X1 U9858 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8391), .S(n9943), .Z(
        P2_U3537) );
  INV_X1 U9859 ( .A(n8359), .ZN(n8364) );
  AOI22_X1 U9860 ( .A1(n8361), .A2(n9899), .B1(n9898), .B2(n8360), .ZN(n8362)
         );
  OAI211_X1 U9861 ( .C1(n8364), .C2(n9904), .A(n8363), .B(n8362), .ZN(n8392)
         );
  MUX2_X1 U9862 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8392), .S(n9943), .Z(
        P2_U3536) );
  INV_X1 U9863 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8370) );
  OAI21_X1 U9864 ( .B1(n8366), .B2(n9919), .A(n8365), .ZN(n8368) );
  AOI211_X1 U9865 ( .C1(n8369), .C2(n9925), .A(n8368), .B(n8367), .ZN(n8393)
         );
  MUX2_X1 U9866 ( .A(n8370), .B(n8393), .S(n9943), .Z(n8371) );
  INV_X1 U9867 ( .A(n8371), .ZN(P2_U3535) );
  INV_X1 U9868 ( .A(n8372), .ZN(n8377) );
  AOI22_X1 U9869 ( .A1(n8374), .A2(n9899), .B1(n9898), .B2(n8373), .ZN(n8375)
         );
  OAI211_X1 U9870 ( .C1(n9880), .C2(n8377), .A(n8376), .B(n8375), .ZN(n8395)
         );
  MUX2_X1 U9871 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8395), .S(n9943), .Z(
        P2_U3533) );
  MUX2_X1 U9872 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8378), .S(n9912), .Z(
        P2_U3519) );
  MUX2_X1 U9873 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8379), .S(n9912), .Z(
        P2_U3517) );
  MUX2_X1 U9874 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8380), .S(n9912), .Z(
        P2_U3516) );
  MUX2_X1 U9875 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8381), .S(n9912), .Z(
        P2_U3515) );
  MUX2_X1 U9876 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8382), .S(n9912), .Z(
        P2_U3514) );
  MUX2_X1 U9877 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8383), .S(n9912), .Z(
        P2_U3513) );
  MUX2_X1 U9878 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8384), .S(n9912), .Z(
        P2_U3512) );
  MUX2_X1 U9879 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8385), .S(n9912), .Z(
        P2_U3511) );
  MUX2_X1 U9880 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8386), .S(n9912), .Z(
        P2_U3510) );
  MUX2_X1 U9881 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8387), .S(n9912), .Z(
        P2_U3509) );
  MUX2_X1 U9882 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8388), .S(n9912), .Z(
        P2_U3508) );
  MUX2_X1 U9883 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8389), .S(n9912), .Z(
        P2_U3507) );
  MUX2_X1 U9884 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8390), .S(n9912), .Z(
        P2_U3505) );
  MUX2_X1 U9885 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8391), .S(n9912), .Z(
        P2_U3502) );
  MUX2_X1 U9886 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8392), .S(n9912), .Z(
        P2_U3499) );
  MUX2_X1 U9887 ( .A(n5134), .B(n8393), .S(n9912), .Z(n8394) );
  INV_X1 U9888 ( .A(n8394), .ZN(P2_U3496) );
  MUX2_X1 U9889 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8395), .S(n9912), .Z(
        P2_U3490) );
  INV_X1 U9890 ( .A(n8665), .ZN(n9459) );
  NOR4_X1 U9891 ( .A1(n8396), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5069), .A4(
        P2_U3152), .ZN(n8397) );
  AOI21_X1 U9892 ( .B1(n8398), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8397), .ZN(
        n8399) );
  OAI21_X1 U9893 ( .B1(n9459), .B2(n8400), .A(n8399), .ZN(P2_U3327) );
  OAI222_X1 U9894 ( .A1(n8404), .A2(n8403), .B1(n8400), .B2(n8402), .C1(n8401), 
        .C2(P2_U3152), .ZN(P2_U3329) );
  NAND2_X1 U9895 ( .A1(n9460), .A2(n8405), .ZN(n8407) );
  OAI211_X1 U9896 ( .C1(n8404), .C2(n8408), .A(n8407), .B(n8406), .ZN(P2_U3330) );
  MUX2_X1 U9897 ( .A(n8409), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9898 ( .A(n8410), .ZN(n8419) );
  NAND2_X1 U9899 ( .A1(n8534), .A2(n8529), .ZN(n8413) );
  NAND2_X1 U9900 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  AOI21_X1 U9901 ( .B1(n8415), .B2(n8410), .A(n8414), .ZN(n8416) );
  NOR2_X1 U9902 ( .A1(n8416), .A2(n8596), .ZN(n8417) );
  OAI21_X1 U9903 ( .B1(n8419), .B2(n8418), .A(n8417), .ZN(n8424) );
  AOI21_X1 U9904 ( .B1(n8587), .B2(n8879), .A(n8420), .ZN(n8421) );
  OAI21_X1 U9905 ( .B1(n9189), .B2(n8590), .A(n8421), .ZN(n8422) );
  AOI21_X1 U9906 ( .B1(n9192), .B2(n8594), .A(n8422), .ZN(n8423) );
  OAI211_X1 U9907 ( .C1(n9195), .C2(n8591), .A(n8424), .B(n8423), .ZN(P1_U3213) );
  NAND2_X1 U9908 ( .A1(n8425), .A2(n8426), .ZN(n8427) );
  XOR2_X1 U9909 ( .A(n8428), .B(n8427), .Z(n8433) );
  AOI22_X1 U9910 ( .A1(n9077), .A2(n8587), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8430) );
  NAND2_X1 U9911 ( .A1(n9044), .A2(n9573), .ZN(n8429) );
  OAI211_X1 U9912 ( .C1(n8483), .C2(n9037), .A(n8430), .B(n8429), .ZN(n8431)
         );
  AOI21_X1 U9913 ( .B1(n9237), .B2(n9575), .A(n8431), .ZN(n8432) );
  OAI21_X1 U9914 ( .B1(n8433), .B2(n8596), .A(n8432), .ZN(P1_U3214) );
  INV_X1 U9915 ( .A(n8434), .ZN(n8438) );
  NOR3_X1 U9916 ( .A1(n8435), .A2(n8555), .A3(n8436), .ZN(n8437) );
  OAI21_X1 U9917 ( .B1(n8438), .B2(n8437), .A(n9576), .ZN(n8442) );
  NAND2_X1 U9918 ( .A1(n8587), .A2(n9137), .ZN(n8439) );
  NAND2_X1 U9919 ( .A1(n4246), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8961) );
  OAI211_X1 U9920 ( .C1(n9106), .C2(n8590), .A(n8439), .B(n8961), .ZN(n8440)
         );
  AOI21_X1 U9921 ( .B1(n9109), .B2(n8594), .A(n8440), .ZN(n8441) );
  OAI211_X1 U9922 ( .C1(n9112), .C2(n8591), .A(n8442), .B(n8441), .ZN(P1_U3217) );
  NAND2_X1 U9923 ( .A1(n8666), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U9924 ( .A1(n9214), .A2(n8445), .ZN(n8447) );
  INV_X1 U9925 ( .A(n8986), .ZN(n8873) );
  NAND2_X1 U9926 ( .A1(n8873), .A2(n4253), .ZN(n8446) );
  NAND2_X1 U9927 ( .A1(n8447), .A2(n8446), .ZN(n8449) );
  XNOR2_X1 U9928 ( .A(n8449), .B(n8448), .ZN(n8453) );
  NAND2_X1 U9929 ( .A1(n9214), .A2(n4253), .ZN(n8450) );
  OAI21_X1 U9930 ( .B1(n8986), .B2(n8451), .A(n8450), .ZN(n8452) );
  XNOR2_X1 U9931 ( .A(n8453), .B(n8452), .ZN(n8466) );
  NAND3_X1 U9932 ( .A1(n8454), .A2(n9576), .A3(n8466), .ZN(n8469) );
  NOR2_X1 U9933 ( .A1(n9015), .A2(n8483), .ZN(n8464) );
  OR2_X1 U9934 ( .A1(n8993), .A2(n4249), .ZN(n8461) );
  NAND2_X1 U9935 ( .A1(n7471), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U9936 ( .A1(n8455), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U9937 ( .A1(n8456), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8457) );
  AND3_X1 U9938 ( .A1(n8459), .A2(n8458), .A3(n8457), .ZN(n8460) );
  NAND2_X1 U9939 ( .A1(n8461), .A2(n8460), .ZN(n8872) );
  INV_X1 U9940 ( .A(n8872), .ZN(n9012) );
  AOI22_X1 U9941 ( .A1(n8874), .A2(n8587), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8462) );
  OAI21_X1 U9942 ( .B1(n9012), .B2(n8590), .A(n8462), .ZN(n8463) );
  AOI211_X1 U9943 ( .C1(n9214), .C2(n9575), .A(n8464), .B(n8463), .ZN(n8468)
         );
  NAND3_X1 U9944 ( .A1(n8466), .A2(n9576), .A3(n8465), .ZN(n8467) );
  NAND4_X1 U9945 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(
        P1_U3218) );
  AOI21_X1 U9946 ( .B1(n8473), .B2(n8472), .A(n8471), .ZN(n8478) );
  AOI22_X1 U9947 ( .A1(n9077), .A2(n9573), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        n4246), .ZN(n8475) );
  NAND2_X1 U9948 ( .A1(n8594), .A2(n9070), .ZN(n8474) );
  OAI211_X1 U9949 ( .C1(n9106), .C2(n8538), .A(n8475), .B(n8474), .ZN(n8476)
         );
  AOI21_X1 U9950 ( .B1(n9248), .B2(n9575), .A(n8476), .ZN(n8477) );
  OAI21_X1 U9951 ( .B1(n8478), .B2(n8596), .A(n8477), .ZN(P1_U3221) );
  OAI21_X1 U9952 ( .B1(n8480), .B2(n8479), .A(n8574), .ZN(n8481) );
  NAND2_X1 U9953 ( .A1(n8481), .A2(n9576), .ZN(n8488) );
  NOR2_X1 U9954 ( .A1(n8483), .A2(n8482), .ZN(n8486) );
  OAI22_X1 U9955 ( .A1(n8763), .A2(n8590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8484), .ZN(n8485) );
  AOI211_X1 U9956 ( .C1(n8587), .C2(n9044), .A(n8486), .B(n8485), .ZN(n8487)
         );
  OAI211_X1 U9957 ( .C1(n8489), .C2(n8591), .A(n8488), .B(n8487), .ZN(P1_U3223) );
  NAND2_X1 U9958 ( .A1(n8491), .A2(n8584), .ZN(n8496) );
  INV_X1 U9959 ( .A(n8493), .ZN(n8494) );
  AOI21_X1 U9960 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8501) );
  AND2_X1 U9961 ( .A1(n4246), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9645) );
  AOI21_X1 U9962 ( .B1(n9573), .B2(n8877), .A(n9645), .ZN(n8498) );
  NAND2_X1 U9963 ( .A1(n8594), .A2(n9159), .ZN(n8497) );
  OAI211_X1 U9964 ( .C1(n9189), .C2(n8538), .A(n8498), .B(n8497), .ZN(n8499)
         );
  AOI21_X1 U9965 ( .B1(n9276), .B2(n9575), .A(n8499), .ZN(n8500) );
  OAI21_X1 U9966 ( .B1(n8501), .B2(n8596), .A(n8500), .ZN(P1_U3224) );
  OAI21_X1 U9967 ( .B1(n8504), .B2(n8502), .A(n8503), .ZN(n8505) );
  NAND2_X1 U9968 ( .A1(n8505), .A2(n9576), .ZN(n8510) );
  NOR2_X1 U9969 ( .A1(n8506), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9658) );
  AOI21_X1 U9970 ( .B1(n9573), .B2(n9137), .A(n9658), .ZN(n8507) );
  OAI21_X1 U9971 ( .B1(n9171), .B2(n8538), .A(n8507), .ZN(n8508) );
  AOI21_X1 U9972 ( .B1(n9145), .B2(n8594), .A(n8508), .ZN(n8509) );
  OAI211_X1 U9973 ( .C1(n9148), .C2(n8591), .A(n8510), .B(n8509), .ZN(P1_U3226) );
  INV_X1 U9974 ( .A(n8511), .ZN(n8514) );
  OAI21_X1 U9975 ( .B1(n8514), .B2(n8513), .A(n9576), .ZN(n8519) );
  INV_X1 U9976 ( .A(n9030), .ZN(n8517) );
  AOI22_X1 U9977 ( .A1(n8876), .A2(n9573), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        n4246), .ZN(n8515) );
  OAI21_X1 U9978 ( .B1(n9026), .B2(n8538), .A(n8515), .ZN(n8516) );
  AOI21_X1 U9979 ( .B1(n8517), .B2(n8594), .A(n8516), .ZN(n8518) );
  OAI211_X1 U9980 ( .C1(n8520), .C2(n8591), .A(n8519), .B(n8518), .ZN(P1_U3227) );
  AND3_X1 U9981 ( .A1(n8434), .A2(n8522), .A3(n8521), .ZN(n8523) );
  OAI21_X1 U9982 ( .B1(n8524), .B2(n8523), .A(n9576), .ZN(n8528) );
  AOI22_X1 U9983 ( .A1(n9573), .A2(n9095), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8525) );
  OAI21_X1 U9984 ( .B1(n9123), .B2(n8538), .A(n8525), .ZN(n8526) );
  AOI21_X1 U9985 ( .B1(n9088), .B2(n8594), .A(n8526), .ZN(n8527) );
  OAI211_X1 U9986 ( .C1(n9090), .C2(n8591), .A(n8528), .B(n8527), .ZN(P1_U3231) );
  INV_X1 U9987 ( .A(n9522), .ZN(n9549) );
  INV_X1 U9988 ( .A(n8529), .ZN(n8533) );
  OAI21_X1 U9989 ( .B1(n8531), .B2(n8533), .A(n8530), .ZN(n8532) );
  OAI21_X1 U9990 ( .B1(n8534), .B2(n8533), .A(n8532), .ZN(n8535) );
  NAND2_X1 U9991 ( .A1(n8535), .A2(n9576), .ZN(n8541) );
  AOI21_X1 U9992 ( .B1(n9573), .B2(n9518), .A(n8536), .ZN(n8537) );
  OAI21_X1 U9993 ( .B1(n9535), .B2(n8538), .A(n8537), .ZN(n8539) );
  AOI21_X1 U9994 ( .B1(n9521), .B2(n8594), .A(n8539), .ZN(n8540) );
  OAI211_X1 U9995 ( .C1(n9549), .C2(n8591), .A(n8541), .B(n8540), .ZN(P1_U3232) );
  NAND2_X1 U9996 ( .A1(n4302), .A2(n8542), .ZN(n8544) );
  XNOR2_X1 U9997 ( .A(n8544), .B(n8543), .ZN(n8551) );
  NOR2_X1 U9998 ( .A1(n8545), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8546) );
  AOI21_X1 U9999 ( .B1(n8587), .B2(n9095), .A(n8546), .ZN(n8548) );
  NAND2_X1 U10000 ( .A1(n8594), .A2(n9061), .ZN(n8547) );
  OAI211_X1 U10001 ( .C1(n9026), .C2(n8590), .A(n8548), .B(n8547), .ZN(n8549)
         );
  AOI21_X1 U10002 ( .B1(n9244), .B2(n9575), .A(n8549), .ZN(n8550) );
  OAI21_X1 U10003 ( .B1(n8551), .B2(n8596), .A(n8550), .ZN(P1_U3233) );
  INV_X1 U10004 ( .A(n8435), .ZN(n8556) );
  OAI21_X1 U10005 ( .B1(n8553), .B2(n8555), .A(n8552), .ZN(n8554) );
  OAI21_X1 U10006 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8557) );
  NAND2_X1 U10007 ( .A1(n8557), .A2(n9576), .ZN(n8561) );
  NAND2_X1 U10008 ( .A1(n8587), .A2(n8877), .ZN(n8558) );
  NAND2_X1 U10009 ( .A1(n4246), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8922) );
  OAI211_X1 U10010 ( .C1(n9123), .C2(n8590), .A(n8558), .B(n8922), .ZN(n8559)
         );
  AOI21_X1 U10011 ( .B1(n9116), .B2(n8594), .A(n8559), .ZN(n8560) );
  OAI211_X1 U10012 ( .C1(n4460), .C2(n8591), .A(n8561), .B(n8560), .ZN(
        P1_U3236) );
  OAI21_X1 U10013 ( .B1(n8564), .B2(n8562), .A(n8563), .ZN(n8565) );
  NAND2_X1 U10014 ( .A1(n8565), .A2(n9576), .ZN(n8572) );
  AOI21_X1 U10015 ( .B1(n9573), .B2(n8884), .A(n8566), .ZN(n8571) );
  AOI22_X1 U10016 ( .A1(n8567), .A2(n9575), .B1(n8587), .B2(n8886), .ZN(n8570)
         );
  NAND2_X1 U10017 ( .A1(n8594), .A2(n8568), .ZN(n8569) );
  NAND4_X1 U10018 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(
        P1_U3237) );
  AND2_X1 U10019 ( .A1(n8574), .A2(n8573), .ZN(n8577) );
  OAI211_X1 U10020 ( .C1(n8577), .C2(n8576), .A(n9576), .B(n8575), .ZN(n8582)
         );
  AOI22_X1 U10021 ( .A1(n8876), .A2(n8587), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8578) );
  OAI21_X1 U10022 ( .B1(n9011), .B2(n8590), .A(n8578), .ZN(n8579) );
  AOI21_X1 U10023 ( .B1(n8580), .B2(n8594), .A(n8579), .ZN(n8581) );
  OAI211_X1 U10024 ( .C1(n8762), .C2(n8591), .A(n8582), .B(n8581), .ZN(
        P1_U3238) );
  NAND2_X1 U10025 ( .A1(n8584), .A2(n8583), .ZN(n8585) );
  XOR2_X1 U10026 ( .A(n8586), .B(n8585), .Z(n8597) );
  NAND2_X1 U10027 ( .A1(n8587), .A2(n9518), .ZN(n8589) );
  NAND2_X1 U10028 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9631) );
  OAI211_X1 U10029 ( .C1(n9171), .C2(n8590), .A(n8589), .B(n9631), .ZN(n8593)
         );
  NOR2_X1 U10030 ( .A1(n9178), .A2(n8591), .ZN(n8592) );
  AOI211_X1 U10031 ( .C1(n9176), .C2(n8594), .A(n8593), .B(n8592), .ZN(n8595)
         );
  OAI21_X1 U10032 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(P1_U3239) );
  INV_X1 U10033 ( .A(n8776), .ZN(n8599) );
  NAND2_X1 U10034 ( .A1(n9214), .A2(n8986), .ZN(n8779) );
  INV_X1 U10035 ( .A(n8779), .ZN(n8983) );
  INV_X1 U10036 ( .A(n8600), .ZN(n8633) );
  INV_X1 U10037 ( .A(n8802), .ZN(n8601) );
  NAND2_X1 U10038 ( .A1(n8602), .A2(n8601), .ZN(n8757) );
  OR2_X1 U10039 ( .A1(n9234), .A2(n8603), .ZN(n8756) );
  NAND2_X1 U10040 ( .A1(n8757), .A2(n8756), .ZN(n8604) );
  NAND2_X1 U10041 ( .A1(n8605), .A2(n8604), .ZN(n8758) );
  INV_X1 U10042 ( .A(n8758), .ZN(n8631) );
  AND2_X1 U10043 ( .A1(n8721), .A2(n8606), .ZN(n8716) );
  INV_X1 U10044 ( .A(n8716), .ZN(n8617) );
  AND2_X1 U10045 ( .A1(n8687), .A2(n8609), .ZN(n8614) );
  AND2_X1 U10046 ( .A1(n8702), .A2(n8607), .ZN(n8608) );
  NAND2_X1 U10047 ( .A1(n9184), .A2(n8608), .ZN(n8712) );
  INV_X1 U10048 ( .A(n8609), .ZN(n8697) );
  NOR2_X1 U10049 ( .A1(n8610), .A2(n8697), .ZN(n8611) );
  OR2_X1 U10050 ( .A1(n8712), .A2(n8611), .ZN(n8651) );
  INV_X1 U10051 ( .A(n8612), .ZN(n8707) );
  NAND3_X1 U10052 ( .A1(n8707), .A2(n9184), .A3(n8702), .ZN(n8613) );
  OAI211_X1 U10053 ( .C1(n8614), .C2(n8651), .A(n4318), .B(n8613), .ZN(n8615)
         );
  AND3_X1 U10054 ( .A1(n8615), .A2(n8650), .A3(n8708), .ZN(n8616) );
  OAI21_X1 U10055 ( .B1(n8617), .B2(n8616), .A(n8719), .ZN(n8618) );
  NOR2_X1 U10056 ( .A1(n8725), .A2(n8618), .ZN(n8622) );
  NAND2_X1 U10057 ( .A1(n8619), .A2(n8728), .ZN(n8621) );
  AND2_X1 U10058 ( .A1(n8731), .A2(n8724), .ZN(n8620) );
  AND2_X1 U10059 ( .A1(n8750), .A2(n8620), .ZN(n8649) );
  OAI21_X1 U10060 ( .B1(n8622), .B2(n8621), .A(n8649), .ZN(n8629) );
  INV_X1 U10061 ( .A(n8744), .ZN(n8623) );
  NAND2_X1 U10062 ( .A1(n9051), .A2(n8623), .ZN(n8625) );
  AND2_X1 U10063 ( .A1(n8625), .A2(n8624), .ZN(n8746) );
  INV_X1 U10064 ( .A(n8746), .ZN(n8626) );
  NAND2_X1 U10065 ( .A1(n8747), .A2(n8626), .ZN(n8627) );
  NAND4_X1 U10066 ( .A1(n8629), .A2(n8628), .A3(n8756), .A4(n8627), .ZN(n8630)
         );
  NAND2_X1 U10067 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  NAND3_X1 U10068 ( .A1(n9008), .A2(n8633), .A3(n8632), .ZN(n8638) );
  NAND2_X1 U10069 ( .A1(n8634), .A2(n7463), .ZN(n8636) );
  NAND2_X1 U10070 ( .A1(n8666), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8635) );
  NOR2_X1 U10071 ( .A1(n9209), .A2(n9012), .ZN(n8800) );
  INV_X1 U10072 ( .A(n8780), .ZN(n8637) );
  AOI211_X1 U10073 ( .C1(n8648), .C2(n8638), .A(n8800), .B(n8637), .ZN(n8849)
         );
  NAND2_X1 U10074 ( .A1(n5913), .A2(n5973), .ZN(n8639) );
  OAI211_X1 U10075 ( .C1(n8640), .C2(n6076), .A(n5762), .B(n8639), .ZN(n8641)
         );
  NAND2_X1 U10076 ( .A1(n8641), .A2(n9705), .ZN(n8644) );
  OAI22_X1 U10077 ( .A1(n8645), .A2(n8644), .B1(n8643), .B2(n8642), .ZN(n8646)
         );
  AND2_X1 U10078 ( .A1(n8646), .A2(n8838), .ZN(n8659) );
  NAND4_X1 U10079 ( .A1(n8657), .A2(n8680), .A3(n8835), .A4(n8647), .ZN(n8845)
         );
  INV_X1 U10080 ( .A(n8648), .ZN(n8656) );
  INV_X1 U10081 ( .A(n8649), .ZN(n8654) );
  NAND2_X1 U10082 ( .A1(n8719), .A2(n8650), .ZN(n8718) );
  INV_X1 U10083 ( .A(n8651), .ZN(n8652) );
  NAND4_X1 U10084 ( .A1(n8708), .A2(n8652), .A3(n8692), .A4(n8681), .ZN(n8653)
         );
  OR4_X1 U10085 ( .A1(n8654), .A2(n8725), .A3(n8718), .A4(n8653), .ZN(n8655)
         );
  NOR3_X1 U10086 ( .A1(n8656), .A2(n8758), .A3(n8655), .ZN(n8844) );
  OAI211_X1 U10087 ( .C1(n8841), .C2(n4542), .A(n8680), .B(n8657), .ZN(n8658)
         );
  OAI211_X1 U10088 ( .C1(n8659), .C2(n8845), .A(n8844), .B(n8658), .ZN(n8660)
         );
  NOR2_X1 U10089 ( .A1(n8997), .A2(n8872), .ZN(n8847) );
  AOI21_X1 U10090 ( .B1(n8849), .B2(n8660), .A(n8847), .ZN(n8669) );
  NAND2_X1 U10091 ( .A1(n8665), .A2(n7463), .ZN(n8668) );
  NAND2_X1 U10092 ( .A1(n8666), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8667) );
  NOR2_X1 U10093 ( .A1(n9199), .A2(n8966), .ZN(n8795) );
  AOI21_X1 U10094 ( .B1(n8988), .B2(n9203), .A(n8795), .ZN(n8830) );
  OAI21_X1 U10095 ( .B1(n8669), .B2(n8829), .A(n8830), .ZN(n8671) );
  INV_X1 U10096 ( .A(n8828), .ZN(n8670) );
  NAND2_X1 U10097 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U10098 ( .A(n8672), .B(n9679), .ZN(n8864) );
  MUX2_X1 U10099 ( .A(n8674), .B(n8673), .S(n8775), .Z(n8676) );
  NOR2_X1 U10100 ( .A1(n8676), .A2(n8675), .ZN(n8685) );
  NAND2_X1 U10101 ( .A1(n8680), .A2(n8677), .ZN(n8839) );
  NAND2_X1 U10102 ( .A1(n8681), .A2(n8678), .ZN(n8679) );
  MUX2_X1 U10103 ( .A(n8839), .B(n8679), .S(n8785), .Z(n8684) );
  INV_X1 U10104 ( .A(n8812), .ZN(n8683) );
  MUX2_X1 U10105 ( .A(n8681), .B(n8680), .S(n8785), .Z(n8682) );
  OAI211_X1 U10106 ( .C1(n8685), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8691)
         );
  INV_X1 U10107 ( .A(n8693), .ZN(n8686) );
  AOI211_X1 U10108 ( .C1(n8691), .C2(n8687), .A(n8686), .B(n8785), .ZN(n8690)
         );
  OAI22_X1 U10109 ( .A1(n8690), .A2(n8689), .B1(n8688), .B2(n8785), .ZN(n8699)
         );
  INV_X1 U10110 ( .A(n8691), .ZN(n8696) );
  NAND2_X1 U10111 ( .A1(n8693), .A2(n8692), .ZN(n8695) );
  OAI211_X1 U10112 ( .C1(n8696), .C2(n8695), .A(n8694), .B(n8785), .ZN(n8698)
         );
  AOI22_X1 U10113 ( .A1(n8699), .A2(n8698), .B1(n8697), .B2(n8785), .ZN(n8701)
         );
  XNOR2_X1 U10114 ( .A(n9540), .B(n8700), .ZN(n9530) );
  NOR2_X1 U10115 ( .A1(n8701), .A2(n9530), .ZN(n8713) );
  INV_X1 U10116 ( .A(n8702), .ZN(n8705) );
  INV_X1 U10117 ( .A(n8703), .ZN(n8704) );
  MUX2_X1 U10118 ( .A(n8705), .B(n8704), .S(n8775), .Z(n8714) );
  INV_X1 U10119 ( .A(n8714), .ZN(n8706) );
  INV_X1 U10120 ( .A(n8708), .ZN(n8715) );
  OAI22_X1 U10121 ( .A1(n8717), .A2(n9167), .B1(n8716), .B2(n8775), .ZN(n8720)
         );
  AOI22_X1 U10122 ( .A1(n8720), .A2(n8719), .B1(n8775), .B2(n8718), .ZN(n8727)
         );
  INV_X1 U10123 ( .A(n8721), .ZN(n8723) );
  MUX2_X1 U10124 ( .A(n9271), .B(n8775), .S(n9156), .Z(n8722) );
  AOI21_X1 U10125 ( .B1(n9148), .B2(n8785), .A(n8722), .ZN(n8726) );
  INV_X1 U10126 ( .A(n8728), .ZN(n8730) );
  INV_X1 U10127 ( .A(n8731), .ZN(n8743) );
  NAND2_X1 U10128 ( .A1(n9105), .A2(n8785), .ZN(n8736) );
  INV_X1 U10129 ( .A(n8736), .ZN(n8733) );
  NOR2_X1 U10130 ( .A1(n9094), .A2(n8775), .ZN(n8732) );
  AOI21_X1 U10131 ( .B1(n9266), .B2(n8733), .A(n8732), .ZN(n8741) );
  NAND2_X1 U10132 ( .A1(n9137), .A2(n8775), .ZN(n8735) );
  OAI22_X1 U10133 ( .A1(n9266), .A2(n8735), .B1(n9123), .B2(n8785), .ZN(n8734)
         );
  NAND2_X1 U10134 ( .A1(n9112), .A2(n8734), .ZN(n8740) );
  NOR2_X1 U10135 ( .A1(n8735), .A2(n9123), .ZN(n8738) );
  OAI21_X1 U10136 ( .B1(n9094), .B2(n8736), .A(n9266), .ZN(n8737) );
  OAI21_X1 U10137 ( .B1(n8738), .B2(n9266), .A(n8737), .ZN(n8739) );
  OAI211_X1 U10138 ( .C1(n9112), .C2(n8741), .A(n8740), .B(n8739), .ZN(n8742)
         );
  AOI21_X1 U10139 ( .B1(n8744), .B2(n8785), .A(n9093), .ZN(n8745) );
  NAND2_X1 U10140 ( .A1(n8747), .A2(n9040), .ZN(n9050) );
  NAND2_X1 U10141 ( .A1(n9040), .A2(n8746), .ZN(n8748) );
  AND2_X1 U10142 ( .A1(n8748), .A2(n8747), .ZN(n8752) );
  INV_X1 U10143 ( .A(n9040), .ZN(n8749) );
  NOR2_X1 U10144 ( .A1(n8750), .A2(n8749), .ZN(n8751) );
  MUX2_X1 U10145 ( .A(n8752), .B(n8751), .S(n8785), .Z(n8754) );
  NAND2_X1 U10146 ( .A1(n8756), .A2(n8801), .ZN(n8753) );
  NOR4_X1 U10147 ( .A1(n8755), .A2(n8754), .A3(n8757), .A4(n8753), .ZN(n8761)
         );
  OAI211_X1 U10148 ( .C1(n8757), .C2(n8801), .A(n7527), .B(n8756), .ZN(n8759)
         );
  MUX2_X1 U10149 ( .A(n8759), .B(n8758), .S(n8775), .Z(n8760) );
  NOR2_X1 U10150 ( .A1(n8761), .A2(n8760), .ZN(n8771) );
  MUX2_X1 U10151 ( .A(n8763), .B(n8762), .S(n8775), .Z(n8770) );
  NOR3_X1 U10152 ( .A1(n8771), .A2(n8770), .A3(n8766), .ZN(n8774) );
  INV_X1 U10153 ( .A(n8766), .ZN(n8767) );
  NOR2_X1 U10154 ( .A1(n8767), .A2(n8875), .ZN(n8768) );
  AOI21_X1 U10155 ( .B1(n8775), .B2(n8875), .A(n8769), .ZN(n8773) );
  AOI21_X1 U10156 ( .B1(n8771), .B2(n8770), .A(n8975), .ZN(n8772) );
  OAI21_X1 U10157 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8778) );
  MUX2_X1 U10158 ( .A(n9008), .B(n8776), .S(n8775), .Z(n8777) );
  MUX2_X1 U10159 ( .A(n8780), .B(n8779), .S(n8785), .Z(n8781) );
  OAI21_X1 U10160 ( .B1(n8966), .B2(n8988), .A(n9203), .ZN(n8852) );
  OAI211_X1 U10161 ( .C1(n8997), .C2(n8785), .A(n8850), .B(n8852), .ZN(n8782)
         );
  NAND3_X1 U10162 ( .A1(n8850), .A2(n8788), .A3(n9209), .ZN(n8784) );
  NAND3_X1 U10163 ( .A1(n8788), .A2(n8872), .A3(n8852), .ZN(n8789) );
  NAND2_X1 U10164 ( .A1(n8789), .A2(n8850), .ZN(n8790) );
  INV_X1 U10165 ( .A(n8795), .ZN(n8796) );
  NAND2_X1 U10166 ( .A1(n8796), .A2(n5762), .ZN(n8856) );
  INV_X1 U10167 ( .A(n8856), .ZN(n8797) );
  NAND2_X1 U10168 ( .A1(n8797), .A2(n8798), .ZN(n8861) );
  NOR2_X1 U10169 ( .A1(n8856), .A2(n8798), .ZN(n8799) );
  NOR2_X1 U10170 ( .A1(n8847), .A2(n8800), .ZN(n8980) );
  INV_X1 U10171 ( .A(n8980), .ZN(n8984) );
  INV_X1 U10172 ( .A(n8801), .ZN(n8803) );
  INV_X1 U10173 ( .A(n9050), .ZN(n9052) );
  INV_X1 U10174 ( .A(n9153), .ZN(n8819) );
  NOR4_X1 U10175 ( .A1(n8806), .A2(n8805), .A3(n9704), .A4(n8804), .ZN(n8809)
         );
  NAND4_X1 U10176 ( .A1(n8809), .A2(n8808), .A3(n9681), .A4(n8807), .ZN(n8813)
         );
  NOR4_X1 U10177 ( .A1(n8813), .A2(n8812), .A3(n8811), .A4(n8810), .ZN(n8816)
         );
  INV_X1 U10178 ( .A(n9530), .ZN(n9532) );
  NAND4_X1 U10179 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n9532), .ZN(n8817)
         );
  NOR4_X1 U10180 ( .A1(n9167), .A2(n8817), .A3(n9185), .A4(n9511), .ZN(n8818)
         );
  NAND3_X1 U10181 ( .A1(n9135), .A2(n8819), .A3(n8818), .ZN(n8820) );
  NOR4_X1 U10182 ( .A1(n9083), .A2(n9103), .A3(n8820), .A4(n9126), .ZN(n8821)
         );
  NAND3_X1 U10183 ( .A1(n9052), .A2(n9075), .A3(n8821), .ZN(n8822) );
  NOR4_X1 U10184 ( .A1(n8823), .A2(n9024), .A3(n9042), .A4(n8822), .ZN(n8825)
         );
  NAND4_X1 U10185 ( .A1(n9007), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n8827)
         );
  AOI21_X1 U10186 ( .B1(n8831), .B2(n8830), .A(n5762), .ZN(n8854) );
  INV_X1 U10187 ( .A(n8834), .ZN(n8846) );
  AOI211_X1 U10188 ( .C1(n8838), .C2(n8837), .A(n4539), .B(n4538), .ZN(n8842)
         );
  INV_X1 U10189 ( .A(n8839), .ZN(n8840) );
  OAI21_X1 U10190 ( .B1(n8842), .B2(n8841), .A(n8840), .ZN(n8843) );
  OAI211_X1 U10191 ( .C1(n8846), .C2(n8845), .A(n8844), .B(n8843), .ZN(n8848)
         );
  AOI21_X1 U10192 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8853) );
  INV_X1 U10193 ( .A(n8850), .ZN(n8851) );
  AOI21_X1 U10194 ( .B1(n8853), .B2(n8852), .A(n8851), .ZN(n8857) );
  INV_X1 U10195 ( .A(n8854), .ZN(n8855) );
  OAI21_X1 U10196 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8858) );
  INV_X1 U10197 ( .A(n8865), .ZN(n8869) );
  OR3_X1 U10198 ( .A1(n8867), .A2(n8866), .A3(n8964), .ZN(n8868) );
  OAI211_X1 U10199 ( .C1(n5764), .C2(n8869), .A(n8868), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8870) );
  NAND2_X1 U10200 ( .A1(n8871), .A2(n8870), .ZN(P1_U3240) );
  MUX2_X1 U10201 ( .A(n8872), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8888), .Z(
        P1_U3584) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8873), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10203 ( .A(n8874), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8888), .Z(
        P1_U3582) );
  MUX2_X1 U10204 ( .A(n8875), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8888), .Z(
        P1_U3581) );
  MUX2_X1 U10205 ( .A(n8876), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8888), .Z(
        P1_U3580) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9044), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10207 ( .A(n9055), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8888), .Z(
        P1_U3578) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9077), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10209 ( .A(n9095), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8888), .Z(
        P1_U3576) );
  MUX2_X1 U10210 ( .A(n9076), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8888), .Z(
        P1_U3575) );
  MUX2_X1 U10211 ( .A(n9094), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8888), .Z(
        P1_U3574) );
  MUX2_X1 U10212 ( .A(n9137), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8888), .Z(
        P1_U3573) );
  MUX2_X1 U10213 ( .A(n8877), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8888), .Z(
        P1_U3572) );
  MUX2_X1 U10214 ( .A(n9138), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8888), .Z(
        P1_U3571) );
  MUX2_X1 U10215 ( .A(n8878), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8888), .Z(
        P1_U3570) );
  MUX2_X1 U10216 ( .A(n9518), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8888), .Z(
        P1_U3569) );
  MUX2_X1 U10217 ( .A(n8879), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8888), .Z(
        P1_U3568) );
  MUX2_X1 U10218 ( .A(n9517), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8888), .Z(
        P1_U3567) );
  MUX2_X1 U10219 ( .A(n8880), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8888), .Z(
        P1_U3566) );
  MUX2_X1 U10220 ( .A(n8881), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8888), .Z(
        P1_U3565) );
  MUX2_X1 U10221 ( .A(n8882), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8888), .Z(
        P1_U3564) );
  MUX2_X1 U10222 ( .A(n8883), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8888), .Z(
        P1_U3563) );
  MUX2_X1 U10223 ( .A(n8884), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8888), .Z(
        P1_U3562) );
  MUX2_X1 U10224 ( .A(n8885), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8888), .Z(
        P1_U3561) );
  MUX2_X1 U10225 ( .A(n8886), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8888), .Z(
        P1_U3560) );
  MUX2_X1 U10226 ( .A(n9701), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8888), .Z(
        P1_U3559) );
  MUX2_X1 U10227 ( .A(n8887), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8888), .Z(
        P1_U3558) );
  MUX2_X1 U10228 ( .A(n4250), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8888), .Z(
        P1_U3557) );
  MUX2_X1 U10229 ( .A(n6414), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8888), .Z(
        P1_U3556) );
  NAND2_X1 U10230 ( .A1(n9659), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n8901) );
  AOI22_X1 U10231 ( .A1(n9634), .A2(n8889), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n8900) );
  OAI211_X1 U10232 ( .C1(n8892), .C2(n8891), .A(n9665), .B(n8890), .ZN(n8899)
         );
  INV_X1 U10233 ( .A(n8893), .ZN(n8895) );
  NAND2_X1 U10234 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8894) );
  NAND2_X1 U10235 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  NAND3_X1 U10236 ( .A1(n9661), .A2(n8897), .A3(n8896), .ZN(n8898) );
  NAND4_X1 U10237 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(
        P1_U3242) );
  NAND2_X1 U10238 ( .A1(n9659), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8913) );
  AOI22_X1 U10239 ( .A1(n9634), .A2(n8902), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n4246), .ZN(n8912) );
  OAI211_X1 U10240 ( .C1(n8905), .C2(n8904), .A(n9665), .B(n8903), .ZN(n8911)
         );
  INV_X1 U10241 ( .A(n8906), .ZN(n8907) );
  OAI211_X1 U10242 ( .C1(n8909), .C2(n8908), .A(n9661), .B(n8907), .ZN(n8910)
         );
  NAND4_X1 U10243 ( .A1(n8913), .A2(n8912), .A3(n8911), .A4(n8910), .ZN(
        P1_U3244) );
  INV_X1 U10244 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8950) );
  AOI22_X1 U10245 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n8951), .B1(n8940), .B2(
        n8950), .ZN(n8921) );
  INV_X1 U10246 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9414) );
  XNOR2_X1 U10247 ( .A(n9655), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9663) );
  INV_X1 U10248 ( .A(n8929), .ZN(n9643) );
  INV_X1 U10249 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8919) );
  XOR2_X1 U10250 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n8929), .Z(n9647) );
  NAND2_X1 U10251 ( .A1(n9633), .A2(n8917), .ZN(n8918) );
  XOR2_X1 U10252 ( .A(n9633), .B(n8917), .Z(n9636) );
  NAND2_X1 U10253 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9636), .ZN(n9635) );
  NAND2_X1 U10254 ( .A1(n8918), .A2(n9635), .ZN(n9648) );
  NAND2_X1 U10255 ( .A1(n9647), .A2(n9648), .ZN(n9646) );
  OAI21_X1 U10256 ( .B1(n9643), .B2(n8919), .A(n9646), .ZN(n9662) );
  NAND2_X1 U10257 ( .A1(n9663), .A2(n9662), .ZN(n9660) );
  OAI21_X1 U10258 ( .B1(n9414), .B2(n9655), .A(n9660), .ZN(n8920) );
  NOR2_X1 U10259 ( .A1(n8921), .A2(n8920), .ZN(n8949) );
  AOI21_X1 U10260 ( .B1(n8921), .B2(n8920), .A(n8949), .ZN(n8945) );
  INV_X1 U10261 ( .A(n8922), .ZN(n8923) );
  AOI21_X1 U10262 ( .B1(n9634), .B2(n8940), .A(n8923), .ZN(n8924) );
  OAI21_X1 U10263 ( .B1(n9605), .B2(n9981), .A(n8924), .ZN(n8925) );
  INV_X1 U10264 ( .A(n8925), .ZN(n8944) );
  NAND2_X1 U10265 ( .A1(n8926), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8939) );
  INV_X1 U10266 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8927) );
  MUX2_X1 U10267 ( .A(n8927), .B(P1_REG2_REG_17__SCAN_IN), .S(n8926), .Z(n8928) );
  INV_X1 U10268 ( .A(n8928), .ZN(n9666) );
  NAND2_X1 U10269 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8929), .ZN(n8938) );
  INV_X1 U10270 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U10271 ( .A(n8930), .B(P1_REG2_REG_16__SCAN_IN), .S(n8929), .Z(n8931) );
  INV_X1 U10272 ( .A(n8931), .ZN(n9650) );
  NOR2_X1 U10273 ( .A1(n8933), .A2(n8932), .ZN(n8935) );
  NOR2_X1 U10274 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND2_X1 U10275 ( .A1(n9633), .A2(n8936), .ZN(n8937) );
  XOR2_X1 U10276 ( .A(n9633), .B(n8936), .Z(n9638) );
  NAND2_X1 U10277 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9638), .ZN(n9637) );
  NAND2_X1 U10278 ( .A1(n8937), .A2(n9637), .ZN(n9651) );
  NAND2_X1 U10279 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  NAND2_X1 U10280 ( .A1(n8938), .A2(n9649), .ZN(n9667) );
  NAND2_X1 U10281 ( .A1(n9666), .A2(n9667), .ZN(n9664) );
  NAND2_X1 U10282 ( .A1(n8939), .A2(n9664), .ZN(n8942) );
  INV_X1 U10283 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U10284 ( .A(n8940), .B(n8947), .ZN(n8941) );
  NAND2_X1 U10285 ( .A1(n8941), .A2(n8942), .ZN(n8946) );
  OAI211_X1 U10286 ( .C1(n8942), .C2(n8941), .A(n9665), .B(n8946), .ZN(n8943)
         );
  OAI211_X1 U10287 ( .C1(n8945), .C2(n9622), .A(n8944), .B(n8943), .ZN(
        P1_U3259) );
  OAI21_X1 U10288 ( .B1(n8951), .B2(n8947), .A(n8946), .ZN(n8948) );
  XNOR2_X1 U10289 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8948), .ZN(n8957) );
  INV_X1 U10290 ( .A(n8957), .ZN(n8955) );
  INV_X1 U10291 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8952) );
  XOR2_X1 U10292 ( .A(n8953), .B(n8952), .Z(n8958) );
  NAND2_X1 U10293 ( .A1(n8958), .A2(n9661), .ZN(n8954) );
  OAI211_X1 U10294 ( .C1(n8956), .C2(n8955), .A(n8954), .B(n9656), .ZN(n8960)
         );
  OAI22_X1 U10295 ( .A1(n8958), .A2(n9622), .B1(n8957), .B2(n8956), .ZN(n8959)
         );
  INV_X1 U10296 ( .A(n9203), .ZN(n8970) );
  NAND2_X1 U10297 ( .A1(n8970), .A2(n8991), .ZN(n8962) );
  XNOR2_X1 U10298 ( .A(n8962), .B(n9199), .ZN(n9201) );
  INV_X1 U10299 ( .A(P1_B_REG_SCAN_IN), .ZN(n8963) );
  NOR2_X1 U10300 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  OR2_X1 U10301 ( .A1(n9687), .A2(n8965), .ZN(n8987) );
  NOR2_X1 U10302 ( .A1(n8966), .A2(n8987), .ZN(n9202) );
  INV_X1 U10303 ( .A(n9202), .ZN(n8967) );
  NOR2_X1 U10304 ( .A1(n8967), .A2(n9715), .ZN(n8972) );
  AOI21_X1 U10305 ( .B1(n9715), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8972), .ZN(
        n8969) );
  NAND2_X1 U10306 ( .A1(n9199), .A2(n9539), .ZN(n8968) );
  OAI211_X1 U10307 ( .C1(n9201), .C2(n8974), .A(n8969), .B(n8968), .ZN(
        P1_U3261) );
  XNOR2_X1 U10308 ( .A(n8970), .B(n8991), .ZN(n9205) );
  NOR2_X1 U10309 ( .A1(n8970), .A2(n9717), .ZN(n8971) );
  AOI211_X1 U10310 ( .C1(n9715), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8972), .B(
        n8971), .ZN(n8973) );
  OAI21_X1 U10311 ( .B1(n9205), .B2(n8974), .A(n8973), .ZN(P1_U3262) );
  NAND2_X1 U10312 ( .A1(n8978), .A2(n9011), .ZN(n9001) );
  AND2_X1 U10313 ( .A1(n9004), .A2(n9001), .ZN(n8979) );
  NAND2_X1 U10314 ( .A1(n9002), .A2(n8979), .ZN(n9003) );
  INV_X1 U10315 ( .A(n9214), .ZN(n9019) );
  NAND2_X1 U10316 ( .A1(n9003), .A2(n4805), .ZN(n8981) );
  XNOR2_X1 U10317 ( .A(n8981), .B(n8980), .ZN(n9206) );
  INV_X1 U10318 ( .A(n9206), .ZN(n9000) );
  INV_X1 U10319 ( .A(n9008), .ZN(n8982) );
  AOI21_X1 U10320 ( .B1(n8873), .B2(n9700), .A(n8989), .ZN(n8990) );
  INV_X1 U10321 ( .A(n9013), .ZN(n8992) );
  AOI211_X1 U10322 ( .C1(n9209), .C2(n8992), .A(n9786), .B(n8991), .ZN(n9208)
         );
  NAND2_X1 U10323 ( .A1(n9208), .A2(n9144), .ZN(n8996) );
  INV_X1 U10324 ( .A(n8993), .ZN(n8994) );
  AOI22_X1 U10325 ( .A1(n8994), .A2(n9714), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9715), .ZN(n8995) );
  OAI211_X1 U10326 ( .C1(n8997), .C2(n9717), .A(n8996), .B(n8995), .ZN(n8998)
         );
  AOI21_X1 U10327 ( .B1(n9207), .B2(n9719), .A(n8998), .ZN(n8999) );
  OAI21_X1 U10328 ( .B1(n9000), .B2(n9198), .A(n8999), .ZN(P1_U3355) );
  AND2_X1 U10329 ( .A1(n9002), .A2(n9001), .ZN(n9005) );
  OAI21_X1 U10330 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9216) );
  AOI21_X1 U10331 ( .B1(n4664), .B2(n9008), .A(n9007), .ZN(n9009) );
  NOR2_X1 U10332 ( .A1(n4282), .A2(n9009), .ZN(n9010) );
  OAI222_X1 U10333 ( .A1(n9687), .A2(n9012), .B1(n9685), .B2(n9011), .C1(n9682), .C2(n9010), .ZN(n9212) );
  AOI211_X1 U10334 ( .C1(n9214), .C2(n9014), .A(n9786), .B(n9013), .ZN(n9213)
         );
  NAND2_X1 U10335 ( .A1(n9213), .A2(n9144), .ZN(n9018) );
  INV_X1 U10336 ( .A(n9015), .ZN(n9016) );
  AOI22_X1 U10337 ( .A1(n9016), .A2(n9714), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9715), .ZN(n9017) );
  OAI211_X1 U10338 ( .C1(n9019), .C2(n9717), .A(n9018), .B(n9017), .ZN(n9020)
         );
  AOI21_X1 U10339 ( .B1(n9212), .B2(n9719), .A(n9020), .ZN(n9021) );
  OAI21_X1 U10340 ( .B1(n9216), .B2(n9198), .A(n9021), .ZN(P1_U3263) );
  XOR2_X1 U10341 ( .A(n9024), .B(n9022), .Z(n9236) );
  AOI22_X1 U10342 ( .A1(n9234), .A2(n9539), .B1(n9715), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9034) );
  XOR2_X1 U10343 ( .A(n9024), .B(n9023), .Z(n9025) );
  OAI222_X1 U10344 ( .A1(n9687), .A2(n9027), .B1(n9685), .B2(n9026), .C1(n9682), .C2(n9025), .ZN(n9232) );
  INV_X1 U10345 ( .A(n9036), .ZN(n9029) );
  AOI211_X1 U10346 ( .C1(n9234), .C2(n9029), .A(n9786), .B(n9028), .ZN(n9233)
         );
  INV_X1 U10347 ( .A(n9233), .ZN(n9031) );
  OAI22_X1 U10348 ( .A1(n9031), .A2(n9679), .B1(n9118), .B2(n9030), .ZN(n9032)
         );
  OAI21_X1 U10349 ( .B1(n9232), .B2(n9032), .A(n9719), .ZN(n9033) );
  OAI211_X1 U10350 ( .C1(n9236), .C2(n9198), .A(n9034), .B(n9033), .ZN(
        P1_U3267) );
  XNOR2_X1 U10351 ( .A(n9035), .B(n9042), .ZN(n9241) );
  AOI21_X1 U10352 ( .B1(n9237), .B2(n9059), .A(n9036), .ZN(n9238) );
  INV_X1 U10353 ( .A(n9037), .ZN(n9038) );
  AOI22_X1 U10354 ( .A1(n9038), .A2(n9714), .B1(n9715), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9039) );
  OAI21_X1 U10355 ( .B1(n4461), .B2(n9717), .A(n9039), .ZN(n9047) );
  NAND2_X1 U10356 ( .A1(n9041), .A2(n9040), .ZN(n9043) );
  XNOR2_X1 U10357 ( .A(n9043), .B(n9042), .ZN(n9045) );
  AOI222_X1 U10358 ( .A1(n9707), .A2(n9045), .B1(n9044), .B2(n9702), .C1(n9077), .C2(n9700), .ZN(n9240) );
  NOR2_X1 U10359 ( .A1(n9240), .A2(n9715), .ZN(n9046) );
  AOI211_X1 U10360 ( .C1(n9238), .C2(n9698), .A(n9047), .B(n9046), .ZN(n9048)
         );
  OAI21_X1 U10361 ( .B1(n9241), .B2(n9198), .A(n9048), .ZN(P1_U3268) );
  XNOR2_X1 U10362 ( .A(n9049), .B(n9050), .ZN(n9246) );
  NAND2_X1 U10363 ( .A1(n9073), .A2(n9051), .ZN(n9053) );
  XNOR2_X1 U10364 ( .A(n9053), .B(n9052), .ZN(n9054) );
  NAND2_X1 U10365 ( .A1(n9054), .A2(n9707), .ZN(n9057) );
  AOI22_X1 U10366 ( .A1(n9055), .A2(n9702), .B1(n9700), .B2(n9095), .ZN(n9056)
         );
  NAND2_X1 U10367 ( .A1(n9057), .A2(n9056), .ZN(n9242) );
  INV_X1 U10368 ( .A(n9059), .ZN(n9060) );
  AOI211_X1 U10369 ( .C1(n9244), .C2(n4465), .A(n9786), .B(n9060), .ZN(n9243)
         );
  NAND2_X1 U10370 ( .A1(n9243), .A2(n9144), .ZN(n9063) );
  AOI22_X1 U10371 ( .A1(n9715), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9061), .B2(
        n9714), .ZN(n9062) );
  OAI211_X1 U10372 ( .C1(n9064), .C2(n9717), .A(n9063), .B(n9062), .ZN(n9065)
         );
  AOI21_X1 U10373 ( .B1(n9242), .B2(n9719), .A(n9065), .ZN(n9066) );
  OAI21_X1 U10374 ( .B1(n9246), .B2(n9198), .A(n9066), .ZN(P1_U3269) );
  OAI21_X1 U10375 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9251) );
  AOI211_X1 U10376 ( .C1(n9248), .C2(n9085), .A(n9786), .B(n9058), .ZN(n9247)
         );
  AOI22_X1 U10377 ( .A1(n9715), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9070), .B2(
        n9714), .ZN(n9071) );
  OAI21_X1 U10378 ( .B1(n9072), .B2(n9717), .A(n9071), .ZN(n9080) );
  OAI21_X1 U10379 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9078) );
  AOI222_X1 U10380 ( .A1(n9707), .A2(n9078), .B1(n9077), .B2(n9702), .C1(n9076), .C2(n9700), .ZN(n9250) );
  NOR2_X1 U10381 ( .A1(n9250), .A2(n9715), .ZN(n9079) );
  AOI211_X1 U10382 ( .C1(n9247), .C2(n9144), .A(n9080), .B(n9079), .ZN(n9081)
         );
  OAI21_X1 U10383 ( .B1(n9251), .B2(n9198), .A(n9081), .ZN(P1_U3270) );
  OAI21_X1 U10384 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9256) );
  INV_X1 U10385 ( .A(n9107), .ZN(n9087) );
  INV_X1 U10386 ( .A(n9085), .ZN(n9086) );
  AOI211_X1 U10387 ( .C1(n9253), .C2(n9087), .A(n9786), .B(n9086), .ZN(n9252)
         );
  AOI22_X1 U10388 ( .A1(n9715), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9088), .B2(
        n9714), .ZN(n9089) );
  OAI21_X1 U10389 ( .B1(n9090), .B2(n9717), .A(n9089), .ZN(n9098) );
  OAI21_X1 U10390 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9096) );
  AOI222_X1 U10391 ( .A1(n9707), .A2(n9096), .B1(n9095), .B2(n9702), .C1(n9094), .C2(n9700), .ZN(n9255) );
  NOR2_X1 U10392 ( .A1(n9255), .A2(n9715), .ZN(n9097) );
  AOI211_X1 U10393 ( .C1(n9252), .C2(n9144), .A(n9098), .B(n9097), .ZN(n9099)
         );
  OAI21_X1 U10394 ( .B1(n9256), .B2(n9198), .A(n9099), .ZN(P1_U3271) );
  OAI21_X1 U10395 ( .B1(n9101), .B2(n9103), .A(n9100), .ZN(n9261) );
  AOI21_X1 U10396 ( .B1(n9103), .B2(n9102), .A(n4298), .ZN(n9104) );
  OAI222_X1 U10397 ( .A1(n9687), .A2(n9106), .B1(n9685), .B2(n9105), .C1(n9682), .C2(n9104), .ZN(n9257) );
  INV_X1 U10398 ( .A(n9115), .ZN(n9108) );
  AOI211_X1 U10399 ( .C1(n9259), .C2(n9108), .A(n9786), .B(n9107), .ZN(n9258)
         );
  NAND2_X1 U10400 ( .A1(n9258), .A2(n9144), .ZN(n9111) );
  AOI22_X1 U10401 ( .A1(n9715), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9109), .B2(
        n9714), .ZN(n9110) );
  OAI211_X1 U10402 ( .C1(n9112), .C2(n9717), .A(n9111), .B(n9110), .ZN(n9113)
         );
  AOI21_X1 U10403 ( .B1(n9257), .B2(n9719), .A(n9113), .ZN(n9114) );
  OAI21_X1 U10404 ( .B1(n9261), .B2(n9198), .A(n9114), .ZN(P1_U3272) );
  AOI211_X1 U10405 ( .C1(n9266), .C2(n9142), .A(n9786), .B(n9115), .ZN(n9265)
         );
  INV_X1 U10406 ( .A(n9116), .ZN(n9117) );
  NOR2_X1 U10407 ( .A1(n9118), .A2(n9117), .ZN(n9124) );
  INV_X1 U10408 ( .A(n9135), .ZN(n9119) );
  NOR2_X1 U10409 ( .A1(n9134), .A2(n9119), .ZN(n9140) );
  NOR2_X1 U10410 ( .A1(n9140), .A2(n9120), .ZN(n9121) );
  XNOR2_X1 U10411 ( .A(n9121), .B(n9126), .ZN(n9122) );
  OAI222_X1 U10412 ( .A1(n9687), .A2(n9123), .B1(n9685), .B2(n9156), .C1(n9682), .C2(n9122), .ZN(n9264) );
  AOI211_X1 U10413 ( .C1(n9265), .C2(n9125), .A(n9124), .B(n9264), .ZN(n9131)
         );
  OR2_X1 U10414 ( .A1(n9127), .A2(n9126), .ZN(n9263) );
  NAND3_X1 U10415 ( .A1(n9263), .A2(n9262), .A3(n9128), .ZN(n9130) );
  AOI22_X1 U10416 ( .A1(n9266), .A2(n9539), .B1(n9715), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9129) );
  OAI211_X1 U10417 ( .C1(n9715), .C2(n9131), .A(n9130), .B(n9129), .ZN(
        P1_U3273) );
  AOI21_X1 U10418 ( .B1(n9135), .B2(n9133), .A(n9132), .ZN(n9273) );
  INV_X1 U10419 ( .A(n9134), .ZN(n9136) );
  OAI21_X1 U10420 ( .B1(n9136), .B2(n9135), .A(n9707), .ZN(n9141) );
  AOI22_X1 U10421 ( .A1(n9700), .A2(n9138), .B1(n9137), .B2(n9702), .ZN(n9139)
         );
  OAI21_X1 U10422 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9269) );
  INV_X1 U10423 ( .A(n9142), .ZN(n9143) );
  AOI211_X1 U10424 ( .C1(n9271), .C2(n9157), .A(n9786), .B(n9143), .ZN(n9270)
         );
  NAND2_X1 U10425 ( .A1(n9270), .A2(n9144), .ZN(n9147) );
  AOI22_X1 U10426 ( .A1(n9715), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9145), .B2(
        n9714), .ZN(n9146) );
  OAI211_X1 U10427 ( .C1(n9148), .C2(n9717), .A(n9147), .B(n9146), .ZN(n9149)
         );
  AOI21_X1 U10428 ( .B1(n9269), .B2(n9719), .A(n9149), .ZN(n9150) );
  OAI21_X1 U10429 ( .B1(n9273), .B2(n9198), .A(n9150), .ZN(P1_U3274) );
  OAI21_X1 U10430 ( .B1(n9152), .B2(n9153), .A(n9151), .ZN(n9278) );
  XNOR2_X1 U10431 ( .A(n9154), .B(n9153), .ZN(n9155) );
  OAI222_X1 U10432 ( .A1(n9687), .A2(n9156), .B1(n9685), .B2(n9189), .C1(n9155), .C2(n9682), .ZN(n9274) );
  INV_X1 U10433 ( .A(n9157), .ZN(n9158) );
  AOI211_X1 U10434 ( .C1(n9276), .C2(n4319), .A(n9786), .B(n9158), .ZN(n9275)
         );
  NAND2_X1 U10435 ( .A1(n9275), .A2(n9191), .ZN(n9161) );
  AOI22_X1 U10436 ( .A1(n9715), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9159), .B2(
        n9714), .ZN(n9160) );
  OAI211_X1 U10437 ( .C1(n9162), .C2(n9717), .A(n9161), .B(n9160), .ZN(n9163)
         );
  AOI21_X1 U10438 ( .B1(n9274), .B2(n9719), .A(n9163), .ZN(n9164) );
  OAI21_X1 U10439 ( .B1(n9278), .B2(n9198), .A(n9164), .ZN(P1_U3275) );
  OAI21_X1 U10440 ( .B1(n9166), .B2(n9167), .A(n9165), .ZN(n9283) );
  INV_X1 U10441 ( .A(n9283), .ZN(n9175) );
  NAND2_X1 U10442 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  AOI21_X1 U10443 ( .B1(n9170), .B2(n9169), .A(n9682), .ZN(n9174) );
  OAI22_X1 U10444 ( .A1(n9172), .A2(n9685), .B1(n9171), .B2(n9687), .ZN(n9173)
         );
  AOI211_X1 U10445 ( .C1(n9175), .C2(n9537), .A(n9174), .B(n9173), .ZN(n9282)
         );
  XNOR2_X1 U10446 ( .A(n9190), .B(n9279), .ZN(n9280) );
  AOI22_X1 U10447 ( .A1(n9715), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9176), .B2(
        n9714), .ZN(n9177) );
  OAI21_X1 U10448 ( .B1(n9178), .B2(n9717), .A(n9177), .ZN(n9181) );
  NOR2_X1 U10449 ( .A1(n9283), .A2(n9179), .ZN(n9180) );
  AOI211_X1 U10450 ( .C1(n9280), .C2(n9698), .A(n9181), .B(n9180), .ZN(n9182)
         );
  OAI21_X1 U10451 ( .B1(n9715), .B2(n9282), .A(n9182), .ZN(P1_U3276) );
  XOR2_X1 U10452 ( .A(n9183), .B(n9185), .Z(n9289) );
  NAND2_X1 U10453 ( .A1(n9513), .A2(n9184), .ZN(n9186) );
  XNOR2_X1 U10454 ( .A(n9186), .B(n9185), .ZN(n9187) );
  OAI222_X1 U10455 ( .A1(n9687), .A2(n9189), .B1(n9685), .B2(n9188), .C1(n9187), .C2(n9682), .ZN(n9284) );
  AOI211_X1 U10456 ( .C1(n9286), .C2(n9524), .A(n9786), .B(n9190), .ZN(n9285)
         );
  NAND2_X1 U10457 ( .A1(n9285), .A2(n9191), .ZN(n9194) );
  AOI22_X1 U10458 ( .A1(n9715), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9192), .B2(
        n9714), .ZN(n9193) );
  OAI211_X1 U10459 ( .C1(n9195), .C2(n9717), .A(n9194), .B(n9193), .ZN(n9196)
         );
  AOI21_X1 U10460 ( .B1(n9284), .B2(n9719), .A(n9196), .ZN(n9197) );
  OAI21_X1 U10461 ( .B1(n9289), .B2(n9198), .A(n9197), .ZN(P1_U3277) );
  AOI21_X1 U10462 ( .B1(n9199), .B2(n9777), .A(n9202), .ZN(n9200) );
  OAI21_X1 U10463 ( .B1(n9201), .B2(n9786), .A(n9200), .ZN(n9291) );
  MUX2_X1 U10464 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9291), .S(n9811), .Z(
        P1_U3554) );
  AOI21_X1 U10465 ( .B1(n9203), .B2(n9777), .A(n9202), .ZN(n9204) );
  OAI21_X1 U10466 ( .B1(n9205), .B2(n9786), .A(n9204), .ZN(n9292) );
  MUX2_X1 U10467 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9292), .S(n9811), .Z(
        P1_U3553) );
  NAND2_X1 U10468 ( .A1(n9206), .A2(n9790), .ZN(n9211) );
  NAND2_X1 U10469 ( .A1(n9211), .A2(n9210), .ZN(n9293) );
  MUX2_X1 U10470 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9293), .S(n9811), .Z(
        P1_U3552) );
  OAI21_X1 U10471 ( .B1(n9216), .B2(n9288), .A(n9215), .ZN(n9294) );
  MUX2_X1 U10472 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9294), .S(n9811), .Z(
        P1_U3551) );
  AOI22_X1 U10473 ( .A1(n9218), .A2(n9778), .B1(n9777), .B2(n9217), .ZN(n9219)
         );
  OAI211_X1 U10474 ( .C1(n9221), .C2(n9288), .A(n9220), .B(n9219), .ZN(n9295)
         );
  MUX2_X1 U10475 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9295), .S(n9811), .Z(
        P1_U3550) );
  AOI22_X1 U10476 ( .A1(n9223), .A2(n9778), .B1(n9777), .B2(n9222), .ZN(n9224)
         );
  OAI211_X1 U10477 ( .C1(n9226), .C2(n9288), .A(n9225), .B(n9224), .ZN(n9296)
         );
  MUX2_X1 U10478 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9296), .S(n9811), .Z(
        P1_U3549) );
  AOI22_X1 U10479 ( .A1(n9228), .A2(n9778), .B1(n9777), .B2(n9227), .ZN(n9229)
         );
  OAI211_X1 U10480 ( .C1(n9231), .C2(n9288), .A(n9230), .B(n9229), .ZN(n9297)
         );
  MUX2_X1 U10481 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9297), .S(n9811), .Z(
        P1_U3548) );
  AOI211_X1 U10482 ( .C1(n9777), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9235)
         );
  OAI21_X1 U10483 ( .B1(n9236), .B2(n9288), .A(n9235), .ZN(n9298) );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9298), .S(n9811), .Z(
        P1_U3547) );
  AOI22_X1 U10485 ( .A1(n9238), .A2(n9778), .B1(n9777), .B2(n9237), .ZN(n9239)
         );
  OAI211_X1 U10486 ( .C1(n9241), .C2(n9288), .A(n9240), .B(n9239), .ZN(n9299)
         );
  MUX2_X1 U10487 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9299), .S(n9811), .Z(
        P1_U3546) );
  AOI211_X1 U10488 ( .C1(n9777), .C2(n9244), .A(n9243), .B(n9242), .ZN(n9245)
         );
  OAI21_X1 U10489 ( .B1(n9246), .B2(n9288), .A(n9245), .ZN(n9300) );
  MUX2_X1 U10490 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9300), .S(n9811), .Z(
        P1_U3545) );
  AOI21_X1 U10491 ( .B1(n9777), .B2(n9248), .A(n9247), .ZN(n9249) );
  OAI211_X1 U10492 ( .C1(n9251), .C2(n9288), .A(n9250), .B(n9249), .ZN(n9449)
         );
  MUX2_X1 U10493 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9449), .S(n9811), .Z(
        P1_U3544) );
  AOI21_X1 U10494 ( .B1(n9777), .B2(n9253), .A(n9252), .ZN(n9254) );
  OAI211_X1 U10495 ( .C1(n9256), .C2(n9288), .A(n9255), .B(n9254), .ZN(n9450)
         );
  MUX2_X1 U10496 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9450), .S(n9811), .Z(
        P1_U3543) );
  AOI211_X1 U10497 ( .C1(n9777), .C2(n9259), .A(n9258), .B(n9257), .ZN(n9260)
         );
  OAI21_X1 U10498 ( .B1(n9261), .B2(n9288), .A(n9260), .ZN(n9451) );
  MUX2_X1 U10499 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9451), .S(n9811), .Z(
        P1_U3542) );
  NAND3_X1 U10500 ( .A1(n9263), .A2(n9262), .A3(n9790), .ZN(n9268) );
  AOI211_X1 U10501 ( .C1(n9777), .C2(n9266), .A(n9265), .B(n9264), .ZN(n9267)
         );
  NAND2_X1 U10502 ( .A1(n9268), .A2(n9267), .ZN(n9452) );
  MUX2_X1 U10503 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9452), .S(n9811), .Z(
        P1_U3541) );
  AOI211_X1 U10504 ( .C1(n9777), .C2(n9271), .A(n9270), .B(n9269), .ZN(n9272)
         );
  OAI21_X1 U10505 ( .B1(n9273), .B2(n9288), .A(n9272), .ZN(n9453) );
  MUX2_X1 U10506 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9453), .S(n9811), .Z(
        P1_U3540) );
  AOI211_X1 U10507 ( .C1(n9777), .C2(n9276), .A(n9275), .B(n9274), .ZN(n9277)
         );
  OAI21_X1 U10508 ( .B1(n9278), .B2(n9288), .A(n9277), .ZN(n9454) );
  MUX2_X1 U10509 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9454), .S(n9811), .Z(
        P1_U3539) );
  AOI22_X1 U10510 ( .A1(n9280), .A2(n9778), .B1(n9777), .B2(n9279), .ZN(n9281)
         );
  OAI211_X1 U10511 ( .C1(n9730), .C2(n9283), .A(n9282), .B(n9281), .ZN(n9455)
         );
  MUX2_X1 U10512 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9455), .S(n9811), .Z(
        P1_U3538) );
  AOI211_X1 U10513 ( .C1(n9777), .C2(n9286), .A(n9285), .B(n9284), .ZN(n9287)
         );
  OAI21_X1 U10514 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9456) );
  MUX2_X1 U10515 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9456), .S(n9811), .Z(
        P1_U3537) );
  MUX2_X1 U10516 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9290), .S(n9811), .Z(
        P1_U3523) );
  MUX2_X1 U10517 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9291), .S(n9794), .Z(
        P1_U3522) );
  MUX2_X1 U10518 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9292), .S(n9794), .Z(
        P1_U3521) );
  MUX2_X1 U10519 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9293), .S(n9794), .Z(
        P1_U3520) );
  MUX2_X1 U10520 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9294), .S(n9794), .Z(
        P1_U3519) );
  MUX2_X1 U10521 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9295), .S(n9794), .Z(
        P1_U3518) );
  MUX2_X1 U10522 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9296), .S(n9794), .Z(
        P1_U3517) );
  MUX2_X1 U10523 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9297), .S(n9794), .Z(
        P1_U3516) );
  MUX2_X1 U10524 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9298), .S(n9794), .Z(
        P1_U3515) );
  MUX2_X1 U10525 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9299), .S(n9794), .Z(
        P1_U3514) );
  MUX2_X1 U10526 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9300), .S(n9794), .Z(n9448) );
  INV_X1 U10527 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U10528 ( .A1(n9856), .A2(keyinput36), .B1(keyinput63), .B2(n9302), 
        .ZN(n9301) );
  OAI221_X1 U10529 ( .B1(n9856), .B2(keyinput36), .C1(n9302), .C2(keyinput63), 
        .A(n9301), .ZN(n9312) );
  INV_X1 U10530 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9852) );
  INV_X1 U10531 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9304) );
  AOI22_X1 U10532 ( .A1(n9852), .A2(keyinput60), .B1(keyinput44), .B2(n9304), 
        .ZN(n9303) );
  OAI221_X1 U10533 ( .B1(n9852), .B2(keyinput60), .C1(n9304), .C2(keyinput44), 
        .A(n9303), .ZN(n9311) );
  INV_X1 U10534 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9306) );
  AOI22_X1 U10535 ( .A1(n9307), .A2(keyinput3), .B1(n9306), .B2(keyinput17), 
        .ZN(n9305) );
  OAI221_X1 U10536 ( .B1(n9307), .B2(keyinput3), .C1(n9306), .C2(keyinput17), 
        .A(n9305), .ZN(n9310) );
  INV_X1 U10537 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9722) );
  AOI22_X1 U10538 ( .A1(n9722), .A2(keyinput7), .B1(keyinput25), .B2(n9805), 
        .ZN(n9308) );
  OAI221_X1 U10539 ( .B1(n9722), .B2(keyinput7), .C1(n9805), .C2(keyinput25), 
        .A(n9308), .ZN(n9309) );
  NOR4_X1 U10540 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9341)
         );
  INV_X1 U10541 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9723) );
  AOI22_X1 U10542 ( .A1(n9813), .A2(keyinput15), .B1(n9723), .B2(keyinput49), 
        .ZN(n9313) );
  OAI221_X1 U10543 ( .B1(n9813), .B2(keyinput15), .C1(n9723), .C2(keyinput49), 
        .A(n9313), .ZN(n9325) );
  INV_X1 U10544 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9854) );
  INV_X1 U10545 ( .A(keyinput57), .ZN(n9315) );
  AOI22_X1 U10546 ( .A1(n9854), .A2(keyinput37), .B1(P1_ADDR_REG_8__SCAN_IN), 
        .B2(n9315), .ZN(n9314) );
  OAI221_X1 U10547 ( .B1(n9854), .B2(keyinput37), .C1(n9315), .C2(
        P1_ADDR_REG_8__SCAN_IN), .A(n9314), .ZN(n9324) );
  INV_X1 U10548 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9317) );
  AOI22_X1 U10549 ( .A1(n9318), .A2(keyinput0), .B1(keyinput61), .B2(n9317), 
        .ZN(n9316) );
  OAI221_X1 U10550 ( .B1(n9318), .B2(keyinput0), .C1(n9317), .C2(keyinput61), 
        .A(n9316), .ZN(n9323) );
  AOI22_X1 U10551 ( .A1(n9321), .A2(keyinput4), .B1(n9320), .B2(keyinput21), 
        .ZN(n9319) );
  OAI221_X1 U10552 ( .B1(n9321), .B2(keyinput4), .C1(n9320), .C2(keyinput21), 
        .A(n9319), .ZN(n9322) );
  NOR4_X1 U10553 ( .A1(n9325), .A2(n9324), .A3(n9323), .A4(n9322), .ZN(n9340)
         );
  INV_X1 U10554 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10555 ( .A1(n9851), .A2(keyinput53), .B1(n9327), .B2(keyinput55), 
        .ZN(n9326) );
  OAI221_X1 U10556 ( .B1(n9851), .B2(keyinput53), .C1(n9327), .C2(keyinput55), 
        .A(n9326), .ZN(n9338) );
  INV_X1 U10557 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9329) );
  AOI22_X1 U10558 ( .A1(n9330), .A2(keyinput1), .B1(keyinput18), .B2(n9329), 
        .ZN(n9328) );
  OAI221_X1 U10559 ( .B1(n9330), .B2(keyinput1), .C1(n9329), .C2(keyinput18), 
        .A(n9328), .ZN(n9337) );
  INV_X1 U10560 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9333) );
  AOI22_X1 U10561 ( .A1(n9333), .A2(keyinput11), .B1(keyinput43), .B2(n9332), 
        .ZN(n9331) );
  OAI221_X1 U10562 ( .B1(n9333), .B2(keyinput11), .C1(n9332), .C2(keyinput43), 
        .A(n9331), .ZN(n9336) );
  INV_X1 U10563 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10564 ( .A1(n6605), .A2(keyinput47), .B1(n9853), .B2(keyinput50), 
        .ZN(n9334) );
  OAI221_X1 U10565 ( .B1(n6605), .B2(keyinput47), .C1(n9853), .C2(keyinput50), 
        .A(n9334), .ZN(n9335) );
  NOR4_X1 U10566 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n9339)
         );
  AND3_X1 U10567 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9446) );
  INV_X1 U10568 ( .A(keyinput54), .ZN(n9343) );
  AOI22_X1 U10569 ( .A1(n4979), .A2(keyinput32), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n9343), .ZN(n9342) );
  OAI221_X1 U10570 ( .B1(n4979), .B2(keyinput32), .C1(n9343), .C2(
        P1_ADDR_REG_18__SCAN_IN), .A(n9342), .ZN(n9355) );
  INV_X1 U10571 ( .A(keyinput9), .ZN(n9345) );
  AOI22_X1 U10572 ( .A1(n9346), .A2(keyinput2), .B1(P1_ADDR_REG_0__SCAN_IN), 
        .B2(n9345), .ZN(n9344) );
  OAI221_X1 U10573 ( .B1(n9346), .B2(keyinput2), .C1(n9345), .C2(
        P1_ADDR_REG_0__SCAN_IN), .A(n9344), .ZN(n9354) );
  INV_X1 U10574 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9349) );
  AOI22_X1 U10575 ( .A1(n9349), .A2(keyinput12), .B1(n9348), .B2(keyinput14), 
        .ZN(n9347) );
  OAI221_X1 U10576 ( .B1(n9349), .B2(keyinput12), .C1(n9348), .C2(keyinput14), 
        .A(n9347), .ZN(n9353) );
  AOI22_X1 U10577 ( .A1(n9351), .A2(keyinput29), .B1(keyinput23), .B2(n6085), 
        .ZN(n9350) );
  OAI221_X1 U10578 ( .B1(n9351), .B2(keyinput29), .C1(n6085), .C2(keyinput23), 
        .A(n9350), .ZN(n9352) );
  NOR4_X1 U10579 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9445)
         );
  INV_X1 U10580 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9358) );
  AOI22_X1 U10581 ( .A1(n9358), .A2(keyinput51), .B1(n9357), .B2(keyinput38), 
        .ZN(n9356) );
  OAI221_X1 U10582 ( .B1(n9358), .B2(keyinput51), .C1(n9357), .C2(keyinput38), 
        .A(n9356), .ZN(n9370) );
  INV_X1 U10583 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9360) );
  AOI22_X1 U10584 ( .A1(n7003), .A2(keyinput20), .B1(n9360), .B2(keyinput48), 
        .ZN(n9359) );
  OAI221_X1 U10585 ( .B1(n7003), .B2(keyinput20), .C1(n9360), .C2(keyinput48), 
        .A(n9359), .ZN(n9369) );
  INV_X1 U10586 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9363) );
  AOI22_X1 U10587 ( .A1(n9363), .A2(keyinput31), .B1(keyinput19), .B2(n9362), 
        .ZN(n9361) );
  OAI221_X1 U10588 ( .B1(n9363), .B2(keyinput31), .C1(n9362), .C2(keyinput19), 
        .A(n9361), .ZN(n9368) );
  AOI22_X1 U10589 ( .A1(n9366), .A2(keyinput62), .B1(keyinput24), .B2(n9365), 
        .ZN(n9364) );
  OAI221_X1 U10590 ( .B1(n9366), .B2(keyinput62), .C1(n9365), .C2(keyinput24), 
        .A(n9364), .ZN(n9367) );
  NOR4_X1 U10591 ( .A1(n9370), .A2(n9369), .A3(n9368), .A4(n9367), .ZN(n9444)
         );
  NOR2_X1 U10592 ( .A1(keyinput61), .A2(keyinput4), .ZN(n9374) );
  NAND3_X1 U10593 ( .A1(keyinput36), .A2(keyinput63), .A3(keyinput60), .ZN(
        n9372) );
  NAND3_X1 U10594 ( .A1(keyinput17), .A2(keyinput7), .A3(keyinput25), .ZN(
        n9371) );
  NOR4_X1 U10595 ( .A1(keyinput44), .A2(keyinput3), .A3(n9372), .A4(n9371), 
        .ZN(n9373) );
  NAND4_X1 U10596 ( .A1(keyinput0), .A2(keyinput21), .A3(n9374), .A4(n9373), 
        .ZN(n9384) );
  NOR2_X1 U10597 ( .A1(keyinput35), .A2(keyinput41), .ZN(n9376) );
  NOR4_X1 U10598 ( .A1(keyinput1), .A2(keyinput18), .A3(keyinput53), .A4(
        keyinput55), .ZN(n9375) );
  NAND4_X1 U10599 ( .A1(keyinput45), .A2(keyinput28), .A3(n9376), .A4(n9375), 
        .ZN(n9383) );
  NOR2_X1 U10600 ( .A1(keyinput15), .A2(keyinput49), .ZN(n9377) );
  NAND3_X1 U10601 ( .A1(keyinput57), .A2(keyinput37), .A3(n9377), .ZN(n9381)
         );
  INV_X1 U10602 ( .A(keyinput50), .ZN(n9378) );
  NAND4_X1 U10603 ( .A1(keyinput47), .A2(keyinput11), .A3(keyinput43), .A4(
        n9378), .ZN(n9380) );
  NAND3_X1 U10604 ( .A1(keyinput27), .A2(keyinput16), .A3(keyinput10), .ZN(
        n9379) );
  OR4_X1 U10605 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(keyinput8), .ZN(
        n9382) );
  NOR3_X1 U10606 ( .A1(n9384), .A2(n9383), .A3(n9382), .ZN(n9442) );
  NOR2_X1 U10607 ( .A1(keyinput33), .A2(keyinput13), .ZN(n9389) );
  NAND3_X1 U10608 ( .A1(keyinput46), .A2(keyinput56), .A3(keyinput5), .ZN(
        n9387) );
  NAND4_X1 U10609 ( .A1(keyinput54), .A2(keyinput32), .A3(keyinput9), .A4(
        keyinput2), .ZN(n9386) );
  NAND4_X1 U10610 ( .A1(keyinput12), .A2(keyinput14), .A3(keyinput29), .A4(
        keyinput23), .ZN(n9385) );
  NOR4_X1 U10611 ( .A1(keyinput59), .A2(n9387), .A3(n9386), .A4(n9385), .ZN(
        n9388) );
  NAND4_X1 U10612 ( .A1(keyinput52), .A2(keyinput6), .A3(n9389), .A4(n9388), 
        .ZN(n9397) );
  NOR3_X1 U10613 ( .A1(keyinput62), .A2(keyinput24), .A3(keyinput19), .ZN(
        n9395) );
  NAND2_X1 U10614 ( .A1(keyinput26), .A2(keyinput39), .ZN(n9390) );
  NOR3_X1 U10615 ( .A1(keyinput58), .A2(keyinput34), .A3(n9390), .ZN(n9394) );
  NAND3_X1 U10616 ( .A1(keyinput20), .A2(keyinput48), .A3(keyinput51), .ZN(
        n9392) );
  NAND3_X1 U10617 ( .A1(keyinput22), .A2(keyinput40), .A3(keyinput42), .ZN(
        n9391) );
  NOR4_X1 U10618 ( .A1(keyinput38), .A2(keyinput30), .A3(n9392), .A4(n9391), 
        .ZN(n9393) );
  NAND4_X1 U10619 ( .A1(keyinput31), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(
        n9396) );
  NOR2_X1 U10620 ( .A1(n9397), .A2(n9396), .ZN(n9441) );
  INV_X1 U10621 ( .A(SI_17_), .ZN(n9399) );
  AOI22_X1 U10622 ( .A1(n9399), .A2(keyinput30), .B1(keyinput42), .B2(n6222), 
        .ZN(n9398) );
  OAI221_X1 U10623 ( .B1(n9399), .B2(keyinput30), .C1(n6222), .C2(keyinput42), 
        .A(n9398), .ZN(n9407) );
  INV_X1 U10624 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9855) );
  INV_X1 U10625 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9401) );
  AOI22_X1 U10626 ( .A1(n9855), .A2(keyinput58), .B1(keyinput39), .B2(n9401), 
        .ZN(n9400) );
  OAI221_X1 U10627 ( .B1(n9855), .B2(keyinput58), .C1(n9401), .C2(keyinput39), 
        .A(n9400), .ZN(n9406) );
  AOI22_X1 U10628 ( .A1(n9404), .A2(keyinput45), .B1(n9403), .B2(keyinput35), 
        .ZN(n9402) );
  OAI221_X1 U10629 ( .B1(n9404), .B2(keyinput45), .C1(n9403), .C2(keyinput35), 
        .A(n9402), .ZN(n9405) );
  NOR3_X1 U10630 ( .A1(n9407), .A2(n9406), .A3(n9405), .ZN(n9439) );
  AOI22_X1 U10631 ( .A1(n9409), .A2(keyinput16), .B1(keyinput10), .B2(n5078), 
        .ZN(n9408) );
  OAI221_X1 U10632 ( .B1(n9409), .B2(keyinput16), .C1(n5078), .C2(keyinput10), 
        .A(n9408), .ZN(n9418) );
  AOI22_X1 U10633 ( .A1(n9412), .A2(keyinput26), .B1(n9411), .B2(keyinput34), 
        .ZN(n9410) );
  OAI221_X1 U10634 ( .B1(n9412), .B2(keyinput26), .C1(n9411), .C2(keyinput34), 
        .A(n9410), .ZN(n9417) );
  AOI22_X1 U10635 ( .A1(n9415), .A2(keyinput8), .B1(n9414), .B2(keyinput27), 
        .ZN(n9413) );
  OAI221_X1 U10636 ( .B1(n9415), .B2(keyinput8), .C1(n9414), .C2(keyinput27), 
        .A(n9413), .ZN(n9416) );
  NOR3_X1 U10637 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9438) );
  XNOR2_X1 U10638 ( .A(SI_2_), .B(keyinput56), .ZN(n9422) );
  XNOR2_X1 U10639 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput5), .ZN(n9421) );
  XNOR2_X1 U10640 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput33), .ZN(n9420) );
  XNOR2_X1 U10641 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput40), .ZN(n9419) );
  NAND4_X1 U10642 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n9428)
         );
  XNOR2_X1 U10643 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput13), .ZN(n9426) );
  XNOR2_X1 U10644 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput41), .ZN(n9425) );
  XNOR2_X1 U10645 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput22), .ZN(n9424) );
  XNOR2_X1 U10646 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput28), .ZN(n9423) );
  NAND4_X1 U10647 ( .A1(n9426), .A2(n9425), .A3(n9424), .A4(n9423), .ZN(n9427)
         );
  NOR2_X1 U10648 ( .A1(n9428), .A2(n9427), .ZN(n9437) );
  AOI22_X1 U10649 ( .A1(n9431), .A2(keyinput46), .B1(keyinput59), .B2(n9430), 
        .ZN(n9429) );
  OAI221_X1 U10650 ( .B1(n9431), .B2(keyinput46), .C1(n9430), .C2(keyinput59), 
        .A(n9429), .ZN(n9435) );
  AOI22_X1 U10651 ( .A1(n5816), .A2(keyinput52), .B1(n9433), .B2(keyinput6), 
        .ZN(n9432) );
  OAI221_X1 U10652 ( .B1(n5816), .B2(keyinput52), .C1(n9433), .C2(keyinput6), 
        .A(n9432), .ZN(n9434) );
  NOR2_X1 U10653 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  NAND4_X1 U10654 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n9440)
         );
  AOI21_X1 U10655 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9443) );
  NAND4_X1 U10656 ( .A1(n9446), .A2(n9445), .A3(n9444), .A4(n9443), .ZN(n9447)
         );
  XNOR2_X1 U10657 ( .A(n9448), .B(n9447), .ZN(P1_U3513) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9449), .S(n9794), .Z(
        P1_U3512) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9450), .S(n9794), .Z(
        P1_U3511) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9451), .S(n9794), .Z(
        P1_U3510) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9452), .S(n9794), .Z(
        P1_U3508) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9453), .S(n9794), .Z(
        P1_U3505) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9454), .S(n9794), .Z(
        P1_U3502) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9455), .S(n9794), .Z(
        P1_U3499) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9456), .S(n9794), .Z(
        P1_U3496) );
  NOR4_X1 U10666 ( .A1(n5654), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n6206), .ZN(n9457) );
  AOI21_X1 U10667 ( .B1(n4244), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9457), .ZN(
        n9458) );
  OAI21_X1 U10668 ( .B1(n9459), .B2(n9464), .A(n9458), .ZN(P1_U3322) );
  INV_X1 U10669 ( .A(n9460), .ZN(n9465) );
  AOI21_X1 U10670 ( .B1(n4244), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9461), .ZN(
        n9463) );
  OAI21_X1 U10671 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(P1_U3325) );
  INV_X1 U10672 ( .A(n9466), .ZN(n9467) );
  MUX2_X1 U10673 ( .A(n9467), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NAND2_X1 U10674 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9469) );
  AOI21_X1 U10675 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(n9471) );
  NAND2_X1 U10676 ( .A1(n9814), .A2(n9471), .ZN(n9475) );
  OAI22_X1 U10677 ( .A1(n9472), .A2(n9948), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4872), .ZN(n9473) );
  INV_X1 U10678 ( .A(n9473), .ZN(n9474) );
  OAI211_X1 U10679 ( .C1(n9815), .C2(n9476), .A(n9475), .B(n9474), .ZN(n9477)
         );
  INV_X1 U10680 ( .A(n9477), .ZN(n9482) );
  INV_X1 U10681 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U10682 ( .A1(n9823), .A2(n9928), .ZN(n9480) );
  OAI211_X1 U10683 ( .C1(n9480), .C2(n9479), .A(n9812), .B(n9478), .ZN(n9481)
         );
  NAND2_X1 U10684 ( .A1(n9482), .A2(n9481), .ZN(P2_U3246) );
  AOI22_X1 U10685 ( .A1(n9820), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9495) );
  AOI211_X1 U10686 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9487)
         );
  AOI21_X1 U10687 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9494) );
  OAI211_X1 U10688 ( .C1(n9492), .C2(n9491), .A(n9812), .B(n9490), .ZN(n9493)
         );
  NAND3_X1 U10689 ( .A1(n9495), .A2(n9494), .A3(n9493), .ZN(P2_U3247) );
  OAI21_X1 U10690 ( .B1(n9497), .B2(n9919), .A(n9496), .ZN(n9498) );
  AOI21_X1 U10691 ( .B1(n9499), .B2(n9899), .A(n9498), .ZN(n9507) );
  AOI22_X1 U10692 ( .A1(n9943), .A2(n9507), .B1(n5412), .B2(n9940), .ZN(
        P2_U3550) );
  OAI22_X1 U10693 ( .A1(n9501), .A2(n9921), .B1(n9500), .B2(n9919), .ZN(n9503)
         );
  AOI211_X1 U10694 ( .C1(n9925), .C2(n9504), .A(n9503), .B(n9502), .ZN(n9509)
         );
  AOI22_X1 U10695 ( .A1(n9943), .A2(n9509), .B1(n9505), .B2(n9940), .ZN(
        P2_U3534) );
  INV_X1 U10696 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U10697 ( .A1(n9912), .A2(n9507), .B1(n9506), .B2(n9927), .ZN(
        P2_U3518) );
  INV_X1 U10698 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U10699 ( .A1(n9912), .A2(n9509), .B1(n9508), .B2(n9927), .ZN(
        P2_U3493) );
  OAI21_X1 U10700 ( .B1(n9512), .B2(n9511), .A(n9510), .ZN(n9553) );
  OAI21_X1 U10701 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(n9516) );
  NAND2_X1 U10702 ( .A1(n9516), .A2(n9707), .ZN(n9520) );
  AOI22_X1 U10703 ( .A1(n9702), .A2(n9518), .B1(n9517), .B2(n9700), .ZN(n9519)
         );
  NAND2_X1 U10704 ( .A1(n9520), .A2(n9519), .ZN(n9552) );
  AOI21_X1 U10705 ( .B1(n9553), .B2(n9537), .A(n9552), .ZN(n9529) );
  AOI222_X1 U10706 ( .A1(n9522), .A2(n9539), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9715), .C1(n9714), .C2(n9521), .ZN(n9528) );
  INV_X1 U10707 ( .A(n9523), .ZN(n9525) );
  INV_X1 U10708 ( .A(n9550), .ZN(n9526) );
  AOI22_X1 U10709 ( .A1(n9553), .A2(n9699), .B1(n9698), .B2(n9526), .ZN(n9527)
         );
  OAI211_X1 U10710 ( .C1(n9715), .C2(n9529), .A(n9528), .B(n9527), .ZN(
        P1_U3278) );
  XNOR2_X1 U10711 ( .A(n9531), .B(n9530), .ZN(n9565) );
  XNOR2_X1 U10712 ( .A(n9533), .B(n9532), .ZN(n9534) );
  OAI222_X1 U10713 ( .A1(n9685), .A2(n9536), .B1(n9687), .B2(n9535), .C1(n9534), .C2(n9682), .ZN(n9564) );
  AOI21_X1 U10714 ( .B1(n9565), .B2(n9537), .A(n9564), .ZN(n9548) );
  AOI222_X1 U10715 ( .A1(n9540), .A2(n9539), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9715), .C1(n9714), .C2(n9538), .ZN(n9547) );
  INV_X1 U10716 ( .A(n9541), .ZN(n9544) );
  INV_X1 U10717 ( .A(n9542), .ZN(n9543) );
  OAI21_X1 U10718 ( .B1(n9561), .B2(n9544), .A(n9543), .ZN(n9562) );
  INV_X1 U10719 ( .A(n9562), .ZN(n9545) );
  AOI22_X1 U10720 ( .A1(n9565), .A2(n9699), .B1(n9698), .B2(n9545), .ZN(n9546)
         );
  OAI211_X1 U10721 ( .C1(n9715), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3280) );
  OAI22_X1 U10722 ( .A1(n9550), .A2(n9786), .B1(n9549), .B2(n9784), .ZN(n9551)
         );
  AOI211_X1 U10723 ( .C1(n9553), .C2(n9790), .A(n9552), .B(n9551), .ZN(n9568)
         );
  AOI22_X1 U10724 ( .A1(n9811), .A2(n9568), .B1(n9554), .B2(n9809), .ZN(
        P1_U3536) );
  OAI211_X1 U10725 ( .C1(n9557), .C2(n9784), .A(n9556), .B(n9555), .ZN(n9558)
         );
  AOI21_X1 U10726 ( .B1(n9559), .B2(n9790), .A(n9558), .ZN(n9570) );
  AOI22_X1 U10727 ( .A1(n9811), .A2(n9570), .B1(n9560), .B2(n9809), .ZN(
        P1_U3535) );
  OAI22_X1 U10728 ( .A1(n9562), .A2(n9786), .B1(n9561), .B2(n9784), .ZN(n9563)
         );
  AOI211_X1 U10729 ( .C1(n9565), .C2(n9790), .A(n9564), .B(n9563), .ZN(n9572)
         );
  AOI22_X1 U10730 ( .A1(n9811), .A2(n9572), .B1(n9566), .B2(n9809), .ZN(
        P1_U3534) );
  INV_X1 U10731 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9567) );
  AOI22_X1 U10732 ( .A1(n9794), .A2(n9568), .B1(n9567), .B2(n9792), .ZN(
        P1_U3493) );
  INV_X1 U10733 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9569) );
  AOI22_X1 U10734 ( .A1(n9794), .A2(n9570), .B1(n9569), .B2(n9792), .ZN(
        P1_U3490) );
  INV_X1 U10735 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9571) );
  AOI22_X1 U10736 ( .A1(n9794), .A2(n9572), .B1(n9571), .B2(n9792), .ZN(
        P1_U3487) );
  XNOR2_X1 U10737 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10738 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI222_X1 U10739 ( .A1(n9577), .A2(n9576), .B1(n9575), .B2(n9574), .C1(n6414), .C2(n9573), .ZN(n9578) );
  OAI21_X1 U10740 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(P1_U3230) );
  INV_X1 U10741 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9949) );
  INV_X1 U10742 ( .A(n9581), .ZN(n9585) );
  OAI21_X1 U10743 ( .B1(n9582), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9587), .ZN(
        n9584) );
  AOI21_X1 U10744 ( .B1(n9585), .B2(n9584), .A(n9583), .ZN(n9586) );
  MUX2_X1 U10745 ( .A(P1_REG3_REG_0__SCAN_IN), .B(n9586), .S(
        P1_STATE_REG_SCAN_IN), .Z(n9589) );
  NOR3_X1 U10746 ( .A1(n9622), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9587), .ZN(
        n9588) );
  AOI21_X1 U10747 ( .B1(n9589), .B2(P1_U3083), .A(n9588), .ZN(n9590) );
  OAI21_X1 U10748 ( .B1(n9949), .B2(n9605), .A(n9590), .ZN(P1_U3241) );
  OAI21_X1 U10749 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9594) );
  AOI22_X1 U10750 ( .A1(n9595), .A2(n9634), .B1(n9661), .B2(n9594), .ZN(n9603)
         );
  XNOR2_X1 U10751 ( .A(n9597), .B(n9596), .ZN(n9599) );
  AOI21_X1 U10752 ( .B1(n9665), .B2(n9599), .A(n9598), .ZN(n9600) );
  AND2_X1 U10753 ( .A1(n9601), .A2(n9600), .ZN(n9602) );
  OAI211_X1 U10754 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(
        P1_U3245) );
  AOI22_X1 U10755 ( .A1(n9659), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9606), .B2(
        n9634), .ZN(n9617) );
  AOI21_X1 U10756 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9610) );
  OR2_X1 U10757 ( .A1(n9610), .A2(n9622), .ZN(n9615) );
  OAI211_X1 U10758 ( .C1(n9613), .C2(n9612), .A(n9665), .B(n9611), .ZN(n9614)
         );
  NAND4_X1 U10759 ( .A1(n9617), .A2(n9616), .A3(n9615), .A4(n9614), .ZN(
        P1_U3250) );
  AOI22_X1 U10760 ( .A1(n9659), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9618), .B2(
        n9634), .ZN(n9630) );
  AOI21_X1 U10761 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9623) );
  OR2_X1 U10762 ( .A1(n9623), .A2(n9622), .ZN(n9628) );
  OAI211_X1 U10763 ( .C1(n9626), .C2(n9625), .A(n9665), .B(n9624), .ZN(n9627)
         );
  NAND4_X1 U10764 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(
        P1_U3251) );
  INV_X1 U10765 ( .A(n9631), .ZN(n9632) );
  AOI21_X1 U10766 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9642) );
  OAI211_X1 U10767 ( .C1(n9636), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9661), .B(
        n9635), .ZN(n9641) );
  NAND2_X1 U10768 ( .A1(n9659), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9640) );
  OAI211_X1 U10769 ( .C1(n9638), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9665), .B(
        n9637), .ZN(n9639) );
  NAND4_X1 U10770 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(
        P1_U3256) );
  NOR2_X1 U10771 ( .A1(n9656), .A2(n9643), .ZN(n9644) );
  AOI211_X1 U10772 ( .C1(n9659), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9645), .B(
        n9644), .ZN(n9654) );
  OAI211_X1 U10773 ( .C1(n9648), .C2(n9647), .A(n9661), .B(n9646), .ZN(n9653)
         );
  OAI211_X1 U10774 ( .C1(n9651), .C2(n9650), .A(n9665), .B(n9649), .ZN(n9652)
         );
  NAND3_X1 U10775 ( .A1(n9654), .A2(n9653), .A3(n9652), .ZN(P1_U3257) );
  NOR2_X1 U10776 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  AOI211_X1 U10777 ( .C1(n9659), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9658), .B(
        n9657), .ZN(n9670) );
  OAI211_X1 U10778 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9669)
         );
  OAI211_X1 U10779 ( .C1(n9667), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9668)
         );
  NAND3_X1 U10780 ( .A1(n9670), .A2(n9669), .A3(n9668), .ZN(P1_U3258) );
  INV_X1 U10781 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9690) );
  XOR2_X1 U10782 ( .A(n9671), .B(n9681), .Z(n9760) );
  AOI21_X1 U10783 ( .B1(n9672), .B2(n9676), .A(n9786), .ZN(n9674) );
  NAND2_X1 U10784 ( .A1(n9674), .A2(n9673), .ZN(n9756) );
  AOI22_X1 U10785 ( .A1(n9714), .A2(n9677), .B1(n9676), .B2(n9675), .ZN(n9678)
         );
  OAI21_X1 U10786 ( .B1(n9756), .B2(n9679), .A(n9678), .ZN(n9688) );
  XOR2_X1 U10787 ( .A(n9681), .B(n9680), .Z(n9683) );
  OAI222_X1 U10788 ( .A1(n9687), .A2(n9686), .B1(n9685), .B2(n9684), .C1(n9683), .C2(n9682), .ZN(n9758) );
  AOI211_X1 U10789 ( .C1(n4814), .C2(n9760), .A(n9688), .B(n9758), .ZN(n9689)
         );
  AOI22_X1 U10790 ( .A1(n9715), .A2(n9690), .B1(n9689), .B2(n9719), .ZN(
        P1_U3286) );
  XNOR2_X1 U10791 ( .A(n9692), .B(n9691), .ZN(n9712) );
  INV_X1 U10792 ( .A(n9712), .ZN(n9748) );
  AND2_X1 U10793 ( .A1(n9694), .A2(n9693), .ZN(n9696) );
  OR2_X1 U10794 ( .A1(n9696), .A2(n9695), .ZN(n9745) );
  INV_X1 U10795 ( .A(n9745), .ZN(n9697) );
  AOI22_X1 U10796 ( .A1(n9748), .A2(n9699), .B1(n9698), .B2(n9697), .ZN(n9721)
         );
  AOI22_X1 U10797 ( .A1(n9702), .A2(n9701), .B1(n4250), .B2(n9700), .ZN(n9711)
         );
  INV_X1 U10798 ( .A(n9703), .ZN(n9709) );
  AND3_X1 U10799 ( .A1(n9706), .A2(n9705), .A3(n9704), .ZN(n9708) );
  OAI21_X1 U10800 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(n9710) );
  OAI211_X1 U10801 ( .C1(n9712), .C2(n9726), .A(n9711), .B(n9710), .ZN(n9746)
         );
  AOI22_X1 U10802 ( .A1(n9715), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9714), .B2(
        n9713), .ZN(n9716) );
  OAI21_X1 U10803 ( .B1(n9744), .B2(n9717), .A(n9716), .ZN(n9718) );
  AOI21_X1 U10804 ( .B1(n9746), .B2(n9719), .A(n9718), .ZN(n9720) );
  NAND2_X1 U10805 ( .A1(n9721), .A2(n9720), .ZN(P1_U3288) );
  AND2_X1 U10806 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9725), .ZN(P1_U3292) );
  AND2_X1 U10807 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9725), .ZN(P1_U3293) );
  AND2_X1 U10808 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9725), .ZN(P1_U3294) );
  AND2_X1 U10809 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9725), .ZN(P1_U3295) );
  AND2_X1 U10810 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9725), .ZN(P1_U3296) );
  AND2_X1 U10811 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9725), .ZN(P1_U3297) );
  AND2_X1 U10812 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9725), .ZN(P1_U3298) );
  AND2_X1 U10813 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9725), .ZN(P1_U3299) );
  AND2_X1 U10814 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9725), .ZN(P1_U3300) );
  AND2_X1 U10815 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9725), .ZN(P1_U3301) );
  AND2_X1 U10816 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9725), .ZN(P1_U3302) );
  AND2_X1 U10817 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9725), .ZN(P1_U3303) );
  AND2_X1 U10818 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9725), .ZN(P1_U3304) );
  AND2_X1 U10819 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9725), .ZN(P1_U3305) );
  AND2_X1 U10820 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9725), .ZN(P1_U3306) );
  AND2_X1 U10821 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9725), .ZN(P1_U3307) );
  AND2_X1 U10822 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9725), .ZN(P1_U3308) );
  AND2_X1 U10823 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9725), .ZN(P1_U3309) );
  AND2_X1 U10824 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9725), .ZN(P1_U3310) );
  AND2_X1 U10825 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9725), .ZN(P1_U3311) );
  AND2_X1 U10826 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9725), .ZN(P1_U3312) );
  INV_X1 U10827 ( .A(n9725), .ZN(n9724) );
  NOR2_X1 U10828 ( .A1(n9724), .A2(n9722), .ZN(P1_U3313) );
  AND2_X1 U10829 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9725), .ZN(P1_U3314) );
  NOR2_X1 U10830 ( .A1(n9724), .A2(n9723), .ZN(P1_U3315) );
  AND2_X1 U10831 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9725), .ZN(P1_U3316) );
  AND2_X1 U10832 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9725), .ZN(P1_U3317) );
  AND2_X1 U10833 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9725), .ZN(P1_U3318) );
  AND2_X1 U10834 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9725), .ZN(P1_U3319) );
  AND2_X1 U10835 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9725), .ZN(P1_U3320) );
  AND2_X1 U10836 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9725), .ZN(P1_U3321) );
  NOR2_X1 U10837 ( .A1(n9729), .A2(n9726), .ZN(n9728) );
  NOR2_X1 U10838 ( .A1(n9728), .A2(n9727), .ZN(n9736) );
  INV_X1 U10839 ( .A(n9729), .ZN(n9734) );
  INV_X1 U10840 ( .A(n9730), .ZN(n9767) );
  OAI21_X1 U10841 ( .B1(n9732), .B2(n9784), .A(n9731), .ZN(n9733) );
  AOI21_X1 U10842 ( .B1(n9734), .B2(n9767), .A(n9733), .ZN(n9735) );
  AND2_X1 U10843 ( .A1(n9736), .A2(n9735), .ZN(n9796) );
  INV_X1 U10844 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9737) );
  AOI22_X1 U10845 ( .A1(n9794), .A2(n9796), .B1(n9737), .B2(n9792), .ZN(
        P1_U3457) );
  OAI22_X1 U10846 ( .A1(n9739), .A2(n9786), .B1(n9738), .B2(n9784), .ZN(n9741)
         );
  AOI211_X1 U10847 ( .C1(n9767), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9798)
         );
  INV_X1 U10848 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U10849 ( .A1(n9794), .A2(n9798), .B1(n9743), .B2(n9792), .ZN(
        P1_U3460) );
  OAI22_X1 U10850 ( .A1(n9745), .A2(n9786), .B1(n9744), .B2(n9784), .ZN(n9747)
         );
  AOI211_X1 U10851 ( .C1(n9767), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9799)
         );
  INV_X1 U10852 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9749) );
  AOI22_X1 U10853 ( .A1(n9794), .A2(n9799), .B1(n9749), .B2(n9792), .ZN(
        P1_U3463) );
  OAI22_X1 U10854 ( .A1(n9751), .A2(n9786), .B1(n9750), .B2(n9784), .ZN(n9753)
         );
  AOI211_X1 U10855 ( .C1(n9767), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9800)
         );
  INV_X1 U10856 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9755) );
  AOI22_X1 U10857 ( .A1(n9794), .A2(n9800), .B1(n9755), .B2(n9792), .ZN(
        P1_U3466) );
  OAI21_X1 U10858 ( .B1(n9757), .B2(n9784), .A(n9756), .ZN(n9759) );
  AOI211_X1 U10859 ( .C1(n9790), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9802)
         );
  INV_X1 U10860 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U10861 ( .A1(n9794), .A2(n9802), .B1(n9761), .B2(n9792), .ZN(
        P1_U3469) );
  OAI22_X1 U10862 ( .A1(n9763), .A2(n9786), .B1(n9762), .B2(n9784), .ZN(n9765)
         );
  AOI211_X1 U10863 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9804)
         );
  INV_X1 U10864 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10865 ( .A1(n9794), .A2(n9804), .B1(n9768), .B2(n9792), .ZN(
        P1_U3472) );
  OAI21_X1 U10866 ( .B1(n9770), .B2(n9784), .A(n9769), .ZN(n9772) );
  AOI211_X1 U10867 ( .C1(n9790), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9806)
         );
  INV_X1 U10868 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10869 ( .A1(n9794), .A2(n9806), .B1(n9774), .B2(n9792), .ZN(
        P1_U3475) );
  NAND2_X1 U10870 ( .A1(n9775), .A2(n9790), .ZN(n9782) );
  AOI22_X1 U10871 ( .A1(n9779), .A2(n9778), .B1(n9777), .B2(n9776), .ZN(n9780)
         );
  INV_X1 U10872 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10873 ( .A1(n9794), .A2(n9808), .B1(n9783), .B2(n9792), .ZN(
        P1_U3478) );
  OAI22_X1 U10874 ( .A1(n9787), .A2(n9786), .B1(n9785), .B2(n9784), .ZN(n9789)
         );
  AOI211_X1 U10875 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9810)
         );
  INV_X1 U10876 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10877 ( .A1(n9794), .A2(n9810), .B1(n9793), .B2(n9792), .ZN(
        P1_U3481) );
  INV_X1 U10878 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U10879 ( .A1(n9811), .A2(n9796), .B1(n9795), .B2(n9809), .ZN(
        P1_U3524) );
  AOI22_X1 U10880 ( .A1(n9811), .A2(n9798), .B1(n9797), .B2(n9809), .ZN(
        P1_U3525) );
  AOI22_X1 U10881 ( .A1(n9811), .A2(n9799), .B1(n5815), .B2(n9809), .ZN(
        P1_U3526) );
  AOI22_X1 U10882 ( .A1(n9811), .A2(n9800), .B1(n5816), .B2(n9809), .ZN(
        P1_U3527) );
  INV_X1 U10883 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U10884 ( .A1(n9811), .A2(n9802), .B1(n9801), .B2(n9809), .ZN(
        P1_U3528) );
  AOI22_X1 U10885 ( .A1(n9811), .A2(n9804), .B1(n9803), .B2(n9809), .ZN(
        P1_U3529) );
  AOI22_X1 U10886 ( .A1(n9811), .A2(n9806), .B1(n9805), .B2(n9809), .ZN(
        P1_U3530) );
  AOI22_X1 U10887 ( .A1(n9811), .A2(n9808), .B1(n9807), .B2(n9809), .ZN(
        P1_U3531) );
  AOI22_X1 U10888 ( .A1(n9811), .A2(n9810), .B1(n5937), .B2(n9809), .ZN(
        P1_U3532) );
  AOI22_X1 U10889 ( .A1(n9814), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9812), .ZN(n9824) );
  NAND2_X1 U10890 ( .A1(n9814), .A2(n9813), .ZN(n9816) );
  OAI211_X1 U10891 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9817), .A(n9816), .B(
        n9815), .ZN(n9818) );
  INV_X1 U10892 ( .A(n9818), .ZN(n9822) );
  AOI22_X1 U10893 ( .A1(n9820), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9821) );
  OAI221_X1 U10894 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9824), .C1(n9823), .C2(
        n9822), .A(n9821), .ZN(P2_U3245) );
  NAND2_X1 U10895 ( .A1(n6562), .A2(n9825), .ZN(n9827) );
  NAND2_X1 U10896 ( .A1(n9827), .A2(n9826), .ZN(n9828) );
  XNOR2_X1 U10897 ( .A(n9828), .B(n9840), .ZN(n9896) );
  OAI21_X1 U10898 ( .B1(n9830), .B2(n9829), .A(n9836), .ZN(n9832) );
  NAND3_X1 U10899 ( .A1(n9832), .A2(n9899), .A3(n9831), .ZN(n9892) );
  AOI22_X1 U10900 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(n9833), .ZN(n9837)
         );
  OAI21_X1 U10901 ( .B1(n9892), .B2(n9838), .A(n9837), .ZN(n9844) );
  XOR2_X1 U10902 ( .A(n9840), .B(n9839), .Z(n9843) );
  OAI21_X1 U10903 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9894) );
  AOI211_X1 U10904 ( .C1(n9845), .C2(n9896), .A(n9844), .B(n9894), .ZN(n9847)
         );
  AOI22_X1 U10905 ( .A1(n9848), .A2(n4926), .B1(n9847), .B2(n9846), .ZN(
        P2_U3291) );
  NOR2_X1 U10906 ( .A1(n9857), .A2(n9851), .ZN(P2_U3297) );
  NOR2_X1 U10907 ( .A1(n9857), .A2(n9852), .ZN(P2_U3298) );
  AND2_X1 U10908 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9860), .ZN(P2_U3299) );
  AND2_X1 U10909 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9860), .ZN(P2_U3300) );
  AND2_X1 U10910 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9860), .ZN(P2_U3301) );
  NOR2_X1 U10911 ( .A1(n9857), .A2(n9853), .ZN(P2_U3302) );
  AND2_X1 U10912 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9860), .ZN(P2_U3303) );
  AND2_X1 U10913 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9860), .ZN(P2_U3304) );
  AND2_X1 U10914 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9860), .ZN(P2_U3305) );
  AND2_X1 U10915 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9860), .ZN(P2_U3306) );
  AND2_X1 U10916 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9860), .ZN(P2_U3307) );
  AND2_X1 U10917 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9860), .ZN(P2_U3308) );
  AND2_X1 U10918 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9860), .ZN(P2_U3309) );
  AND2_X1 U10919 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9860), .ZN(P2_U3310) );
  AND2_X1 U10920 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9860), .ZN(P2_U3311) );
  NOR2_X1 U10921 ( .A1(n9857), .A2(n9854), .ZN(P2_U3312) );
  AND2_X1 U10922 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9860), .ZN(P2_U3313) );
  AND2_X1 U10923 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9860), .ZN(P2_U3314) );
  AND2_X1 U10924 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9860), .ZN(P2_U3315) );
  AND2_X1 U10925 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9860), .ZN(P2_U3316) );
  NOR2_X1 U10926 ( .A1(n9857), .A2(n9855), .ZN(P2_U3317) );
  AND2_X1 U10927 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9860), .ZN(P2_U3318) );
  AND2_X1 U10928 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9860), .ZN(P2_U3319) );
  AND2_X1 U10929 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9860), .ZN(P2_U3320) );
  AND2_X1 U10930 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9860), .ZN(P2_U3321) );
  AND2_X1 U10931 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9860), .ZN(P2_U3322) );
  AND2_X1 U10932 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9860), .ZN(P2_U3323) );
  AND2_X1 U10933 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9860), .ZN(P2_U3324) );
  AND2_X1 U10934 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9860), .ZN(P2_U3325) );
  NOR2_X1 U10935 ( .A1(n9857), .A2(n9856), .ZN(P2_U3326) );
  AOI22_X1 U10936 ( .A1(n9863), .A2(n9859), .B1(n9858), .B2(n9860), .ZN(
        P2_U3437) );
  AOI22_X1 U10937 ( .A1(n9863), .A2(n9862), .B1(n9861), .B2(n9860), .ZN(
        P2_U3438) );
  AOI22_X1 U10938 ( .A1(n9866), .A2(n9925), .B1(n9865), .B2(n9864), .ZN(n9867)
         );
  AND2_X1 U10939 ( .A1(n9868), .A2(n9867), .ZN(n9929) );
  AOI22_X1 U10940 ( .A1(n9912), .A2(n9929), .B1(n4792), .B2(n9927), .ZN(
        P2_U3451) );
  NAND3_X1 U10941 ( .A1(n9870), .A2(n9869), .A3(n9899), .ZN(n9871) );
  OAI21_X1 U10942 ( .B1(n6346), .B2(n9919), .A(n9871), .ZN(n9874) );
  INV_X1 U10943 ( .A(n9872), .ZN(n9873) );
  AOI211_X1 U10944 ( .C1(n9925), .C2(n9875), .A(n9874), .B(n9873), .ZN(n9930)
         );
  AOI22_X1 U10945 ( .A1(n9912), .A2(n9930), .B1(n4875), .B2(n9927), .ZN(
        P2_U3454) );
  OAI22_X1 U10946 ( .A1(n9876), .A2(n9921), .B1(n6349), .B2(n9919), .ZN(n9878)
         );
  AOI211_X1 U10947 ( .C1(n9925), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9931)
         );
  AOI22_X1 U10948 ( .A1(n9912), .A2(n9931), .B1(n4847), .B2(n9927), .ZN(
        P2_U3457) );
  INV_X1 U10949 ( .A(n9880), .ZN(n9917) );
  OAI22_X1 U10950 ( .A1(n9881), .A2(n9921), .B1(n6257), .B2(n9919), .ZN(n9882)
         );
  AOI21_X1 U10951 ( .B1(n9883), .B2(n9917), .A(n9882), .ZN(n9884) );
  INV_X1 U10952 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9886) );
  AOI22_X1 U10953 ( .A1(n9912), .A2(n9932), .B1(n9886), .B2(n9927), .ZN(
        P2_U3460) );
  OAI22_X1 U10954 ( .A1(n9888), .A2(n9921), .B1(n9887), .B2(n9919), .ZN(n9890)
         );
  AOI211_X1 U10955 ( .C1(n9925), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9934)
         );
  AOI22_X1 U10956 ( .A1(n9912), .A2(n9934), .B1(n4906), .B2(n9927), .ZN(
        P2_U3463) );
  OAI21_X1 U10957 ( .B1(n9893), .B2(n9919), .A(n9892), .ZN(n9895) );
  AOI211_X1 U10958 ( .C1(n9925), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9935)
         );
  AOI22_X1 U10959 ( .A1(n9912), .A2(n9935), .B1(n4925), .B2(n9927), .ZN(
        P2_U3466) );
  AOI22_X1 U10960 ( .A1(n9900), .A2(n9899), .B1(n9898), .B2(n9897), .ZN(n9901)
         );
  OAI211_X1 U10961 ( .C1(n9904), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9905)
         );
  INV_X1 U10962 ( .A(n9905), .ZN(n9937) );
  INV_X1 U10963 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9906) );
  AOI22_X1 U10964 ( .A1(n9912), .A2(n9937), .B1(n9906), .B2(n9927), .ZN(
        P2_U3469) );
  OAI22_X1 U10965 ( .A1(n9908), .A2(n9921), .B1(n9907), .B2(n9919), .ZN(n9910)
         );
  AOI211_X1 U10966 ( .C1(n9917), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9938)
         );
  AOI22_X1 U10967 ( .A1(n9912), .A2(n9938), .B1(n4979), .B2(n9927), .ZN(
        P2_U3475) );
  OAI22_X1 U10968 ( .A1(n9913), .A2(n9921), .B1(n6802), .B2(n9919), .ZN(n9915)
         );
  AOI211_X1 U10969 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9939)
         );
  INV_X1 U10970 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U10971 ( .A1(n9912), .A2(n9939), .B1(n9918), .B2(n9927), .ZN(
        P2_U3481) );
  OAI22_X1 U10972 ( .A1(n9922), .A2(n9921), .B1(n9920), .B2(n9919), .ZN(n9924)
         );
  AOI211_X1 U10973 ( .C1(n9926), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9942)
         );
  AOI22_X1 U10974 ( .A1(n9912), .A2(n9942), .B1(n5077), .B2(n9927), .ZN(
        P2_U3487) );
  AOI22_X1 U10975 ( .A1(n9943), .A2(n9929), .B1(n9928), .B2(n9940), .ZN(
        P2_U3520) );
  AOI22_X1 U10976 ( .A1(n9943), .A2(n9930), .B1(n6106), .B2(n9940), .ZN(
        P2_U3521) );
  AOI22_X1 U10977 ( .A1(n9943), .A2(n9931), .B1(n6104), .B2(n9940), .ZN(
        P2_U3522) );
  AOI22_X1 U10978 ( .A1(n9943), .A2(n9932), .B1(n6103), .B2(n9940), .ZN(
        P2_U3523) );
  AOI22_X1 U10979 ( .A1(n9943), .A2(n9934), .B1(n9933), .B2(n9940), .ZN(
        P2_U3524) );
  AOI22_X1 U10980 ( .A1(n9943), .A2(n9935), .B1(n6101), .B2(n9940), .ZN(
        P2_U3525) );
  AOI22_X1 U10981 ( .A1(n9943), .A2(n9937), .B1(n9936), .B2(n9940), .ZN(
        P2_U3526) );
  AOI22_X1 U10982 ( .A1(n9943), .A2(n9938), .B1(n6111), .B2(n9940), .ZN(
        P2_U3528) );
  AOI22_X1 U10983 ( .A1(n9943), .A2(n9939), .B1(n6222), .B2(n9940), .ZN(
        P2_U3530) );
  AOI22_X1 U10984 ( .A1(n9943), .A2(n9942), .B1(n9941), .B2(n9940), .ZN(
        P2_U3532) );
  INV_X1 U10985 ( .A(n9944), .ZN(n9945) );
  NAND2_X1 U10986 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  XOR2_X1 U10987 ( .A(n9948), .B(n9947), .Z(ADD_1071_U5) );
  INV_X1 U10988 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U10989 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9950), .B2(n9949), .ZN(ADD_1071_U46) );
  OAI21_X1 U10990 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(ADD_1071_U56) );
  OAI21_X1 U10991 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(ADD_1071_U57) );
  OAI21_X1 U10992 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(ADD_1071_U58) );
  OAI21_X1 U10993 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(ADD_1071_U59) );
  OAI21_X1 U10994 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(ADD_1071_U60) );
  OAI21_X1 U10995 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(ADD_1071_U61) );
  AOI21_X1 U10996 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(ADD_1071_U62) );
  AOI21_X1 U10997 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(ADD_1071_U63) );
  XOR2_X1 U10998 ( .A(n9975), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10999 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  XOR2_X1 U11000 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9978), .Z(ADD_1071_U51) );
  OAI21_X1 U11001 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9982) );
  XNOR2_X1 U11002 ( .A(n9982), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11003 ( .B1(n9985), .B2(n9984), .A(n9983), .ZN(ADD_1071_U47) );
  XOR2_X1 U11004 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9986), .Z(ADD_1071_U48) );
  XOR2_X1 U11005 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9987), .Z(ADD_1071_U49) );
  XOR2_X1 U11006 ( .A(n9989), .B(n9988), .Z(ADD_1071_U54) );
  XOR2_X1 U11007 ( .A(n9991), .B(n9990), .Z(ADD_1071_U53) );
  XNOR2_X1 U11008 ( .A(n9993), .B(n9992), .ZN(ADD_1071_U52) );
  AND2_X1 U5988 ( .A1(n4523), .A2(n4522), .ZN(n5633) );
  NAND4_X2 U4788 ( .A1(n5661), .A2(n5660), .A3(n5659), .A4(n5658), .ZN(n5913)
         );
  OAI21_X1 U4750 ( .B1(n9525), .B2(n9549), .A(n9524), .ZN(n9550) );
  CLKBUF_X1 U4769 ( .A(n4882), .Z(n5396) );
  NOR3_X1 U4855 ( .A1(n5916), .A2(P1_IR_REG_19__SCAN_IN), .A3(n5667), .ZN(
        n4520) );
  CLKBUF_X1 U4918 ( .A(n9846), .Z(n8253) );
  XNOR2_X1 U4919 ( .A(n5607), .B(n5606), .ZN(n7050) );
endmodule

