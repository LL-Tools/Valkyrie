

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910;

  XNOR2_X1 U11030 ( .A(n14363), .B(n14362), .ZN(n19127) );
  OR2_X1 U11031 ( .A1(n9985), .A2(n15002), .ZN(n9983) );
  INV_X2 U11032 ( .A(n19111), .ZN(n19089) );
  NOR2_X1 U11033 ( .A1(n15813), .A2(n17839), .ZN(n18121) );
  NOR2_X1 U11034 ( .A1(n17840), .A2(n18161), .ZN(n17839) );
  NAND2_X1 U11035 ( .A1(n16328), .A2(n12619), .ZN(n14493) );
  CLKBUF_X2 U11036 ( .A(n14319), .Z(n9591) );
  INV_X2 U11037 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n10675) );
  OR2_X1 U11038 ( .A1(n11377), .A2(n11368), .ZN(n15480) );
  AND2_X1 U11039 ( .A1(n11355), .A2(n11352), .ZN(n16368) );
  AND2_X1 U11040 ( .A1(n13425), .A2(n11392), .ZN(n12600) );
  AND2_X1 U11041 ( .A1(n13421), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12597) );
  AND2_X1 U11042 ( .A1(n9601), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12598) );
  CLKBUF_X2 U11043 ( .A(n13601), .Z(n11105) );
  CLKBUF_X2 U11044 ( .A(n13332), .Z(n13382) );
  INV_X1 U11045 ( .A(n12722), .ZN(n13230) );
  BUF_X2 U11046 ( .A(n15752), .Z(n17239) );
  CLKBUF_X2 U11047 ( .A(n15738), .Z(n17242) );
  INV_X1 U11048 ( .A(n10232), .ZN(n17020) );
  CLKBUF_X1 U11049 ( .A(n15739), .Z(n17243) );
  CLKBUF_X1 U11050 ( .A(n14891), .Z(n9606) );
  INV_X1 U11051 ( .A(n11279), .ZN(n11301) );
  NOR2_X2 U11052 ( .A1(n11813), .A2(n16983), .ZN(n15740) );
  NAND2_X2 U11053 ( .A1(n9856), .A2(n9855), .ZN(n16408) );
  NAND4_X1 U11054 ( .A1(n9857), .A2(n11259), .A3(n11257), .A4(n11256), .ZN(
        n9855) );
  NAND2_X1 U11055 ( .A1(n12508), .A2(n12658), .ZN(n13593) );
  INV_X1 U11056 ( .A(n12959), .ZN(n10345) );
  BUF_X1 U11057 ( .A(n10414), .Z(n10474) );
  BUF_X1 U11058 ( .A(n10350), .Z(n14281) );
  INV_X1 U11059 ( .A(n12978), .ZN(n20101) );
  NAND2_X1 U11060 ( .A1(n12012), .A2(n12500), .ZN(n12162) );
  BUF_X2 U11061 ( .A(n13417), .Z(n9599) );
  INV_X1 U11062 ( .A(n13429), .ZN(n13417) );
  OR2_X1 U11063 ( .A1(n10299), .A2(n10298), .ZN(n10524) );
  BUF_X1 U11064 ( .A(n10816), .Z(n11131) );
  AND2_X2 U11065 ( .A1(n12425), .A2(n14286), .ZN(n10436) );
  AND2_X1 U11066 ( .A1(n12425), .A2(n10242), .ZN(n10315) );
  AND2_X1 U11067 ( .A1(n10243), .A2(n10245), .ZN(n10383) );
  AND2_X1 U11068 ( .A1(n10245), .A2(n14286), .ZN(n13601) );
  CLKBUF_X2 U11069 ( .A(n10816), .Z(n13602) );
  AND2_X1 U11070 ( .A1(n10029), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10243) );
  INV_X4 U11071 ( .A(n18181), .ZN(n9593) );
  BUF_X1 U11072 ( .A(n10314), .Z(n11089) );
  NAND3_X2 U11073 ( .A1(n15449), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n10171), .ZN(n13242) );
  AND2_X1 U11074 ( .A1(n11383), .A2(n11392), .ZN(n13236) );
  AND2_X1 U11075 ( .A1(n9598), .A2(n11392), .ZN(n11415) );
  INV_X1 U11076 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11392) );
  NOR2_X1 U11077 ( .A1(n12162), .A2(n20101), .ZN(n11993) );
  NAND2_X1 U11078 ( .A1(n11255), .A2(n11254), .ZN(n11293) );
  BUF_X1 U11079 ( .A(n11330), .Z(n14307) );
  AND3_X1 U11080 ( .A1(n16421), .A2(n9590), .A3(n12070), .ZN(n12903) );
  CLKBUF_X2 U11081 ( .A(n12508), .Z(n12501) );
  NOR2_X1 U11082 ( .A1(n12978), .A2(n12959), .ZN(n12131) );
  INV_X1 U11083 ( .A(n12501), .ZN(n13646) );
  NOR2_X2 U11084 ( .A1(n13628), .A2(n13653), .ZN(n13652) );
  AND2_X1 U11085 ( .A1(n13792), .A2(n9697), .ZN(n13720) );
  NAND2_X1 U11087 ( .A1(n11280), .A2(n11279), .ZN(n11556) );
  INV_X1 U11088 ( .A(n11329), .ZN(n13536) );
  OAI21_X1 U11089 ( .B1(n12464), .B2(n12463), .A(n12462), .ZN(n12567) );
  CLKBUF_X3 U11090 ( .A(n15559), .Z(n9603) );
  NAND2_X1 U11091 ( .A1(n11345), .A2(n11352), .ZN(n11344) );
  AND2_X1 U11092 ( .A1(n9751), .A2(n9681), .ZN(n9790) );
  NAND2_X1 U11093 ( .A1(n10066), .A2(n10064), .ZN(n10063) );
  OAI211_X1 U11094 ( .C1(n10063), .C2(n9789), .A(n9818), .B(n9817), .ZN(n12763) );
  INV_X1 U11096 ( .A(n19948), .ZN(n19879) );
  AOI21_X1 U11097 ( .B1(n13628), .B2(n13653), .A(n13652), .ZN(n13936) );
  XNOR2_X1 U11098 ( .A(n13341), .B(n13342), .ZN(n14599) );
  AND2_X1 U11099 ( .A1(n11280), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19149) );
  NOR2_X1 U11101 ( .A1(n14327), .A2(n16285), .ZN(n14330) );
  XNOR2_X1 U11102 ( .A(n9748), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15001) );
  INV_X1 U11103 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16435) );
  OAI21_X1 U11105 ( .B1(n11151), .B2(n11152), .A(n13628), .ZN(n13857) );
  AND4_X1 U11106 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n9586) );
  NAND2_X2 U11107 ( .A1(n10401), .A2(n10400), .ZN(n10402) );
  NAND2_X2 U11108 ( .A1(n12486), .A2(n10544), .ZN(n10553) );
  XNOR2_X1 U11110 ( .A(n10682), .B(n10533), .ZN(n12446) );
  NOR2_X2 U11111 ( .A1(n10610), .A2(n16031), .ZN(n14029) );
  AND2_X2 U11112 ( .A1(n12291), .A2(n12568), .ZN(n12464) );
  NOR2_X2 U11113 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15461) );
  AOI211_X2 U11114 ( .C1(n18120), .C2(n17946), .A(n17960), .B(n17945), .ZN(
        n17954) );
  NOR2_X1 U11115 ( .A1(n16445), .A2(n16617), .ZN(n17924) );
  INV_X2 U11116 ( .A(n9606), .ZN(n9590) );
  INV_X1 U11117 ( .A(n11293), .ZN(n14891) );
  OAI21_X1 U11118 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n14918), .A(n14305), 
        .ZN(n14319) );
  AND2_X4 U11119 ( .A1(n12428), .A2(n10242), .ZN(n10441) );
  AOI211_X1 U11120 ( .C1(n19227), .C2(n15180), .A(n14966), .B(n14965), .ZN(
        n14967) );
  OR2_X1 U11121 ( .A1(n14972), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10167) );
  AOI21_X1 U11122 ( .B1(n10073), .B2(n10070), .A(n9695), .ZN(n15357) );
  NOR2_X1 U11123 ( .A1(n15334), .A2(n15341), .ZN(n15323) );
  NOR2_X2 U11124 ( .A1(n15003), .A2(n15225), .ZN(n14995) );
  NAND2_X1 U11125 ( .A1(n15032), .A2(n9638), .ZN(n15259) );
  NAND2_X1 U11126 ( .A1(n14902), .A2(n14901), .ZN(n16281) );
  INV_X1 U11127 ( .A(n14000), .ZN(n9595) );
  AND2_X1 U11128 ( .A1(n12298), .A2(n12297), .ZN(n19803) );
  NAND2_X1 U11129 ( .A1(n9742), .A2(n9741), .ZN(n19502) );
  NAND2_X1 U11130 ( .A1(n9742), .A2(n11357), .ZN(n12825) );
  OR2_X1 U11131 ( .A1(n11366), .A2(n11368), .ZN(n19554) );
  BUF_X2 U11132 ( .A(n12186), .Z(n9592) );
  NOR2_X1 U11133 ( .A1(n18767), .A2(n11918), .ZN(n16971) );
  AND2_X1 U11134 ( .A1(n13017), .A2(n13016), .ZN(n14251) );
  NOR2_X1 U11135 ( .A1(n14796), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14804) );
  INV_X2 U11136 ( .A(n9591), .ZN(n19094) );
  NAND2_X1 U11137 ( .A1(n12164), .A2(n12132), .ZN(n10357) );
  INV_X4 U11138 ( .A(n16986), .ZN(n9694) );
  INV_X4 U11139 ( .A(n11720), .ZN(n14828) );
  NAND2_X1 U11141 ( .A1(n12628), .A2(n12501), .ZN(n12004) );
  NOR3_X2 U11142 ( .A1(n17571), .A2(n17592), .A3(n17572), .ZN(n16482) );
  CLKBUF_X2 U11143 ( .A(n10352), .Z(n12015) );
  INV_X4 U11144 ( .A(n15526), .ZN(n16421) );
  CLKBUF_X2 U11145 ( .A(n12604), .Z(n13222) );
  BUF_X1 U11146 ( .A(n10320), .Z(n10419) );
  CLKBUF_X2 U11147 ( .A(n10436), .Z(n10993) );
  BUF_X4 U11148 ( .A(n10305), .Z(n9594) );
  CLKBUF_X2 U11149 ( .A(n13122), .Z(n13229) );
  INV_X2 U11150 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10171) );
  OAI21_X1 U11151 ( .B1(n13929), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10143), .ZN(n10142) );
  NAND2_X1 U11152 ( .A1(n13947), .A2(n14074), .ZN(n13923) );
  NOR2_X1 U11153 ( .A1(n15328), .A2(n9779), .ZN(n9778) );
  AOI211_X1 U11154 ( .C1(n16369), .C2(n16189), .A(n15152), .B(n15151), .ZN(
        n15153) );
  OR2_X1 U11155 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  AOI211_X1 U11156 ( .C1(n19227), .C2(n16189), .A(n14930), .B(n14929), .ZN(
        n14931) );
  AND2_X1 U11157 ( .A1(n9897), .A2(n9895), .ZN(n9894) );
  AND2_X1 U11158 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  OR2_X1 U11159 ( .A1(n13857), .A2(n20098), .ZN(n11160) );
  NAND2_X1 U11160 ( .A1(n10167), .A2(n10166), .ZN(n15150) );
  OR2_X1 U11161 ( .A1(n15086), .A2(n10082), .ZN(n10076) );
  OAI21_X1 U11162 ( .B1(n9782), .B2(n9781), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9780) );
  OR2_X1 U11163 ( .A1(n15086), .A2(n15023), .ZN(n10085) );
  NAND2_X1 U11164 ( .A1(n15359), .A2(n15355), .ZN(n15086) );
  OR2_X1 U11165 ( .A1(n15361), .A2(n15362), .ZN(n16238) );
  NAND2_X1 U11166 ( .A1(n13991), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13968) );
  OR2_X1 U11167 ( .A1(n15320), .A2(n9783), .ZN(n9782) );
  OR2_X1 U11168 ( .A1(n16256), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16258) );
  NAND2_X1 U11169 ( .A1(n9793), .A2(n9791), .ZN(n15002) );
  OR2_X1 U11170 ( .A1(n15386), .A2(n15397), .ZN(n9743) );
  CLKBUF_X1 U11171 ( .A(n13720), .Z(n13721) );
  NAND2_X1 U11172 ( .A1(n14599), .A2(n14598), .ZN(n14597) );
  NAND2_X1 U11173 ( .A1(n15362), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15334) );
  NAND2_X1 U11174 ( .A1(n9656), .A2(n9914), .ZN(n9913) );
  XNOR2_X1 U11175 ( .A(n14314), .B(n14313), .ZN(n15140) );
  NAND2_X1 U11176 ( .A1(n9732), .A2(n9730), .ZN(n9729) );
  XNOR2_X1 U11177 ( .A(n9653), .B(n14303), .ZN(n16189) );
  NAND2_X1 U11178 ( .A1(n9785), .A2(n10235), .ZN(n10075) );
  NAND2_X1 U11179 ( .A1(n9947), .A2(n9946), .ZN(n16449) );
  AOI21_X1 U11180 ( .B1(n14782), .B2(n14783), .A(n9654), .ZN(n9785) );
  NOR2_X1 U11181 ( .A1(n14388), .A2(n10103), .ZN(n14314) );
  OR2_X1 U11182 ( .A1(n9644), .A2(n14386), .ZN(n14388) );
  OR2_X1 U11183 ( .A1(n9890), .A2(n9728), .ZN(n9727) );
  NOR2_X1 U11184 ( .A1(n14046), .A2(n14044), .ZN(n16051) );
  NOR2_X1 U11185 ( .A1(n14621), .A2(n14620), .ZN(n14622) );
  OR2_X1 U11186 ( .A1(n14462), .A2(n14463), .ZN(n14621) );
  NAND2_X1 U11187 ( .A1(n16053), .A2(n9621), .ZN(n14046) );
  AOI21_X1 U11188 ( .B1(n9892), .B2(n14908), .A(n9891), .ZN(n9890) );
  AND2_X1 U11189 ( .A1(n9767), .A2(n10724), .ZN(n12846) );
  INV_X1 U11190 ( .A(n14913), .ZN(n9728) );
  NOR2_X1 U11191 ( .A1(n14649), .A2(n14638), .ZN(n14640) );
  AND2_X1 U11192 ( .A1(n10723), .A2(n9768), .ZN(n9767) );
  NOR2_X1 U11193 ( .A1(n11546), .A2(n9775), .ZN(n9774) );
  XNOR2_X1 U11194 ( .A(n14910), .B(n11643), .ZN(n16279) );
  OR2_X1 U11195 ( .A1(n14905), .A2(n14904), .ZN(n14910) );
  NAND2_X1 U11196 ( .A1(n9912), .A2(n10519), .ZN(n10587) );
  INV_X1 U11197 ( .A(n10576), .ZN(n9912) );
  AND2_X1 U11198 ( .A1(n14490), .A2(n14489), .ZN(n14492) );
  NAND2_X1 U11199 ( .A1(n9744), .A2(n11509), .ZN(n14905) );
  NOR2_X2 U11200 ( .A1(n19470), .A2(n19659), .ZN(n19707) );
  XNOR2_X1 U11201 ( .A(n10565), .B(n10564), .ZN(n10722) );
  XNOR2_X1 U11202 ( .A(n11508), .B(n11509), .ZN(n11677) );
  NOR2_X1 U11203 ( .A1(n12709), .A2(n12710), .ZN(n14489) );
  NAND2_X1 U11204 ( .A1(n14455), .A2(n14868), .ZN(n14871) );
  OR2_X1 U11205 ( .A1(n19803), .A2(n15477), .ZN(n19368) );
  AND2_X2 U11206 ( .A1(n12695), .A2(n12694), .ZN(n12704) );
  AND2_X1 U11207 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  AND2_X1 U11208 ( .A1(n11543), .A2(n11542), .ZN(n14903) );
  NAND2_X1 U11209 ( .A1(n9646), .A2(n14819), .ZN(n14455) );
  NOR2_X1 U11210 ( .A1(n18082), .A2(n18081), .ZN(n18080) );
  NAND2_X1 U11211 ( .A1(n13725), .A2(n13714), .ZN(n13716) );
  NAND2_X1 U11212 ( .A1(n12472), .A2(n12471), .ZN(n12544) );
  AND2_X1 U11213 ( .A1(n13086), .A2(n11793), .ZN(n12472) );
  NAND2_X1 U11214 ( .A1(n14760), .A2(n14749), .ZN(n14750) );
  AND2_X1 U11215 ( .A1(n13085), .A2(n13084), .ZN(n13086) );
  OR2_X2 U11216 ( .A1(n11372), .A2(n11376), .ZN(n19341) );
  NAND2_X1 U11217 ( .A1(n11354), .A2(n9741), .ZN(n19609) );
  CLKBUF_X1 U11218 ( .A(n13849), .Z(n13910) );
  CLKBUF_X1 U11219 ( .A(n13845), .Z(n13908) );
  OR2_X1 U11220 ( .A1(n11366), .A2(n11376), .ZN(n12813) );
  NOR2_X1 U11221 ( .A1(n20103), .A2(n20348), .ZN(n20104) );
  OR2_X1 U11222 ( .A1(n11369), .A2(n11376), .ZN(n19460) );
  OR2_X1 U11223 ( .A1(n13005), .A2(n12984), .ZN(n14085) );
  OR2_X1 U11224 ( .A1(n11366), .A2(n11375), .ZN(n19648) );
  NOR2_X1 U11225 ( .A1(n13098), .A2(n13097), .ZN(n13085) );
  OR2_X1 U11226 ( .A1(n12293), .A2(n12292), .ZN(n12461) );
  OAI211_X1 U11227 ( .C1(n9592), .C2(n9867), .A(n9861), .B(n9859), .ZN(n12293)
         );
  NAND2_X1 U11228 ( .A1(n10483), .A2(n10482), .ZN(n14273) );
  INV_X1 U11229 ( .A(n17931), .ZN(n17903) );
  NAND2_X1 U11230 ( .A1(n13839), .A2(n20136), .ZN(n19954) );
  NAND2_X1 U11231 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17850), .ZN(
        n15811) );
  NAND2_X1 U11232 ( .A1(n10434), .A2(n10520), .ZN(n10456) );
  NAND2_X1 U11233 ( .A1(n9750), .A2(n9707), .ZN(n14838) );
  OAI21_X1 U11234 ( .B1(n10533), .B2(n10345), .A(n10532), .ZN(n10534) );
  NOR2_X1 U11235 ( .A1(n18308), .A2(n17449), .ZN(n17387) );
  AND2_X1 U11236 ( .A1(n10108), .A2(n10109), .ZN(n14439) );
  OR2_X1 U11237 ( .A1(n15448), .A2(n16368), .ZN(n11368) );
  XNOR2_X1 U11238 ( .A(n9881), .B(n11343), .ZN(n12186) );
  OAI21_X1 U11239 ( .B1(n9803), .B2(n9801), .A(n11343), .ZN(n9800) );
  NAND2_X2 U11240 ( .A1(n15915), .A2(n17424), .ZN(n17449) );
  NOR2_X1 U11241 ( .A1(n17860), .A2(n17859), .ZN(n17858) );
  NAND2_X1 U11242 ( .A1(n10162), .A2(n10452), .ZN(n20511) );
  NAND2_X1 U11243 ( .A1(n11344), .A2(n9805), .ZN(n9804) );
  AND2_X2 U11244 ( .A1(n10670), .A2(n10669), .ZN(n12973) );
  NAND2_X1 U11245 ( .A1(n9807), .A2(n11336), .ZN(n9806) );
  AND2_X1 U11246 ( .A1(n14251), .A2(n9702), .ZN(n13835) );
  NAND2_X1 U11247 ( .A1(n11351), .A2(n11350), .ZN(n11355) );
  AND2_X1 U11248 ( .A1(n11325), .A2(n9808), .ZN(n9805) );
  OAI211_X1 U11249 ( .C1(n20109), .C2(n11156), .A(n10380), .B(n10379), .ZN(
        n10381) );
  NAND2_X1 U11250 ( .A1(n12033), .A2(n12032), .ZN(n12031) );
  XNOR2_X1 U11251 ( .A(n11774), .B(n11775), .ZN(n11773) );
  NAND2_X1 U11252 ( .A1(n10201), .A2(n10202), .ZN(n11325) );
  NOR2_X1 U11253 ( .A1(n12948), .A2(n12949), .ZN(n13017) );
  NAND2_X1 U11254 ( .A1(n11348), .A2(n11349), .ZN(n11352) );
  CLKBUF_X1 U11255 ( .A(n10378), .Z(n10462) );
  NAND2_X1 U11256 ( .A1(n11341), .A2(n11340), .ZN(n11774) );
  NAND2_X1 U11257 ( .A1(n11320), .A2(n11319), .ZN(n11348) );
  XNOR2_X1 U11258 ( .A(n11740), .B(n11737), .ZN(n12033) );
  OAI211_X1 U11259 ( .C1(n14299), .C2(n19836), .A(n11324), .B(n11323), .ZN(
        n11349) );
  NAND2_X1 U11260 ( .A1(n12125), .A2(n11733), .ZN(n11740) );
  AOI21_X1 U11261 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11334), .ZN(n11343) );
  OR2_X1 U11262 ( .A1(n12123), .A2(n12122), .ZN(n12125) );
  NOR2_X1 U11263 ( .A1(n9610), .A2(n12786), .ZN(n11292) );
  OR2_X1 U11264 ( .A1(n9609), .A2(n12087), .ZN(n11319) );
  NAND2_X2 U11265 ( .A1(n11770), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11329) );
  OAI21_X1 U11266 ( .B1(n10357), .B2(n10359), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10373) );
  OAI211_X1 U11267 ( .C1(n9604), .C2(n14557), .A(n11290), .B(n11289), .ZN(
        n11291) );
  NOR2_X1 U11268 ( .A1(n14315), .A2(n14928), .ZN(n12785) );
  OR2_X2 U11269 ( .A1(n11321), .A2(n16435), .ZN(n13534) );
  AND2_X1 U11270 ( .A1(n11728), .A2(n11727), .ZN(n11732) );
  NAND2_X1 U11271 ( .A1(n11330), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11290) );
  NAND2_X2 U11272 ( .A1(n17500), .A2(n17501), .ZN(n17567) );
  AND2_X1 U11273 ( .A1(n11767), .A2(n11288), .ZN(n11330) );
  NAND2_X1 U11274 ( .A1(n9738), .A2(n11311), .ZN(n9736) );
  AOI21_X1 U11275 ( .B1(n9866), .B2(n9864), .A(n9624), .ZN(n9861) );
  INV_X1 U11276 ( .A(n14361), .ZN(n11738) );
  NOR3_X1 U11277 ( .A1(n14323), .A2(n14316), .A3(n10121), .ZN(n14317) );
  AND2_X1 U11278 ( .A1(n11604), .A2(n19149), .ZN(n9738) );
  AOI21_X1 U11279 ( .B1(n11706), .B2(n11707), .A(n16435), .ZN(n11309) );
  NAND2_X1 U11280 ( .A1(n9657), .A2(n11310), .ZN(n16407) );
  AND2_X1 U11281 ( .A1(n14340), .A2(n10113), .ZN(n14324) );
  NOR2_X1 U11282 ( .A1(n12015), .A2(n12978), .ZN(n10353) );
  AND2_X1 U11283 ( .A1(n12979), .A2(n10312), .ZN(n12161) );
  AND2_X1 U11284 ( .A1(n10313), .A2(n13593), .ZN(n12018) );
  AND2_X1 U11285 ( .A1(n10349), .A2(n10362), .ZN(n12152) );
  INV_X2 U11286 ( .A(n9606), .ZN(n11720) );
  AND3_X1 U11287 ( .A1(n18281), .A2(n18308), .A3(n18293), .ZN(n11894) );
  OR2_X1 U11288 ( .A1(n10352), .A2(n12508), .ZN(n12979) );
  AND2_X1 U11289 ( .A1(n10347), .A2(n10672), .ZN(n12012) );
  INV_X1 U11290 ( .A(n11298), .ZN(n11310) );
  BUF_X4 U11291 ( .A(n11279), .Z(n15526) );
  OR2_X1 U11292 ( .A1(n11424), .A2(n11423), .ZN(n11736) );
  NAND2_X1 U11293 ( .A1(n15728), .A2(n10176), .ZN(n15817) );
  NAND3_X1 U11294 ( .A1(n11891), .A2(n11890), .A3(n11889), .ZN(n16445) );
  INV_X2 U11295 ( .A(n12145), .ZN(n10344) );
  NAND2_X2 U11296 ( .A1(n11220), .A2(n11219), .ZN(n15543) );
  CLKBUF_X2 U11297 ( .A(n10346), .Z(n12208) );
  INV_X1 U11298 ( .A(n13848), .ZN(n20128) );
  INV_X1 U11299 ( .A(n10524), .ZN(n20120) );
  NAND4_X1 U11300 ( .A1(n9858), .A2(n11264), .A3(n11261), .A4(n11262), .ZN(
        n9856) );
  NOR2_X1 U11301 ( .A1(n11868), .A2(n9754), .ZN(n9753) );
  OR2_X1 U11302 ( .A1(n10413), .A2(n10412), .ZN(n10591) );
  AND4_X1 U11303 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10271) );
  NOR2_X2 U11304 ( .A1(n20095), .A2(n20098), .ZN(n20096) );
  AND2_X1 U11305 ( .A1(n11263), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9858) );
  AND4_X1 U11306 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  INV_X2 U11307 ( .A(U214), .ZN(n16565) );
  BUF_X2 U11308 ( .A(n10383), .Z(n13608) );
  NAND2_X2 U11309 ( .A1(n18935), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18861) );
  NAND2_X2 U11310 ( .A1(n18935), .A2(n18801), .ZN(n18857) );
  CLKBUF_X2 U11311 ( .A(n10475), .Z(n10407) );
  BUF_X2 U11312 ( .A(n10305), .Z(n13607) );
  NAND2_X2 U11313 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19783), .ZN(n19787) );
  BUF_X2 U11314 ( .A(n10300), .Z(n13611) );
  BUF_X4 U11315 ( .A(n10300), .Z(n11136) );
  BUF_X2 U11316 ( .A(n15738), .Z(n17259) );
  BUF_X2 U11317 ( .A(n15739), .Z(n17268) );
  CLKBUF_X3 U11318 ( .A(n15751), .Z(n17260) );
  OR2_X1 U11319 ( .A1(n16983), .A2(n11814), .ZN(n10232) );
  NOR2_X4 U11320 ( .A1(n11813), .A2(n11815), .ZN(n15648) );
  NOR2_X1 U11321 ( .A1(n18885), .A2(n17932), .ZN(n18920) );
  OR2_X1 U11322 ( .A1(n11815), .A2(n11814), .ZN(n15605) );
  BUF_X4 U11323 ( .A(n15742), .Z(n9596) );
  NOR2_X1 U11324 ( .A1(n11812), .A2(n11811), .ZN(n15729) );
  INV_X2 U11325 ( .A(n16603), .ZN(n16605) );
  OR3_X2 U11326 ( .A1(n18884), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18181) );
  OR2_X2 U11327 ( .A1(n11156), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20068) );
  AND2_X1 U11328 ( .A1(n12425), .A2(n14287), .ZN(n10305) );
  AND2_X1 U11329 ( .A1(n10242), .A2(n10245), .ZN(n10816) );
  INV_X1 U11330 ( .A(n13383), .ZN(n9597) );
  AND2_X2 U11331 ( .A1(n12425), .A2(n10243), .ZN(n10475) );
  NAND2_X1 U11332 ( .A1(n18905), .A2(n18899), .ZN(n16983) );
  NAND2_X1 U11333 ( .A1(n18892), .A2(n18880), .ZN(n11814) );
  NOR2_X2 U11334 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U11335 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18740) );
  INV_X1 U11336 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18899) );
  INV_X2 U11337 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18892) );
  INV_X1 U11338 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18880) );
  INV_X1 U11339 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10237) );
  AND2_X1 U11340 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12304) );
  INV_X4 U11341 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U11342 ( .A1(n12567), .A2(n10221), .ZN(n10217) );
  NAND2_X1 U11343 ( .A1(n9911), .A2(n10461), .ZN(n10546) );
  NOR2_X4 U11344 ( .A1(n16329), .A2(n16330), .ZN(n16328) );
  NAND2_X2 U11345 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12308) );
  AND2_X1 U11346 ( .A1(n11258), .A2(n11392), .ZN(n9857) );
  BUF_X2 U11347 ( .A(n13417), .Z(n9598) );
  INV_X2 U11348 ( .A(n13242), .ZN(n9600) );
  NAND2_X2 U11349 ( .A1(n9883), .A2(n9882), .ZN(n15494) );
  AND3_X1 U11350 ( .A1(n11550), .A2(n15449), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U11351 ( .A1(n12978), .A2(n12959), .ZN(n13544) );
  XNOR2_X2 U11352 ( .A(n10397), .B(n10396), .ZN(n10461) );
  OAI22_X2 U11353 ( .A1(n12171), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n10547), 
        .B2(n10469), .ZN(n10397) );
  NAND2_X1 U11355 ( .A1(n9885), .A2(n9884), .ZN(n15559) );
  AND2_X2 U11356 ( .A1(n15559), .A2(n15537), .ZN(n11307) );
  OR2_X1 U11357 ( .A1(n11321), .A2(n16435), .ZN(n9604) );
  OR2_X1 U11358 ( .A1(n11321), .A2(n16435), .ZN(n9605) );
  NAND2_X2 U11359 ( .A1(n11556), .A2(n12044), .ZN(n11700) );
  OR2_X2 U11360 ( .A1(n12299), .A2(n9592), .ZN(n11377) );
  NAND2_X1 U11361 ( .A1(n11344), .A2(n11347), .ZN(n15448) );
  AND2_X2 U11362 ( .A1(n12704), .A2(n10218), .ZN(n14662) );
  NAND2_X2 U11363 ( .A1(n11363), .A2(n9592), .ZN(n11372) );
  NAND4_X2 U11364 ( .A1(n11436), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n10067) );
  XNOR2_X2 U11365 ( .A(n11474), .B(n11475), .ZN(n15119) );
  NAND2_X2 U11366 ( .A1(n14602), .A2(n14603), .ZN(n10210) );
  XNOR2_X2 U11367 ( .A(n13314), .B(n13311), .ZN(n14602) );
  NOR2_X2 U11368 ( .A1(n11283), .A2(n11282), .ZN(n11766) );
  INV_X4 U11369 ( .A(n13249), .ZN(n9607) );
  OR2_X4 U11370 ( .A1(n12308), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13249) );
  NAND2_X2 U11371 ( .A1(n11322), .A2(n9870), .ZN(n11770) );
  INV_X2 U11372 ( .A(n16408), .ZN(n11280) );
  NAND2_X1 U11373 ( .A1(n11301), .A2(n16408), .ZN(n12044) );
  NAND2_X2 U11374 ( .A1(n13133), .A2(n13132), .ZN(n14643) );
  INV_X4 U11375 ( .A(n13429), .ZN(n9608) );
  NAND2_X1 U11376 ( .A1(n11770), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U11377 ( .A1(n11770), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9610) );
  AOI211_X1 U11378 ( .C1(n9592), .C2(n19115), .A(n12841), .B(n12840), .ZN(
        n12842) );
  INV_X2 U11379 ( .A(n19021), .ZN(n19115) );
  CLKBUF_X1 U11380 ( .A(n10419), .Z(n13600) );
  INV_X1 U11381 ( .A(n9806), .ZN(n9801) );
  AND3_X1 U11382 ( .A1(n11300), .A2(n16408), .A3(n11607), .ZN(n11703) );
  NAND4_X1 U11383 ( .A1(n10170), .A2(n11382), .A3(n10169), .A4(n11381), .ZN(
        n10065) );
  NOR2_X1 U11384 ( .A1(n11362), .A2(n11358), .ZN(n10169) );
  NOR2_X1 U11385 ( .A1(n11814), .A2(n18740), .ZN(n15742) );
  NAND2_X1 U11386 ( .A1(n10354), .A2(n9622), .ZN(n9821) );
  CLKBUF_X2 U11388 ( .A(n10315), .Z(n10988) );
  OAI21_X1 U11389 ( .B1(n10660), .B2(n10507), .A(n10506), .ZN(n10564) );
  OAI21_X1 U11390 ( .B1(n10660), .B2(n10495), .A(n10494), .ZN(n10555) );
  AND2_X1 U11391 ( .A1(n10339), .A2(n12978), .ZN(n10429) );
  NOR2_X1 U11392 ( .A1(n14838), .A2(n14347), .ZN(n9933) );
  NAND2_X1 U11393 ( .A1(n11326), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11313) );
  AND2_X1 U11394 ( .A1(n10062), .A2(n11748), .ZN(n9788) );
  NAND2_X1 U11395 ( .A1(n9887), .A2(n16408), .ZN(n9886) );
  AOI21_X1 U11396 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19809), .A(
        n11575), .ZN(n11571) );
  AOI21_X1 U11397 ( .B1(n18750), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11905), .ZN(n11911) );
  NOR2_X1 U11398 ( .A1(n13063), .A2(n13062), .ZN(n11905) );
  NAND2_X1 U11399 ( .A1(n17315), .A2(n15683), .ZN(n11896) );
  AND2_X1 U11400 ( .A1(n10158), .A2(n11152), .ZN(n9766) );
  NAND2_X1 U11401 ( .A1(n13985), .A2(n9945), .ZN(n9944) );
  NAND2_X1 U11402 ( .A1(n16055), .A2(n14089), .ZN(n9945) );
  NOR2_X1 U11403 ( .A1(n10393), .A2(n10392), .ZN(n10547) );
  OR2_X1 U11405 ( .A1(n14507), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14796) );
  AOI211_X1 U11406 ( .C1(n13364), .C2(n13366), .A(n13363), .B(n13407), .ZN(
        n13365) );
  AND2_X1 U11407 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  INV_X1 U11408 ( .A(n14645), .ZN(n9877) );
  AND2_X1 U11409 ( .A1(n9690), .A2(n9879), .ZN(n9878) );
  INV_X1 U11410 ( .A(n14619), .ZN(n9879) );
  NAND3_X1 U11411 ( .A1(n12100), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n15526), 
        .ZN(n13363) );
  AND2_X1 U11412 ( .A1(n19004), .A2(n14896), .ZN(n14856) );
  AOI21_X1 U11413 ( .B1(n11544), .B2(n9774), .A(n9675), .ZN(n9773) );
  INV_X1 U11414 ( .A(n16299), .ZN(n9775) );
  NAND2_X1 U11415 ( .A1(n11326), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11328) );
  AND2_X1 U11416 ( .A1(n14395), .A2(n9916), .ZN(n14890) );
  NOR2_X1 U11417 ( .A1(n14879), .A2(n9917), .ZN(n9916) );
  INV_X1 U11418 ( .A(n14372), .ZN(n9917) );
  NOR2_X1 U11419 ( .A1(n15104), .A2(n10011), .ZN(n10010) );
  INV_X1 U11420 ( .A(n10074), .ZN(n10011) );
  NAND2_X1 U11421 ( .A1(n9777), .A2(n11685), .ZN(n14901) );
  NAND2_X1 U11422 ( .A1(n11544), .A2(n16299), .ZN(n9777) );
  NAND2_X1 U11423 ( .A1(n11766), .A2(n11284), .ZN(n11322) );
  AND4_X1 U11424 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11641) );
  AND4_X1 U11425 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11642) );
  AND2_X1 U11426 ( .A1(n11425), .A2(n11451), .ZN(n10062) );
  NAND2_X1 U11427 ( .A1(n9949), .A2(n9950), .ZN(n15838) );
  AND2_X1 U11428 ( .A1(n18041), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U11429 ( .A(n15831), .ZN(n9949) );
  NOR2_X1 U11430 ( .A1(n17445), .A2(n15819), .ZN(n15821) );
  AND2_X1 U11431 ( .A1(n9703), .A2(n12942), .ZN(n9770) );
  INV_X1 U11432 ( .A(n13043), .ZN(n10155) );
  NAND2_X1 U11433 ( .A1(n12977), .A2(n12976), .ZN(n13005) );
  AOI21_X1 U11434 ( .B1(n10111), .B2(n9591), .A(n15007), .ZN(n10109) );
  NAND2_X1 U11435 ( .A1(n10208), .A2(n10207), .ZN(n10206) );
  INV_X1 U11436 ( .A(n14615), .ZN(n10207) );
  NAND2_X1 U11437 ( .A1(n11191), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9884) );
  NAND2_X1 U11438 ( .A1(n11196), .A2(n11392), .ZN(n9885) );
  NAND2_X1 U11439 ( .A1(n11742), .A2(n9708), .ZN(n10188) );
  OR2_X1 U11440 ( .A1(n10083), .A2(n15025), .ZN(n10081) );
  NAND2_X1 U11441 ( .A1(n15024), .A2(n15085), .ZN(n10082) );
  NAND2_X1 U11442 ( .A1(n11676), .A2(n11675), .ZN(n16296) );
  INV_X1 U11443 ( .A(n15113), .ZN(n10087) );
  NAND2_X1 U11444 ( .A1(n14951), .A2(n9662), .ZN(n9749) );
  NOR2_X1 U11445 ( .A1(n9651), .A2(n14887), .ZN(n14888) );
  AOI21_X1 U11446 ( .B1(n9795), .B2(n9615), .A(n9792), .ZN(n9791) );
  NAND2_X1 U11447 ( .A1(n15094), .A2(n9794), .ZN(n9793) );
  INV_X1 U11448 ( .A(n15013), .ZN(n9792) );
  NOR2_X1 U11449 ( .A1(n15077), .A2(n10084), .ZN(n10083) );
  INV_X1 U11450 ( .A(n15084), .ZN(n10084) );
  AND2_X1 U11451 ( .A1(n9632), .A2(n16245), .ZN(n10070) );
  NAND2_X1 U11452 ( .A1(n10065), .A2(n11425), .ZN(n10064) );
  AND2_X1 U11453 ( .A1(n11622), .A2(n12098), .ZN(n11771) );
  NAND2_X1 U11454 ( .A1(n12060), .A2(n12059), .ZN(n12195) );
  NAND2_X1 U11455 ( .A1(n16368), .A2(n12284), .ZN(n12060) );
  AOI211_X1 U11456 ( .C1(n17269), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n11888), .B(n11887), .ZN(n11889) );
  NOR2_X1 U11457 ( .A1(n17929), .A2(n17921), .ZN(n17919) );
  NAND2_X1 U11458 ( .A1(n17725), .A2(n17829), .ZN(n17683) );
  NAND2_X1 U11459 ( .A1(n10172), .A2(n17829), .ZN(n15837) );
  AND2_X1 U11460 ( .A1(n9719), .A2(n18161), .ZN(n10173) );
  INV_X1 U11461 ( .A(n20083), .ZN(n20071) );
  NOR2_X2 U11462 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19799) );
  NAND2_X1 U11463 ( .A1(n10036), .A2(n10035), .ZN(n10576) );
  NOR2_X1 U11464 ( .A1(n10508), .A2(n10562), .ZN(n10035) );
  INV_X1 U11465 ( .A(n10563), .ZN(n10036) );
  INV_X1 U11466 ( .A(n12162), .ZN(n12965) );
  AND2_X1 U11467 ( .A1(n11549), .A2(n11548), .ZN(n11559) );
  OR2_X1 U11468 ( .A1(n11584), .A2(n11563), .ZN(n11549) );
  NAND2_X1 U11469 ( .A1(n11560), .A2(n11554), .ZN(n11573) );
  NAND2_X1 U11470 ( .A1(n11309), .A2(n16408), .ZN(n9740) );
  AOI21_X1 U11471 ( .B1(n9989), .B2(n9991), .A(n14992), .ZN(n9988) );
  NOR2_X1 U11472 ( .A1(n9991), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9986) );
  INV_X1 U11473 ( .A(n11508), .ZN(n9744) );
  NAND3_X1 U11474 ( .A1(n11285), .A2(n11302), .A3(n9887), .ZN(n11308) );
  AND2_X1 U11475 ( .A1(n11303), .A2(n11301), .ZN(n11707) );
  NOR2_X1 U11476 ( .A1(n15543), .A2(n11297), .ZN(n11233) );
  AND2_X1 U11477 ( .A1(n17441), .A2(n15799), .ZN(n15784) );
  AND2_X1 U11478 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n9754) );
  INV_X1 U11479 ( .A(n12173), .ZN(n12211) );
  AND2_X1 U11480 ( .A1(n11127), .A2(n9692), .ZN(n10158) );
  NOR2_X1 U11481 ( .A1(n13695), .A2(n10161), .ZN(n10160) );
  INV_X1 U11482 ( .A(n13708), .ZN(n10161) );
  NOR2_X1 U11483 ( .A1(n13739), .A2(n9762), .ZN(n9761) );
  INV_X1 U11484 ( .A(n13793), .ZN(n9762) );
  NAND2_X1 U11485 ( .A1(n10151), .A2(n13887), .ZN(n10150) );
  INV_X1 U11486 ( .A(n10153), .ZN(n10151) );
  INV_X1 U11487 ( .A(n13625), .ZN(n11144) );
  NAND2_X1 U11488 ( .A1(n12166), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13625) );
  XNOR2_X1 U11489 ( .A(n10587), .B(n10586), .ZN(n10733) );
  INV_X1 U11490 ( .A(n12655), .ZN(n10723) );
  INV_X1 U11491 ( .A(n13947), .ZN(n10032) );
  NOR2_X1 U11492 ( .A1(n9910), .A2(n9903), .ZN(n10616) );
  NAND2_X1 U11493 ( .A1(n13990), .A2(n9904), .ZN(n9903) );
  INV_X1 U11494 ( .A(n13938), .ZN(n9904) );
  INV_X1 U11495 ( .A(n9837), .ZN(n9835) );
  NAND2_X1 U11496 ( .A1(n9838), .A2(n14021), .ZN(n9837) );
  INV_X1 U11497 ( .A(n10144), .ZN(n9838) );
  NAND2_X1 U11498 ( .A1(n14029), .A2(n16027), .ZN(n9914) );
  NOR2_X1 U11499 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  INV_X1 U11500 ( .A(n12868), .ZN(n10018) );
  OR2_X1 U11501 ( .A1(n12853), .A2(n10020), .ZN(n10019) );
  INV_X1 U11502 ( .A(n12859), .ZN(n10020) );
  AND2_X1 U11503 ( .A1(n12144), .A2(n12143), .ZN(n12971) );
  NAND2_X1 U11504 ( .A1(n10138), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10136) );
  INV_X1 U11505 ( .A(n10522), .ZN(n10141) );
  NAND2_X1 U11506 ( .A1(n20101), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10468) );
  NAND2_X1 U11507 ( .A1(n20124), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U11508 ( .A1(n10429), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10660) );
  OR2_X1 U11509 ( .A1(n10481), .A2(n10480), .ZN(n10566) );
  NAND2_X2 U11510 ( .A1(n10469), .A2(n10468), .ZN(n10665) );
  AOI221_X1 U11511 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10664), 
        .C1(n16173), .C2(n10664), .A(n10663), .ZN(n12000) );
  OR2_X1 U11512 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  MUX2_X1 U11513 ( .A(n10340), .B(n10339), .S(n20132), .Z(n10342) );
  NAND2_X1 U11514 ( .A1(n10467), .A2(n10466), .ZN(n20234) );
  NOR2_X1 U11515 ( .A1(n20349), .A2(n20348), .ZN(n20442) );
  AND2_X1 U11516 ( .A1(n11615), .A2(n11614), .ZN(n11694) );
  NAND2_X1 U11517 ( .A1(n19827), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11548) );
  AND3_X1 U11518 ( .A1(n11588), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11571), .ZN(n11671) );
  NAND2_X1 U11519 ( .A1(n10112), .A2(n15850), .ZN(n10111) );
  NAND2_X1 U11520 ( .A1(n14350), .A2(n14842), .ZN(n14846) );
  INV_X1 U11521 ( .A(n14844), .ZN(n14350) );
  INV_X1 U11522 ( .A(n9933), .ZN(n14834) );
  INV_X1 U11523 ( .A(n14812), .ZN(n9750) );
  NAND2_X1 U11524 ( .A1(n9674), .A2(n11682), .ZN(n14507) );
  AND2_X1 U11525 ( .A1(n11682), .A2(n9926), .ZN(n14787) );
  INV_X1 U11526 ( .A(n11680), .ZN(n11681) );
  AND2_X2 U11527 ( .A1(n11679), .A2(n11678), .ZN(n11682) );
  NAND2_X1 U11528 ( .A1(n11682), .A2(n11681), .ZN(n11687) );
  NAND2_X1 U11529 ( .A1(n9925), .A2(n9924), .ZN(n11649) );
  OAI21_X1 U11530 ( .B1(n11743), .B2(n11646), .A(n9590), .ZN(n9925) );
  AND2_X1 U11531 ( .A1(n9635), .A2(n14445), .ZN(n10195) );
  OR2_X1 U11532 ( .A1(n10199), .A2(n9700), .ZN(n10198) );
  NAND2_X1 U11533 ( .A1(n10102), .A2(n12552), .ZN(n10101) );
  INV_X1 U11534 ( .A(n12543), .ZN(n10102) );
  NAND2_X1 U11535 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  INV_X1 U11536 ( .A(n14575), .ZN(n10105) );
  INV_X1 U11537 ( .A(n14370), .ZN(n10106) );
  INV_X1 U11538 ( .A(n14582), .ZN(n10107) );
  AND2_X1 U11539 ( .A1(n14979), .A2(n14886), .ZN(n14946) );
  NAND2_X1 U11540 ( .A1(n10100), .A2(n12696), .ZN(n10099) );
  INV_X1 U11541 ( .A(n10101), .ZN(n10100) );
  OR2_X1 U11542 ( .A1(n10193), .A2(n12354), .ZN(n10192) );
  INV_X1 U11543 ( .A(n14307), .ZN(n13540) );
  NAND2_X1 U11544 ( .A1(n11677), .A2(n11643), .ZN(n9982) );
  NAND2_X1 U11545 ( .A1(n11335), .A2(n9808), .ZN(n9747) );
  NAND2_X1 U11546 ( .A1(n9746), .A2(n11343), .ZN(n9745) );
  NAND2_X1 U11547 ( .A1(n11287), .A2(n11278), .ZN(n12306) );
  NOR2_X1 U11548 ( .A1(n9886), .A2(n13480), .ZN(n11277) );
  NAND2_X1 U11549 ( .A1(n10215), .A2(n9887), .ZN(n10214) );
  NAND2_X1 U11550 ( .A1(n12058), .A2(n12070), .ZN(n12287) );
  AOI221_X1 U11551 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11571), 
        .C1(n11588), .C2(n11571), .A(n11555), .ZN(n11579) );
  AOI22_X1 U11552 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11229) );
  INV_X1 U11553 ( .A(n19831), .ZN(n15477) );
  NOR2_X1 U11554 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  INV_X1 U11555 ( .A(n15731), .ZN(n9972) );
  NAND2_X1 U11556 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18892), .ZN(
        n11811) );
  NAND2_X1 U11557 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18905), .ZN(
        n11812) );
  NOR2_X1 U11558 ( .A1(n11811), .A2(n16983), .ZN(n15738) );
  NOR2_X1 U11559 ( .A1(n16667), .A2(n17927), .ZN(n10060) );
  NOR2_X1 U11560 ( .A1(n16448), .A2(n17818), .ZN(n16452) );
  NOR2_X1 U11561 ( .A1(n17433), .A2(n15826), .ZN(n15827) );
  AND2_X1 U11562 ( .A1(n9959), .A2(n9841), .ZN(n15842) );
  INV_X1 U11563 ( .A(n17642), .ZN(n9959) );
  AND2_X1 U11564 ( .A1(n17623), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9841) );
  NOR2_X1 U11565 ( .A1(n15825), .A2(n17858), .ZN(n15828) );
  AND2_X1 U11566 ( .A1(n9951), .A2(n9678), .ZN(n15820) );
  NOR2_X1 U11567 ( .A1(n18316), .A2(n18287), .ZN(n15676) );
  XNOR2_X1 U11568 ( .A(n17455), .B(n15817), .ZN(n15818) );
  OAI22_X1 U11569 ( .A1(n18899), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18750), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13063) );
  AOI21_X1 U11570 ( .B1(n11911), .B2(n11910), .A(n11909), .ZN(n15684) );
  INV_X1 U11571 ( .A(n11896), .ZN(n11881) );
  AND2_X1 U11572 ( .A1(n13075), .A2(n18721), .ZN(n13067) );
  NOR2_X1 U11573 ( .A1(n16616), .A2(n15673), .ZN(n15677) );
  INV_X1 U11574 ( .A(n18729), .ZN(n18732) );
  NAND2_X1 U11575 ( .A1(n12137), .A2(n12136), .ZN(n12207) );
  OR2_X1 U11576 ( .A1(n12973), .A2(n12134), .ZN(n12137) );
  AND4_X1 U11577 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10269) );
  AND4_X1 U11578 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10270) );
  AND2_X1 U11579 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n10949), .ZN(
        n10950) );
  INV_X1 U11580 ( .A(n10948), .ZN(n10949) );
  NAND2_X1 U11581 ( .A1(n10950), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10983) );
  NOR2_X1 U11582 ( .A1(n12929), .A2(n10165), .ZN(n10164) );
  INV_X1 U11583 ( .A(n10224), .ZN(n10165) );
  NAND2_X1 U11584 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U11585 ( .A1(n9827), .A2(n10542), .ZN(n12484) );
  INV_X1 U11586 ( .A(n13662), .ZN(n10021) );
  NAND2_X1 U11587 ( .A1(n10032), .A2(n9840), .ZN(n9839) );
  AND2_X1 U11588 ( .A1(n10030), .A2(n14115), .ZN(n9840) );
  NOR2_X1 U11589 ( .A1(n9634), .A2(n14094), .ZN(n9901) );
  NAND2_X1 U11590 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U11591 ( .A1(n9944), .A2(n9940), .ZN(n9939) );
  NOR3_X1 U11592 ( .A1(n13938), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U11593 ( .A1(n13025), .A2(n10601), .ZN(n10603) );
  AOI21_X1 U11594 ( .B1(n9936), .B2(n10583), .A(n9669), .ZN(n9935) );
  XNOR2_X1 U11595 ( .A(n10456), .B(n10457), .ZN(n10680) );
  INV_X1 U11596 ( .A(n19849), .ZN(n12976) );
  INV_X1 U11597 ( .A(n20208), .ZN(n20205) );
  OR2_X1 U11598 ( .A1(n20595), .A2(n9587), .ZN(n20515) );
  INV_X1 U11599 ( .A(n10688), .ZN(n20507) );
  NOR2_X1 U11600 ( .A1(n9919), .A2(n14879), .ZN(n9918) );
  NAND2_X1 U11601 ( .A1(n14889), .A2(n14372), .ZN(n9919) );
  NOR3_X1 U11602 ( .A1(n14871), .A2(n9921), .A3(n14436), .ZN(n14371) );
  NAND2_X1 U11603 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  NAND2_X1 U11604 ( .A1(n14395), .A2(n14372), .ZN(n14881) );
  OR2_X1 U11605 ( .A1(n14473), .A2(n10111), .ZN(n10110) );
  NAND2_X1 U11606 ( .A1(n14787), .A2(n11720), .ZN(n14819) );
  INV_X1 U11607 ( .A(n14653), .ZN(n10091) );
  AND2_X1 U11608 ( .A1(n13426), .A2(n11392), .ZN(n13224) );
  AND2_X1 U11609 ( .A1(n9691), .A2(n9633), .ZN(n9869) );
  NAND2_X1 U11610 ( .A1(n14597), .A2(n9645), .ZN(n10211) );
  INV_X1 U11611 ( .A(n13266), .ZN(n10205) );
  OR2_X1 U11612 ( .A1(n9876), .A2(n9875), .ZN(n9873) );
  NAND2_X1 U11613 ( .A1(n9876), .A2(n9875), .ZN(n9874) );
  OR2_X1 U11614 ( .A1(n14613), .A2(n14615), .ZN(n10209) );
  AND2_X1 U11615 ( .A1(n10219), .A2(n12902), .ZN(n10218) );
  NOR2_X1 U11616 ( .A1(n10188), .A2(n10186), .ZN(n10185) );
  INV_X1 U11617 ( .A(n12563), .ZN(n10186) );
  XNOR2_X1 U11618 ( .A(n12785), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14918) );
  OR3_X1 U11619 ( .A1(n10093), .A2(n10095), .A3(n14404), .ZN(n10092) );
  AND2_X1 U11620 ( .A1(n9630), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10113) );
  NAND2_X1 U11621 ( .A1(n14340), .A2(n9630), .ZN(n14341) );
  NAND2_X1 U11622 ( .A1(n14492), .A2(n12923), .ZN(n14672) );
  AND2_X1 U11623 ( .A1(n9977), .A2(n9980), .ZN(n9976) );
  NAND2_X1 U11624 ( .A1(n11677), .A2(n9975), .ZN(n9974) );
  NAND2_X1 U11625 ( .A1(n9978), .A2(n14896), .ZN(n9977) );
  NAND2_X1 U11626 ( .A1(n14971), .A2(n14946), .ZN(n14949) );
  NAND2_X1 U11627 ( .A1(n14873), .A2(n14896), .ZN(n9748) );
  NOR2_X1 U11628 ( .A1(n9647), .A2(n9797), .ZN(n9796) );
  INV_X1 U11629 ( .A(n10230), .ZN(n9797) );
  AND2_X1 U11630 ( .A1(n9632), .A2(n10007), .ZN(n10006) );
  NAND2_X1 U11631 ( .A1(n10008), .A2(n16254), .ZN(n10007) );
  NAND2_X1 U11632 ( .A1(n10075), .A2(n10010), .ZN(n9799) );
  NAND2_X1 U11633 ( .A1(n14900), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14902) );
  INV_X1 U11634 ( .A(n9819), .ZN(n9818) );
  OAI21_X1 U11635 ( .B1(n9789), .B2(n11643), .A(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U11636 ( .A1(n11667), .A2(n11666), .ZN(n12764) );
  OAI21_X1 U11637 ( .B1(n9816), .B2(n9815), .A(n14543), .ZN(n11665) );
  INV_X1 U11638 ( .A(n9973), .ZN(n9815) );
  INV_X2 U11639 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U11640 ( .A1(n12198), .A2(n12197), .ZN(n12292) );
  NOR2_X1 U11641 ( .A1(n15543), .A2(n12046), .ZN(n11299) );
  OR2_X1 U11642 ( .A1(n19803), .A2(n19831), .ZN(n19406) );
  NAND2_X1 U11643 ( .A1(n19803), .A2(n19831), .ZN(n19598) );
  NAND2_X1 U11644 ( .A1(n19812), .A2(n19823), .ZN(n19659) );
  INV_X1 U11645 ( .A(n19463), .ZN(n19655) );
  NOR2_X1 U11646 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16426) );
  INV_X1 U11647 ( .A(n17600), .ZN(n10040) );
  NOR2_X1 U11648 ( .A1(n16707), .A2(n9694), .ZN(n10038) );
  NAND2_X1 U11649 ( .A1(n9854), .A2(n9851), .ZN(n9850) );
  AOI21_X1 U11650 ( .B1(n17237), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(n9852), .ZN(n9851) );
  NAND2_X1 U11651 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9854) );
  OAI21_X1 U11652 ( .B1(n9642), .B2(n20791), .A(n9853), .ZN(n9852) );
  NOR2_X1 U11653 ( .A1(n9637), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9846) );
  OR2_X1 U11654 ( .A1(n17601), .A2(n10180), .ZN(n10179) );
  NAND2_X1 U11655 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  NAND2_X1 U11656 ( .A1(n17818), .A2(n17941), .ZN(n10181) );
  INV_X1 U11657 ( .A(n17622), .ZN(n10182) );
  NAND2_X1 U11658 ( .A1(n9948), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17586) );
  INV_X1 U11659 ( .A(n10179), .ZN(n9948) );
  NOR2_X1 U11660 ( .A1(n17602), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17601) );
  NAND2_X1 U11661 ( .A1(n10184), .A2(n9689), .ZN(n10183) );
  NAND2_X1 U11662 ( .A1(n17730), .A2(n17633), .ZN(n10184) );
  NAND2_X1 U11663 ( .A1(n9842), .A2(n17683), .ZN(n17623) );
  AND2_X1 U11664 ( .A1(n10183), .A2(n17938), .ZN(n9842) );
  NOR2_X1 U11665 ( .A1(n9844), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9843) );
  INV_X1 U11666 ( .A(n15836), .ZN(n9844) );
  NOR2_X1 U11667 ( .A1(n18121), .A2(n18092), .ZN(n17757) );
  AOI21_X1 U11668 ( .B1(n18721), .B2(n18729), .A(n18720), .ZN(n18731) );
  NAND3_X1 U11669 ( .A1(n15783), .A2(n15782), .A3(n15781), .ZN(n16505) );
  NOR2_X1 U11670 ( .A1(n15831), .A2(n18161), .ZN(n17747) );
  NAND2_X1 U11671 ( .A1(n9845), .A2(n17870), .ZN(n17860) );
  OAI21_X1 U11672 ( .B1(n17871), .B2(n17872), .A(n18198), .ZN(n9845) );
  AND2_X1 U11673 ( .A1(n9956), .A2(n9957), .ZN(n17871) );
  INV_X1 U11674 ( .A(n15822), .ZN(n9956) );
  AOI21_X1 U11675 ( .B1(n10175), .B2(n9649), .A(n18206), .ZN(n15822) );
  OR2_X1 U11676 ( .A1(n9649), .A2(n18206), .ZN(n9954) );
  OR2_X1 U11677 ( .A1(n10175), .A2(n18206), .ZN(n9952) );
  XNOR2_X1 U11678 ( .A(n15820), .B(n18187), .ZN(n17897) );
  NAND2_X1 U11679 ( .A1(n9848), .A2(n9847), .ZN(n10175) );
  INV_X1 U11680 ( .A(n17898), .ZN(n9847) );
  INV_X1 U11681 ( .A(n17897), .ZN(n9848) );
  NOR2_X1 U11682 ( .A1(n17919), .A2(n15816), .ZN(n17911) );
  XNOR2_X1 U11683 ( .A(n15818), .B(n18234), .ZN(n17910) );
  OR2_X1 U11684 ( .A1(n17911), .A2(n17910), .ZN(n9951) );
  INV_X1 U11685 ( .A(n12500), .ZN(n20136) );
  INV_X1 U11686 ( .A(n13917), .ZN(n13906) );
  XNOR2_X1 U11687 ( .A(n13651), .B(n13650), .ZN(n14104) );
  OR2_X1 U11688 ( .A1(n13005), .A2(n13004), .ZN(n20083) );
  NAND2_X1 U11689 ( .A1(n20511), .A2(n10453), .ZN(n20540) );
  CLKBUF_X1 U11690 ( .A(n12171), .Z(n20479) );
  NOR2_X1 U11691 ( .A1(n11287), .A2(n12834), .ZN(n18946) );
  NAND2_X1 U11692 ( .A1(n10076), .A2(n10081), .ZN(n15071) );
  OAI21_X1 U11693 ( .B1(n19224), .B2(n19043), .A(n16240), .ZN(n9896) );
  INV_X1 U11694 ( .A(n19216), .ZN(n16287) );
  NAND2_X1 U11695 ( .A1(n12079), .A2(n12078), .ZN(n16305) );
  AND2_X1 U11696 ( .A1(n12074), .A2(n16421), .ZN(n19216) );
  OR2_X1 U11697 ( .A1(n14934), .A2(n9997), .ZN(n9994) );
  NAND2_X1 U11698 ( .A1(n10001), .A2(n9998), .ZN(n9997) );
  INV_X1 U11699 ( .A(n14899), .ZN(n9998) );
  NAND2_X1 U11700 ( .A1(n9992), .A2(n9650), .ZN(n9995) );
  OR2_X1 U11701 ( .A1(n14899), .A2(n9999), .ZN(n9993) );
  NAND2_X1 U11702 ( .A1(n14934), .A2(n14932), .ZN(n14923) );
  INV_X1 U11703 ( .A(n9784), .ZN(n9783) );
  AOI21_X1 U11704 ( .B1(n15322), .B2(n15321), .A(n15346), .ZN(n9784) );
  NAND2_X1 U11705 ( .A1(n10085), .A2(n15084), .ZN(n15078) );
  NAND2_X1 U11706 ( .A1(n15319), .A2(n15316), .ZN(n16376) );
  INV_X1 U11707 ( .A(n16652), .ZN(n10054) );
  NOR2_X1 U11708 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  NOR2_X1 U11709 ( .A1(n16987), .A2(n16654), .ZN(n10053) );
  INV_X1 U11710 ( .A(n16653), .ZN(n10052) );
  NAND2_X1 U11711 ( .A1(n17320), .A2(n17449), .ZN(n17319) );
  NAND2_X1 U11712 ( .A1(n17325), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17320) );
  NOR2_X1 U11713 ( .A1(n15727), .A2(n15726), .ZN(n17445) );
  AOI22_X1 U11714 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U11715 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U11716 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10409) );
  INV_X1 U11717 ( .A(n13209), .ZN(n13233) );
  OAI22_X1 U11718 ( .A1(n19307), .A2(n13369), .B1(n13196), .B2(n19502), .ZN(
        n11486) );
  AND2_X1 U11719 ( .A1(n14891), .A2(n15494), .ZN(n11302) );
  NOR2_X1 U11720 ( .A1(n15543), .A2(n9603), .ZN(n11285) );
  NAND2_X1 U11721 ( .A1(n11610), .A2(n11701), .ZN(n11305) );
  NAND2_X1 U11722 ( .A1(n11303), .A2(n15543), .ZN(n11306) );
  AOI22_X1 U11724 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U11725 ( .A1(n10331), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10898) );
  AOI21_X1 U11726 ( .B1(n10994), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n10129), .ZN(n10742) );
  AND2_X1 U11727 ( .A1(n13600), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10129) );
  AOI22_X1 U11728 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10514) );
  OR2_X1 U11729 ( .A1(n10493), .A2(n10492), .ZN(n10567) );
  OR2_X1 U11730 ( .A1(n10447), .A2(n10446), .ZN(n10529) );
  AOI22_X1 U11731 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11732 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10477) );
  AOI21_X1 U11733 ( .B1(n20474), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10629), .ZN(n10664) );
  AOI22_X1 U11734 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n10331), .ZN(n10295) );
  AOI22_X1 U11735 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10239) );
  NAND2_X1 U11736 ( .A1(n9826), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U11737 ( .A1(n9821), .A2(n20101), .ZN(n9820) );
  NOR2_X1 U11738 ( .A1(n9825), .A2(n12018), .ZN(n9824) );
  NOR2_X1 U11739 ( .A1(n15494), .A2(n11293), .ZN(n11281) );
  AND2_X1 U11740 ( .A1(n9927), .A2(n14519), .ZN(n9926) );
  AND2_X1 U11741 ( .A1(n11681), .A2(n9928), .ZN(n9927) );
  INV_X1 U11742 ( .A(n11686), .ZN(n9928) );
  NAND2_X1 U11743 ( .A1(n14828), .A2(n14542), .ZN(n9924) );
  AOI22_X1 U11744 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n9607), .ZN(n11194) );
  NOR2_X1 U11745 ( .A1(n11505), .A2(n11504), .ZN(n11752) );
  INV_X1 U11746 ( .A(n15494), .ZN(n12100) );
  INV_X1 U11747 ( .A(n9804), .ZN(n9746) );
  INV_X1 U11748 ( .A(n9802), .ZN(n9803) );
  OAI22_X1 U11749 ( .A1(n20842), .A2(n15480), .B1(n11523), .B2(n11433), .ZN(
        n11435) );
  NOR2_X1 U11750 ( .A1(n11364), .A2(n11359), .ZN(n10170) );
  NAND2_X1 U11751 ( .A1(n11285), .A2(n11302), .ZN(n11706) );
  NAND2_X1 U11752 ( .A1(n11305), .A2(n11306), .ZN(n11697) );
  OR2_X1 U11753 ( .A1(n17437), .A2(n15823), .ZN(n15826) );
  INV_X1 U11754 ( .A(n13686), .ZN(n10159) );
  INV_X1 U11755 ( .A(n13785), .ZN(n9760) );
  NAND2_X1 U11756 ( .A1(n10154), .A2(n10918), .ZN(n10153) );
  INV_X1 U11757 ( .A(n13802), .ZN(n10154) );
  AOI22_X1 U11758 ( .A1(n13609), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10806) );
  AND2_X1 U11759 ( .A1(n10829), .A2(n10157), .ZN(n10156) );
  OR2_X1 U11760 ( .A1(n13011), .A2(n13033), .ZN(n10157) );
  NOR2_X1 U11761 ( .A1(n10781), .A2(n19876), .ZN(n10785) );
  AND2_X1 U11762 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n10725), .ZN(
        n10734) );
  NOR2_X1 U11763 ( .A1(n20862), .A2(n10717), .ZN(n10725) );
  INV_X1 U11764 ( .A(n12656), .ZN(n10724) );
  NOR2_X1 U11765 ( .A1(n9595), .A2(n10031), .ZN(n10030) );
  NAND2_X1 U11766 ( .A1(n10619), .A2(n10620), .ZN(n10031) );
  NAND2_X1 U11767 ( .A1(n10024), .A2(n13592), .ZN(n10023) );
  NOR2_X1 U11768 ( .A1(n13696), .A2(n13681), .ZN(n10024) );
  NOR2_X1 U11769 ( .A1(n14188), .A2(n14187), .ZN(n10026) );
  AND2_X1 U11770 ( .A1(n10148), .A2(n10145), .ZN(n10144) );
  NAND2_X1 U11771 ( .A1(n14000), .A2(n9718), .ZN(n10145) );
  INV_X1 U11772 ( .A(n16028), .ZN(n10148) );
  INV_X1 U11773 ( .A(n13054), .ZN(n10012) );
  NOR2_X1 U11774 ( .A1(n10014), .A2(n13757), .ZN(n10013) );
  INV_X1 U11775 ( .A(n14250), .ZN(n10014) );
  INV_X1 U11776 ( .A(n10591), .ZN(n10598) );
  INV_X1 U11777 ( .A(n10574), .ZN(n9936) );
  NAND2_X1 U11778 ( .A1(n13646), .A2(n13585), .ZN(n13596) );
  INV_X1 U11779 ( .A(n13590), .ZN(n13044) );
  OR2_X1 U11780 ( .A1(n10426), .A2(n10425), .ZN(n10528) );
  NAND2_X1 U11781 ( .A1(n10524), .A2(n12959), .ZN(n12508) );
  NOR2_X1 U11782 ( .A1(n10660), .A2(n10628), .ZN(n10668) );
  NAND2_X1 U11783 ( .A1(n10344), .A2(n20120), .ZN(n12173) );
  AND2_X1 U11784 ( .A1(n10464), .A2(n20590), .ZN(n20350) );
  AOI21_X1 U11785 ( .B1(n16176), .B2(n16180), .A(n14285), .ZN(n20100) );
  AND2_X1 U11786 ( .A1(n12151), .A2(n12150), .ZN(n12442) );
  AND2_X1 U11787 ( .A1(n11561), .A2(n11560), .ZN(n11590) );
  NAND2_X1 U11788 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19836), .ZN(
        n11563) );
  OR2_X1 U11789 ( .A1(n11575), .A2(n11574), .ZN(n11647) );
  NOR2_X1 U11790 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n9923) );
  NOR2_X1 U11791 ( .A1(n14846), .A2(n14825), .ZN(n9931) );
  NAND2_X1 U11792 ( .A1(n9933), .A2(n14349), .ZN(n14844) );
  NAND2_X1 U11793 ( .A1(n14808), .A2(n14344), .ZN(n14812) );
  NAND2_X1 U11794 ( .A1(n14819), .A2(n14810), .ZN(n14808) );
  AND2_X1 U11795 ( .A1(n11673), .A2(n11672), .ZN(n11678) );
  NOR2_X2 U11796 ( .A1(n11656), .A2(n11650), .ZN(n11679) );
  INV_X1 U11797 ( .A(n13236), .ZN(n13211) );
  INV_X1 U11798 ( .A(n13224), .ZN(n13214) );
  OR2_X1 U11799 ( .A1(n11329), .A2(n11666), .ZN(n11341) );
  AOI21_X1 U11800 ( .B1(n11326), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11342), .ZN(n11775) );
  INV_X1 U11801 ( .A(n14608), .ZN(n10208) );
  NAND2_X1 U11802 ( .A1(n9603), .A2(n15494), .ZN(n13480) );
  AND2_X1 U11803 ( .A1(n14637), .A2(n14632), .ZN(n10220) );
  AOI22_X1 U11804 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11190) );
  OR2_X1 U11805 ( .A1(n14494), .A2(n10200), .ZN(n10199) );
  OR2_X1 U11806 ( .A1(n12331), .A2(n10194), .ZN(n10193) );
  INV_X1 U11807 ( .A(n12282), .ZN(n10194) );
  NOR2_X1 U11808 ( .A1(n14325), .A2(n10115), .ZN(n10114) );
  INV_X1 U11809 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U11810 ( .A1(n20861), .A2(n10125), .ZN(n10124) );
  INV_X1 U11811 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U11812 ( .A1(n16269), .A2(n10119), .ZN(n10118) );
  INV_X1 U11813 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U11814 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9975) );
  NAND2_X1 U11815 ( .A1(n9981), .A2(n11783), .ZN(n9980) );
  INV_X1 U11816 ( .A(n14532), .ZN(n9981) );
  NAND2_X1 U11817 ( .A1(n14952), .A2(n14946), .ZN(n14887) );
  AOI22_X1 U11818 ( .A1(n9988), .A2(n9990), .B1(n9984), .B2(n9986), .ZN(n9751)
         );
  INV_X1 U11819 ( .A(n15001), .ZN(n9984) );
  NOR2_X1 U11820 ( .A1(n9988), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U11821 ( .A1(n10094), .A2(n14426), .ZN(n10093) );
  INV_X1 U11822 ( .A(n14620), .ZN(n10094) );
  AND2_X1 U11823 ( .A1(n9796), .A2(n9795), .ZN(n9794) );
  INV_X1 U11824 ( .A(n9773), .ZN(n9733) );
  INV_X1 U11825 ( .A(n14906), .ZN(n9892) );
  INV_X1 U11826 ( .A(n15403), .ZN(n9891) );
  NOR2_X1 U11827 ( .A1(n10230), .A2(n10069), .ZN(n10068) );
  INV_X1 U11828 ( .A(n16245), .ZN(n10069) );
  INV_X1 U11829 ( .A(n14803), .ZN(n10008) );
  NOR2_X1 U11830 ( .A1(n10009), .A2(n10005), .ZN(n10004) );
  INV_X1 U11831 ( .A(n16254), .ZN(n10009) );
  INV_X1 U11832 ( .A(n10010), .ZN(n10005) );
  AND2_X1 U11833 ( .A1(n14791), .A2(n14792), .ZN(n10074) );
  INV_X1 U11834 ( .A(n14903), .ZN(n14904) );
  INV_X1 U11835 ( .A(n13534), .ZN(n14308) );
  NAND2_X1 U11836 ( .A1(n11689), .A2(n12806), .ZN(n14784) );
  NOR2_X1 U11837 ( .A1(n11541), .A2(n11540), .ZN(n11758) );
  NOR2_X1 U11838 ( .A1(n9789), .A2(n9787), .ZN(n9786) );
  INV_X1 U11839 ( .A(n10062), .ZN(n9787) );
  NAND2_X1 U11840 ( .A1(n10063), .A2(n11643), .ZN(n9816) );
  INV_X1 U11841 ( .A(n11308), .ZN(n12047) );
  AOI22_X1 U11842 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12604), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U11843 ( .A1(n9670), .A2(n9616), .ZN(n11727) );
  OR2_X1 U11844 ( .A1(n11411), .A2(n11410), .ZN(n11729) );
  OR2_X1 U11845 ( .A1(n11448), .A2(n11449), .ZN(n11743) );
  NOR2_X1 U11846 ( .A1(n9603), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11719) );
  AND2_X1 U11847 ( .A1(n12192), .A2(n9863), .ZN(n9862) );
  NAND2_X1 U11848 ( .A1(n12190), .A2(n9864), .ZN(n9863) );
  NAND2_X1 U11849 ( .A1(n9860), .A2(n9862), .ZN(n12459) );
  OR2_X1 U11850 ( .A1(n9592), .A2(n9865), .ZN(n9860) );
  OR2_X2 U11851 ( .A1(n11372), .A2(n11375), .ZN(n19397) );
  INV_X1 U11852 ( .A(n11375), .ZN(n11357) );
  NAND2_X1 U11853 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18899), .ZN(
        n11815) );
  NAND2_X1 U11854 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18880), .ZN(
        n11813) );
  NAND3_X1 U11855 ( .A1(n18905), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18719), .ZN(n17207) );
  NOR2_X1 U11856 ( .A1(n11813), .A2(n18740), .ZN(n15737) );
  NAND2_X1 U11857 ( .A1(n15737), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9853) );
  NOR2_X1 U11858 ( .A1(n11813), .A2(n11812), .ZN(n15753) );
  INV_X1 U11859 ( .A(n17207), .ZN(n15752) );
  NOR2_X1 U11860 ( .A1(n11815), .A2(n11811), .ZN(n15751) );
  OR2_X1 U11861 ( .A1(n11815), .A2(n11806), .ZN(n9642) );
  NOR2_X1 U11862 ( .A1(n17655), .A2(n17656), .ZN(n17610) );
  NAND2_X1 U11863 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10048) );
  AND2_X1 U11864 ( .A1(n15788), .A2(n15787), .ZN(n15799) );
  NOR2_X1 U11865 ( .A1(n16500), .A2(n15848), .ZN(n9946) );
  INV_X1 U11866 ( .A(n17586), .ZN(n9947) );
  AND2_X1 U11867 ( .A1(n10179), .A2(n9715), .ZN(n16448) );
  NAND2_X1 U11868 ( .A1(n17683), .A2(n17670), .ZN(n17671) );
  AND2_X1 U11869 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15786), .ZN(
        n15801) );
  AND2_X1 U11870 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18719) );
  OR2_X1 U11871 ( .A1(n11867), .A2(n9752), .ZN(n15683) );
  NOR3_X1 U11872 ( .A1(n18926), .A2(n13073), .A3(n16614), .ZN(n15914) );
  INV_X1 U11873 ( .A(n12961), .ZN(n10034) );
  NOR3_X1 U11874 ( .A1(n10339), .A2(n12208), .A3(n13848), .ZN(n10347) );
  AOI21_X1 U11875 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n11152) );
  AND2_X1 U11876 ( .A1(n13663), .A2(n13622), .ZN(n11148) );
  OR2_X1 U11877 ( .A1(n11126), .A2(n11125), .ZN(n13670) );
  AND2_X1 U11878 ( .A1(n11076), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11077) );
  AND2_X1 U11879 ( .A1(n13967), .A2(n13622), .ZN(n11056) );
  AND2_X1 U11880 ( .A1(n11034), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U11881 ( .A1(n11035), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U11882 ( .A1(n10984), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11033) );
  AND2_X1 U11883 ( .A1(n10968), .A2(n10967), .ZN(n13793) );
  AND2_X1 U11884 ( .A1(n10952), .A2(n10951), .ZN(n13887) );
  NOR2_X1 U11885 ( .A1(n10912), .A2(n15971), .ZN(n10914) );
  NAND2_X1 U11886 ( .A1(n10914), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10948) );
  INV_X1 U11887 ( .A(n13809), .ZN(n10152) );
  NOR2_X1 U11888 ( .A1(n10878), .A2(n10877), .ZN(n10879) );
  NAND2_X1 U11889 ( .A1(n10879), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10912) );
  NAND2_X1 U11890 ( .A1(n10846), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10878) );
  INV_X1 U11891 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U11892 ( .A1(n14034), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16053) );
  NOR2_X1 U11893 ( .A1(n20808), .A2(n10824), .ZN(n10830) );
  INV_X1 U11894 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20808) );
  AND2_X1 U11895 ( .A1(n10785), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10786) );
  AND2_X1 U11896 ( .A1(n10734), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U11897 ( .A1(n10741), .A2(n10740), .ZN(n12845) );
  AOI21_X1 U11898 ( .B1(n10722), .B2(n10855), .A(n10721), .ZN(n12655) );
  NAND2_X1 U11899 ( .A1(n10724), .A2(n10723), .ZN(n9769) );
  NOR2_X1 U11900 ( .A1(n10698), .A2(n10697), .ZN(n10709) );
  NAND2_X1 U11901 ( .A1(n12336), .A2(n10696), .ZN(n12453) );
  INV_X1 U11902 ( .A(n9763), .ZN(n10234) );
  OAI21_X1 U11903 ( .B1(n12454), .B2(n10678), .A(n9764), .ZN(n9763) );
  AOI21_X1 U11904 ( .B1(n10679), .B2(n9765), .A(n10149), .ZN(n9764) );
  INV_X1 U11905 ( .A(n10696), .ZN(n10149) );
  NOR2_X1 U11906 ( .A1(n13716), .A2(n10023), .ZN(n13671) );
  NOR2_X1 U11907 ( .A1(n13716), .A2(n10022), .ZN(n13682) );
  INV_X1 U11908 ( .A(n10024), .ZN(n10022) );
  AND2_X1 U11909 ( .A1(n13787), .A2(n13578), .ZN(n13725) );
  NOR2_X1 U11910 ( .A1(n13796), .A2(n13748), .ZN(n13787) );
  NAND2_X1 U11911 ( .A1(n9835), .A2(n9612), .ZN(n9834) );
  NAND2_X1 U11912 ( .A1(n10026), .A2(n10025), .ZN(n13796) );
  INV_X1 U11913 ( .A(n13794), .ZN(n10025) );
  INV_X1 U11914 ( .A(n10026), .ZN(n14190) );
  NOR2_X1 U11915 ( .A1(n13820), .A2(n13812), .ZN(n13814) );
  NAND2_X1 U11916 ( .A1(n13814), .A2(n13804), .ZN(n14188) );
  OR2_X1 U11917 ( .A1(n20056), .A2(n14235), .ZN(n14157) );
  OR2_X1 U11918 ( .A1(n14228), .A2(n14077), .ZN(n14195) );
  AND2_X1 U11919 ( .A1(n9833), .A2(n9837), .ZN(n13999) );
  OR2_X1 U11920 ( .A1(n13827), .A2(n13818), .ZN(n13820) );
  NAND2_X1 U11921 ( .A1(n13835), .A2(n13825), .ZN(n13827) );
  NAND2_X1 U11922 ( .A1(n14251), .A2(n14250), .ZN(n14253) );
  NAND2_X1 U11923 ( .A1(n14251), .A2(n10013), .ZN(n13759) );
  INV_X1 U11924 ( .A(n12936), .ZN(n10015) );
  NAND2_X1 U11925 ( .A1(n10016), .A2(n10017), .ZN(n12937) );
  NOR2_X1 U11926 ( .A1(n19932), .A2(n10019), .ZN(n12869) );
  NOR2_X1 U11927 ( .A1(n19932), .A2(n12853), .ZN(n16150) );
  INV_X1 U11928 ( .A(n10554), .ZN(n9831) );
  NAND2_X1 U11929 ( .A1(n16089), .A2(n16088), .ZN(n16087) );
  INV_X1 U11930 ( .A(n14263), .ZN(n20058) );
  NAND2_X1 U11931 ( .A1(n12224), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12226) );
  OR2_X1 U11932 ( .A1(n13005), .A2(n12986), .ZN(n20073) );
  OR2_X1 U11933 ( .A1(n12160), .A2(n13844), .ZN(n13001) );
  INV_X1 U11934 ( .A(n10135), .ZN(n10134) );
  NAND2_X1 U11935 ( .A1(n9672), .A2(n10402), .ZN(n10130) );
  NOR2_X1 U11936 ( .A1(n10141), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U11937 ( .A1(n10133), .A2(n10138), .ZN(n10132) );
  INV_X1 U11938 ( .A(n10452), .ZN(n10370) );
  NAND2_X1 U11939 ( .A1(n10460), .A2(n10459), .ZN(n10538) );
  OAI21_X1 U11940 ( .B1(n10382), .B2(n10381), .A(n9759), .ZN(n12171) );
  NAND2_X1 U11941 ( .A1(n20103), .A2(n20650), .ZN(n10483) );
  INV_X1 U11942 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12174) );
  INV_X1 U11943 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U11944 ( .A1(n10033), .A2(n12959), .ZN(n12985) );
  INV_X1 U11945 ( .A(n12144), .ZN(n10033) );
  OR2_X1 U11946 ( .A1(n20515), .A2(n20507), .ZN(n20475) );
  AOI21_X1 U11947 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20509), .A(n20148), 
        .ZN(n20597) );
  OR3_X1 U11948 ( .A1(n20355), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20100), 
        .ZN(n20137) );
  AND2_X1 U11949 ( .A1(n16397), .A2(n16395), .ZN(n12320) );
  AND2_X1 U11950 ( .A1(n11694), .A2(n11693), .ZN(n16398) );
  NAND2_X1 U11951 ( .A1(n11548), .A2(n11547), .ZN(n11584) );
  NOR2_X1 U11952 ( .A1(n11671), .A2(n11647), .ZN(n11591) );
  NAND2_X1 U11953 ( .A1(n14353), .A2(n14819), .ZN(n14395) );
  INV_X1 U11954 ( .A(n9923), .ZN(n9920) );
  AND2_X1 U11955 ( .A1(n14438), .A2(n14611), .ZN(n14419) );
  NAND2_X1 U11956 ( .A1(n9591), .A2(n14459), .ZN(n10112) );
  NAND2_X1 U11957 ( .A1(n9931), .A2(n14633), .ZN(n14456) );
  INV_X1 U11958 ( .A(n9931), .ZN(n14827) );
  NAND2_X1 U11959 ( .A1(n14340), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14339) );
  AND2_X1 U11960 ( .A1(n13448), .A2(n13447), .ZN(n14741) );
  NOR2_X1 U11961 ( .A1(n14337), .A2(n15054), .ZN(n14340) );
  NOR2_X1 U11962 ( .A1(n14821), .A2(n14820), .ZN(n19017) );
  AND2_X1 U11963 ( .A1(n14841), .A2(n14840), .ZN(n19038) );
  AND2_X1 U11964 ( .A1(n12703), .A2(n12911), .ZN(n10219) );
  AND2_X1 U11965 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  NOR2_X1 U11966 ( .A1(n12544), .A2(n12543), .ZN(n12553) );
  AND2_X1 U11967 ( .A1(n12569), .A2(n9716), .ZN(n10216) );
  AND2_X1 U11968 ( .A1(n11782), .A2(n11781), .ZN(n13097) );
  INV_X1 U11969 ( .A(n13365), .ZN(n10212) );
  NAND2_X1 U11970 ( .A1(n13452), .A2(n9693), .ZN(n14428) );
  AND2_X1 U11971 ( .A1(n13452), .A2(n10195), .ZN(n14447) );
  INV_X1 U11972 ( .A(n9876), .ZN(n9872) );
  NAND2_X1 U11973 ( .A1(n13452), .A2(n13451), .ZN(n14719) );
  NOR2_X2 U11974 ( .A1(n14493), .A2(n10196), .ZN(n14760) );
  NAND2_X1 U11975 ( .A1(n10197), .A2(n14758), .ZN(n10196) );
  INV_X1 U11976 ( .A(n10198), .ZN(n10197) );
  CLKBUF_X1 U11977 ( .A(n14643), .Z(n14644) );
  NOR2_X1 U11978 ( .A1(n14493), .A2(n10198), .ZN(n14772) );
  OR2_X1 U11979 ( .A1(n13116), .A2(n13115), .ZN(n14663) );
  CLKBUF_X1 U11980 ( .A(n14654), .Z(n14655) );
  NOR2_X1 U11981 ( .A1(n14493), .A2(n10199), .ZN(n14769) );
  AND2_X1 U11982 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  OR2_X1 U11983 ( .A1(n12332), .A2(n10193), .ZN(n12355) );
  INV_X1 U11984 ( .A(n19146), .ZN(n12098) );
  INV_X1 U11985 ( .A(n11184), .ZN(n13482) );
  NOR3_X1 U11986 ( .A1(n14323), .A2(n14986), .A3(n10122), .ZN(n14320) );
  NAND2_X1 U11987 ( .A1(n14324), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14323) );
  NOR2_X1 U11988 ( .A1(n14323), .A2(n14986), .ZN(n14322) );
  AND2_X1 U11989 ( .A1(n13509), .A2(n13508), .ZN(n14463) );
  OR2_X1 U11990 ( .A1(n14647), .A2(n14646), .ZN(n14649) );
  AND2_X1 U11991 ( .A1(n13502), .A2(n13501), .ZN(n14638) );
  AND2_X1 U11992 ( .A1(n14335), .A2(n10123), .ZN(n14338) );
  AND2_X1 U11993 ( .A1(n9631), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10123) );
  NAND2_X1 U11994 ( .A1(n14335), .A2(n9631), .ZN(n14336) );
  INV_X1 U11995 ( .A(n14671), .ZN(n10090) );
  NAND2_X1 U11996 ( .A1(n14492), .A2(n9611), .ZN(n14667) );
  NAND2_X1 U11997 ( .A1(n14335), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14334) );
  NOR2_X1 U11998 ( .A1(n14332), .A2(n16252), .ZN(n14335) );
  NAND2_X1 U11999 ( .A1(n14333), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14332) );
  AND2_X1 U12000 ( .A1(n14330), .A2(n10117), .ZN(n14333) );
  AND2_X1 U12001 ( .A1(n9617), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10117) );
  NOR2_X1 U12002 ( .A1(n12544), .A2(n10101), .ZN(n12697) );
  NAND2_X1 U12003 ( .A1(n14330), .A2(n9617), .ZN(n14331) );
  NAND2_X1 U12004 ( .A1(n14330), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14329) );
  NOR2_X1 U12005 ( .A1(n16306), .A2(n10127), .ZN(n10126) );
  NAND2_X1 U12006 ( .A1(n9776), .A2(n9773), .ZN(n14900) );
  NAND2_X1 U12007 ( .A1(n11545), .A2(n11546), .ZN(n9776) );
  NAND2_X1 U12008 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12787) );
  NOR2_X1 U12009 ( .A1(n12787), .A2(n14541), .ZN(n12789) );
  INV_X1 U12010 ( .A(n11325), .ZN(n9807) );
  OR3_X1 U12011 ( .A1(n10104), .A2(n10107), .A3(n14304), .ZN(n10103) );
  NOR2_X1 U12012 ( .A1(n14924), .A2(n10000), .ZN(n9999) );
  INV_X1 U12013 ( .A(n14932), .ZN(n10000) );
  INV_X1 U12014 ( .A(n14933), .ZN(n10002) );
  OR2_X1 U12015 ( .A1(n14882), .A2(n14937), .ZN(n14952) );
  XNOR2_X1 U12016 ( .A(n14949), .B(n14947), .ZN(n14960) );
  OR2_X1 U12017 ( .A1(n14884), .A2(n14883), .ZN(n14979) );
  NOR3_X1 U12018 ( .A1(n14621), .A2(n10095), .A3(n14620), .ZN(n14444) );
  NAND2_X1 U12019 ( .A1(n15032), .A2(n15124), .ZN(n15033) );
  CLKBUF_X1 U12020 ( .A(n14465), .Z(n14483) );
  AND2_X1 U12021 ( .A1(n14853), .A2(n15298), .ZN(n15049) );
  AND2_X1 U12022 ( .A1(n14847), .A2(n15310), .ZN(n15060) );
  NOR2_X1 U12023 ( .A1(n15359), .A2(n9619), .ZN(n9813) );
  AOI21_X1 U12024 ( .B1(n10081), .B2(n10079), .A(n10078), .ZN(n10077) );
  INV_X1 U12025 ( .A(n15069), .ZN(n10078) );
  AND2_X1 U12026 ( .A1(n10082), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U12027 ( .A1(n9641), .A2(n15366), .ZN(n9893) );
  INV_X1 U12028 ( .A(n16257), .ZN(n15360) );
  NAND2_X1 U12029 ( .A1(n15385), .A2(n9641), .ZN(n16257) );
  NOR2_X1 U12030 ( .A1(n12544), .A2(n10099), .ZN(n12699) );
  NOR2_X1 U12031 ( .A1(n10099), .A2(n10098), .ZN(n10097) );
  INV_X1 U12032 ( .A(n12679), .ZN(n10098) );
  AND2_X1 U12033 ( .A1(n12618), .A2(n12617), .ZN(n16330) );
  AND2_X1 U12034 ( .A1(n14797), .A2(n15374), .ZN(n15104) );
  NAND2_X1 U12035 ( .A1(n10075), .A2(n10074), .ZN(n15103) );
  OR2_X2 U12036 ( .A1(n12332), .A2(n10190), .ZN(n16329) );
  OR2_X1 U12037 ( .A1(n10192), .A2(n10191), .ZN(n10190) );
  INV_X1 U12038 ( .A(n12389), .ZN(n10191) );
  NAND2_X1 U12039 ( .A1(n12306), .A2(n16421), .ZN(n9870) );
  NAND2_X1 U12040 ( .A1(n9798), .A2(n11684), .ZN(n14783) );
  NAND2_X1 U12041 ( .A1(n9982), .A2(n14532), .ZN(n11683) );
  CLKBUF_X1 U12042 ( .A(n12306), .Z(n12307) );
  XNOR2_X1 U12043 ( .A(n12195), .B(n12196), .ZN(n12194) );
  AOI21_X1 U12044 ( .B1(n15448), .B2(n12284), .A(n12102), .ZN(n12193) );
  AND2_X1 U12045 ( .A1(n11581), .A2(n11580), .ZN(n16401) );
  INV_X1 U12046 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U12047 ( .A1(n9810), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9809) );
  NAND2_X1 U12048 ( .A1(n9812), .A2(n11392), .ZN(n9811) );
  OR2_X1 U12049 ( .A1(n19803), .A2(n18957), .ZN(n19399) );
  NAND2_X1 U12050 ( .A1(n11225), .A2(n11392), .ZN(n11232) );
  NAND2_X1 U12051 ( .A1(n11230), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U12052 ( .A1(n11201), .A2(n11392), .ZN(n11208) );
  OR2_X1 U12053 ( .A1(n19470), .A2(n19338), .ZN(n19599) );
  NAND2_X1 U12054 ( .A1(n19803), .A2(n15477), .ZN(n19470) );
  OR2_X1 U12055 ( .A1(n13482), .A2(n15115), .ZN(n15563) );
  OR2_X1 U12056 ( .A1(n13481), .A2(n15115), .ZN(n15564) );
  AOI21_X1 U12057 ( .B1(n15684), .B2(n11915), .A(n13064), .ZN(n18710) );
  OR2_X1 U12058 ( .A1(n10039), .A2(n16688), .ZN(n10037) );
  NOR2_X1 U12059 ( .A1(n10046), .A2(n16867), .ZN(n10045) );
  OR2_X1 U12060 ( .A1(n10048), .A2(n16873), .ZN(n10046) );
  INV_X1 U12061 ( .A(n17874), .ZN(n10047) );
  NAND2_X1 U12062 ( .A1(n18941), .A2(n17462), .ZN(n11918) );
  AND3_X1 U12063 ( .A1(n9676), .A2(n10177), .A3(n9970), .ZN(n10176) );
  NAND2_X1 U12064 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10177) );
  INV_X1 U12065 ( .A(n17499), .ZN(n17463) );
  NOR2_X1 U12066 ( .A1(n13072), .A2(n18792), .ZN(n17461) );
  NOR2_X1 U12067 ( .A1(n16614), .A2(n18773), .ZN(n17501) );
  NAND2_X1 U12068 ( .A1(n16482), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16479) );
  OR2_X1 U12069 ( .A1(n17686), .A2(n17685), .ZN(n17655) );
  NAND2_X1 U12070 ( .A1(n17758), .A2(n10041), .ZN(n17686) );
  AND2_X1 U12071 ( .A1(n9618), .A2(n10044), .ZN(n10041) );
  INV_X1 U12072 ( .A(n17701), .ZN(n10044) );
  NAND2_X1 U12073 ( .A1(n17758), .A2(n9618), .ZN(n17700) );
  NOR2_X1 U12074 ( .A1(n17734), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U12075 ( .A1(n17758), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17733) );
  NOR2_X1 U12076 ( .A1(n17776), .A2(n17778), .ZN(n17758) );
  AOI21_X1 U12077 ( .B1(n17687), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18653), .ZN(n17777) );
  NAND3_X1 U12078 ( .A1(n10047), .A2(n10045), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17776) );
  OR2_X1 U12079 ( .A1(n17874), .A2(n10048), .ZN(n17833) );
  NAND2_X1 U12080 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17874) );
  AND2_X1 U12081 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17892) );
  NOR2_X1 U12082 ( .A1(n16452), .A2(n9967), .ZN(n9966) );
  INV_X1 U12083 ( .A(n16451), .ZN(n9965) );
  NOR2_X1 U12084 ( .A1(n15899), .A2(n16460), .ZN(n16451) );
  OAI21_X1 U12085 ( .B1(n15842), .B2(n17964), .A(n9958), .ZN(n17602) );
  AND2_X1 U12086 ( .A1(n15841), .A2(n9698), .ZN(n9958) );
  NAND2_X1 U12087 ( .A1(n17671), .A2(n15840), .ZN(n17642) );
  NOR2_X1 U12088 ( .A1(n18119), .A2(n18016), .ZN(n18073) );
  OR2_X1 U12089 ( .A1(n18088), .A2(n17774), .ZN(n18092) );
  NAND2_X1 U12090 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17828), .ZN(
        n18119) );
  AOI21_X1 U12091 ( .B1(n15812), .B2(n15811), .A(n15810), .ZN(n17840) );
  NAND2_X1 U12092 ( .A1(n18165), .A2(n17829), .ZN(n17828) );
  NOR2_X1 U12093 ( .A1(n17869), .A2(n17868), .ZN(n17867) );
  NAND2_X1 U12094 ( .A1(n17871), .A2(n17872), .ZN(n17870) );
  INV_X1 U12095 ( .A(n17887), .ZN(n9953) );
  NOR2_X1 U12096 ( .A1(n18940), .A2(n15674), .ZN(n18717) );
  INV_X1 U12097 ( .A(n18228), .ZN(n18706) );
  INV_X1 U12098 ( .A(n18710), .ZN(n16614) );
  INV_X1 U12099 ( .A(n18225), .ZN(n18712) );
  INV_X1 U12100 ( .A(n18726), .ZN(n18745) );
  NOR2_X1 U12101 ( .A1(n15677), .A2(n9757), .ZN(n18729) );
  OR2_X1 U12102 ( .A1(n9758), .A2(n17502), .ZN(n9757) );
  AND2_X1 U12103 ( .A1(n11904), .A2(n13067), .ZN(n9758) );
  NOR2_X1 U12104 ( .A1(n15675), .A2(n18732), .ZN(n18735) );
  INV_X1 U12105 ( .A(n16445), .ZN(n18274) );
  INV_X1 U12106 ( .A(n15682), .ZN(n18281) );
  NOR2_X1 U12107 ( .A1(n11880), .A2(n11879), .ZN(n18293) );
  NOR2_X1 U12108 ( .A1(n11851), .A2(n11850), .ZN(n18300) );
  OAI22_X1 U12109 ( .A1(n16439), .A2(n18228), .B1(n18705), .B2(n18712), .ZN(
        n18765) );
  NAND2_X1 U12110 ( .A1(n12231), .A2(n12002), .ZN(n20739) );
  NAND2_X1 U12111 ( .A1(n12637), .A2(n12636), .ZN(n19890) );
  INV_X1 U12112 ( .A(n15943), .ZN(n19904) );
  INV_X1 U12113 ( .A(n19934), .ZN(n16011) );
  INV_X1 U12114 ( .A(n19926), .ZN(n19901) );
  NOR2_X1 U12115 ( .A1(n19890), .A2(n19922), .ZN(n19917) );
  AND2_X1 U12116 ( .A1(n19890), .A2(n19889), .ZN(n15982) );
  INV_X1 U12117 ( .A(n19914), .ZN(n19939) );
  INV_X1 U12118 ( .A(n16020), .ZN(n19956) );
  INV_X1 U12119 ( .A(n19954), .ZN(n19950) );
  OR2_X1 U12120 ( .A1(n12496), .A2(n19849), .ZN(n12499) );
  NAND2_X1 U12121 ( .A1(n13839), .A2(n12500), .ZN(n16020) );
  INV_X1 U12122 ( .A(n13890), .ZN(n13907) );
  INV_X1 U12123 ( .A(n13920), .ZN(n13059) );
  NAND2_X1 U12124 ( .A1(n12213), .A2(n12212), .ZN(n13917) );
  NAND2_X1 U12125 ( .A1(n12207), .A2(n12976), .ZN(n12213) );
  OR2_X1 U12126 ( .A1(n13906), .A2(n12215), .ZN(n13920) );
  CLKBUF_X1 U12127 ( .A(n19987), .Z(n20742) );
  INV_X1 U12128 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15971) );
  AND2_X1 U12129 ( .A1(n11153), .A2(n20510), .ZN(n20028) );
  INV_X1 U12130 ( .A(n20022), .ZN(n14062) );
  NOR2_X2 U12131 ( .A1(n20022), .A2(n12222), .ZN(n16064) );
  INV_X1 U12132 ( .A(n20028), .ZN(n20098) );
  AND2_X2 U12133 ( .A1(n16067), .A2(n11154), .ZN(n20022) );
  XNOR2_X1 U12134 ( .A(n10142), .B(n14075), .ZN(n14102) );
  NAND2_X1 U12135 ( .A1(n13930), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10143) );
  NAND2_X1 U12136 ( .A1(n9941), .A2(n9938), .ZN(n13939) );
  NAND2_X1 U12137 ( .A1(n9939), .A2(n14000), .ZN(n9938) );
  NAND2_X1 U12138 ( .A1(n9942), .A2(n9595), .ZN(n9941) );
  AND2_X1 U12139 ( .A1(n14183), .A2(n14072), .ZN(n14162) );
  AND2_X1 U12140 ( .A1(n14195), .A2(n14157), .ZN(n14209) );
  NAND2_X1 U12141 ( .A1(n20058), .A2(n20076), .ZN(n20056) );
  NAND2_X1 U12142 ( .A1(n10603), .A2(n10602), .ZN(n14059) );
  INV_X1 U12143 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20509) );
  NAND2_X1 U12144 ( .A1(n10402), .A2(n10452), .ZN(n13768) );
  INV_X1 U12145 ( .A(n10680), .ZN(n10682) );
  XNOR2_X1 U12146 ( .A(n10546), .B(n14273), .ZN(n20099) );
  INV_X1 U12147 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12170) );
  NOR2_X1 U12148 ( .A1(n20355), .A2(n12973), .ZN(n14285) );
  INV_X1 U12149 ( .A(n20647), .ZN(n20139) );
  OAI21_X1 U12150 ( .B1(n20256), .B2(n20240), .A(n20548), .ZN(n20259) );
  OR2_X1 U12151 ( .A1(n20262), .A2(n10688), .ZN(n20298) );
  INV_X1 U12152 ( .A(n20298), .ZN(n20312) );
  OAI211_X1 U12153 ( .C1(n20370), .C2(n20355), .A(n20408), .B(n20354), .ZN(
        n20373) );
  INV_X1 U12154 ( .A(n20434), .ZN(n20398) );
  INV_X1 U12155 ( .A(n20473), .ZN(n20462) );
  INV_X1 U12156 ( .A(n20475), .ZN(n20534) );
  INV_X1 U12157 ( .A(n20550), .ZN(n20643) );
  INV_X1 U12158 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20649) );
  INV_X1 U12159 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20355) );
  OR2_X1 U12160 ( .A1(n14364), .A2(n12796), .ZN(n19087) );
  AND2_X1 U12161 ( .A1(n10110), .A2(n9591), .ZN(n14440) );
  INV_X1 U12162 ( .A(n10110), .ZN(n15852) );
  AND2_X1 U12163 ( .A1(n12805), .A2(n12804), .ZN(n19104) );
  AND2_X1 U12164 ( .A1(n12795), .A2(n16420), .ZN(n19070) );
  OR2_X1 U12165 ( .A1(n12587), .A2(n12586), .ZN(n12705) );
  AND2_X1 U12166 ( .A1(n9869), .A2(n12351), .ZN(n9868) );
  OR2_X1 U12167 ( .A1(n12386), .A2(n12385), .ZN(n12694) );
  OR2_X1 U12168 ( .A1(n14659), .A2(n12103), .ZN(n14677) );
  AND2_X1 U12169 ( .A1(n14682), .A2(n14681), .ZN(n16215) );
  NAND2_X1 U12170 ( .A1(n10204), .A2(n10203), .ZN(n14607) );
  AND2_X1 U12171 ( .A1(n19144), .A2(n13437), .ZN(n16230) );
  AND2_X1 U12172 ( .A1(n14779), .A2(n14776), .ZN(n19135) );
  AND2_X1 U12173 ( .A1(n12031), .A2(n10187), .ZN(n12564) );
  INV_X1 U12174 ( .A(n10188), .ZN(n10187) );
  INV_X1 U12175 ( .A(n14776), .ZN(n19129) );
  NAND2_X1 U12176 ( .A1(n19144), .A2(n12103), .ZN(n14776) );
  NOR2_X1 U12178 ( .A1(n19180), .A2(n19190), .ZN(n19197) );
  CLKBUF_X1 U12179 ( .A(n19197), .Z(n19209) );
  AND2_X2 U12180 ( .A1(n18946), .A2(n16421), .ZN(n12795) );
  NAND2_X1 U12181 ( .A1(n15094), .A2(n10230), .ZN(n16247) );
  INV_X1 U12182 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16269) );
  INV_X1 U12183 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16285) );
  AND2_X1 U12184 ( .A1(n16305), .A2(n12095), .ZN(n16295) );
  INV_X1 U12185 ( .A(n16305), .ZN(n19215) );
  NAND2_X1 U12186 ( .A1(n15002), .A2(n15001), .ZN(n9987) );
  AOI21_X1 U12187 ( .B1(n15094), .B2(n9796), .A(n9615), .ZN(n15015) );
  NOR2_X1 U12188 ( .A1(n10072), .A2(n10071), .ZN(n15096) );
  INV_X1 U12189 ( .A(n9712), .ZN(n10071) );
  INV_X1 U12190 ( .A(n10073), .ZN(n10072) );
  INV_X1 U12191 ( .A(n9889), .ZN(n15404) );
  AOI21_X1 U12192 ( .B1(n16281), .B2(n14906), .A(n9771), .ZN(n9889) );
  NAND2_X1 U12193 ( .A1(n12764), .A2(n10088), .ZN(n15114) );
  INV_X1 U12194 ( .A(n12774), .ZN(n9888) );
  NAND2_X1 U12195 ( .A1(n9973), .A2(n10063), .ZN(n11653) );
  INV_X1 U12196 ( .A(n16369), .ZN(n16309) );
  INV_X1 U12197 ( .A(n16319), .ZN(n16371) );
  INV_X1 U12198 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19836) );
  OR2_X1 U12199 ( .A1(n12195), .A2(n12064), .ZN(n19831) );
  INV_X1 U12200 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19827) );
  INV_X1 U12201 ( .A(n19823), .ZN(n19820) );
  INV_X1 U12202 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19817) );
  INV_X1 U12203 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19809) );
  NAND2_X1 U12204 ( .A1(n12031), .A2(n11742), .ZN(n12531) );
  XNOR2_X1 U12205 ( .A(n12194), .B(n12193), .ZN(n19823) );
  XNOR2_X1 U12206 ( .A(n12293), .B(n12199), .ZN(n19812) );
  NOR2_X1 U12207 ( .A1(n19659), .A2(n19406), .ZN(n19426) );
  OAI21_X1 U12208 ( .B1(n19452), .B2(n19432), .A(n19655), .ZN(n19454) );
  NAND2_X1 U12209 ( .A1(n19437), .A2(n19436), .ZN(n19453) );
  NOR2_X2 U12210 ( .A1(n19598), .A2(n19469), .ZN(n19489) );
  NOR2_X1 U12211 ( .A1(n19470), .A2(n19469), .ZN(n19500) );
  OAI22_X1 U12212 ( .A1(n18265), .A2(n15563), .B1(n16529), .B2(n15564), .ZN(
        n19605) );
  OAI22_X1 U12213 ( .A1(n18273), .A2(n15563), .B1(n16527), .B2(n15564), .ZN(
        n19615) );
  OAI22_X1 U12214 ( .A1(n18280), .A2(n15563), .B1(n13868), .B2(n15564), .ZN(
        n19619) );
  OAI22_X1 U12215 ( .A1(n16524), .A2(n15564), .B1(n18285), .B2(n15563), .ZN(
        n19623) );
  OAI22_X1 U12216 ( .A1(n13859), .A2(n15564), .B1(n18292), .B2(n15563), .ZN(
        n19627) );
  OAI22_X1 U12217 ( .A1(n16521), .A2(n15564), .B1(n18298), .B2(n15563), .ZN(
        n19631) );
  OAI22_X1 U12218 ( .A1(n18307), .A2(n15563), .B1(n16519), .B2(n15564), .ZN(
        n19635) );
  INV_X1 U12219 ( .A(n19599), .ZN(n19642) );
  OAI22_X1 U12220 ( .A1(n16517), .A2(n15564), .B1(n18312), .B2(n15563), .ZN(
        n19641) );
  INV_X1 U12221 ( .A(n19605), .ZN(n19665) );
  INV_X1 U12222 ( .A(n19615), .ZN(n19671) );
  INV_X1 U12223 ( .A(n19233), .ZN(n19672) );
  INV_X1 U12224 ( .A(n19236), .ZN(n19678) );
  INV_X1 U12225 ( .A(n19623), .ZN(n19683) );
  INV_X1 U12226 ( .A(n19627), .ZN(n19689) );
  INV_X1 U12227 ( .A(n19242), .ZN(n19690) );
  INV_X1 U12228 ( .A(n19631), .ZN(n19695) );
  INV_X1 U12229 ( .A(n19635), .ZN(n19701) );
  INV_X1 U12230 ( .A(n19245), .ZN(n19703) );
  INV_X1 U12231 ( .A(n19646), .ZN(n19704) );
  INV_X1 U12232 ( .A(n19641), .ZN(n19712) );
  NOR3_X1 U12233 ( .A1(n16426), .A2(n16425), .A3(n16424), .ZN(n19719) );
  NOR2_X1 U12234 ( .A1(n17502), .A2(n13079), .ZN(n16616) );
  NOR2_X1 U12235 ( .A1(n16697), .A2(n17600), .ZN(n16696) );
  NOR2_X1 U12236 ( .A1(n16707), .A2(n9694), .ZN(n16697) );
  NOR2_X1 U12237 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16764), .ZN(n16751) );
  NOR2_X1 U12238 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16840), .ZN(n16817) );
  INV_X1 U12239 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16844) );
  NOR2_X1 U12240 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16872), .ZN(n16871) );
  INV_X1 U12241 ( .A(n16963), .ZN(n16987) );
  NOR2_X2 U12242 ( .A1(n18872), .A2(n16969), .ZN(n16963) );
  NAND4_X1 U12243 ( .A1(n18181), .A2(n16947), .A3(n18781), .A4(n18772), .ZN(
        n16999) );
  INV_X1 U12244 ( .A(n16976), .ZN(n16996) );
  INV_X1 U12245 ( .A(n18316), .ZN(n17424) );
  NOR2_X1 U12246 ( .A1(n17330), .A2(n17527), .ZN(n17325) );
  NOR2_X1 U12247 ( .A1(n17523), .A2(n17340), .ZN(n17335) );
  NAND2_X1 U12248 ( .A1(n17341), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17340) );
  AND2_X1 U12249 ( .A1(n17347), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17341) );
  NOR2_X1 U12250 ( .A1(n17350), .A2(n17424), .ZN(n17347) );
  NOR2_X1 U12251 ( .A1(n17389), .A2(n9755), .ZN(n17351) );
  NAND2_X1 U12252 ( .A1(n9720), .A2(n9756), .ZN(n9755) );
  INV_X1 U12253 ( .A(n17355), .ZN(n9756) );
  NOR3_X1 U12254 ( .A1(n17424), .A2(n17389), .A3(n17506), .ZN(n17378) );
  NAND2_X1 U12255 ( .A1(n9652), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17389) );
  NOR2_X1 U12256 ( .A1(n15707), .A2(n15706), .ZN(n17433) );
  NAND2_X1 U12257 ( .A1(n18744), .A2(n15915), .ZN(n17451) );
  INV_X1 U12258 ( .A(n17457), .ZN(n17454) );
  NOR2_X1 U12259 ( .A1(n15747), .A2(n9850), .ZN(n9849) );
  NOR2_X1 U12260 ( .A1(n18744), .A2(n17449), .ZN(n17457) );
  INV_X1 U12261 ( .A(n17451), .ZN(n17456) );
  NOR2_X1 U12262 ( .A1(n18920), .A2(n17463), .ZN(n17489) );
  CLKBUF_X1 U12263 ( .A(n17489), .Z(n17496) );
  CLKBUF_X1 U12264 ( .A(n17565), .Z(n17561) );
  BUF_X1 U12265 ( .A(n17556), .Z(n17564) );
  NOR2_X1 U12266 ( .A1(n18274), .A2(n17564), .ZN(n17565) );
  AOI21_X1 U12267 ( .B1(n9965), .B2(n9961), .A(n9963), .ZN(n9960) );
  AND2_X1 U12268 ( .A1(n9966), .A2(n9969), .ZN(n9961) );
  NOR2_X1 U12269 ( .A1(n9968), .A2(n17824), .ZN(n9963) );
  NAND2_X1 U12270 ( .A1(n16454), .A2(n9964), .ZN(n9962) );
  NOR2_X1 U12271 ( .A1(n9968), .A2(n16453), .ZN(n9964) );
  NAND3_X1 U12272 ( .A1(n10056), .A2(n10055), .A3(n10057), .ZN(n16986) );
  NAND2_X1 U12273 ( .A1(n10059), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10057) );
  OAI22_X1 U12274 ( .A1(n17751), .A2(n18119), .B1(n17937), .B2(n18121), .ZN(
        n17787) );
  NAND2_X1 U12275 ( .A1(n16505), .A2(n17920), .ZN(n17844) );
  NOR2_X1 U12276 ( .A1(n17847), .A2(n17835), .ZN(n17831) );
  INV_X1 U12277 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17835) );
  NOR2_X1 U12278 ( .A1(n16505), .A2(n17935), .ZN(n17841) );
  NOR2_X1 U12279 ( .A1(n17874), .A2(n17875), .ZN(n17876) );
  INV_X1 U12280 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17902) );
  INV_X1 U12281 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17918) );
  INV_X2 U12282 ( .A(n18653), .ZN(n18395) );
  INV_X1 U12283 ( .A(n17935), .ZN(n17920) );
  OAI21_X1 U12284 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18922), .A(n16617), 
        .ZN(n17931) );
  INV_X1 U12285 ( .A(n17924), .ZN(n17937) );
  AOI22_X1 U12286 ( .A1(n9966), .A2(n9965), .B1(n16454), .B2(n9967), .ZN(
        n16495) );
  NAND2_X1 U12287 ( .A1(n10179), .A2(n9846), .ZN(n15897) );
  NAND2_X1 U12288 ( .A1(n17683), .A2(n10183), .ZN(n17635) );
  INV_X1 U12289 ( .A(n17623), .ZN(n17634) );
  AND2_X1 U12290 ( .A1(n9701), .A2(n15839), .ZN(n17726) );
  NAND2_X1 U12291 ( .A1(n18738), .A2(n18745), .ZN(n18126) );
  INV_X1 U12292 ( .A(n9588), .ZN(n18743) );
  NAND2_X1 U12293 ( .A1(n17817), .A2(n10174), .ZN(n17819) );
  INV_X1 U12294 ( .A(n18169), .ZN(n18150) );
  NOR2_X1 U12295 ( .A1(n17747), .A2(n9673), .ZN(n18165) );
  INV_X1 U12296 ( .A(n18251), .ZN(n18236) );
  INV_X1 U12297 ( .A(n10175), .ZN(n17896) );
  NOR2_X1 U12298 ( .A1(n15815), .A2(n15814), .ZN(n18225) );
  INV_X1 U12299 ( .A(n9951), .ZN(n17909) );
  INV_X1 U12300 ( .A(n18248), .ZN(n18231) );
  NOR2_X1 U12301 ( .A1(n18712), .A2(n18248), .ZN(n18247) );
  INV_X1 U12302 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18759) );
  INV_X1 U12303 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18872) );
  NAND2_X1 U12304 ( .A1(n18799), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18936) );
  CLKBUF_X1 U12305 ( .A(n16593), .Z(n20772) );
  OAI211_X1 U12306 ( .C1(n14108), .C2(n20085), .A(n10028), .B(n10027), .ZN(
        P1_U3001) );
  AOI21_X1 U12307 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(n10028) );
  OR2_X1 U12308 ( .A1(n14104), .A2(n20083), .ZN(n10027) );
  AND2_X1 U12309 ( .A1(n9906), .A2(n14114), .ZN(n9905) );
  OR2_X1 U12310 ( .A1(n14116), .A2(n14115), .ZN(n9906) );
  NAND2_X1 U12311 ( .A1(n9932), .A2(n14922), .ZN(P2_U2983) );
  NOR2_X1 U12312 ( .A1(n15150), .A2(n16287), .ZN(n14929) );
  OAI21_X1 U12313 ( .B1(n16238), .B2(n16287), .A(n9894), .ZN(P2_U3000) );
  AOI21_X1 U12314 ( .B1(n19045), .B2(n19227), .A(n9896), .ZN(n9895) );
  OR2_X1 U12315 ( .A1(n16239), .A2(n19218), .ZN(n9897) );
  NAND2_X1 U12316 ( .A1(n9780), .A2(n9778), .ZN(P2_U3029) );
  NOR2_X1 U12317 ( .A1(n15363), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9781) );
  INV_X1 U12318 ( .A(n9782), .ZN(n15342) );
  OAI21_X1 U12319 ( .B1(n16656), .B2(n9711), .A(n10049), .ZN(P3_U2640) );
  AOI21_X1 U12320 ( .B1(n16661), .B2(n17034), .A(n10050), .ZN(n10049) );
  NAND2_X1 U12321 ( .A1(n10054), .A2(n10051), .ZN(n10050) );
  NAND2_X1 U12322 ( .A1(n17319), .A2(n9713), .ZN(n17311) );
  NAND2_X1 U12323 ( .A1(n14635), .A2(n9690), .ZN(n14618) );
  INV_X1 U12324 ( .A(n12787), .ZN(n10128) );
  AND2_X1 U12325 ( .A1(n9620), .A2(n14665), .ZN(n9611) );
  AND2_X1 U12326 ( .A1(n9723), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9612) );
  AND2_X1 U12327 ( .A1(n9600), .A2(n11392), .ZN(n11402) );
  CLKBUF_X3 U12328 ( .A(n15648), .Z(n17263) );
  NAND2_X1 U12329 ( .A1(n16069), .A2(n10605), .ZN(n14027) );
  INV_X1 U12330 ( .A(n11297), .ZN(n12046) );
  INV_X1 U12331 ( .A(n9785), .ZN(n15405) );
  NAND2_X1 U12332 ( .A1(n12941), .A2(n10156), .ZN(n13041) );
  NAND2_X1 U12333 ( .A1(n14635), .A2(n10220), .ZN(n14626) );
  NAND2_X1 U12334 ( .A1(n14873), .A2(n14872), .ZN(n9613) );
  NAND2_X1 U12335 ( .A1(n13707), .A2(n9692), .ZN(n9614) );
  OR2_X1 U12336 ( .A1(n14867), .A2(n15021), .ZN(n9615) );
  AND2_X1 U12337 ( .A1(n16421), .A2(n9664), .ZN(n9616) );
  INV_X1 U12338 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14541) );
  AND2_X1 U12339 ( .A1(n10118), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9617) );
  AND2_X1 U12340 ( .A1(n10042), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9618) );
  NAND2_X1 U12341 ( .A1(n10081), .A2(n10080), .ZN(n9619) );
  AND2_X1 U12342 ( .A1(n10090), .A2(n12923), .ZN(n9620) );
  INV_X2 U12343 ( .A(n14000), .ZN(n16055) );
  NAND2_X1 U12344 ( .A1(n15448), .A2(n12120), .ZN(n11373) );
  INV_X1 U12345 ( .A(n11373), .ZN(n9741) );
  OR2_X1 U12346 ( .A1(n14034), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9621) );
  AND2_X1 U12347 ( .A1(n12173), .A2(n10345), .ZN(n9622) );
  AND2_X1 U12348 ( .A1(n12563), .A2(n12561), .ZN(n9623) );
  AND2_X1 U12349 ( .A1(n9862), .A2(n9865), .ZN(n9624) );
  AND2_X1 U12350 ( .A1(n10013), .A2(n10012), .ZN(n9625) );
  AND2_X1 U12351 ( .A1(n10017), .A2(n10015), .ZN(n9626) );
  AND2_X1 U12352 ( .A1(n10136), .A2(n10140), .ZN(n9627) );
  AND2_X1 U12353 ( .A1(n9623), .A2(n9708), .ZN(n9628) );
  INV_X1 U12354 ( .A(n11739), .ZN(n12888) );
  INV_X1 U12355 ( .A(n12888), .ZN(n13471) );
  NAND2_X1 U12356 ( .A1(n10217), .A2(n12569), .ZN(n12489) );
  NAND2_X1 U12357 ( .A1(n10217), .A2(n9869), .ZN(n12672) );
  AND4_X1 U12358 ( .A1(n10128), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9629) );
  AND2_X1 U12359 ( .A1(n10114), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9630) );
  AND2_X1 U12360 ( .A1(n10124), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9631) );
  INV_X1 U12361 ( .A(n14543), .ZN(n9789) );
  AND2_X1 U12362 ( .A1(n15095), .A2(n9712), .ZN(n9632) );
  OR2_X1 U12363 ( .A1(n12275), .A2(n12274), .ZN(n9633) );
  OR2_X1 U12364 ( .A1(n14000), .A2(n14115), .ZN(n9634) );
  AND2_X1 U12365 ( .A1(n13455), .A2(n13451), .ZN(n9635) );
  NAND2_X1 U12366 ( .A1(n11311), .A2(n11604), .ZN(n9636) );
  AND2_X1 U12367 ( .A1(n13425), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12599) );
  INV_X1 U12368 ( .A(n13289), .ZN(n9875) );
  OR2_X1 U12369 ( .A1(n17818), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9637) );
  AND2_X1 U12370 ( .A1(n15124), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9638) );
  AND2_X1 U12371 ( .A1(n9638), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9639) );
  AND2_X1 U12372 ( .A1(n15145), .A2(n15125), .ZN(n9640) );
  AND2_X1 U12373 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9641) );
  INV_X4 U12374 ( .A(n15605), .ZN(n15780) );
  OR3_X1 U12375 ( .A1(n13716), .A2(n10021), .A3(n10023), .ZN(n9643) );
  XNOR2_X1 U12376 ( .A(n14905), .B(n14903), .ZN(n11685) );
  OR2_X1 U12377 ( .A1(n14621), .A2(n10092), .ZN(n9644) );
  NAND3_X2 U12378 ( .A1(n10171), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13429) );
  OR2_X1 U12379 ( .A1(n13343), .A2(n13342), .ZN(n9645) );
  OR2_X1 U12380 ( .A1(n14456), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n9646) );
  OR4_X1 U12381 ( .A1(n15020), .A2(n15037), .A3(n15077), .A4(n14851), .ZN(
        n9647) );
  NOR2_X1 U12382 ( .A1(n13809), .A2(n10153), .ZN(n13800) );
  NOR2_X1 U12383 ( .A1(n13823), .A2(n13824), .ZN(n13816) );
  AND2_X1 U12384 ( .A1(n13452), .A2(n9635), .ZN(n9648) );
  OR2_X1 U12385 ( .A1(n15820), .A2(n18187), .ZN(n9649) );
  OR2_X1 U12386 ( .A1(n10001), .A2(n14899), .ZN(n9650) );
  NAND2_X1 U12387 ( .A1(n16253), .A2(n16254), .ZN(n10073) );
  NOR2_X1 U12388 ( .A1(n14882), .A2(n15182), .ZN(n9651) );
  NOR2_X1 U12389 ( .A1(n17398), .A2(n17568), .ZN(n9652) );
  OR3_X1 U12390 ( .A1(n14388), .A2(n10107), .A3(n10104), .ZN(n9653) );
  AND2_X1 U12391 ( .A1(n14784), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9654) );
  OR2_X1 U12392 ( .A1(n16055), .A2(n10604), .ZN(n9655) );
  AND2_X1 U12393 ( .A1(n16033), .A2(n16040), .ZN(n9656) );
  AND2_X1 U12394 ( .A1(n11233), .A2(n11307), .ZN(n9657) );
  AND2_X1 U12395 ( .A1(n10279), .A2(n10278), .ZN(n9658) );
  XNOR2_X1 U12396 ( .A(n14784), .B(n9772), .ZN(n14782) );
  NAND2_X1 U12397 ( .A1(n9799), .A2(n14803), .ZN(n16253) );
  NAND2_X1 U12398 ( .A1(n10075), .A2(n14791), .ZN(n15393) );
  AND2_X1 U12399 ( .A1(n12928), .A2(n12942), .ZN(n12941) );
  AND2_X1 U12400 ( .A1(n14021), .A2(n10605), .ZN(n9659) );
  OR2_X1 U12401 ( .A1(n11369), .A2(n11368), .ZN(n11478) );
  NAND2_X1 U12402 ( .A1(n13968), .A2(n13990), .ZN(n13985) );
  NAND2_X1 U12403 ( .A1(n10003), .A2(n10006), .ZN(n15094) );
  NOR3_X1 U12404 ( .A1(n16194), .A2(n11643), .A3(n15125), .ZN(n9660) );
  AND2_X1 U12405 ( .A1(n13707), .A2(n10158), .ZN(n11151) );
  OR3_X1 U12406 ( .A1(n14621), .A2(n10093), .A3(n10095), .ZN(n9661) );
  AND2_X1 U12407 ( .A1(n14587), .A2(n10213), .ZN(n14592) );
  OR2_X1 U12408 ( .A1(n14948), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9662) );
  AND2_X1 U12409 ( .A1(n11742), .A2(n9628), .ZN(n9663) );
  NAND2_X1 U12410 ( .A1(n12289), .A2(n12288), .ZN(n12465) );
  AND2_X1 U12411 ( .A1(n9603), .A2(n12070), .ZN(n9664) );
  OR2_X1 U12412 ( .A1(n13716), .A2(n13696), .ZN(n9665) );
  OAI21_X1 U12413 ( .B1(n9619), .B2(n15355), .A(n10077), .ZN(n9814) );
  INV_X1 U12414 ( .A(n9990), .ZN(n9989) );
  OAI21_X1 U12415 ( .B1(n9991), .B2(n15001), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U12416 ( .A1(n14428), .A2(n14406), .ZN(n14396) );
  AND2_X1 U12417 ( .A1(n14899), .A2(n9999), .ZN(n9666) );
  NAND2_X1 U12418 ( .A1(n12200), .A2(n12299), .ZN(n11369) );
  INV_X1 U12419 ( .A(n11369), .ZN(n9742) );
  AND2_X1 U12420 ( .A1(n9655), .A2(n10602), .ZN(n9667) );
  AND2_X1 U12421 ( .A1(n10561), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9668) );
  AND2_X1 U12422 ( .A1(n16083), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9669) );
  AND2_X1 U12423 ( .A1(n14828), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9670) );
  NAND2_X2 U12424 ( .A1(n11208), .A2(n11207), .ZN(n15537) );
  INV_X1 U12425 ( .A(n15537), .ZN(n9887) );
  NAND2_X1 U12426 ( .A1(n13816), .A2(n13817), .ZN(n13809) );
  AND3_X1 U12427 ( .A1(n11387), .A2(n11386), .A3(n11385), .ZN(n9671) );
  AND2_X1 U12428 ( .A1(n10452), .A2(n10131), .ZN(n9672) );
  NAND2_X1 U12429 ( .A1(n13707), .A2(n10160), .ZN(n13684) );
  NAND2_X1 U12430 ( .A1(n13792), .A2(n9761), .ZN(n13737) );
  NAND2_X1 U12431 ( .A1(n13707), .A2(n13708), .ZN(n13693) );
  NAND2_X1 U12432 ( .A1(n10085), .A2(n10083), .ZN(n10086) );
  NAND2_X1 U12433 ( .A1(n13792), .A2(n13793), .ZN(n13736) );
  AND2_X1 U12434 ( .A1(n15831), .A2(n18161), .ZN(n9673) );
  NAND2_X1 U12435 ( .A1(n12941), .A2(n13011), .ZN(n13010) );
  AND2_X1 U12436 ( .A1(n9926), .A2(n14785), .ZN(n9674) );
  NOR2_X1 U12437 ( .A1(n16299), .A2(n14903), .ZN(n9675) );
  INV_X1 U12438 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17875) );
  AND3_X1 U12439 ( .A1(n15732), .A2(n15735), .A3(n15733), .ZN(n9676) );
  OR2_X1 U12440 ( .A1(n9813), .A2(n9814), .ZN(n9677) );
  NAND2_X1 U12441 ( .A1(n10152), .A2(n10918), .ZN(n13801) );
  OR2_X1 U12442 ( .A1(n18234), .A2(n15818), .ZN(n9678) );
  AND2_X1 U12443 ( .A1(n11546), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9679) );
  OR2_X1 U12444 ( .A1(n17178), .A2(n18284), .ZN(n9680) );
  NOR2_X1 U12445 ( .A1(n9660), .A2(n10002), .ZN(n10001) );
  AND2_X1 U12446 ( .A1(n14878), .A2(n14877), .ZN(n9681) );
  AND2_X1 U12447 ( .A1(n9649), .A2(n18206), .ZN(n9682) );
  INV_X1 U12448 ( .A(n9969), .ZN(n9968) );
  NAND2_X1 U12449 ( .A1(n16494), .A2(n9589), .ZN(n9969) );
  INV_X1 U12450 ( .A(n11336), .ZN(n9808) );
  NAND2_X1 U12451 ( .A1(n11328), .A2(n11327), .ZN(n11336) );
  AND2_X1 U12452 ( .A1(n9954), .A2(n9953), .ZN(n9683) );
  INV_X1 U12453 ( .A(n10139), .ZN(n10138) );
  NAND2_X1 U12454 ( .A1(n10428), .A2(n10141), .ZN(n10139) );
  NOR2_X2 U12455 ( .A1(n20137), .A2(n20132), .ZN(n9684) );
  NAND2_X1 U12456 ( .A1(n20120), .A2(n12978), .ZN(n12658) );
  INV_X1 U12457 ( .A(n9592), .ZN(n12200) );
  NAND2_X1 U12458 ( .A1(n12704), .A2(n12703), .ZN(n12909) );
  AND2_X1 U12459 ( .A1(n10217), .A2(n10216), .ZN(n12546) );
  INV_X1 U12460 ( .A(n12190), .ZN(n9865) );
  NOR2_X1 U12461 ( .A1(n14643), .A2(n14645), .ZN(n14635) );
  AND2_X1 U12462 ( .A1(n14635), .A2(n14637), .ZN(n14631) );
  AND2_X1 U12463 ( .A1(n12928), .A2(n9770), .ZN(n13042) );
  NOR2_X1 U12464 ( .A1(n12332), .A2(n12331), .ZN(n9685) );
  AND2_X1 U12465 ( .A1(n14330), .A2(n10118), .ZN(n9686) );
  AND2_X1 U12466 ( .A1(n14335), .A2(n10124), .ZN(n9687) );
  NAND2_X1 U12467 ( .A1(n12846), .A2(n12845), .ZN(n12844) );
  INV_X1 U12468 ( .A(n12557), .ZN(n10715) );
  NOR2_X1 U12469 ( .A1(n14493), .A2(n14494), .ZN(n9688) );
  OR3_X1 U12470 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17662), .ZN(n9689) );
  INV_X1 U12471 ( .A(n15012), .ZN(n9795) );
  AND2_X1 U12472 ( .A1(n10220), .A2(n13204), .ZN(n9690) );
  AND2_X1 U12473 ( .A1(n10216), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9691) );
  NOR2_X1 U12474 ( .A1(n9694), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U12475 ( .A1(n16087), .A2(n10574), .ZN(n16082) );
  AOI21_X1 U12476 ( .B1(n10732), .B2(n10855), .A(n10731), .ZN(n12714) );
  INV_X1 U12477 ( .A(n12714), .ZN(n9768) );
  AND2_X1 U12478 ( .A1(n10160), .A2(n10159), .ZN(n9692) );
  AND2_X1 U12479 ( .A1(n10205), .A2(n10209), .ZN(n14606) );
  NAND2_X1 U12480 ( .A1(n20132), .A2(n13848), .ZN(n12214) );
  INV_X2 U12481 ( .A(n13978), .ZN(n14000) );
  AND2_X1 U12482 ( .A1(n10195), .A2(n14429), .ZN(n9693) );
  INV_X1 U12483 ( .A(n10628), .ZN(n10137) );
  INV_X1 U12484 ( .A(n13978), .ZN(n14034) );
  AND2_X1 U12486 ( .A1(n14831), .A2(n14830), .ZN(n15068) );
  INV_X1 U12487 ( .A(n15068), .ZN(n10080) );
  NAND2_X1 U12488 ( .A1(n11682), .A2(n9927), .ZN(n9930) );
  NAND2_X1 U12489 ( .A1(n10354), .A2(n10353), .ZN(n12144) );
  AND3_X1 U12490 ( .A1(n12846), .A2(n12845), .A3(n10164), .ZN(n12928) );
  OR2_X1 U12491 ( .A1(n10068), .A2(n15022), .ZN(n9695) );
  INV_X1 U12492 ( .A(n9867), .ZN(n9866) );
  OR2_X1 U12493 ( .A1(n12192), .A2(n9865), .ZN(n9867) );
  AND2_X1 U12494 ( .A1(n14492), .A2(n9620), .ZN(n9696) );
  AND2_X1 U12495 ( .A1(n9761), .A2(n9760), .ZN(n9697) );
  NAND2_X1 U12496 ( .A1(n14340), .A2(n10114), .ZN(n10116) );
  OR2_X1 U12497 ( .A1(n17829), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9698) );
  OR2_X1 U12498 ( .A1(n10038), .A2(n10039), .ZN(n9699) );
  NAND2_X1 U12499 ( .A1(n14770), .A2(n14768), .ZN(n9700) );
  AND2_X1 U12500 ( .A1(n15837), .A2(n15836), .ZN(n9701) );
  AND2_X1 U12501 ( .A1(n9625), .A2(n13833), .ZN(n9702) );
  INV_X1 U12502 ( .A(n9613), .ZN(n9991) );
  AND2_X1 U12503 ( .A1(n10156), .A2(n10155), .ZN(n9703) );
  AND2_X1 U12504 ( .A1(n9611), .A2(n10091), .ZN(n9704) );
  INV_X1 U12505 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16306) );
  INV_X1 U12506 ( .A(n9979), .ZN(n9978) );
  NAND2_X1 U12507 ( .A1(n14532), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9979) );
  AND2_X1 U12508 ( .A1(n16482), .A2(n10060), .ZN(n9705) );
  NAND2_X1 U12509 ( .A1(n12704), .A2(n10219), .ZN(n13103) );
  NOR2_X2 U12510 ( .A1(n12208), .A2(n10675), .ZN(n10855) );
  INV_X1 U12511 ( .A(n10855), .ZN(n9765) );
  NOR2_X2 U12512 ( .A1(n16503), .A2(n17430), .ZN(n17818) );
  INV_X1 U12513 ( .A(n17818), .ZN(n17829) );
  AND2_X1 U12514 ( .A1(n14251), .A2(n9625), .ZN(n9706) );
  INV_X1 U12515 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10043) );
  AOI21_X1 U12516 ( .B1(n14474), .B2(n15042), .A(n19094), .ZN(n14473) );
  OR2_X1 U12517 ( .A1(n9590), .A2(n14345), .ZN(n9707) );
  INV_X1 U12518 ( .A(n14519), .ZN(n9929) );
  NAND4_X1 U12519 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n9708) );
  OR3_X1 U12520 ( .A1(n13289), .A2(n13288), .A3(n14610), .ZN(n9709) );
  AND2_X1 U12521 ( .A1(n10185), .A2(n12031), .ZN(n12559) );
  OR2_X1 U12522 ( .A1(n19931), .A2(n12664), .ZN(n19932) );
  INV_X1 U12523 ( .A(n19932), .ZN(n10016) );
  AND2_X1 U12524 ( .A1(n10217), .A2(n9691), .ZN(n9710) );
  OR2_X1 U12525 ( .A1(n16818), .A2(n16657), .ZN(n9711) );
  INV_X1 U12526 ( .A(n16453), .ZN(n9967) );
  OR2_X1 U12527 ( .A1(n19065), .A2(n14809), .ZN(n9712) );
  OR2_X1 U12528 ( .A1(n17358), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9713) );
  INV_X1 U12529 ( .A(n10189), .ZN(n12390) );
  OR2_X1 U12530 ( .A1(n12332), .A2(n10192), .ZN(n10189) );
  OR2_X1 U12531 ( .A1(n14323), .A2(n10121), .ZN(n9714) );
  INV_X1 U12532 ( .A(n10059), .ZN(n10058) );
  NAND2_X1 U12533 ( .A1(n10060), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10059) );
  AND2_X1 U12534 ( .A1(n13383), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12604) );
  AND2_X1 U12535 ( .A1(n9846), .A2(n15848), .ZN(n9715) );
  AND2_X1 U12536 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9716) );
  AND2_X1 U12537 ( .A1(n14458), .A2(n10112), .ZN(n9717) );
  OR2_X1 U12538 ( .A1(n12079), .A2(n16421), .ZN(n19218) );
  OR3_X1 U12539 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9718) );
  AND4_X1 U12540 ( .A1(n15835), .A2(n18113), .A3(n17774), .A4(n18082), .ZN(
        n9719) );
  INV_X1 U12541 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10122) );
  AND4_X1 U12542 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9720)
         );
  AND2_X1 U12543 ( .A1(n17758), .A2(n10042), .ZN(n9721) );
  NOR2_X1 U12544 ( .A1(n15123), .A2(n15182), .ZN(n10168) );
  AND2_X1 U12545 ( .A1(n14182), .A2(n14008), .ZN(n9722) );
  AND2_X1 U12546 ( .A1(n16435), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12284) );
  INV_X1 U12547 ( .A(n12284), .ZN(n9864) );
  AND2_X1 U12548 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9723) );
  INV_X1 U12549 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n9922) );
  AND2_X1 U12550 ( .A1(n10047), .A2(n10045), .ZN(n9724) );
  INV_X1 U12551 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9772) );
  INV_X1 U12552 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10061) );
  INV_X1 U12553 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10178) );
  INV_X1 U12554 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10120) );
  AND2_X1 U12555 ( .A1(n10168), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9725) );
  INV_X1 U12556 ( .A(n16373), .ZN(n16360) );
  NOR2_X1 U12557 ( .A1(n15329), .A2(n16373), .ZN(n9779) );
  AOI22_X2 U12558 ( .A1(DATAI_23_), .A2(n20096), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20138), .ZN(n20648) );
  CLKBUF_X1 U12559 ( .A(n20609), .Z(n9726) );
  NAND2_X1 U12560 ( .A1(n9679), .A2(n11545), .ZN(n9734) );
  AND2_X4 U12561 ( .A1(n9729), .A2(n9727), .ZN(n15032) );
  INV_X1 U12562 ( .A(n9731), .ZN(n9730) );
  NAND4_X1 U12563 ( .A1(n14908), .A2(n9734), .A3(n14913), .A4(n14901), .ZN(
        n9731) );
  NAND2_X1 U12564 ( .A1(n9733), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9732) );
  NAND4_X2 U12565 ( .A1(n9740), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(n11326) );
  NAND3_X1 U12566 ( .A1(n9739), .A2(n11308), .A3(n11309), .ZN(n9735) );
  NAND2_X1 U12567 ( .A1(n11703), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9737) );
  NAND3_X1 U12568 ( .A1(n11305), .A2(n11306), .A3(n11307), .ZN(n9739) );
  INV_X1 U12569 ( .A(n9743), .ZN(n15385) );
  NOR2_X1 U12570 ( .A1(n9743), .A2(n15374), .ZN(n16256) );
  NOR2_X1 U12571 ( .A1(n9743), .A2(n9893), .ZN(n16242) );
  NAND3_X1 U12572 ( .A1(n10067), .A2(n10065), .A3(n9788), .ZN(n11508) );
  NAND3_X1 U12573 ( .A1(n9800), .A2(n9747), .A3(n9745), .ZN(n11772) );
  NOR2_X2 U12574 ( .A1(n14438), .A2(n14437), .ZN(n14873) );
  NAND2_X1 U12575 ( .A1(n11654), .A2(n11657), .ZN(n11656) );
  OAI21_X2 U12576 ( .B1(n14971), .B2(n9749), .A(n14888), .ZN(n14934) );
  NAND2_X1 U12577 ( .A1(n9983), .A2(n9751), .ZN(n14982) );
  NAND3_X1 U12578 ( .A1(n11870), .A2(n11869), .A3(n9753), .ZN(n9752) );
  NAND4_X1 U12579 ( .A1(n17423), .A2(n17310), .A3(P3_EAX_REG_13__SCAN_IN), 
        .A4(P3_EAX_REG_14__SCAN_IN), .ZN(n17398) );
  INV_X1 U12580 ( .A(n17341), .ZN(n17346) );
  INV_X2 U12581 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18905) );
  NAND2_X2 U12582 ( .A1(n10382), .A2(n10381), .ZN(n9759) );
  OR2_X1 U12583 ( .A1(n9759), .A2(n20478), .ZN(n12440) );
  XNOR2_X1 U12584 ( .A(n9759), .B(n20234), .ZN(n20103) );
  XNOR2_X2 U12585 ( .A(n10461), .B(n10538), .ZN(n12454) );
  NAND2_X2 U12586 ( .A1(n13707), .A2(n9766), .ZN(n13628) );
  AND2_X1 U12588 ( .A1(n9769), .A2(n12657), .ZN(n19918) );
  XNOR2_X1 U12589 ( .A(n9769), .B(n9768), .ZN(n19951) );
  NAND2_X1 U12590 ( .A1(n13042), .A2(n10861), .ZN(n13823) );
  NOR2_X4 U12591 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14287) );
  AND2_X2 U12592 ( .A1(n10244), .A2(n14287), .ZN(n10331) );
  OR2_X2 U12593 ( .A1(n11377), .A2(n11376), .ZN(n19258) );
  XNOR2_X2 U12594 ( .A(n11772), .B(n11773), .ZN(n12299) );
  INV_X1 U12595 ( .A(n14908), .ZN(n9771) );
  NAND3_X1 U12596 ( .A1(n11345), .A2(n11336), .A3(n11352), .ZN(n9802) );
  XNOR2_X2 U12597 ( .A(n9880), .B(n10202), .ZN(n11345) );
  NAND3_X2 U12598 ( .A1(n10063), .A2(n9973), .A3(n9888), .ZN(n12780) );
  NAND2_X2 U12599 ( .A1(n12780), .A2(n11460), .ZN(n11475) );
  INV_X1 U12600 ( .A(n15032), .ZN(n15386) );
  AND2_X1 U12601 ( .A1(n15032), .A2(n15318), .ZN(n15362) );
  INV_X4 U12602 ( .A(n13242), .ZN(n13421) );
  NAND2_X1 U12603 ( .A1(n9902), .A2(n14273), .ZN(n10563) );
  NAND2_X1 U12604 ( .A1(n11218), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11219) );
  AOI211_X2 U12605 ( .C1(n15191), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15190), .B(n15189), .ZN(n15192) );
  OR2_X2 U12606 ( .A1(n14022), .A2(n10146), .ZN(n10613) );
  NOR2_X2 U12607 ( .A1(n11377), .A2(n11373), .ZN(n15503) );
  INV_X1 U12608 ( .A(n10538), .ZN(n9911) );
  INV_X1 U12609 ( .A(n10546), .ZN(n9902) );
  NAND2_X1 U12610 ( .A1(n9934), .A2(n9935), .ZN(n12990) );
  NAND2_X1 U12611 ( .A1(n13956), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13958) );
  NAND2_X1 U12612 ( .A1(n9915), .A2(n10428), .ZN(n10523) );
  NAND2_X1 U12613 ( .A1(n9836), .A2(n10144), .ZN(n14022) );
  NAND2_X1 U12614 ( .A1(n9830), .A2(n9828), .ZN(n16089) );
  NAND2_X1 U12615 ( .A1(n10067), .A2(n11451), .ZN(n10066) );
  NAND2_X1 U12616 ( .A1(n11265), .A2(n11293), .ZN(n11276) );
  NAND2_X1 U12617 ( .A1(n11243), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9883) );
  NAND3_X1 U12618 ( .A1(n10065), .A2(n10067), .A3(n10062), .ZN(n9973) );
  NAND3_X1 U12619 ( .A1(n10065), .A2(n10067), .A3(n9786), .ZN(n9817) );
  NAND2_X1 U12620 ( .A1(n9973), .A2(n11668), .ZN(n11473) );
  NAND2_X2 U12621 ( .A1(n9983), .A2(n9790), .ZN(n14971) );
  NAND2_X1 U12622 ( .A1(n16296), .A2(n16297), .ZN(n9798) );
  NAND2_X1 U12623 ( .A1(n11344), .A2(n11325), .ZN(n11335) );
  NAND3_X1 U12624 ( .A1(n9802), .A2(n9804), .A3(n9806), .ZN(n9881) );
  NAND2_X2 U12625 ( .A1(n9811), .A2(n9809), .ZN(n11279) );
  NAND4_X1 U12626 ( .A1(n11270), .A2(n11272), .A3(n11271), .A4(n11273), .ZN(
        n9810) );
  NAND4_X1 U12627 ( .A1(n11266), .A2(n11267), .A3(n11269), .A4(n11268), .ZN(
        n9812) );
  NOR3_X1 U12628 ( .A1(n9813), .A2(n15059), .A3(n9814), .ZN(n15048) );
  NAND4_X1 U12629 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9820), .ZN(n9826)
         );
  INV_X1 U12630 ( .A(n10357), .ZN(n9822) );
  INV_X1 U12631 ( .A(n10367), .ZN(n9823) );
  NAND2_X1 U12632 ( .A1(n10358), .A2(n10351), .ZN(n9825) );
  OAI21_X2 U12633 ( .B1(n10378), .B2(n12170), .A(n10361), .ZN(n10398) );
  NAND2_X1 U12634 ( .A1(n12454), .A2(n10137), .ZN(n9827) );
  NAND2_X1 U12635 ( .A1(n12484), .A2(n12485), .ZN(n12486) );
  NAND3_X1 U12636 ( .A1(n10583), .A2(n16088), .A3(n16089), .ZN(n9934) );
  NAND2_X1 U12637 ( .A1(n9829), .A2(n20024), .ZN(n9828) );
  INV_X1 U12638 ( .A(n12754), .ZN(n9829) );
  AOI21_X1 U12639 ( .B1(n20024), .B2(n9831), .A(n9668), .ZN(n9830) );
  NAND2_X1 U12640 ( .A1(n20025), .A2(n20024), .ZN(n20023) );
  NAND2_X1 U12641 ( .A1(n12754), .A2(n10554), .ZN(n20025) );
  NAND3_X1 U12642 ( .A1(n9832), .A2(n16055), .A3(n9834), .ZN(n13991) );
  NAND4_X1 U12643 ( .A1(n16069), .A2(n9898), .A3(n9659), .A4(n9612), .ZN(n9832) );
  NAND3_X1 U12644 ( .A1(n16069), .A2(n9898), .A3(n9659), .ZN(n9833) );
  NAND3_X1 U12645 ( .A1(n16069), .A2(n9898), .A3(n10605), .ZN(n9836) );
  NAND2_X1 U12646 ( .A1(n10032), .A2(n10030), .ZN(n13922) );
  INV_X1 U12647 ( .A(n9839), .ZN(n13929) );
  NAND2_X1 U12648 ( .A1(n9839), .A2(n13930), .ZN(n13931) );
  NAND3_X1 U12649 ( .A1(n15839), .A2(n15837), .A3(n9843), .ZN(n17725) );
  AND2_X1 U12650 ( .A1(n10179), .A2(n10178), .ZN(n17585) );
  NAND3_X1 U12651 ( .A1(n15749), .A2(n9849), .A3(n15748), .ZN(n17455) );
  NAND2_X1 U12652 ( .A1(n9592), .A2(n9862), .ZN(n9859) );
  AND2_X2 U12653 ( .A1(n10217), .A2(n9868), .ZN(n12695) );
  NAND2_X1 U12654 ( .A1(n14643), .A2(n13289), .ZN(n9871) );
  NOR2_X1 U12655 ( .A1(n14643), .A2(n9872), .ZN(n13265) );
  OAI211_X1 U12656 ( .C1(n14643), .C2(n9874), .A(n9873), .B(n9871), .ZN(n14613) );
  INV_X1 U12657 ( .A(n9880), .ZN(n10201) );
  OR2_X2 U12658 ( .A1(n11291), .A2(n11292), .ZN(n9880) );
  NAND2_X1 U12659 ( .A1(n11238), .A2(n11392), .ZN(n9882) );
  OAI21_X1 U12660 ( .B1(n9913), .B2(n13553), .A(n16055), .ZN(n9898) );
  NAND2_X2 U12661 ( .A1(n10603), .A2(n9667), .ZN(n16069) );
  INV_X1 U12662 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9899) );
  INV_X1 U12663 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9900) );
  AND2_X2 U12664 ( .A1(n9899), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10242) );
  AND2_X2 U12665 ( .A1(n9900), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12428) );
  NAND2_X1 U12666 ( .A1(n13947), .A2(n9901), .ZN(n13930) );
  INV_X2 U12667 ( .A(n14034), .ZN(n16070) );
  NAND2_X2 U12668 ( .A1(n10453), .A2(n10374), .ZN(n10382) );
  NAND2_X2 U12669 ( .A1(n10370), .A2(n20206), .ZN(n10453) );
  NAND2_X2 U12670 ( .A1(n10613), .A2(n14000), .ZN(n13990) );
  NAND2_X1 U12671 ( .A1(n9907), .A2(n9905), .ZN(P1_U3002) );
  NAND2_X1 U12672 ( .A1(n14109), .A2(n20075), .ZN(n9907) );
  XNOR2_X2 U12673 ( .A(n9908), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14109) );
  OAI21_X2 U12674 ( .B1(n13923), .B2(n9595), .A(n9909), .ZN(n9908) );
  NAND2_X1 U12675 ( .A1(n13923), .A2(n13922), .ZN(n9909) );
  INV_X1 U12676 ( .A(n13968), .ZN(n9910) );
  NAND2_X2 U12677 ( .A1(n10587), .A2(n10521), .ZN(n13978) );
  INV_X1 U12678 ( .A(n9913), .ZN(n14030) );
  NAND3_X1 U12679 ( .A1(n10402), .A2(n20650), .A3(n10452), .ZN(n9915) );
  NAND2_X1 U12680 ( .A1(n14395), .A2(n9918), .ZN(n14893) );
  NOR2_X1 U12681 ( .A1(n14871), .A2(n14436), .ZN(n14438) );
  OR3_X1 U12682 ( .A1(n14871), .A2(n9920), .A3(n14436), .ZN(n14392) );
  INV_X1 U12683 ( .A(n9930), .ZN(n14520) );
  AND2_X2 U12684 ( .A1(n11388), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13209) );
  NAND4_X1 U12685 ( .A1(n9995), .A2(n9996), .A3(n9994), .A4(n16302), .ZN(n9932) );
  XNOR2_X2 U12686 ( .A(n9937), .B(n10373), .ZN(n20206) );
  OAI21_X2 U12687 ( .B1(n10378), .B2(n10029), .A(n10356), .ZN(n9937) );
  NAND4_X4 U12688 ( .A1(n10276), .A2(n10277), .A3(n9658), .A4(n9586), .ZN(
        n12978) );
  INV_X1 U12689 ( .A(n13544), .ZN(n12848) );
  NAND2_X1 U12690 ( .A1(n15838), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15839) );
  NOR2_X2 U12691 ( .A1(n17848), .A2(n15830), .ZN(n15831) );
  NAND3_X1 U12692 ( .A1(n9955), .A2(n9954), .A3(n9952), .ZN(n17888) );
  NAND3_X1 U12693 ( .A1(n9955), .A2(n9683), .A3(n9952), .ZN(n9957) );
  NAND2_X1 U12694 ( .A1(n10175), .A2(n9682), .ZN(n9955) );
  INV_X1 U12695 ( .A(n9957), .ZN(n17886) );
  NAND2_X1 U12696 ( .A1(n9962), .A2(n9960), .ZN(n16455) );
  NAND3_X1 U12697 ( .A1(n15734), .A2(n15730), .A3(n9680), .ZN(n9971) );
  AND3_X2 U12698 ( .A1(n11233), .A2(n11307), .A3(n11281), .ZN(n11616) );
  OAI211_X1 U12699 ( .C1(n11677), .C2(n9979), .A(n9974), .B(n9976), .ZN(n16297) );
  AND2_X1 U12700 ( .A1(n9987), .A2(n9613), .ZN(n14994) );
  NAND2_X1 U12701 ( .A1(n14934), .A2(n9666), .ZN(n9996) );
  NAND2_X1 U12702 ( .A1(n9993), .A2(n10001), .ZN(n9992) );
  NAND3_X1 U12703 ( .A1(n9996), .A2(n9995), .A3(n9994), .ZN(n15144) );
  NAND2_X1 U12704 ( .A1(n10075), .A2(n10004), .ZN(n10003) );
  NAND2_X1 U12705 ( .A1(n10016), .A2(n9626), .ZN(n12948) );
  INV_X1 U12706 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10029) );
  NAND2_X2 U12707 ( .A1(n13958), .A2(n10618), .ZN(n13947) );
  NAND3_X1 U12708 ( .A1(n10354), .A2(n10345), .A3(n10353), .ZN(n12164) );
  NOR2_X1 U12709 ( .A1(n12144), .A2(n10034), .ZN(n12135) );
  NOR2_X1 U12710 ( .A1(n10038), .A2(n10037), .ZN(n16687) );
  NOR2_X1 U12711 ( .A1(n16664), .A2(n9694), .ZN(n16656) );
  NAND3_X1 U12712 ( .A1(n16482), .A2(n16654), .A3(n10058), .ZN(n10055) );
  OR2_X1 U12713 ( .A1(n16482), .A2(n16654), .ZN(n10056) );
  INV_X1 U12714 ( .A(n10086), .ZN(n15330) );
  NAND2_X1 U12715 ( .A1(n12763), .A2(n12765), .ZN(n10088) );
  NAND3_X1 U12716 ( .A1(n12764), .A2(n10088), .A3(n10087), .ZN(n11676) );
  AND2_X4 U12717 ( .A1(n12304), .A2(n11550), .ZN(n13425) );
  NAND2_X1 U12718 ( .A1(n10089), .A2(n11777), .ZN(n13098) );
  NAND2_X1 U12719 ( .A1(n11772), .A2(n11773), .ZN(n10089) );
  NAND2_X1 U12720 ( .A1(n14492), .A2(n9704), .ZN(n14647) );
  INV_X1 U12721 ( .A(n14442), .ZN(n10095) );
  INV_X1 U12722 ( .A(n12544), .ZN(n10096) );
  NAND2_X1 U12723 ( .A1(n10096), .A2(n10097), .ZN(n12709) );
  NOR2_X1 U12724 ( .A1(n14388), .A2(n14370), .ZN(n14583) );
  OR3_X1 U12725 ( .A1(n14388), .A2(n14370), .A3(n10107), .ZN(n14585) );
  NAND2_X1 U12726 ( .A1(n14473), .A2(n9591), .ZN(n10108) );
  INV_X1 U12727 ( .A(n10116), .ZN(n14342) );
  NAND3_X1 U12728 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12729 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10127) );
  NAND3_X1 U12730 ( .A1(n10128), .A2(n10126), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14327) );
  NAND3_X1 U12731 ( .A1(n10128), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U12732 ( .A1(n12393), .A2(n10536), .ZN(n10543) );
  NAND2_X1 U12733 ( .A1(n12394), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12393) );
  XNOR2_X1 U12734 ( .A(n12226), .B(n10534), .ZN(n12394) );
  NAND4_X1 U12735 ( .A1(n10134), .A2(n10137), .A3(n10132), .A4(n10130), .ZN(
        n10527) );
  NAND3_X1 U12736 ( .A1(n10130), .A2(n10134), .A3(n10132), .ZN(n10688) );
  INV_X1 U12737 ( .A(n10402), .ZN(n10133) );
  OAI21_X1 U12738 ( .B1(n10452), .B2(n10139), .A(n9627), .ZN(n10135) );
  NAND2_X1 U12739 ( .A1(n10427), .A2(n10522), .ZN(n10140) );
  NAND2_X1 U12740 ( .A1(n9722), .A2(n10147), .ZN(n10146) );
  NOR2_X1 U12741 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10147) );
  NOR2_X2 U12742 ( .A1(n13809), .A2(n10150), .ZN(n13792) );
  INV_X1 U12743 ( .A(n20206), .ZN(n10162) );
  NAND3_X1 U12744 ( .A1(n20511), .A2(n20650), .A3(n10453), .ZN(n10163) );
  NAND2_X2 U12745 ( .A1(n10163), .A2(n10455), .ZN(n10533) );
  NAND3_X1 U12746 ( .A1(n12846), .A2(n12845), .A3(n10224), .ZN(n12862) );
  AOI21_X1 U12747 ( .B1(n14972), .B2(n9725), .A(n9640), .ZN(n10166) );
  NAND2_X1 U12748 ( .A1(n14972), .A2(n10168), .ZN(n14938) );
  NAND2_X1 U12749 ( .A1(n14972), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14964) );
  NAND2_X2 U12750 ( .A1(n15032), .A2(n9639), .ZN(n15003) );
  NAND2_X1 U12751 ( .A1(n15831), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U12752 ( .A1(n9673), .A2(n17829), .ZN(n10174) );
  NAND2_X1 U12753 ( .A1(n12031), .A2(n9663), .ZN(n12560) );
  NAND2_X2 U12754 ( .A1(n9616), .A2(n14828), .ZN(n14361) );
  INV_X1 U12755 ( .A(n12750), .ZN(n10200) );
  AND2_X2 U12756 ( .A1(n11313), .A2(n11312), .ZN(n10202) );
  NAND2_X1 U12757 ( .A1(n13266), .A2(n10208), .ZN(n10204) );
  AND3_X2 U12758 ( .A1(n10204), .A2(n9709), .A3(n10203), .ZN(n13314) );
  OR2_X2 U12759 ( .A1(n14613), .A2(n10206), .ZN(n10203) );
  INV_X1 U12760 ( .A(n10209), .ZN(n14614) );
  NAND2_X2 U12761 ( .A1(n10210), .A2(n13317), .ZN(n13341) );
  OAI21_X1 U12762 ( .B1(n14602), .B2(n14603), .A(n10210), .ZN(n14712) );
  NAND2_X2 U12763 ( .A1(n10211), .A2(n13365), .ZN(n14587) );
  NAND3_X1 U12764 ( .A1(n14597), .A2(n9645), .A3(n10212), .ZN(n10213) );
  NAND2_X1 U12765 ( .A1(n10214), .A2(n11296), .ZN(n11282) );
  NAND2_X1 U12766 ( .A1(n11303), .A2(n15537), .ZN(n11296) );
  NAND2_X2 U12767 ( .A1(n12100), .A2(n11293), .ZN(n11303) );
  NAND2_X1 U12768 ( .A1(n11281), .A2(n11301), .ZN(n10215) );
  AND3_X4 U12769 ( .A1(n11550), .A2(n15450), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13332) );
  CLKBUF_X1 U12770 ( .A(n11993), .Z(n13000) );
  NAND2_X1 U12771 ( .A1(n11993), .A2(n12007), .ZN(n10358) );
  NAND2_X1 U12772 ( .A1(n10338), .A2(n10236), .ZN(n10350) );
  NOR2_X1 U12773 ( .A1(n20137), .A2(n10344), .ZN(n20609) );
  AND2_X1 U12774 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  NAND2_X1 U12775 ( .A1(n14640), .A2(n14478), .ZN(n14462) );
  AOI221_X1 U12776 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18730), 
        .C1(n18729), .C2(n18730), .A(n18892), .ZN(n18741) );
  OAI21_X1 U12777 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18892), .A(
        n11906), .ZN(n11907) );
  NAND2_X1 U12778 ( .A1(n11274), .A2(n9606), .ZN(n11275) );
  AOI21_X1 U12779 ( .B1(n16191), .B2(n16190), .A(n19717), .ZN(n16200) );
  NOR2_X2 U12780 ( .A1(n13968), .A2(n14089), .ZN(n13946) );
  INV_X1 U12781 ( .A(n14396), .ZN(n14408) );
  INV_X1 U12782 ( .A(n11665), .ZN(n11667) );
  OR2_X1 U12783 ( .A1(n12465), .A2(n12290), .ZN(n12291) );
  OAI211_X1 U12784 ( .C1(n13534), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        n11334) );
  CLKBUF_X1 U12785 ( .A(n12299), .Z(n14546) );
  NAND2_X1 U12786 ( .A1(n12299), .A2(n12284), .ZN(n12289) );
  NAND2_X1 U12787 ( .A1(n12299), .A2(n9592), .ZN(n11366) );
  INV_X1 U12788 ( .A(n17687), .ZN(n17613) );
  NAND2_X2 U12789 ( .A1(n12499), .A2(n12498), .ZN(n13839) );
  NAND2_X1 U12790 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10221) );
  AND3_X1 U12791 ( .A1(n11536), .A2(n11535), .A3(n11534), .ZN(n10222) );
  AND3_X1 U12792 ( .A1(n11500), .A2(n11499), .A3(n11498), .ZN(n10223) );
  NAND3_X1 U12793 ( .A1(n10754), .A2(n10753), .A3(n10752), .ZN(n10224) );
  AND3_X1 U12794 ( .A1(n11467), .A2(n11466), .A3(n11465), .ZN(n10225) );
  AND3_X1 U12795 ( .A1(n11414), .A2(n11413), .A3(n11412), .ZN(n10226) );
  OR4_X1 U12796 ( .A1(n15145), .A2(n15125), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n15170), .ZN(n10227) );
  NOR2_X1 U12797 ( .A1(n20440), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10228) );
  OR2_X1 U12798 ( .A1(n13593), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10229) );
  OR2_X1 U12799 ( .A1(n14813), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10230) );
  OR2_X1 U12800 ( .A1(n13593), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10231) );
  INV_X1 U12801 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19876) );
  AND3_X1 U12802 ( .A1(n11401), .A2(n11400), .A3(n11399), .ZN(n10233) );
  INV_X1 U12803 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n16425) );
  INV_X1 U12804 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10625) );
  INV_X1 U12805 ( .A(n13465), .ZN(n14397) );
  INV_X1 U12806 ( .A(n13042), .ZN(n13831) );
  INV_X1 U12807 ( .A(n15741), .ZN(n17241) );
  INV_X1 U12808 ( .A(n11719), .ZN(n11751) );
  INV_X1 U12809 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n12070) );
  AND2_X1 U12810 ( .A1(n15407), .A2(n16277), .ZN(n10235) );
  INV_X1 U12811 ( .A(n15394), .ZN(n14801) );
  INV_X1 U12812 ( .A(n11685), .ZN(n11546) );
  INV_X1 U12813 ( .A(n10690), .ZN(n11118) );
  AND2_X1 U12814 ( .A1(n10339), .A2(n12500), .ZN(n10236) );
  INV_X1 U12815 ( .A(n15503), .ZN(n11523) );
  INV_X1 U12816 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10622) );
  INV_X1 U12817 ( .A(n10665), .ZN(n10654) );
  AOI21_X1 U12818 ( .B1(n10665), .B2(n12959), .A(n10633), .ZN(n10642) );
  NAND2_X1 U12819 ( .A1(n19817), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11554) );
  OR3_X1 U12820 ( .A1(n10654), .A2(n10653), .A3(n11996), .ZN(n10655) );
  OR2_X1 U12821 ( .A1(n10505), .A2(n10504), .ZN(n10578) );
  INV_X1 U12822 ( .A(n11559), .ZN(n11553) );
  NOR2_X1 U12823 ( .A1(n11429), .A2(n11428), .ZN(n11438) );
  NAND2_X1 U12824 ( .A1(n11304), .A2(n11303), .ZN(n11610) );
  INV_X1 U12825 ( .A(n10555), .ZN(n10562) );
  OR2_X1 U12826 ( .A1(n10518), .A2(n10517), .ZN(n10589) );
  NOR2_X1 U12827 ( .A1(n10469), .A2(n10598), .ZN(n10433) );
  NAND2_X1 U12828 ( .A1(n11553), .A2(n11552), .ZN(n11560) );
  NAND2_X1 U12829 ( .A1(n19068), .A2(n14804), .ZN(n14810) );
  INV_X1 U12830 ( .A(n15543), .ZN(n11701) );
  AND2_X1 U12831 ( .A1(n11573), .A2(n11572), .ZN(n11575) );
  AND2_X1 U12832 ( .A1(n10631), .A2(n10632), .ZN(n10629) );
  AOI21_X1 U12833 ( .B1(n10352), .B2(n12145), .A(n20136), .ZN(n10341) );
  NOR2_X1 U12834 ( .A1(n11556), .A2(n11297), .ZN(n11286) );
  INV_X1 U12835 ( .A(n14657), .ZN(n13132) );
  AND2_X1 U12836 ( .A1(n15526), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11288) );
  OR2_X1 U12837 ( .A1(n11910), .A2(n11911), .ZN(n11906) );
  NOR2_X1 U12838 ( .A1(n16983), .A2(n11806), .ZN(n15741) );
  AND2_X1 U12839 ( .A1(n12172), .A2(n12133), .ZN(n12134) );
  OR2_X1 U12840 ( .A1(n11121), .A2(n13952), .ZN(n11123) );
  INV_X1 U12841 ( .A(n11033), .ZN(n11034) );
  INV_X1 U12842 ( .A(n13810), .ZN(n10918) );
  AND2_X1 U12843 ( .A1(n13752), .A2(n13036), .ZN(n10829) );
  NAND2_X1 U12844 ( .A1(n10733), .A2(n10855), .ZN(n10741) );
  OR2_X1 U12845 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n10823) );
  NAND2_X1 U12846 ( .A1(n12965), .A2(n12848), .ZN(n12132) );
  INV_X1 U12847 ( .A(n10528), .ZN(n10432) );
  INV_X1 U12848 ( .A(n10660), .ZN(n10648) );
  NOR2_X1 U12849 ( .A1(n14675), .A2(n12910), .ZN(n12911) );
  NAND2_X1 U12850 ( .A1(n14396), .A2(n14398), .ZN(n13465) );
  BUF_X1 U12851 ( .A(n13314), .Z(n13316) );
  AND2_X1 U12852 ( .A1(n13265), .A2(n9875), .ZN(n13266) );
  INV_X1 U12853 ( .A(n14981), .ZN(n14877) );
  NOR2_X1 U12854 ( .A1(n14802), .A2(n14801), .ZN(n14803) );
  AND4_X1 U12855 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11640) );
  NOR2_X1 U12856 ( .A1(n11811), .A2(n18740), .ZN(n15739) );
  INV_X1 U12857 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20791) );
  NAND2_X1 U12858 ( .A1(n17818), .A2(n18070), .ZN(n15836) );
  NOR2_X1 U12859 ( .A1(n17315), .A2(n18308), .ZN(n13075) );
  AOI21_X1 U12860 ( .B1(n17502), .B2(n16445), .A(n18735), .ZN(n13073) );
  INV_X1 U12861 ( .A(n13596), .ZN(n13584) );
  OR2_X1 U12862 ( .A1(n11123), .A2(n11122), .ZN(n12623) );
  NAND2_X1 U12863 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11121) );
  NOR2_X1 U12864 ( .A1(n10983), .A2(n15927), .ZN(n10984) );
  AND2_X1 U12865 ( .A1(n10675), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13629) );
  NAND2_X1 U12866 ( .A1(n13946), .A2(n9595), .ZN(n10614) );
  AND2_X1 U12867 ( .A1(n20440), .A2(n10377), .ZN(n20109) );
  INV_X1 U12868 ( .A(n11751), .ZN(n14358) );
  NOR2_X1 U12869 ( .A1(n14781), .A2(n11643), .ZN(n14948) );
  NOR2_X1 U12870 ( .A1(n19050), .A2(n11643), .ZN(n14813) );
  INV_X1 U12871 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11666) );
  OR2_X1 U12872 ( .A1(n11398), .A2(n11397), .ZN(n11721) );
  INV_X1 U12873 ( .A(n11741), .ZN(n11737) );
  AND2_X1 U12874 ( .A1(n11912), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U12875 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11806) );
  NOR2_X1 U12876 ( .A1(n11812), .A2(n11814), .ZN(n15736) );
  NOR2_X1 U12877 ( .A1(n17932), .A2(n17903), .ZN(n17687) );
  INV_X1 U12878 ( .A(n18072), .ZN(n18120) );
  NOR2_X1 U12879 ( .A1(n15801), .A2(n17867), .ZN(n15803) );
  INV_X1 U12880 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n20811) );
  NAND2_X1 U12881 ( .A1(n10755), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10781) );
  INV_X1 U12882 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20862) );
  INV_X1 U12883 ( .A(n20739), .ZN(n12635) );
  OR2_X1 U12884 ( .A1(n11081), .A2(n11080), .ZN(n13695) );
  AND2_X1 U12885 ( .A1(n10830), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10846) );
  INV_X1 U12886 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10697) );
  INV_X1 U12887 ( .A(n12335), .ZN(n10695) );
  AND2_X1 U12888 ( .A1(n14091), .A2(n14090), .ZN(n14147) );
  AND2_X1 U12889 ( .A1(n14070), .A2(n14069), .ZN(n14228) );
  AND2_X1 U12890 ( .A1(n14085), .A2(n14232), .ZN(n14263) );
  NOR2_X1 U12891 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20100), .ZN(n20239) );
  OR2_X1 U12892 ( .A1(n20099), .A2(n12454), .ZN(n20208) );
  INV_X1 U12893 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20474) );
  AND2_X1 U12894 ( .A1(n11595), .A2(n11594), .ZN(n16395) );
  OR2_X1 U12895 ( .A1(n19840), .A2(n11623), .ZN(n11603) );
  NAND2_X1 U12896 ( .A1(n19087), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16196) );
  INV_X1 U12897 ( .A(n19087), .ZN(n19109) );
  INV_X1 U12898 ( .A(n12292), .ZN(n12199) );
  INV_X1 U12899 ( .A(n14948), .ZN(n14947) );
  OR3_X1 U12900 ( .A1(n14859), .A2(n11643), .A3(n16244), .ZN(n16245) );
  INV_X1 U12901 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12087) );
  AND2_X1 U12902 ( .A1(n12326), .A2(n12325), .ZN(n16413) );
  NOR2_X1 U12903 ( .A1(n15519), .A2(n15518), .ZN(n15561) );
  AND2_X1 U12904 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15511) );
  AND3_X1 U12905 ( .A1(n19397), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19431), 
        .ZN(n19403) );
  NAND2_X1 U12906 ( .A1(n15476), .A2(n19820), .ZN(n19469) );
  OR2_X1 U12907 ( .A1(n19812), .A2(n19820), .ZN(n19800) );
  NAND2_X1 U12908 ( .A1(n19812), .A2(n19820), .ZN(n19338) );
  INV_X1 U12909 ( .A(n15493), .ZN(n15558) );
  NOR2_X1 U12910 ( .A1(n18281), .A2(n11892), .ZN(n13079) );
  NOR2_X1 U12911 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16790), .ZN(n16772) );
  INV_X1 U12912 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16873) );
  NOR2_X1 U12913 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16907), .ZN(n16886) );
  NOR2_X1 U12914 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16936), .ZN(n16915) );
  INV_X1 U12915 ( .A(n16971), .ZN(n16989) );
  INV_X1 U12916 ( .A(n18300), .ZN(n17315) );
  AND4_X1 U12917 ( .A1(n17462), .A2(n15676), .A3(n18300), .A4(n11894), .ZN(
        n17502) );
  NOR2_X1 U12918 ( .A1(n17609), .A2(n17941), .ZN(n16471) );
  INV_X1 U12919 ( .A(n15827), .ZN(n16503) );
  AOI211_X1 U12920 ( .C1(n18073), .C2(n18120), .A(n15844), .B(n17962), .ZN(
        n17986) );
  NOR2_X1 U12921 ( .A1(n18188), .A2(n17862), .ZN(n17861) );
  INV_X1 U12922 ( .A(n18717), .ZN(n18738) );
  NOR2_X1 U12923 ( .A1(n18126), .A2(n18743), .ZN(n18158) );
  NOR2_X1 U12924 ( .A1(n11821), .A2(n11820), .ZN(n18925) );
  NOR2_X1 U12925 ( .A1(n11841), .A2(n11840), .ZN(n18287) );
  NAND2_X1 U12926 ( .A1(n18274), .A2(n18158), .ZN(n18228) );
  NOR3_X1 U12927 ( .A1(n20877), .A2(n19874), .A3(n19873), .ZN(n16016) );
  AND2_X1 U12928 ( .A1(n12637), .A2(n12630), .ZN(n19934) );
  OR2_X1 U12929 ( .A1(n20739), .A2(n12622), .ZN(n19889) );
  INV_X1 U12930 ( .A(n13839), .ZN(n13828) );
  OR2_X1 U12931 ( .A1(n12497), .A2(n12628), .ZN(n12212) );
  AND2_X1 U12932 ( .A1(n12107), .A2(n12629), .ZN(n19959) );
  INV_X1 U12933 ( .A(n12261), .ZN(n20003) );
  NAND2_X1 U12934 ( .A1(n10786), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10824) );
  NAND2_X1 U12935 ( .A1(n10709), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10717) );
  INV_X1 U12936 ( .A(n16067), .ZN(n20029) );
  AND2_X1 U12937 ( .A1(n14162), .A2(n14073), .ZN(n14143) );
  AND2_X1 U12938 ( .A1(n12995), .A2(n12994), .ZN(n20072) );
  OAI21_X1 U12939 ( .B1(n20052), .B2(n20056), .A(n20073), .ZN(n16120) );
  INV_X1 U12940 ( .A(n20085), .ZN(n20075) );
  INV_X1 U12941 ( .A(n20239), .ZN(n20148) );
  NOR2_X1 U12942 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16170) );
  OAI22_X1 U12943 ( .A1(n20111), .A2(n20110), .B1(n20410), .B2(n20236), .ZN(
        n20142) );
  NOR2_X1 U12944 ( .A1(n20208), .A2(n9587), .ZN(n20146) );
  INV_X1 U12945 ( .A(n20228), .ZN(n20229) );
  INV_X1 U12946 ( .A(n20287), .ZN(n20279) );
  OR2_X1 U12947 ( .A1(n20325), .A2(n9587), .ZN(n20262) );
  NAND2_X1 U12948 ( .A1(n12454), .A2(n14272), .ZN(n20325) );
  INV_X1 U12949 ( .A(n20347), .ZN(n20372) );
  NOR2_X1 U12950 ( .A1(n20451), .A2(n9587), .ZN(n20381) );
  NAND2_X1 U12951 ( .A1(n14275), .A2(n20099), .ZN(n20451) );
  OAI211_X1 U12952 ( .C1(n20579), .C2(n20549), .A(n20548), .B(n20547), .ZN(
        n20582) );
  INV_X1 U12953 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20670) );
  INV_X1 U12954 ( .A(n19091), .ZN(n19112) );
  INV_X1 U12955 ( .A(n14677), .ZN(n14658) );
  INV_X1 U12956 ( .A(n14769), .ZN(n12751) );
  INV_X1 U12957 ( .A(n19144), .ZN(n19131) );
  INV_X1 U12958 ( .A(n11980), .ZN(n11988) );
  INV_X1 U12959 ( .A(n19218), .ZN(n16302) );
  AOI21_X1 U12960 ( .B1(n14960), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14950), .ZN(n14954) );
  OR2_X1 U12961 ( .A1(n12768), .A2(n12772), .ZN(n16355) );
  AND2_X1 U12962 ( .A1(n11771), .A2(n19839), .ZN(n16358) );
  INV_X1 U12963 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15450) );
  NOR2_X1 U12964 ( .A1(n16401), .A2(n12070), .ZN(n16428) );
  OAI21_X1 U12965 ( .B1(n15482), .B2(n15485), .A(n15481), .ZN(n19247) );
  NOR2_X1 U12966 ( .A1(n19469), .A2(n19368), .ZN(n19252) );
  NOR2_X2 U12967 ( .A1(n19469), .A2(n19406), .ZN(n19298) );
  NOR2_X2 U12968 ( .A1(n19368), .A2(n19800), .ZN(n19299) );
  NOR2_X2 U12969 ( .A1(n19406), .A2(n19800), .ZN(n19330) );
  NOR2_X2 U12970 ( .A1(n19368), .A2(n19338), .ZN(n19360) );
  NOR2_X1 U12971 ( .A1(n19406), .A2(n19338), .ZN(n19369) );
  NOR2_X1 U12972 ( .A1(n19659), .A2(n19368), .ZN(n19396) );
  OAI21_X1 U12973 ( .B1(n19468), .B2(n19467), .A(n19466), .ZN(n19488) );
  OAI21_X1 U12974 ( .B1(n19503), .B2(n19518), .A(n19655), .ZN(n19520) );
  NOR2_X2 U12975 ( .A1(n19598), .A2(n19800), .ZN(n19539) );
  NOR2_X1 U12976 ( .A1(n19470), .A2(n19800), .ZN(n19549) );
  AND2_X1 U12977 ( .A1(n12817), .A2(n12816), .ZN(n19592) );
  INV_X1 U12978 ( .A(n19711), .ZN(n19640) );
  INV_X1 U12979 ( .A(n19230), .ZN(n19666) );
  INV_X1 U12980 ( .A(n19239), .ZN(n19684) );
  INV_X1 U12981 ( .A(n19661), .ZN(n19708) );
  INV_X1 U12982 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20815) );
  NAND2_X1 U12983 ( .A1(n18925), .A2(n16445), .ZN(n15673) );
  NOR3_X1 U12984 ( .A1(n17502), .A2(n15677), .A3(n18735), .ZN(n18709) );
  NOR2_X1 U12985 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16750), .ZN(n16738) );
  INV_X1 U12986 ( .A(n16965), .ZN(n16995) );
  NOR2_X1 U12987 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16810), .ZN(n16795) );
  NOR2_X1 U12988 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16862), .ZN(n16845) );
  INV_X1 U12989 ( .A(n16999), .ZN(n16969) );
  AND2_X1 U12990 ( .A1(n17305), .A2(n17424), .ZN(n17303) );
  NOR2_X1 U12991 ( .A1(n17508), .A2(n17382), .ZN(n17373) );
  NOR3_X1 U12992 ( .A1(n17309), .A2(n17429), .A3(n17308), .ZN(n17423) );
  NOR2_X2 U12993 ( .A1(n11831), .A2(n11830), .ZN(n18316) );
  INV_X1 U12994 ( .A(n18925), .ZN(n17462) );
  INV_X1 U12995 ( .A(n17741), .ZN(n17666) );
  INV_X1 U12996 ( .A(n18080), .ZN(n18002) );
  INV_X1 U12997 ( .A(n17797), .ZN(n17772) );
  INV_X1 U12998 ( .A(n17844), .ZN(n17824) );
  NOR2_X2 U12999 ( .A1(n18394), .A2(n18620), .ZN(n18653) );
  NAND2_X1 U13000 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17757), .ZN(
        n18081) );
  INV_X1 U13001 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18137) );
  INV_X1 U13002 ( .A(n18233), .ZN(n18239) );
  NAND2_X1 U13003 ( .A1(n18928), .A2(n18266), .ZN(n18394) );
  NOR2_X1 U13004 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18872), .ZN(
        n18900) );
  INV_X1 U13005 ( .A(n18773), .ZN(n18923) );
  INV_X1 U13006 ( .A(n18371), .ZN(n18435) );
  INV_X1 U13007 ( .A(n18393), .ZN(n18458) );
  INV_X1 U13008 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18748) );
  INV_X1 U13009 ( .A(n18552), .ZN(n18614) );
  INV_X1 U13010 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18885) );
  INV_X1 U13011 ( .A(n13482), .ZN(n13481) );
  INV_X1 U13012 ( .A(U212), .ZN(n16556) );
  OR2_X1 U13013 ( .A1(n12973), .A2(n11994), .ZN(n12231) );
  INV_X1 U13014 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20650) );
  NAND2_X1 U13015 ( .A1(n19889), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19926) );
  NAND2_X1 U13016 ( .A1(n19889), .A2(n12627), .ZN(n15943) );
  NAND2_X1 U13017 ( .A1(n19889), .A2(n12633), .ZN(n19948) );
  INV_X1 U13018 ( .A(n19959), .ZN(n19989) );
  NOR2_X1 U13019 ( .A1(n12231), .A2(n12230), .ZN(n12259) );
  OR2_X1 U13020 ( .A1(n12973), .A2(n10673), .ZN(n16067) );
  INV_X1 U13021 ( .A(n16064), .ZN(n20033) );
  OR2_X1 U13022 ( .A1(n13005), .A2(n12993), .ZN(n20085) );
  INV_X1 U13023 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16173) );
  NAND2_X1 U13024 ( .A1(n20146), .A2(n10688), .ZN(n20167) );
  NAND2_X1 U13025 ( .A1(n20146), .A2(n20507), .ZN(n20198) );
  NAND2_X1 U13026 ( .A1(n20205), .A2(n20174), .ZN(n20228) );
  NAND2_X1 U13027 ( .A1(n20205), .A2(n20204), .ZN(n20255) );
  OR2_X1 U13028 ( .A1(n20262), .A2(n20507), .ZN(n20287) );
  OR2_X1 U13029 ( .A1(n20325), .A2(n20541), .ZN(n20336) );
  OR2_X1 U13030 ( .A1(n20325), .A2(n20450), .ZN(n20347) );
  NAND2_X1 U13031 ( .A1(n20381), .A2(n10688), .ZN(n20402) );
  NAND2_X1 U13032 ( .A1(n20381), .A2(n20507), .ZN(n20434) );
  OR2_X1 U13033 ( .A1(n20451), .A2(n20541), .ZN(n20473) );
  OR2_X1 U13034 ( .A1(n20451), .A2(n20450), .ZN(n20506) );
  NAND2_X1 U13035 ( .A1(n20508), .A2(n20507), .ZN(n20585) );
  OR2_X1 U13036 ( .A1(n20595), .A2(n20450), .ZN(n20647) );
  INV_X1 U13037 ( .A(n20721), .ZN(n20654) );
  INV_X1 U13038 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20668) );
  INV_X1 U13039 ( .A(n20736), .ZN(n20738) );
  INV_X1 U13040 ( .A(n19799), .ZN(n19552) );
  AND2_X1 U13041 ( .A1(n12320), .A2(n12098), .ZN(n18951) );
  AOI21_X1 U13042 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(n16201) );
  OR2_X1 U13043 ( .A1(n18951), .A2(n12798), .ZN(n19091) );
  INV_X1 U13044 ( .A(n19104), .ZN(n19075) );
  OR2_X1 U13045 ( .A1(n12793), .A2(n12802), .ZN(n19021) );
  INV_X1 U13046 ( .A(n19070), .ZN(n19107) );
  INV_X1 U13047 ( .A(n19812), .ZN(n15476) );
  INV_X1 U13048 ( .A(n14652), .ZN(n14659) );
  NAND2_X1 U13049 ( .A1(n12051), .A2(n12050), .ZN(n19144) );
  NAND2_X1 U13050 ( .A1(n19144), .A2(n12065), .ZN(n14779) );
  INV_X1 U13051 ( .A(n19180), .ZN(n19212) );
  INV_X1 U13052 ( .A(n12795), .ZN(n19145) );
  INV_X1 U13053 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16262) );
  INV_X1 U13054 ( .A(n16295), .ZN(n19224) );
  NAND3_X1 U13055 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19799), .A3(n19655), 
        .ZN(n15115) );
  OR2_X1 U13056 ( .A1(n11691), .A2(n19844), .ZN(n16373) );
  INV_X1 U13057 ( .A(n16358), .ZN(n16383) );
  AOI211_X2 U13058 ( .C1(n15486), .C2(n15485), .A(n19463), .B(n15484), .ZN(
        n19251) );
  INV_X1 U13059 ( .A(n19252), .ZN(n19280) );
  NOR2_X1 U13060 ( .A1(n15502), .A2(n19463), .ZN(n19303) );
  AOI211_X2 U13061 ( .C1(n15560), .C2(n15515), .A(n19463), .B(n15514), .ZN(
        n15568) );
  AOI211_X2 U13062 ( .C1(n19312), .C2(n19309), .A(n19463), .B(n19308), .ZN(
        n19334) );
  AOI21_X1 U13063 ( .B1(n19339), .B2(n19343), .A(n19337), .ZN(n19364) );
  INV_X1 U13064 ( .A(n19369), .ZN(n19395) );
  INV_X1 U13065 ( .A(n19396), .ZN(n19425) );
  INV_X1 U13066 ( .A(n19426), .ZN(n19457) );
  AOI211_X2 U13067 ( .C1(n19464), .C2(n19467), .A(n19463), .B(n19462), .ZN(
        n19493) );
  INV_X1 U13068 ( .A(n19500), .ZN(n19523) );
  AOI21_X1 U13069 ( .B1(n12827), .B2(n12828), .A(n12826), .ZN(n19543) );
  INV_X1 U13070 ( .A(n19549), .ZN(n19576) );
  AND4_X1 U13071 ( .A1(n12815), .A2(n19655), .A3(n12817), .A4(n12814), .ZN(
        n19597) );
  AOI21_X1 U13072 ( .B1(n19607), .B2(n19604), .A(n19603), .ZN(n19647) );
  INV_X1 U13073 ( .A(n19619), .ZN(n19677) );
  OR2_X1 U13074 ( .A1(n19598), .A2(n19659), .ZN(n19711) );
  INV_X1 U13075 ( .A(n19796), .ZN(n19720) );
  NOR2_X1 U13076 ( .A1(n18709), .A2(n16607), .ZN(n18941) );
  NAND2_X1 U13077 ( .A1(n18923), .A2(n18765), .ZN(n16617) );
  INV_X1 U13078 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17847) );
  INV_X2 U13079 ( .A(n17303), .ZN(n17300) );
  AND3_X1 U13080 ( .A1(n17462), .A2(n15912), .A3(n16440), .ZN(n17305) );
  AND2_X1 U13081 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17406), .ZN(n17409) );
  INV_X1 U13082 ( .A(n16505), .ZN(n17430) );
  NOR2_X1 U13083 ( .A1(n15772), .A2(n15771), .ZN(n17437) );
  OR2_X1 U13084 ( .A1(n17533), .A2(n17358), .ZN(n17460) );
  NAND2_X1 U13085 ( .A1(n17501), .A2(n17461), .ZN(n17499) );
  INV_X1 U13086 ( .A(n17841), .ZN(n17751) );
  NAND2_X1 U13087 ( .A1(n17787), .A2(n18041), .ZN(n17741) );
  NAND2_X1 U13088 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17928), .ZN(n17797) );
  INV_X1 U13089 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18144) );
  INV_X1 U13090 ( .A(n17923), .ZN(n17915) );
  NOR2_X1 U13091 ( .A1(n17903), .A2(n17834), .ZN(n17928) );
  NAND2_X1 U13092 ( .A1(n15693), .A2(n18923), .ZN(n18248) );
  INV_X1 U13093 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18750) );
  INV_X1 U13094 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18284) );
  INV_X1 U13095 ( .A(n18322), .ZN(n18657) );
  INV_X1 U13096 ( .A(n18335), .ZN(n18681) );
  INV_X1 U13097 ( .A(n16951), .ZN(n18781) );
  INV_X1 U13098 ( .A(n18869), .ZN(n18785) );
  INV_X1 U13099 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18799) );
  INV_X1 U13100 ( .A(n16567), .ZN(n16558) );
  AND2_X2 U13101 ( .A1(n12428), .A2(n14287), .ZN(n10314) );
  AOI22_X1 U13102 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10241) );
  NOR2_X2 U13103 ( .A1(n10237), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12425) );
  AND2_X2 U13104 ( .A1(n12428), .A2(n10243), .ZN(n10320) );
  AOI22_X1 U13105 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10320), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10240) );
  AND2_X2 U13106 ( .A1(n10242), .A2(n10244), .ZN(n10300) );
  AND2_X4 U13107 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14286) );
  AND2_X4 U13108 ( .A1(n10244), .A2(n14286), .ZN(n13610) );
  AND2_X4 U13109 ( .A1(n12428), .A2(n14286), .ZN(n10420) );
  AOI22_X1 U13110 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10238) );
  NAND4_X1 U13111 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10251) );
  AOI22_X1 U13112 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10249) );
  AND2_X2 U13113 ( .A1(n10243), .A2(n10244), .ZN(n10414) );
  AOI22_X1 U13114 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13115 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10247) );
  AND2_X4 U13116 ( .A1(n14287), .A2(n10245), .ZN(n10994) );
  AOI22_X1 U13117 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10246) );
  NAND4_X1 U13118 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10250) );
  OR2_X2 U13119 ( .A1(n10251), .A2(n10250), .ZN(n10339) );
  INV_X4 U13120 ( .A(n10339), .ZN(n20124) );
  NAND2_X1 U13121 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10255) );
  NAND2_X1 U13122 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10254) );
  NAND2_X1 U13123 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10253) );
  NAND2_X1 U13124 ( .A1(n13601), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10252) );
  NAND2_X1 U13125 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10259) );
  NAND2_X1 U13126 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10258) );
  NAND2_X1 U13127 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10257) );
  NAND2_X1 U13128 ( .A1(n10994), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U13129 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U13130 ( .A1(n10300), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U13131 ( .A1(n10383), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U13132 ( .A1(n13610), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10260) );
  NAND2_X1 U13133 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10267) );
  BUF_X4 U13134 ( .A(n10320), .Z(n11137) );
  NAND2_X1 U13135 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10266) );
  NAND2_X1 U13136 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U13137 ( .A1(n10331), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10264) );
  NAND4_X4 U13138 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n12959) );
  AOI22_X1 U13139 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13140 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13141 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13142 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13143 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13144 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10278) );
  CLKBUF_X3 U13145 ( .A(n10331), .Z(n13609) );
  AOI22_X1 U13146 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13147 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U13148 ( .A1(n10345), .A2(n12978), .ZN(n20744) );
  AOI22_X1 U13149 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13150 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13151 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13152 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10280) );
  NAND4_X1 U13153 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10289) );
  AOI22_X1 U13154 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13155 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13156 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13157 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10284) );
  NAND4_X1 U13158 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10288) );
  OR2_X4 U13159 ( .A1(n10289), .A2(n10288), .ZN(n13848) );
  NAND2_X1 U13160 ( .A1(n20124), .A2(n13848), .ZN(n10352) );
  AOI22_X1 U13161 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13162 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13163 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13164 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10290) );
  NAND4_X1 U13165 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10299) );
  AOI22_X1 U13166 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13167 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13168 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10294) );
  NAND4_X1 U13169 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  AOI22_X1 U13170 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13171 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10300), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13172 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13173 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10301) );
  NAND4_X1 U13174 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10311) );
  AOI22_X1 U13175 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13176 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13177 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13178 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U13179 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  OR2_X2 U13180 ( .A1(n10311), .A2(n10310), .ZN(n12145) );
  NAND2_X1 U13181 ( .A1(n12145), .A2(n12978), .ZN(n10312) );
  OAI21_X1 U13182 ( .B1(n20124), .B2(n20744), .A(n12161), .ZN(n10367) );
  AND2_X2 U13183 ( .A1(n10344), .A2(n10524), .ZN(n10672) );
  INV_X1 U13184 ( .A(n10672), .ZN(n10313) );
  AOI22_X1 U13185 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13186 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13187 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13188 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10316) );
  NAND4_X1 U13189 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10326) );
  AOI22_X1 U13190 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13191 ( .A1(n10320), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13192 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13193 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U13194 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  OR2_X2 U13195 ( .A1(n10326), .A2(n10325), .ZN(n10346) );
  INV_X2 U13196 ( .A(n10346), .ZN(n20132) );
  INV_X1 U13197 ( .A(n12214), .ZN(n10338) );
  AOI22_X1 U13198 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13199 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13200 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13201 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10327) );
  NAND4_X1 U13202 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10337) );
  AOI22_X1 U13203 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13204 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10383), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13205 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13206 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10332) );
  NAND4_X1 U13207 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10336) );
  OR2_X4 U13208 ( .A1(n10337), .A2(n10336), .ZN(n12500) );
  NAND2_X1 U13209 ( .A1(n10350), .A2(n10524), .ZN(n10343) );
  NAND2_X1 U13210 ( .A1(n10344), .A2(n13848), .ZN(n10340) );
  AND3_X2 U13211 ( .A1(n10343), .A2(n10342), .A3(n10341), .ZN(n10354) );
  INV_X1 U13212 ( .A(n10354), .ZN(n10366) );
  XNOR2_X1 U13213 ( .A(n20670), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12007) );
  OR2_X1 U13214 ( .A1(n12214), .A2(n10339), .ZN(n10349) );
  NAND2_X1 U13215 ( .A1(n20128), .A2(n12208), .ZN(n10348) );
  AND2_X1 U13216 ( .A1(n10348), .A2(n12500), .ZN(n10362) );
  NAND2_X1 U13217 ( .A1(n12152), .A2(n20124), .ZN(n12141) );
  NAND2_X1 U13218 ( .A1(n12141), .A2(n14281), .ZN(n10351) );
  INV_X4 U13219 ( .A(n13544), .ZN(n13585) );
  NAND2_X1 U13220 ( .A1(n16170), .A2(n20650), .ZN(n11156) );
  NAND2_X1 U13221 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10376) );
  OAI21_X1 U13222 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10376), .ZN(n20406) );
  NAND2_X1 U13223 ( .A1(n20649), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15887) );
  NAND2_X1 U13224 ( .A1(n15887), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10371) );
  OAI21_X1 U13225 ( .B1(n11156), .B2(n20406), .A(n10371), .ZN(n10355) );
  INV_X1 U13226 ( .A(n10355), .ZN(n10356) );
  NAND3_X1 U13227 ( .A1(n12211), .A2(n12131), .A3(n20128), .ZN(n12160) );
  NAND2_X1 U13228 ( .A1(n12208), .A2(n12500), .ZN(n13844) );
  NAND2_X1 U13229 ( .A1(n10358), .A2(n13001), .ZN(n10359) );
  INV_X1 U13230 ( .A(n15887), .ZN(n10360) );
  MUX2_X1 U13231 ( .A(n10360), .B(n11156), .S(n20509), .Z(n10361) );
  AND2_X1 U13232 ( .A1(n12214), .A2(n10524), .ZN(n10363) );
  INV_X1 U13233 ( .A(n12131), .ZN(n12628) );
  OAI22_X1 U13234 ( .A1(n10363), .A2(n12004), .B1(n10362), .B2(n20744), .ZN(
        n10365) );
  NAND2_X1 U13235 ( .A1(n12211), .A2(n20132), .ZN(n12980) );
  NAND2_X1 U13236 ( .A1(n20101), .A2(n12959), .ZN(n12634) );
  NAND4_X1 U13237 ( .A1(n12980), .A2(n16170), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n12634), .ZN(n10364) );
  NOR2_X1 U13238 ( .A1(n10365), .A2(n10364), .ZN(n10369) );
  NAND3_X1 U13239 ( .A1(n12141), .A2(n12959), .A3(n14281), .ZN(n10368) );
  NAND2_X1 U13240 ( .A1(n10366), .A2(n12131), .ZN(n12157) );
  NAND4_X1 U13241 ( .A1(n10369), .A2(n10368), .A3(n12157), .A4(n9823), .ZN(
        n10399) );
  NAND2_X2 U13242 ( .A1(n10398), .A2(n10399), .ZN(n10452) );
  AND2_X1 U13243 ( .A1(n10371), .A2(n10029), .ZN(n10372) );
  INV_X1 U13244 ( .A(n10376), .ZN(n10375) );
  NAND2_X1 U13245 ( .A1(n10375), .A2(n10625), .ZN(n20440) );
  NAND2_X1 U13246 ( .A1(n10376), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10377) );
  OR2_X1 U13247 ( .A1(n10462), .A2(n12174), .ZN(n10380) );
  NAND2_X1 U13248 ( .A1(n15887), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10379) );
  AOI22_X1 U13249 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13250 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13251 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13252 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10384) );
  NAND4_X1 U13253 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10393) );
  AOI22_X1 U13254 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13255 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10390) );
  INV_X1 U13256 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20797) );
  AOI22_X1 U13257 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13258 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10392) );
  INV_X1 U13259 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10394) );
  OAI22_X1 U13260 ( .A1(n10660), .A2(n10394), .B1(n10468), .B2(n10547), .ZN(
        n10395) );
  INV_X1 U13261 ( .A(n10395), .ZN(n10396) );
  INV_X1 U13262 ( .A(n10398), .ZN(n10401) );
  INV_X1 U13263 ( .A(n10399), .ZN(n10400) );
  AOI22_X1 U13264 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13265 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13266 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13267 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10403) );
  NAND4_X1 U13268 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10413) );
  AOI22_X1 U13269 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13270 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10410) );
  INV_X1 U13271 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U13272 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10408) );
  NAND4_X1 U13273 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10412) );
  NOR2_X1 U13274 ( .A1(n10469), .A2(n10591), .ZN(n10435) );
  AOI22_X1 U13275 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U13276 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13277 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13278 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10415) );
  NAND4_X1 U13279 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10426) );
  AOI22_X1 U13280 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13281 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13282 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13283 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10421) );
  NAND4_X1 U13284 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  MUX2_X1 U13285 ( .A(n10435), .B(n10433), .S(n10432), .Z(n10427) );
  INV_X1 U13286 ( .A(n10427), .ZN(n10428) );
  AOI21_X1 U13287 ( .B1(n20124), .B2(n10591), .A(n20650), .ZN(n10431) );
  NAND2_X1 U13288 ( .A1(n10429), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10430) );
  OAI211_X1 U13289 ( .C1(n10432), .C2(n12978), .A(n10431), .B(n10430), .ZN(
        n10522) );
  NAND2_X1 U13290 ( .A1(n10523), .A2(n10522), .ZN(n10434) );
  INV_X1 U13291 ( .A(n10433), .ZN(n10520) );
  INV_X1 U13292 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10450) );
  INV_X1 U13293 ( .A(n10435), .ZN(n10449) );
  AOI22_X1 U13294 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13295 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10407), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13296 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13297 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13298 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10447) );
  AOI22_X1 U13299 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13300 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13301 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13302 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13601), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10442) );
  NAND4_X1 U13303 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10446) );
  INV_X1 U13304 ( .A(n10529), .ZN(n10454) );
  OR2_X1 U13305 ( .A1(n10468), .A2(n10454), .ZN(n10448) );
  OAI211_X1 U13306 ( .C1(n10660), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10451) );
  INV_X1 U13307 ( .A(n10451), .ZN(n10457) );
  OR2_X1 U13308 ( .A1(n10469), .A2(n10454), .ZN(n10455) );
  INV_X1 U13309 ( .A(n10533), .ZN(n10681) );
  NAND2_X1 U13310 ( .A1(n10680), .A2(n10681), .ZN(n10460) );
  INV_X1 U13311 ( .A(n10456), .ZN(n10458) );
  NAND2_X1 U13312 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  OR2_X1 U13313 ( .A1(n10462), .A2(n12424), .ZN(n10467) );
  INV_X1 U13314 ( .A(n11156), .ZN(n10465) );
  NAND3_X1 U13315 ( .A1(n20474), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20319) );
  INV_X1 U13316 ( .A(n20319), .ZN(n20324) );
  NAND2_X1 U13317 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20324), .ZN(
        n20317) );
  NAND2_X1 U13318 ( .A1(n20474), .A2(n20317), .ZN(n10464) );
  NAND3_X1 U13319 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20594) );
  INV_X1 U13320 ( .A(n20594), .ZN(n10463) );
  NAND2_X1 U13321 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10463), .ZN(
        n20590) );
  AOI22_X1 U13322 ( .A1(n10465), .A2(n20350), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15887), .ZN(n10466) );
  AOI22_X1 U13323 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13324 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13325 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13326 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10470) );
  NAND4_X1 U13327 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10481) );
  AOI22_X1 U13328 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13329 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13330 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10476) );
  NAND4_X1 U13331 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  AOI22_X1 U13332 ( .A1(n10648), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10665), .B2(n10566), .ZN(n10482) );
  INV_X1 U13333 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13334 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13335 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13336 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13337 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13338 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10493) );
  AOI22_X1 U13339 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13340 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13341 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11137), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13342 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10407), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10488) );
  NAND4_X1 U13343 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  NAND2_X1 U13344 ( .A1(n10665), .A2(n10567), .ZN(n10494) );
  INV_X1 U13345 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13346 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13347 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13348 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13349 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10496) );
  NAND4_X1 U13350 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10505) );
  AOI22_X1 U13351 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13352 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13353 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10500) );
  NAND4_X1 U13354 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  NAND2_X1 U13355 ( .A1(n10665), .A2(n10578), .ZN(n10506) );
  INV_X1 U13356 ( .A(n10564), .ZN(n10508) );
  AOI22_X1 U13357 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13358 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13359 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13360 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10509) );
  NAND4_X1 U13361 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10518) );
  AOI22_X1 U13362 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13363 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13364 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10513) );
  NAND4_X1 U13365 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10517) );
  AOI22_X1 U13366 ( .A1(n10648), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10665), .B2(n10589), .ZN(n10575) );
  INV_X1 U13367 ( .A(n10575), .ZN(n10519) );
  NAND2_X1 U13368 ( .A1(n13848), .A2(n12959), .ZN(n10628) );
  NOR2_X1 U13369 ( .A1(n10520), .A2(n10628), .ZN(n10521) );
  NAND2_X1 U13370 ( .A1(n20101), .A2(n10524), .ZN(n10539) );
  OAI21_X1 U13371 ( .B1(n20744), .B2(n10528), .A(n10539), .ZN(n10525) );
  INV_X1 U13372 ( .A(n10525), .ZN(n10526) );
  NAND2_X1 U13373 ( .A1(n10527), .A2(n10526), .ZN(n12224) );
  NAND2_X1 U13374 ( .A1(n10528), .A2(n10529), .ZN(n10548) );
  OAI21_X1 U13375 ( .B1(n10529), .B2(n10528), .A(n10548), .ZN(n10530) );
  OAI211_X1 U13376 ( .C1(n10530), .C2(n20744), .A(n10672), .B(n13848), .ZN(
        n10531) );
  INV_X1 U13377 ( .A(n10531), .ZN(n10532) );
  INV_X1 U13378 ( .A(n10534), .ZN(n10535) );
  OR2_X1 U13379 ( .A1(n12226), .A2(n10535), .ZN(n10536) );
  INV_X1 U13380 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10537) );
  XNOR2_X1 U13381 ( .A(n10543), .B(n10537), .ZN(n12485) );
  XNOR2_X1 U13382 ( .A(n10548), .B(n10547), .ZN(n10541) );
  INV_X1 U13383 ( .A(n20744), .ZN(n10592) );
  INV_X1 U13384 ( .A(n10539), .ZN(n10540) );
  AOI21_X1 U13385 ( .B1(n10541), .B2(n10592), .A(n10540), .ZN(n10542) );
  NAND2_X1 U13386 ( .A1(n10543), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10544) );
  INV_X1 U13387 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10545) );
  XNOR2_X1 U13388 ( .A(n10553), .B(n10545), .ZN(n12756) );
  NAND2_X1 U13389 ( .A1(n20099), .A2(n10137), .ZN(n10552) );
  NAND2_X1 U13390 ( .A1(n10548), .A2(n10547), .ZN(n10569) );
  INV_X1 U13391 ( .A(n10566), .ZN(n10549) );
  XNOR2_X1 U13392 ( .A(n10569), .B(n10549), .ZN(n10550) );
  NAND2_X1 U13393 ( .A1(n10550), .A2(n10592), .ZN(n10551) );
  NAND2_X1 U13394 ( .A1(n10552), .A2(n10551), .ZN(n12755) );
  NAND2_X1 U13395 ( .A1(n12756), .A2(n12755), .ZN(n12754) );
  NAND2_X1 U13396 ( .A1(n10553), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10554) );
  XNOR2_X1 U13397 ( .A(n10563), .B(n10555), .ZN(n10714) );
  NAND2_X1 U13398 ( .A1(n10714), .A2(n10137), .ZN(n10559) );
  NAND2_X1 U13399 ( .A1(n10569), .A2(n10566), .ZN(n10556) );
  XNOR2_X1 U13400 ( .A(n10556), .B(n10567), .ZN(n10557) );
  NAND2_X1 U13401 ( .A1(n10557), .A2(n10592), .ZN(n10558) );
  NAND2_X1 U13402 ( .A1(n10559), .A2(n10558), .ZN(n10561) );
  INV_X1 U13403 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10560) );
  XNOR2_X1 U13404 ( .A(n10561), .B(n10560), .ZN(n20024) );
  OR2_X1 U13405 ( .A1(n10563), .A2(n10562), .ZN(n10565) );
  NAND2_X1 U13406 ( .A1(n10722), .A2(n10137), .ZN(n10572) );
  AND2_X1 U13407 ( .A1(n10567), .A2(n10566), .ZN(n10568) );
  NAND2_X1 U13408 ( .A1(n10569), .A2(n10568), .ZN(n10577) );
  XNOR2_X1 U13409 ( .A(n10577), .B(n10578), .ZN(n10570) );
  NAND2_X1 U13410 ( .A1(n10570), .A2(n10592), .ZN(n10571) );
  NAND2_X1 U13411 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  INV_X1 U13412 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16168) );
  XNOR2_X1 U13413 ( .A(n10573), .B(n16168), .ZN(n16088) );
  NAND2_X1 U13414 ( .A1(n10573), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13415 ( .A1(n10576), .A2(n10575), .ZN(n10732) );
  NAND3_X1 U13416 ( .A1(n10587), .A2(n10137), .A3(n10732), .ZN(n10582) );
  INV_X1 U13417 ( .A(n10577), .ZN(n10579) );
  NAND2_X1 U13418 ( .A1(n10579), .A2(n10578), .ZN(n10588) );
  XNOR2_X1 U13419 ( .A(n10588), .B(n10589), .ZN(n10580) );
  NAND2_X1 U13420 ( .A1(n10580), .A2(n10592), .ZN(n10581) );
  NAND2_X1 U13421 ( .A1(n10582), .A2(n10581), .ZN(n16083) );
  OR2_X1 U13422 ( .A1(n16083), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10583) );
  INV_X1 U13423 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13424 ( .A1(n10665), .A2(n10591), .ZN(n10584) );
  OAI21_X1 U13425 ( .B1(n10585), .B2(n10660), .A(n10584), .ZN(n10586) );
  NAND2_X1 U13426 ( .A1(n10733), .A2(n10137), .ZN(n10595) );
  INV_X1 U13427 ( .A(n10588), .ZN(n10590) );
  NAND2_X1 U13428 ( .A1(n10590), .A2(n10589), .ZN(n10599) );
  XNOR2_X1 U13429 ( .A(n10599), .B(n10591), .ZN(n10593) );
  NAND2_X1 U13430 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NAND2_X1 U13431 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  OR2_X1 U13432 ( .A1(n10596), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12988) );
  NAND2_X1 U13433 ( .A1(n12990), .A2(n12988), .ZN(n10597) );
  NAND2_X1 U13434 ( .A1(n10596), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12987) );
  NAND2_X1 U13435 ( .A1(n10597), .A2(n12987), .ZN(n13025) );
  OR3_X1 U13436 ( .A1(n10599), .A2(n10598), .A3(n20744), .ZN(n10600) );
  NAND2_X1 U13437 ( .A1(n16070), .A2(n10600), .ZN(n13026) );
  OR2_X1 U13438 ( .A1(n13026), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10601) );
  NAND2_X1 U13439 ( .A1(n13026), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10602) );
  INV_X1 U13440 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U13441 ( .A1(n16070), .A2(n10604), .ZN(n10605) );
  INV_X1 U13442 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14077) );
  INV_X1 U13443 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14248) );
  AND2_X1 U13444 ( .A1(n13978), .A2(n14248), .ZN(n14044) );
  NAND3_X1 U13445 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13446 ( .A1(n16070), .A2(n10606), .ZN(n10607) );
  NAND2_X1 U13447 ( .A1(n16051), .A2(n10607), .ZN(n16027) );
  INV_X1 U13448 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16114) );
  OR2_X1 U13449 ( .A1(n13978), .A2(n16114), .ZN(n10608) );
  NAND2_X1 U13450 ( .A1(n16053), .A2(n10608), .ZN(n10610) );
  INV_X1 U13451 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13547) );
  NOR2_X1 U13452 ( .A1(n9595), .A2(n13547), .ZN(n16031) );
  OR2_X1 U13453 ( .A1(n13978), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14033) );
  NAND2_X1 U13454 ( .A1(n9595), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13455 ( .A1(n14033), .A2(n10609), .ZN(n16033) );
  NAND2_X1 U13456 ( .A1(n16055), .A2(n13547), .ZN(n16040) );
  INV_X1 U13457 ( .A(n10610), .ZN(n10612) );
  NOR2_X1 U13458 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14041) );
  AND2_X1 U13459 ( .A1(n14041), .A2(n14248), .ZN(n10611) );
  OR2_X1 U13460 ( .A1(n13978), .A2(n10611), .ZN(n14028) );
  NAND2_X1 U13461 ( .A1(n10612), .A2(n14028), .ZN(n16028) );
  XNOR2_X1 U13462 ( .A(n16055), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14021) );
  INV_X1 U13463 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14182) );
  INV_X1 U13464 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14008) );
  INV_X1 U13465 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14146) );
  INV_X1 U13466 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14165) );
  INV_X1 U13467 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14086) );
  NAND3_X1 U13468 ( .A1(n14146), .A2(n14165), .A3(n14086), .ZN(n13938) );
  NAND2_X1 U13469 ( .A1(n10616), .A2(n14000), .ZN(n10615) );
  AND2_X1 U13470 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U13471 ( .A1(n14073), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14089) );
  NAND2_X1 U13472 ( .A1(n10615), .A2(n10614), .ZN(n13956) );
  INV_X1 U13473 ( .A(n10616), .ZN(n10617) );
  NAND2_X1 U13474 ( .A1(n10617), .A2(n14000), .ZN(n10618) );
  INV_X1 U13475 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10620) );
  INV_X1 U13476 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10619) );
  AND2_X1 U13477 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14074) );
  MUX2_X1 U13478 ( .A(n10622), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10639) );
  NAND2_X1 U13479 ( .A1(n20509), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10640) );
  INV_X1 U13480 ( .A(n10640), .ZN(n10621) );
  NAND2_X1 U13481 ( .A1(n10639), .A2(n10621), .ZN(n10624) );
  NAND2_X1 U13482 ( .A1(n10622), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13483 ( .A1(n10624), .A2(n10623), .ZN(n10647) );
  MUX2_X1 U13484 ( .A(n10625), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10646) );
  NAND2_X1 U13485 ( .A1(n10647), .A2(n10646), .ZN(n10627) );
  NAND2_X1 U13486 ( .A1(n10625), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13487 ( .A1(n10627), .A2(n10626), .ZN(n10631) );
  XNOR2_X1 U13488 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10632) );
  NAND3_X1 U13489 ( .A1(n16173), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10664), .ZN(n11998) );
  INV_X1 U13490 ( .A(n11998), .ZN(n10661) );
  INV_X1 U13491 ( .A(n10629), .ZN(n10630) );
  OAI21_X1 U13492 ( .B1(n10632), .B2(n10631), .A(n10630), .ZN(n11995) );
  NOR2_X1 U13493 ( .A1(n13848), .A2(n20650), .ZN(n10633) );
  NAND2_X1 U13494 ( .A1(n10642), .A2(n12959), .ZN(n10641) );
  NOR2_X1 U13495 ( .A1(n10641), .A2(n11998), .ZN(n10658) );
  OAI21_X1 U13496 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20509), .A(
        n10640), .ZN(n10635) );
  NOR2_X1 U13497 ( .A1(n10654), .A2(n10635), .ZN(n10638) );
  NAND2_X1 U13498 ( .A1(n20128), .A2(n12978), .ZN(n10634) );
  NAND2_X1 U13499 ( .A1(n10634), .A2(n10345), .ZN(n10653) );
  INV_X1 U13500 ( .A(n10635), .ZN(n10636) );
  OAI211_X1 U13501 ( .C1(n12015), .C2(n20101), .A(n10653), .B(n10636), .ZN(
        n10637) );
  OAI21_X1 U13502 ( .B1(n10638), .B2(n10668), .A(n10637), .ZN(n10644) );
  XOR2_X1 U13503 ( .A(n10640), .B(n10639), .Z(n11997) );
  OAI211_X1 U13504 ( .C1(n10644), .C2(n10642), .A(n11997), .B(n10641), .ZN(
        n10652) );
  INV_X1 U13505 ( .A(n10642), .ZN(n10643) );
  NOR2_X1 U13506 ( .A1(n11997), .A2(n10643), .ZN(n10645) );
  NAND2_X1 U13507 ( .A1(n10645), .A2(n10644), .ZN(n10651) );
  XNOR2_X1 U13508 ( .A(n10647), .B(n10646), .ZN(n11996) );
  NAND2_X1 U13509 ( .A1(n10648), .A2(n11996), .ZN(n10649) );
  OAI211_X1 U13510 ( .C1(n10654), .C2(n11996), .A(n10649), .B(n10653), .ZN(
        n10650) );
  NAND3_X1 U13511 ( .A1(n10652), .A2(n10651), .A3(n10650), .ZN(n10656) );
  AOI22_X1 U13512 ( .A1(n10656), .A2(n10655), .B1(n10660), .B2(n11995), .ZN(
        n10657) );
  AOI211_X1 U13513 ( .C1(n10668), .C2(n11995), .A(n10658), .B(n10657), .ZN(
        n10659) );
  AOI21_X1 U13514 ( .B1(n10661), .B2(n10660), .A(n10659), .ZN(n10662) );
  AOI21_X1 U13515 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20650), .A(
        n10662), .ZN(n10667) );
  INV_X1 U13516 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20094) );
  NOR2_X1 U13517 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20094), .ZN(
        n10663) );
  NAND2_X1 U13518 ( .A1(n12000), .A2(n10665), .ZN(n10666) );
  NAND2_X1 U13519 ( .A1(n10667), .A2(n10666), .ZN(n10670) );
  NAND2_X1 U13520 ( .A1(n12000), .A2(n10668), .ZN(n10669) );
  NAND2_X1 U13521 ( .A1(n14281), .A2(n20101), .ZN(n10671) );
  NAND3_X1 U13522 ( .A1(n12152), .A2(n10672), .A3(n10671), .ZN(n12009) );
  NOR2_X1 U13523 ( .A1(n12009), .A2(n12015), .ZN(n15875) );
  OR2_X1 U13524 ( .A1(n15887), .A2(n20650), .ZN(n19849) );
  NAND2_X1 U13525 ( .A1(n15875), .A2(n12976), .ZN(n10673) );
  NAND2_X1 U13526 ( .A1(n14109), .A2(n20029), .ZN(n11162) );
  INV_X1 U13527 ( .A(n13844), .ZN(n10674) );
  NAND2_X1 U13528 ( .A1(n10674), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10706) );
  INV_X2 U13529 ( .A(n10823), .ZN(n13622) );
  XNOR2_X1 U13530 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12481) );
  AOI21_X1 U13531 ( .B1(n13622), .B2(n12481), .A(n13629), .ZN(n10677) );
  NOR2_X2 U13532 ( .A1(n12500), .A2(n10675), .ZN(n10690) );
  INV_X1 U13533 ( .A(n11118), .ZN(n10874) );
  NAND2_X1 U13534 ( .A1(n10874), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10676) );
  OAI211_X1 U13535 ( .C1(n10706), .C2(n12174), .A(n10677), .B(n10676), .ZN(
        n10678) );
  INV_X1 U13536 ( .A(n10678), .ZN(n10679) );
  NAND2_X1 U13537 ( .A1(n13629), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10696) );
  NAND2_X1 U13538 ( .A1(n12446), .A2(n10855), .ZN(n10687) );
  NAND2_X1 U13539 ( .A1(n10874), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U13540 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10683) );
  OAI211_X1 U13541 ( .C1(n10706), .C2(n10029), .A(n10684), .B(n10683), .ZN(
        n10685) );
  INV_X1 U13542 ( .A(n10685), .ZN(n10686) );
  NAND2_X1 U13543 ( .A1(n10687), .A2(n10686), .ZN(n12219) );
  NAND2_X1 U13544 ( .A1(n10688), .A2(n20132), .ZN(n10689) );
  NAND2_X1 U13545 ( .A1(n10689), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12204) );
  INV_X1 U13546 ( .A(n13768), .ZN(n20207) );
  NAND2_X1 U13547 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10692) );
  NAND2_X1 U13548 ( .A1(n10690), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10691) );
  OAI211_X1 U13549 ( .C1(n10706), .C2(n12170), .A(n10692), .B(n10691), .ZN(
        n10693) );
  AOI21_X1 U13550 ( .B1(n20207), .B2(n10855), .A(n10693), .ZN(n12203) );
  OR2_X1 U13551 ( .A1(n12204), .A2(n12203), .ZN(n12206) );
  NAND2_X1 U13552 ( .A1(n12203), .A2(n13622), .ZN(n10694) );
  NAND2_X1 U13553 ( .A1(n12206), .A2(n10694), .ZN(n12218) );
  NAND2_X1 U13554 ( .A1(n12219), .A2(n12218), .ZN(n12335) );
  NAND2_X1 U13555 ( .A1(n10234), .A2(n10695), .ZN(n12336) );
  NAND2_X1 U13556 ( .A1(n20099), .A2(n10855), .ZN(n10705) );
  INV_X1 U13557 ( .A(n10698), .ZN(n10700) );
  INV_X1 U13558 ( .A(n10709), .ZN(n10699) );
  OAI21_X1 U13559 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10700), .A(
        n10699), .ZN(n12758) );
  AOI22_X1 U13560 ( .A1(n13622), .A2(n12758), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U13561 ( .A1(n10874), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10701) );
  OAI211_X1 U13562 ( .C1(n10706), .C2(n12424), .A(n10702), .B(n10701), .ZN(
        n10703) );
  INV_X1 U13563 ( .A(n10703), .ZN(n10704) );
  NAND2_X1 U13564 ( .A1(n10705), .A2(n10704), .ZN(n12452) );
  NAND2_X1 U13565 ( .A1(n12453), .A2(n12452), .ZN(n12451) );
  INV_X1 U13566 ( .A(n12451), .ZN(n10716) );
  INV_X1 U13567 ( .A(n10706), .ZN(n10707) );
  NAND2_X1 U13568 ( .A1(n10707), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10712) );
  INV_X1 U13569 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19927) );
  AOI21_X1 U13570 ( .B1(n19927), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10708) );
  AOI21_X1 U13571 ( .B1(n10874), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10708), .ZN(
        n10711) );
  OAI21_X1 U13572 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10709), .A(
        n10717), .ZN(n20032) );
  INV_X1 U13573 ( .A(n20032), .ZN(n10710) );
  AOI22_X1 U13574 ( .A1(n10712), .A2(n10711), .B1(n13622), .B2(n10710), .ZN(
        n10713) );
  AOI21_X1 U13575 ( .B1(n10714), .B2(n10855), .A(n10713), .ZN(n12557) );
  NAND2_X1 U13576 ( .A1(n10716), .A2(n10715), .ZN(n12656) );
  INV_X1 U13577 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10720) );
  INV_X1 U13578 ( .A(n10717), .ZN(n10718) );
  INV_X1 U13579 ( .A(n10725), .ZN(n10726) );
  OAI21_X1 U13580 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10718), .A(
        n10726), .ZN(n19921) );
  AOI22_X1 U13581 ( .A1(n13622), .A2(n19921), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10719) );
  OAI21_X1 U13582 ( .B1(n11118), .B2(n10720), .A(n10719), .ZN(n10721) );
  INV_X1 U13583 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10730) );
  INV_X1 U13584 ( .A(n10734), .ZN(n10735) );
  INV_X1 U13585 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13586 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  NAND2_X1 U13587 ( .A1(n10735), .A2(n10728), .ZN(n19907) );
  AOI22_X1 U13588 ( .A1(n19907), .A2(n13622), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10729) );
  OAI21_X1 U13589 ( .B1(n11118), .B2(n10730), .A(n10729), .ZN(n10731) );
  INV_X1 U13590 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19886) );
  INV_X1 U13591 ( .A(n13629), .ZN(n10894) );
  INV_X1 U13592 ( .A(n10755), .ZN(n10737) );
  NAND2_X1 U13593 ( .A1(n10735), .A2(n19886), .ZN(n10736) );
  NAND2_X1 U13594 ( .A1(n10737), .A2(n10736), .ZN(n19896) );
  NAND2_X1 U13595 ( .A1(n19896), .A2(n13622), .ZN(n10738) );
  OAI21_X1 U13596 ( .B1(n19886), .B2(n10894), .A(n10738), .ZN(n10739) );
  AOI21_X1 U13597 ( .B1(n10874), .B2(P1_EAX_REG_7__SCAN_IN), .A(n10739), .ZN(
        n10740) );
  AOI22_X1 U13598 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13599 ( .A1(n13608), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13600 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13601 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10751) );
  AOI22_X1 U13602 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13603 ( .A1(n13607), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10407), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13604 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13605 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U13606 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10750) );
  OAI21_X1 U13607 ( .B1(n10751), .B2(n10750), .A(n10855), .ZN(n10754) );
  XNOR2_X1 U13608 ( .A(n10755), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13028) );
  AOI22_X1 U13609 ( .A1(n13028), .A2(n13622), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13610 ( .A1(n10690), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10752) );
  XOR2_X1 U13611 ( .A(n19876), .B(n10781), .Z(n19878) );
  INV_X1 U13612 ( .A(n19878), .ZN(n10770) );
  AOI22_X1 U13613 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13614 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13615 ( .A1(n13608), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13616 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10756) );
  NAND4_X1 U13617 ( .A1(n10759), .A2(n10758), .A3(n10757), .A4(n10756), .ZN(
        n10765) );
  AOI22_X1 U13618 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13619 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13620 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13621 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10760) );
  NAND4_X1 U13622 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  OAI21_X1 U13623 ( .B1(n10765), .B2(n10764), .A(n10855), .ZN(n10768) );
  NAND2_X1 U13624 ( .A1(n10874), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13625 ( .A1(n13629), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10766) );
  NAND3_X1 U13626 ( .A1(n10768), .A2(n10767), .A3(n10766), .ZN(n10769) );
  AOI21_X1 U13627 ( .B1(n10770), .B2(n13622), .A(n10769), .ZN(n12929) );
  AOI22_X1 U13628 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10407), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13629 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13630 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13631 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13632 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10780) );
  AOI22_X1 U13633 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13634 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13635 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13636 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10775) );
  NAND4_X1 U13637 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  NOR2_X1 U13638 ( .A1(n10780), .A2(n10779), .ZN(n10784) );
  XNOR2_X1 U13639 ( .A(n10785), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U13640 ( .A1(n12953), .A2(n13622), .ZN(n10783) );
  AOI22_X1 U13641 ( .A1(n10690), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13629), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10782) );
  OAI211_X1 U13642 ( .C1(n10784), .C2(n9765), .A(n10783), .B(n10782), .ZN(
        n12942) );
  NAND2_X1 U13643 ( .A1(n10690), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10788) );
  OAI21_X1 U13644 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10786), .A(
        n10824), .ZN(n16078) );
  AOI22_X1 U13645 ( .A1(n13622), .A2(n16078), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13646 ( .A1(n10788), .A2(n10787), .ZN(n13011) );
  AOI22_X1 U13647 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13648 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13649 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13650 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10789) );
  NAND4_X1 U13651 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10798) );
  AOI22_X1 U13652 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13653 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13654 ( .A1(n13608), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13655 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10793) );
  NAND4_X1 U13656 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10797) );
  OR2_X1 U13657 ( .A1(n10798), .A2(n10797), .ZN(n10799) );
  AND2_X1 U13658 ( .A1(n10855), .A2(n10799), .ZN(n13033) );
  INV_X1 U13659 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U13660 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13661 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10407), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13662 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13663 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U13664 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10809) );
  AOI22_X1 U13665 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13666 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13667 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10804) );
  NAND4_X1 U13668 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10808) );
  OAI21_X1 U13669 ( .B1(n10809), .B2(n10808), .A(n10855), .ZN(n10811) );
  XNOR2_X1 U13670 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10830), .ZN(
        n14048) );
  AOI22_X1 U13671 ( .A1(n13622), .A2(n14048), .B1(n13629), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10810) );
  OAI211_X1 U13672 ( .C1(n11118), .C2(n13918), .A(n10811), .B(n10810), .ZN(
        n13752) );
  AOI22_X1 U13673 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13674 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9594), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13675 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11089), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13676 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10407), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13677 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10822) );
  AOI22_X1 U13678 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13679 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13680 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10993), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13681 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10817) );
  NAND4_X1 U13682 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        n10821) );
  NOR2_X1 U13683 ( .A1(n10822), .A2(n10821), .ZN(n10828) );
  AOI21_X1 U13684 ( .B1(n20808), .B2(n10824), .A(n10830), .ZN(n16063) );
  OAI22_X1 U13685 ( .A1(n10823), .A2(n16063), .B1(n10894), .B2(n20808), .ZN(
        n10825) );
  INV_X1 U13686 ( .A(n10825), .ZN(n10827) );
  NAND2_X1 U13687 ( .A1(n10690), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10826) );
  OAI211_X1 U13688 ( .C1(n9765), .C2(n10828), .A(n10827), .B(n10826), .ZN(
        n13036) );
  XOR2_X1 U13689 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10846), .Z(
        n16058) );
  INV_X1 U13690 ( .A(n16058), .ZN(n10845) );
  AOI22_X1 U13691 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13692 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13693 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13694 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10831) );
  NAND4_X1 U13695 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n10840) );
  AOI22_X1 U13696 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13697 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13698 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13699 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10835) );
  NAND4_X1 U13700 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10839) );
  OAI21_X1 U13701 ( .B1(n10840), .B2(n10839), .A(n10855), .ZN(n10843) );
  NAND2_X1 U13702 ( .A1(n10690), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10842) );
  NAND2_X1 U13703 ( .A1(n13629), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10841) );
  NAND3_X1 U13704 ( .A1(n10843), .A2(n10842), .A3(n10841), .ZN(n10844) );
  AOI21_X1 U13705 ( .B1(n10845), .B2(n13622), .A(n10844), .ZN(n13043) );
  XNOR2_X1 U13706 ( .A(n10878), .B(n10877), .ZN(n16045) );
  AOI22_X1 U13707 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13708 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13709 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13710 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10847) );
  NAND4_X1 U13711 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n10857) );
  AOI22_X1 U13712 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13713 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13714 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13715 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13716 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10856) );
  OAI21_X1 U13717 ( .B1(n10857), .B2(n10856), .A(n10855), .ZN(n10859) );
  NAND2_X1 U13718 ( .A1(n10690), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10858) );
  OAI211_X1 U13719 ( .C1(n10894), .C2(n10877), .A(n10859), .B(n10858), .ZN(
        n10860) );
  AOI21_X1 U13720 ( .B1(n16045), .B2(n13622), .A(n10860), .ZN(n13832) );
  INV_X1 U13721 ( .A(n13832), .ZN(n10861) );
  INV_X1 U13722 ( .A(n14281), .ZN(n12166) );
  AOI22_X1 U13723 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13724 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13725 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13726 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10862) );
  NAND4_X1 U13727 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n10871) );
  AOI22_X1 U13728 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11131), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13729 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13730 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13731 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10866) );
  NAND4_X1 U13732 ( .A1(n10869), .A2(n10868), .A3(n10867), .A4(n10866), .ZN(
        n10870) );
  NOR2_X1 U13733 ( .A1(n10871), .A2(n10870), .ZN(n10876) );
  NAND2_X1 U13734 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10872) );
  NAND2_X1 U13735 ( .A1(n10823), .A2(n10872), .ZN(n10873) );
  AOI21_X1 U13736 ( .B1(n10874), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10873), .ZN(
        n10875) );
  OAI21_X1 U13737 ( .B1(n13625), .B2(n10876), .A(n10875), .ZN(n10882) );
  OAI21_X1 U13738 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10879), .A(
        n10912), .ZN(n16038) );
  INV_X1 U13739 ( .A(n16038), .ZN(n10880) );
  NAND2_X1 U13740 ( .A1(n10880), .A2(n13622), .ZN(n10881) );
  NAND2_X1 U13741 ( .A1(n10882), .A2(n10881), .ZN(n13824) );
  AOI22_X1 U13742 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13743 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13744 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13745 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10883) );
  NAND4_X1 U13746 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(
        n10892) );
  AOI22_X1 U13747 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13748 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13749 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13750 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10887) );
  NAND4_X1 U13751 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10891) );
  OR2_X1 U13752 ( .A1(n10892), .A2(n10891), .ZN(n10893) );
  NAND2_X1 U13753 ( .A1(n11144), .A2(n10893), .ZN(n10897) );
  XNOR2_X1 U13754 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10912), .ZN(
        n15973) );
  OAI22_X1 U13755 ( .A1(n10823), .A2(n15973), .B1(n15971), .B2(n10894), .ZN(
        n10895) );
  AOI21_X1 U13756 ( .B1(n10690), .B2(P1_EAX_REG_17__SCAN_IN), .A(n10895), .ZN(
        n10896) );
  NAND2_X1 U13757 ( .A1(n10897), .A2(n10896), .ZN(n13817) );
  AOI22_X1 U13758 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13759 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13760 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10899) );
  NAND4_X1 U13761 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n10907) );
  AOI22_X1 U13762 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13763 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13764 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13765 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10902) );
  NAND4_X1 U13766 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n10906) );
  NOR2_X1 U13767 ( .A1(n10907), .A2(n10906), .ZN(n10911) );
  INV_X1 U13768 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20542) );
  OAI21_X1 U13769 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20542), .A(
        n10675), .ZN(n10908) );
  INV_X1 U13770 ( .A(n10908), .ZN(n10909) );
  AOI21_X1 U13771 ( .B1(n10690), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10909), .ZN(
        n10910) );
  OAI21_X1 U13772 ( .B1(n13625), .B2(n10911), .A(n10910), .ZN(n10917) );
  INV_X1 U13773 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14024) );
  INV_X1 U13774 ( .A(n10914), .ZN(n10913) );
  NAND2_X1 U13775 ( .A1(n14024), .A2(n10913), .ZN(n10915) );
  AND2_X1 U13776 ( .A1(n10915), .A2(n10948), .ZN(n15962) );
  NAND2_X1 U13777 ( .A1(n15962), .A2(n13622), .ZN(n10916) );
  NAND2_X1 U13778 ( .A1(n10917), .A2(n10916), .ZN(n13810) );
  AOI22_X1 U13779 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13780 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13781 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13782 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10919) );
  NAND4_X1 U13783 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n10928) );
  AOI22_X1 U13784 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13785 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13786 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13787 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10923) );
  NAND4_X1 U13788 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n10927) );
  NOR2_X1 U13789 ( .A1(n10928), .A2(n10927), .ZN(n10932) );
  NAND2_X1 U13790 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10929) );
  NAND2_X1 U13791 ( .A1(n10823), .A2(n10929), .ZN(n10930) );
  AOI21_X1 U13792 ( .B1(n10690), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10930), .ZN(
        n10931) );
  OAI21_X1 U13793 ( .B1(n13625), .B2(n10932), .A(n10931), .ZN(n10934) );
  XNOR2_X1 U13794 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n10948), .ZN(
        n15949) );
  NAND2_X1 U13795 ( .A1(n13622), .A2(n15949), .ZN(n10933) );
  NAND2_X1 U13796 ( .A1(n10934), .A2(n10933), .ZN(n13802) );
  AOI22_X1 U13797 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13798 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9594), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13799 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13800 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13801 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10944) );
  AOI22_X1 U13802 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10988), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13803 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13804 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10475), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U13805 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10943) );
  NOR2_X1 U13806 ( .A1(n10944), .A2(n10943), .ZN(n10947) );
  INV_X1 U13807 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15939) );
  OAI21_X1 U13808 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15939), .A(n10823), 
        .ZN(n10945) );
  AOI21_X1 U13809 ( .B1(n10690), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10945), .ZN(
        n10946) );
  OAI21_X1 U13810 ( .B1(n13625), .B2(n10947), .A(n10946), .ZN(n10952) );
  OAI21_X1 U13811 ( .B1(n10950), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n10983), .ZN(n15947) );
  OR2_X1 U13812 ( .A1(n15947), .A2(n10823), .ZN(n10951) );
  AOI22_X1 U13813 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13814 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13815 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U13816 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10953) );
  NAND4_X1 U13817 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10962) );
  AOI22_X1 U13818 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13819 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13820 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13821 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10957) );
  NAND4_X1 U13822 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10961) );
  NOR2_X1 U13823 ( .A1(n10962), .A2(n10961), .ZN(n10966) );
  INV_X1 U13824 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15927) );
  NOR2_X1 U13825 ( .A1(n15927), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10963) );
  OR2_X1 U13826 ( .A1(n13622), .A2(n10963), .ZN(n10964) );
  AOI21_X1 U13827 ( .B1(n10690), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10964), .ZN(
        n10965) );
  OAI21_X1 U13828 ( .B1(n13625), .B2(n10966), .A(n10965), .ZN(n10968) );
  XNOR2_X1 U13829 ( .A(n10983), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15935) );
  NAND2_X1 U13830 ( .A1(n15935), .A2(n13622), .ZN(n10967) );
  AOI22_X1 U13831 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13832 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U13833 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13834 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U13835 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10978) );
  AOI22_X1 U13836 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13837 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13838 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13839 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10973) );
  NAND4_X1 U13840 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10977) );
  NOR2_X1 U13841 ( .A1(n10978), .A2(n10977), .ZN(n10982) );
  NAND2_X1 U13842 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10979) );
  NAND2_X1 U13843 ( .A1(n10823), .A2(n10979), .ZN(n10980) );
  AOI21_X1 U13844 ( .B1(n10690), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10980), .ZN(
        n10981) );
  OAI21_X1 U13845 ( .B1(n13625), .B2(n10982), .A(n10981), .ZN(n10987) );
  OR2_X1 U13846 ( .A1(n10984), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10985) );
  AND2_X1 U13847 ( .A1(n11033), .A2(n10985), .ZN(n13996) );
  NAND2_X1 U13848 ( .A1(n13996), .A2(n13622), .ZN(n10986) );
  NAND2_X1 U13849 ( .A1(n10987), .A2(n10986), .ZN(n13739) );
  AOI22_X1 U13850 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13851 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13852 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13853 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10989) );
  NAND4_X1 U13854 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n11000) );
  AOI22_X1 U13855 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13856 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13857 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10331), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13858 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10995) );
  NAND4_X1 U13859 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n10999) );
  NOR2_X1 U13860 ( .A1(n11000), .A2(n10999), .ZN(n11017) );
  AOI22_X1 U13861 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13862 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U13863 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13864 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11001) );
  NAND4_X1 U13865 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11010) );
  AOI22_X1 U13866 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U13867 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U13868 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13869 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11005) );
  NAND4_X1 U13870 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n11009) );
  NOR2_X1 U13871 ( .A1(n11010), .A2(n11009), .ZN(n11018) );
  XOR2_X1 U13872 ( .A(n11017), .B(n11018), .Z(n11011) );
  NAND2_X1 U13873 ( .A1(n11011), .A2(n11144), .ZN(n11014) );
  INV_X1 U13874 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15926) );
  OAI21_X1 U13875 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15926), .A(n10823), 
        .ZN(n11012) );
  AOI21_X1 U13876 ( .B1(n10690), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11012), .ZN(
        n11013) );
  NAND2_X1 U13877 ( .A1(n11014), .A2(n11013), .ZN(n11016) );
  XNOR2_X1 U13878 ( .A(n11033), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15917) );
  NAND2_X1 U13879 ( .A1(n15917), .A2(n13622), .ZN(n11015) );
  NAND2_X1 U13880 ( .A1(n11016), .A2(n11015), .ZN(n13785) );
  NOR2_X1 U13881 ( .A1(n11018), .A2(n11017), .ZN(n11042) );
  AOI22_X1 U13882 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U13883 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U13884 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U13885 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11019) );
  NAND4_X1 U13886 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(
        n11028) );
  AOI22_X1 U13887 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13888 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13889 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U13890 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11023) );
  NAND4_X1 U13891 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n11027) );
  OR2_X1 U13892 ( .A1(n11028), .A2(n11027), .ZN(n11041) );
  INV_X1 U13893 ( .A(n11041), .ZN(n11029) );
  XNOR2_X1 U13894 ( .A(n11042), .B(n11029), .ZN(n11030) );
  NAND2_X1 U13895 ( .A1(n11030), .A2(n11144), .ZN(n11040) );
  NAND2_X1 U13896 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U13897 ( .A1(n10823), .A2(n11031), .ZN(n11032) );
  AOI21_X1 U13898 ( .B1(n10690), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11032), .ZN(
        n11039) );
  INV_X1 U13899 ( .A(n11035), .ZN(n11036) );
  INV_X1 U13900 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U13901 ( .A1(n11036), .A2(n13729), .ZN(n11037) );
  NAND2_X1 U13902 ( .A1(n11075), .A2(n11037), .ZN(n13975) );
  NOR2_X1 U13903 ( .A1(n13975), .A2(n10823), .ZN(n11038) );
  AOI21_X1 U13904 ( .B1(n11040), .B2(n11039), .A(n11038), .ZN(n13723) );
  AND2_X2 U13905 ( .A1(n13720), .A2(n13723), .ZN(n13707) );
  NAND2_X1 U13906 ( .A1(n11042), .A2(n11041), .ZN(n11059) );
  AOI22_X1 U13907 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13908 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13909 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U13910 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11043) );
  NAND4_X1 U13911 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11052) );
  AOI22_X1 U13912 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10441), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U13913 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U13914 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13915 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11047) );
  NAND4_X1 U13916 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(
        n11051) );
  NOR2_X1 U13917 ( .A1(n11052), .A2(n11051), .ZN(n11060) );
  XOR2_X1 U13918 ( .A(n11059), .B(n11060), .Z(n11053) );
  NAND2_X1 U13919 ( .A1(n11053), .A2(n11144), .ZN(n11058) );
  NAND2_X1 U13920 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U13921 ( .A1(n10823), .A2(n11054), .ZN(n11055) );
  AOI21_X1 U13922 ( .B1(n10690), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11055), .ZN(
        n11057) );
  XNOR2_X1 U13923 ( .A(n11075), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13967) );
  AOI21_X1 U13924 ( .B1(n11058), .B2(n11057), .A(n11056), .ZN(n13708) );
  NOR2_X1 U13925 ( .A1(n11060), .A2(n11059), .ZN(n11083) );
  AOI22_X1 U13926 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U13927 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U13928 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U13929 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11061) );
  NAND4_X1 U13930 ( .A1(n11064), .A2(n11063), .A3(n11062), .A4(n11061), .ZN(
        n11070) );
  AOI22_X1 U13931 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U13932 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U13933 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13934 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U13935 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11069) );
  OR2_X1 U13936 ( .A1(n11070), .A2(n11069), .ZN(n11082) );
  INV_X1 U13937 ( .A(n11082), .ZN(n11071) );
  XNOR2_X1 U13938 ( .A(n11083), .B(n11071), .ZN(n11074) );
  INV_X1 U13939 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13867) );
  NAND2_X1 U13940 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11072) );
  OAI211_X1 U13941 ( .C1(n11118), .C2(n13867), .A(n10823), .B(n11072), .ZN(
        n11073) );
  AOI21_X1 U13942 ( .B1(n11074), .B2(n11144), .A(n11073), .ZN(n11081) );
  INV_X1 U13943 ( .A(n11075), .ZN(n11076) );
  INV_X1 U13944 ( .A(n11077), .ZN(n11078) );
  INV_X1 U13945 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U13946 ( .A1(n11078), .A2(n13698), .ZN(n11079) );
  NAND2_X1 U13947 ( .A1(n11121), .A2(n11079), .ZN(n13960) );
  NOR2_X1 U13948 ( .A1(n13960), .A2(n10823), .ZN(n11080) );
  NAND2_X1 U13949 ( .A1(n11083), .A2(n11082), .ZN(n11103) );
  AOI22_X1 U13950 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10441), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U13951 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11084), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U13952 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U13953 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11095) );
  AOI22_X1 U13954 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11089), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U13955 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U13956 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U13957 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11090) );
  NAND4_X1 U13958 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11090), .ZN(
        n11094) );
  NOR2_X1 U13959 ( .A1(n11095), .A2(n11094), .ZN(n11104) );
  XOR2_X1 U13960 ( .A(n11103), .B(n11104), .Z(n11096) );
  NAND2_X1 U13961 ( .A1(n11096), .A2(n11144), .ZN(n11100) );
  NAND2_X1 U13962 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U13963 ( .A1(n10823), .A2(n11097), .ZN(n11098) );
  AOI21_X1 U13964 ( .B1(n10690), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11098), .ZN(
        n11099) );
  NAND2_X1 U13965 ( .A1(n11100), .A2(n11099), .ZN(n11102) );
  XNOR2_X1 U13966 ( .A(n11121), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13950) );
  NAND2_X1 U13967 ( .A1(n13950), .A2(n13622), .ZN(n11101) );
  NAND2_X1 U13968 ( .A1(n11102), .A2(n11101), .ZN(n13686) );
  NOR2_X1 U13969 ( .A1(n11104), .A2(n11103), .ZN(n11129) );
  AOI22_X1 U13970 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U13971 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U13972 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U13973 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11106) );
  NAND4_X1 U13974 ( .A1(n11109), .A2(n11108), .A3(n11107), .A4(n11106), .ZN(
        n11115) );
  AOI22_X1 U13975 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U13976 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U13977 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U13978 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11110) );
  NAND4_X1 U13979 ( .A1(n11113), .A2(n11112), .A3(n11111), .A4(n11110), .ZN(
        n11114) );
  OR2_X1 U13980 ( .A1(n11115), .A2(n11114), .ZN(n11128) );
  INV_X1 U13981 ( .A(n11128), .ZN(n11116) );
  XNOR2_X1 U13982 ( .A(n11129), .B(n11116), .ZN(n11120) );
  INV_X1 U13983 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13858) );
  NAND2_X1 U13984 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11117) );
  OAI211_X1 U13985 ( .C1(n11118), .C2(n13858), .A(n10823), .B(n11117), .ZN(
        n11119) );
  AOI21_X1 U13986 ( .B1(n11120), .B2(n11144), .A(n11119), .ZN(n11126) );
  INV_X1 U13987 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13952) );
  INV_X1 U13988 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U13989 ( .A1(n11123), .A2(n11122), .ZN(n11124) );
  NAND2_X1 U13990 ( .A1(n12623), .A2(n11124), .ZN(n13942) );
  NOR2_X1 U13991 ( .A1(n13942), .A2(n10823), .ZN(n11125) );
  INV_X1 U13992 ( .A(n13670), .ZN(n11127) );
  NAND2_X1 U13993 ( .A1(n11129), .A2(n11128), .ZN(n13618) );
  AOI22_X1 U13994 ( .A1(n10436), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10314), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U13995 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U13996 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10474), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U13997 ( .A1(n10420), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11132) );
  NAND4_X1 U13998 ( .A1(n11135), .A2(n11134), .A3(n11133), .A4(n11132), .ZN(
        n11143) );
  AOI22_X1 U13999 ( .A1(n10988), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14000 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14001 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14002 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11138) );
  NAND4_X1 U14003 ( .A1(n11141), .A2(n11140), .A3(n11139), .A4(n11138), .ZN(
        n11142) );
  NOR2_X1 U14004 ( .A1(n11143), .A2(n11142), .ZN(n13619) );
  XOR2_X1 U14005 ( .A(n13618), .B(n13619), .Z(n11145) );
  NAND2_X1 U14006 ( .A1(n11145), .A2(n11144), .ZN(n11150) );
  NAND2_X1 U14007 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14008 ( .A1(n10823), .A2(n11146), .ZN(n11147) );
  AOI21_X1 U14009 ( .B1(n10690), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11147), .ZN(
        n11149) );
  XNOR2_X1 U14010 ( .A(n12623), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13663) );
  NAND3_X1 U14011 ( .A1(n20650), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16178) );
  INV_X1 U14012 ( .A(n16178), .ZN(n11153) );
  NOR2_X2 U14013 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20510) );
  INV_X1 U14014 ( .A(n20510), .ZN(n20587) );
  NAND2_X1 U14015 ( .A1(n20587), .A2(n11156), .ZN(n20740) );
  NAND2_X1 U14016 ( .A1(n20740), .A2(n20650), .ZN(n11154) );
  NAND2_X1 U14017 ( .A1(n20650), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15888) );
  NAND2_X1 U14018 ( .A1(n20542), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11155) );
  AND2_X1 U14019 ( .A1(n15888), .A2(n11155), .ZN(n12222) );
  INV_X1 U14020 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11157) );
  INV_X2 U14021 ( .A(n20068), .ZN(n20021) );
  NAND2_X1 U14022 ( .A1(n20021), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U14023 ( .B1(n14062), .B2(n11157), .A(n14110), .ZN(n11158) );
  AOI21_X1 U14024 ( .B1(n13663), .B2(n16064), .A(n11158), .ZN(n11159) );
  NAND2_X1 U14025 ( .A1(n11162), .A2(n11161), .ZN(P1_U2970) );
  NOR4_X1 U14026 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11166) );
  NOR4_X1 U14027 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n11165) );
  NOR4_X1 U14028 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11164) );
  NOR4_X1 U14029 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11163) );
  AND4_X1 U14030 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n11171) );
  NOR4_X1 U14031 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n11169) );
  NOR4_X1 U14032 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n11168) );
  NOR4_X1 U14033 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n11167) );
  INV_X1 U14034 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20674) );
  AND4_X1 U14035 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n20674), .ZN(
        n11170) );
  NAND2_X1 U14036 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  AND2_X2 U14037 ( .A1(n11172), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20095)
         );
  INV_X1 U14038 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20737) );
  NOR3_X1 U14039 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20737), .ZN(n11174) );
  NOR4_X1 U14040 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n11173) );
  NAND4_X1 U14041 ( .A1(n20095), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n11174), .A4(
        n11173), .ZN(U214) );
  NOR4_X1 U14042 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n11178) );
  NOR4_X1 U14043 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n11177) );
  NOR4_X1 U14044 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11176) );
  NOR4_X1 U14045 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11175) );
  NAND4_X1 U14046 ( .A1(n11178), .A2(n11177), .A3(n11176), .A4(n11175), .ZN(
        n11183) );
  NOR4_X1 U14047 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n11181) );
  NOR4_X1 U14048 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n11180) );
  NOR4_X1 U14049 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n11179) );
  INV_X1 U14050 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19744) );
  NAND4_X1 U14051 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n19744), .ZN(
        n11182) );
  OAI21_X1 U14052 ( .B1(n11183), .B2(n11182), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11184) );
  NOR2_X1 U14053 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .ZN(n11186) );
  NOR4_X1 U14054 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n11185) );
  NAND4_X1 U14055 ( .A1(n11186), .A2(P2_W_R_N_REG_SCAN_IN), .A3(
        P2_M_IO_N_REG_SCAN_IN), .A4(n11185), .ZN(n11802) );
  NOR2_X1 U14056 ( .A1(n13481), .A2(n11802), .ZN(n16516) );
  NAND2_X1 U14057 ( .A1(n16516), .A2(U214), .ZN(U212) );
  INV_X1 U14058 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13278) );
  AND2_X4 U14059 ( .A1(n15461), .A2(n15449), .ZN(n11388) );
  AND3_X4 U14060 ( .A1(n11550), .A2(n15449), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14061 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11189) );
  INV_X2 U14062 ( .A(n13242), .ZN(n11260) );
  AOI22_X1 U14063 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11188) );
  AND2_X4 U14064 ( .A1(n12304), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13426) );
  AOI22_X1 U14065 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11187) );
  NAND4_X1 U14066 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11191) );
  AOI22_X1 U14067 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14068 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14069 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11192) );
  NAND4_X1 U14070 ( .A1(n11195), .A2(n11194), .A3(n11193), .A4(n11192), .ZN(
        n11196) );
  AOI22_X1 U14071 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14072 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14073 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11198) );
  INV_X2 U14074 ( .A(n13249), .ZN(n13383) );
  AOI22_X1 U14075 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11197) );
  NAND4_X1 U14076 ( .A1(n11200), .A2(n11199), .A3(n11198), .A4(n11197), .ZN(
        n11201) );
  AOI22_X1 U14077 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14078 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14079 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14080 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11202) );
  NAND4_X1 U14081 ( .A1(n11205), .A2(n11204), .A3(n11203), .A4(n11202), .ZN(
        n11206) );
  NAND2_X1 U14082 ( .A1(n11206), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11207) );
  AOI22_X1 U14083 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14084 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14085 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14086 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14087 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  NAND2_X1 U14088 ( .A1(n11213), .A2(n11392), .ZN(n11220) );
  AOI22_X1 U14089 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14090 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14091 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14092 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14093 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  AOI22_X1 U14094 ( .A1(n11383), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11388), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14095 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14096 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14097 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11221) );
  NAND4_X1 U14098 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .ZN(
        n11225) );
  AOI22_X1 U14099 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14100 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14101 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11226) );
  NAND4_X1 U14102 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n11226), .ZN(
        n11230) );
  NAND2_X2 U14103 ( .A1(n11232), .A2(n11231), .ZN(n11297) );
  AOI22_X1 U14104 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11237) );
  AOI22_X1 U14105 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9607), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14106 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14107 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11234) );
  NAND4_X1 U14108 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(
        n11238) );
  AOI22_X1 U14109 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14110 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14111 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14112 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U14113 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11243) );
  AOI22_X1 U14114 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14115 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14116 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14117 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11244) );
  NAND4_X1 U14118 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11248) );
  NAND2_X1 U14119 ( .A1(n11248), .A2(n11392), .ZN(n11255) );
  AOI22_X1 U14120 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14121 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14122 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14123 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11249) );
  NAND4_X1 U14124 ( .A1(n11252), .A2(n11251), .A3(n11250), .A4(n11249), .ZN(
        n11253) );
  NAND2_X1 U14125 ( .A1(n11253), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11254) );
  AOI22_X1 U14126 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14127 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14128 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14129 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14130 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14131 ( .A1(n13417), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14132 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14133 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14134 ( .A1(n11616), .A2(n11280), .ZN(n11287) );
  NAND2_X1 U14135 ( .A1(n11701), .A2(n11297), .ZN(n11265) );
  AOI22_X1 U14136 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14137 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14138 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14139 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14140 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14141 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13332), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14142 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14143 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11270) );
  NAND2_X1 U14144 ( .A1(n11301), .A2(n12046), .ZN(n11274) );
  NAND3_X1 U14145 ( .A1(n11277), .A2(n11276), .A3(n11275), .ZN(n11278) );
  NAND3_X1 U14146 ( .A1(n11700), .A2(n15543), .A3(n9603), .ZN(n11283) );
  NOR2_X1 U14147 ( .A1(n15537), .A2(n11297), .ZN(n11284) );
  NAND2_X1 U14148 ( .A1(n12047), .A2(n11286), .ZN(n11321) );
  INV_X1 U14149 ( .A(n11287), .ZN(n11767) );
  NAND2_X1 U14150 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11289) );
  MUX2_X1 U14151 ( .A(n15494), .B(n9603), .S(n15543), .Z(n11295) );
  NAND2_X1 U14152 ( .A1(n11293), .A2(n15494), .ZN(n11298) );
  AND2_X1 U14153 ( .A1(n11298), .A2(n12046), .ZN(n11294) );
  NAND3_X1 U14154 ( .A1(n11296), .A2(n11295), .A3(n11294), .ZN(n11300) );
  NAND4_X1 U14155 ( .A1(n11299), .A2(n9887), .A3(n11310), .A4(n9603), .ZN(
        n11607) );
  INV_X1 U14156 ( .A(n11302), .ZN(n11304) );
  INV_X1 U14157 ( .A(n11616), .ZN(n11604) );
  NAND3_X1 U14158 ( .A1(n16407), .A2(n12046), .A3(n15526), .ZN(n11311) );
  AOI22_X1 U14159 ( .A1(n12306), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16426), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11312) );
  INV_X1 U14160 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U14161 ( .A1(n11330), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11316) );
  AND2_X1 U14162 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11314) );
  NOR2_X1 U14163 ( .A1(n16426), .A2(n11314), .ZN(n11315) );
  OAI211_X1 U14164 ( .C1(n9605), .C2(n11317), .A(n11316), .B(n11315), .ZN(
        n11318) );
  NOR2_X1 U14165 ( .A1(n11318), .A2(n11326), .ZN(n11320) );
  INV_X1 U14166 ( .A(n16426), .ZN(n14299) );
  NAND2_X1 U14167 ( .A1(n11326), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11324) );
  NAND2_X1 U14168 ( .A1(n11322), .A2(n11321), .ZN(n12311) );
  NAND2_X1 U14169 ( .A1(n12311), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11323) );
  AOI21_X1 U14170 ( .B1(n16435), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11327) );
  INV_X1 U14171 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U14172 ( .A1(n14307), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14173 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11331) );
  INV_X1 U14174 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U14175 ( .A1(n14307), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U14176 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11337) );
  OAI211_X1 U14177 ( .C1(n13534), .C2(n14542), .A(n11338), .B(n11337), .ZN(
        n11339) );
  INV_X1 U14178 ( .A(n11339), .ZN(n11340) );
  AND2_X1 U14179 ( .A1(n16426), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11342) );
  INV_X1 U14180 ( .A(n11345), .ZN(n11365) );
  INV_X1 U14181 ( .A(n11352), .ZN(n11346) );
  NAND2_X1 U14182 ( .A1(n11365), .A2(n11346), .ZN(n11347) );
  INV_X1 U14183 ( .A(n11348), .ZN(n11351) );
  INV_X1 U14184 ( .A(n11349), .ZN(n11350) );
  INV_X1 U14185 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11353) );
  OAI22_X1 U14186 ( .A1(n13278), .A2(n19554), .B1(n11478), .B2(n11353), .ZN(
        n11359) );
  INV_X1 U14187 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13277) );
  INV_X1 U14188 ( .A(n11366), .ZN(n11354) );
  INV_X1 U14189 ( .A(n16368), .ZN(n12120) );
  INV_X1 U14190 ( .A(n11355), .ZN(n11356) );
  OR2_X1 U14191 ( .A1(n11344), .A2(n11356), .ZN(n11375) );
  INV_X1 U14192 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n19526) );
  OAI22_X1 U14193 ( .A1(n13277), .A2(n19609), .B1(n12825), .B2(n19526), .ZN(
        n11358) );
  INV_X1 U14194 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11361) );
  INV_X1 U14195 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11360) );
  OAI22_X1 U14196 ( .A1(n11361), .A2(n15480), .B1(n19502), .B2(n11360), .ZN(
        n11362) );
  INV_X1 U14197 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13268) );
  INV_X1 U14198 ( .A(n12299), .ZN(n11363) );
  INV_X1 U14199 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13276) );
  OAI22_X1 U14200 ( .A1(n13268), .A2(n19397), .B1(n19648), .B2(n13276), .ZN(
        n11364) );
  INV_X1 U14201 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13269) );
  OR2_X2 U14202 ( .A1(n11372), .A2(n11373), .ZN(n19365) );
  NAND2_X1 U14203 ( .A1(n11365), .A2(n16368), .ZN(n11376) );
  INV_X1 U14204 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11367) );
  OAI22_X1 U14205 ( .A1(n13269), .A2(n19365), .B1(n12813), .B2(n11367), .ZN(
        n11371) );
  INV_X1 U14206 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13270) );
  OR2_X2 U14207 ( .A1(n11372), .A2(n11368), .ZN(n19307) );
  INV_X1 U14208 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12343) );
  OAI22_X1 U14209 ( .A1(n13270), .A2(n19307), .B1(n19460), .B2(n12343), .ZN(
        n11370) );
  NOR2_X1 U14210 ( .A1(n11371), .A2(n11370), .ZN(n11382) );
  INV_X1 U14211 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U14212 ( .A1(n15503), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11374) );
  OAI211_X1 U14213 ( .C1(n13121), .C2(n19341), .A(n11374), .B(n15526), .ZN(
        n11380) );
  INV_X1 U14214 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15530) );
  OR2_X2 U14215 ( .A1(n11377), .A2(n11375), .ZN(n15516) );
  INV_X1 U14216 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11378) );
  OAI22_X1 U14217 ( .A1(n15530), .A2(n15516), .B1(n19258), .B2(n11378), .ZN(
        n11379) );
  NOR2_X1 U14218 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  NAND2_X1 U14219 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U14220 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11386) );
  NAND3_X1 U14221 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11587) );
  INV_X1 U14222 ( .A(n11587), .ZN(n11384) );
  NAND2_X1 U14223 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11384), .ZN(
        n12722) );
  NOR4_X2 U14224 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U14225 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n13229), .ZN(n11385) );
  NAND2_X1 U14226 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U14227 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11389) );
  NAND4_X1 U14228 ( .A1(n9671), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(
        n11398) );
  AND2_X2 U14229 ( .A1(n13382), .A2(n11392), .ZN(n13223) );
  AND2_X2 U14230 ( .A1(n13382), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12594) );
  AOI22_X1 U14231 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11396) );
  AND2_X2 U14232 ( .A1(n9599), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12592) );
  AND2_X2 U14233 ( .A1(n13383), .A2(n11392), .ZN(n13235) );
  AOI22_X1 U14234 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__0__SCAN_IN), .B2(n13235), .ZN(n11395) );
  AOI22_X1 U14235 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14236 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12600), .B1(
        n12599), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11393) );
  NAND4_X1 U14237 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n11397) );
  AND2_X1 U14238 ( .A1(n11721), .A2(n16421), .ZN(n12088) );
  NAND2_X1 U14239 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11401) );
  NAND2_X1 U14240 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11400) );
  AOI22_X1 U14241 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14242 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12604), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U14243 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14244 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11403) );
  NAND4_X1 U14245 ( .A1(n10233), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11411) );
  AOI22_X1 U14246 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14247 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14248 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14249 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11406) );
  NAND4_X1 U14250 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11410) );
  NAND2_X1 U14251 ( .A1(n12088), .A2(n11729), .ZN(n11456) );
  NAND2_X1 U14252 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11414) );
  NAND2_X1 U14253 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11413) );
  AOI22_X1 U14254 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11412) );
  INV_X1 U14255 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U14256 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12604), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14257 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11417) );
  NAND2_X1 U14258 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11416) );
  NAND4_X1 U14259 ( .A1(n10226), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11424) );
  AOI22_X1 U14260 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14261 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14262 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14263 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11419) );
  NAND4_X1 U14264 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(
        n11423) );
  INV_X1 U14265 ( .A(n11736), .ZN(n11455) );
  NAND2_X1 U14266 ( .A1(n11456), .A2(n11455), .ZN(n11425) );
  INV_X1 U14267 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13320) );
  INV_X1 U14268 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13152) );
  OAI22_X1 U14269 ( .A1(n13320), .A2(n19307), .B1(n19502), .B2(n13152), .ZN(
        n11427) );
  INV_X1 U14270 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13318) );
  INV_X1 U14271 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12593) );
  OAI22_X1 U14272 ( .A1(n13318), .A2(n19397), .B1(n11478), .B2(n12593), .ZN(
        n11426) );
  NOR2_X1 U14273 ( .A1(n11427), .A2(n11426), .ZN(n11439) );
  INV_X1 U14274 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13319) );
  INV_X1 U14275 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13149) );
  OAI22_X1 U14276 ( .A1(n13319), .A2(n19365), .B1(n19341), .B2(n13149), .ZN(
        n11429) );
  INV_X1 U14277 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12601) );
  INV_X1 U14278 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13158) );
  OAI22_X1 U14279 ( .A1(n12601), .A2(n12813), .B1(n19460), .B2(n13158), .ZN(
        n11428) );
  INV_X1 U14280 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13327) );
  INV_X1 U14281 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13326) );
  OAI22_X1 U14282 ( .A1(n13327), .A2(n12825), .B1(n19648), .B2(n13326), .ZN(
        n11432) );
  INV_X1 U14283 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11430) );
  INV_X1 U14284 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13329) );
  OAI22_X1 U14285 ( .A1(n11430), .A2(n19258), .B1(n19554), .B2(n13329), .ZN(
        n11431) );
  NOR2_X1 U14286 ( .A1(n11432), .A2(n11431), .ZN(n11437) );
  INV_X1 U14287 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11433) );
  INV_X1 U14288 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15541) );
  INV_X1 U14289 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13328) );
  OAI22_X1 U14290 ( .A1(n15541), .A2(n15516), .B1(n19609), .B2(n13328), .ZN(
        n11434) );
  NOR2_X1 U14291 ( .A1(n11435), .A2(n11434), .ZN(n11436) );
  AOI22_X1 U14292 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13223), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14293 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14294 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14295 ( .A1(n12598), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11440) );
  NAND4_X1 U14296 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11449) );
  AOI22_X1 U14297 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14298 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13230), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14299 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14300 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11444) );
  NAND4_X1 U14301 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11448) );
  INV_X1 U14302 ( .A(n11743), .ZN(n11450) );
  NAND2_X1 U14303 ( .A1(n11450), .A2(n16421), .ZN(n11451) );
  INV_X1 U14304 ( .A(n12088), .ZN(n11452) );
  NAND2_X1 U14305 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12090) );
  XNOR2_X1 U14306 ( .A(n11721), .B(n11729), .ZN(n11453) );
  NOR2_X1 U14307 ( .A1(n12090), .A2(n11453), .ZN(n11454) );
  INV_X1 U14308 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12786) );
  XNOR2_X1 U14309 ( .A(n12090), .B(n11453), .ZN(n12073) );
  NOR2_X1 U14310 ( .A1(n12786), .A2(n12073), .ZN(n12072) );
  NOR2_X1 U14311 ( .A1(n11454), .A2(n12072), .ZN(n11457) );
  XNOR2_X1 U14312 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11457), .ZN(
        n12036) );
  XNOR2_X1 U14313 ( .A(n11456), .B(n11455), .ZN(n12035) );
  NAND2_X1 U14314 ( .A1(n12036), .A2(n12035), .ZN(n12034) );
  INV_X1 U14315 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12027) );
  OR2_X1 U14316 ( .A1(n11457), .A2(n12027), .ZN(n11458) );
  NAND2_X1 U14317 ( .A1(n12034), .A2(n11458), .ZN(n11459) );
  XNOR2_X1 U14318 ( .A(n11459), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12774) );
  NAND2_X1 U14319 ( .A1(n11459), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11460) );
  AOI22_X1 U14320 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14321 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14322 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14323 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14324 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11472) );
  NAND2_X1 U14325 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U14326 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11466) );
  AOI22_X1 U14327 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11465) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19483) );
  AOI22_X1 U14329 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14330 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U14331 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11468) );
  NAND4_X1 U14332 ( .A1(n10225), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11471) );
  NOR2_X1 U14333 ( .A1(n11472), .A2(n11471), .ZN(n11668) );
  INV_X1 U14334 ( .A(n11668), .ZN(n11748) );
  NAND2_X1 U14335 ( .A1(n11508), .A2(n11473), .ZN(n11474) );
  INV_X1 U14336 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15118) );
  INV_X1 U14337 ( .A(n11474), .ZN(n11476) );
  NOR2_X1 U14338 ( .A1(n11476), .A2(n11475), .ZN(n11477) );
  AOI21_X2 U14339 ( .B1(n15119), .B2(n15118), .A(n11477), .ZN(n16301) );
  INV_X1 U14340 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12739) );
  OAI22_X1 U14341 ( .A1(n19588), .A2(n12813), .B1(n19460), .B2(n12739), .ZN(
        n11481) );
  INV_X1 U14342 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13367) );
  INV_X1 U14343 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11479) );
  OAI22_X1 U14344 ( .A1(n13367), .A2(n19397), .B1(n11478), .B2(n11479), .ZN(
        n11480) );
  NOR2_X1 U14345 ( .A1(n11481), .A2(n11480), .ZN(n11493) );
  INV_X1 U14346 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12490) );
  INV_X1 U14347 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11482) );
  OAI22_X1 U14348 ( .A1(n12490), .A2(n15480), .B1(n11523), .B2(n11482), .ZN(
        n11485) );
  INV_X1 U14349 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11483) );
  INV_X1 U14350 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13376) );
  OAI22_X1 U14351 ( .A1(n11483), .A2(n19258), .B1(n12825), .B2(n13376), .ZN(
        n11484) );
  NOR2_X1 U14352 ( .A1(n11485), .A2(n11484), .ZN(n11492) );
  INV_X1 U14353 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13368) );
  INV_X1 U14354 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13193) );
  OAI22_X1 U14355 ( .A1(n13368), .A2(n19365), .B1(n19341), .B2(n13193), .ZN(
        n11487) );
  INV_X1 U14356 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13369) );
  INV_X1 U14357 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13196) );
  NOR2_X1 U14358 ( .A1(n11487), .A2(n11486), .ZN(n11491) );
  INV_X1 U14359 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13379) );
  INV_X1 U14360 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13375) );
  OAI22_X1 U14361 ( .A1(n13379), .A2(n19554), .B1(n19648), .B2(n13375), .ZN(
        n11489) );
  INV_X1 U14362 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15552) );
  INV_X1 U14363 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13377) );
  OAI22_X1 U14364 ( .A1(n15552), .A2(n15516), .B1(n19609), .B2(n13377), .ZN(
        n11488) );
  NOR2_X1 U14365 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  NAND4_X1 U14366 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11507) );
  AOI22_X1 U14367 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14368 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14369 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14370 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11494) );
  NAND4_X1 U14371 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n11505) );
  NAND2_X1 U14372 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14373 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11499) );
  AOI22_X1 U14374 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14375 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14376 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14377 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11501) );
  NAND4_X1 U14378 ( .A1(n10223), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11504) );
  NAND2_X1 U14379 ( .A1(n11752), .A2(n16421), .ZN(n11506) );
  OR2_X1 U14380 ( .A1(n11677), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16298) );
  NAND2_X1 U14381 ( .A1(n16301), .A2(n16298), .ZN(n11544) );
  NAND2_X1 U14382 ( .A1(n11677), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16299) );
  INV_X1 U14383 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13210) );
  INV_X1 U14384 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11510) );
  OAI22_X1 U14385 ( .A1(n13210), .A2(n19341), .B1(n19365), .B2(n11510), .ZN(
        n11514) );
  INV_X1 U14386 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11512) );
  INV_X1 U14387 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11511) );
  OAI22_X1 U14388 ( .A1(n11512), .A2(n19307), .B1(n12813), .B2(n11511), .ZN(
        n11513) );
  NOR2_X1 U14389 ( .A1(n11514), .A2(n11513), .ZN(n11529) );
  INV_X1 U14390 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13397) );
  INV_X1 U14391 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11515) );
  OAI22_X1 U14392 ( .A1(n13397), .A2(n19648), .B1(n19554), .B2(n11515), .ZN(
        n11518) );
  INV_X1 U14393 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15557) );
  INV_X1 U14394 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11516) );
  OAI22_X1 U14395 ( .A1(n15557), .A2(n15516), .B1(n19609), .B2(n11516), .ZN(
        n11517) );
  NOR2_X1 U14396 ( .A1(n11518), .A2(n11517), .ZN(n11528) );
  INV_X1 U14397 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13395) );
  INV_X1 U14398 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11519) );
  OAI22_X1 U14399 ( .A1(n13395), .A2(n19502), .B1(n19460), .B2(n11519), .ZN(
        n11521) );
  INV_X1 U14400 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13389) );
  INV_X1 U14401 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13396) );
  OAI22_X1 U14402 ( .A1(n13389), .A2(n19397), .B1(n11478), .B2(n13396), .ZN(
        n11520) );
  NOR2_X1 U14403 ( .A1(n11521), .A2(n11520), .ZN(n11527) );
  INV_X1 U14404 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15497) );
  INV_X1 U14405 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11522) );
  OAI22_X1 U14406 ( .A1(n15497), .A2(n15480), .B1(n11523), .B2(n11522), .ZN(
        n11525) );
  INV_X1 U14407 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12721) );
  INV_X1 U14408 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13399) );
  OAI22_X1 U14409 ( .A1(n12721), .A2(n19258), .B1(n12825), .B2(n13399), .ZN(
        n11524) );
  NOR2_X1 U14410 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  NAND4_X1 U14411 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11543) );
  AOI22_X1 U14412 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12594), .B1(
        n13223), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14413 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n13235), .ZN(n11532) );
  AOI22_X1 U14414 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14415 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12600), .B1(
        n12599), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14416 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11541) );
  NAND2_X1 U14417 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14418 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11535) );
  AOI22_X1 U14419 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13229), .ZN(n11534) );
  AOI22_X1 U14420 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14421 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U14422 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11537) );
  NAND4_X1 U14423 ( .A1(n10222), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11540) );
  NAND2_X1 U14424 ( .A1(n11758), .A2(n16421), .ZN(n11542) );
  INV_X1 U14425 ( .A(n11544), .ZN(n11545) );
  XNOR2_X1 U14426 ( .A(n14900), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16288) );
  NAND2_X1 U14427 ( .A1(n15450), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14428 ( .A1(n11550), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U14429 ( .A1(n11554), .A2(n11551), .ZN(n11558) );
  INV_X1 U14430 ( .A(n11558), .ZN(n11552) );
  MUX2_X1 U14431 ( .A(n19809), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11572) );
  INV_X1 U14432 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15911) );
  NOR2_X1 U14433 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15911), .ZN(
        n11555) );
  INV_X1 U14434 ( .A(n11579), .ZN(n11594) );
  INV_X1 U14435 ( .A(n19149), .ZN(n11557) );
  NAND2_X1 U14436 ( .A1(n11557), .A2(n15526), .ZN(n11562) );
  NAND2_X1 U14437 ( .A1(n11559), .A2(n11558), .ZN(n11561) );
  MUX2_X1 U14438 ( .A(n11562), .B(n11646), .S(n11590), .Z(n11570) );
  INV_X1 U14439 ( .A(n11590), .ZN(n11568) );
  OAI21_X1 U14440 ( .B1(n19836), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11563), .ZN(n11597) );
  INV_X1 U14441 ( .A(n11646), .ZN(n12792) );
  OAI21_X1 U14442 ( .B1(n11597), .B2(n11584), .A(n12792), .ZN(n11567) );
  INV_X1 U14443 ( .A(n11597), .ZN(n11565) );
  INV_X1 U14444 ( .A(n11563), .ZN(n11564) );
  XNOR2_X1 U14445 ( .A(n11584), .B(n11564), .ZN(n11593) );
  OAI211_X1 U14446 ( .C1(n15526), .C2(n11565), .A(n16408), .B(n11593), .ZN(
        n11566) );
  OAI211_X1 U14447 ( .C1(n12044), .C2(n11568), .A(n11567), .B(n11566), .ZN(
        n11569) );
  NAND2_X1 U14448 ( .A1(n11570), .A2(n11569), .ZN(n11576) );
  NOR2_X1 U14449 ( .A1(n11573), .A2(n11572), .ZN(n11574) );
  MUX2_X1 U14450 ( .A(n11646), .B(n11576), .S(n11591), .Z(n11577) );
  NAND2_X1 U14451 ( .A1(n11594), .A2(n11577), .ZN(n11578) );
  MUX2_X1 U14452 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11578), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11581) );
  NAND2_X1 U14453 ( .A1(n11579), .A2(n19149), .ZN(n11580) );
  NOR2_X1 U14454 ( .A1(n16401), .A2(n16421), .ZN(n12317) );
  NAND2_X1 U14455 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19714) );
  INV_X1 U14456 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18949) );
  NOR2_X1 U14457 ( .A1(n20815), .A2(n18949), .ZN(n19734) );
  NOR2_X1 U14458 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19721) );
  NOR3_X1 U14459 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19734), .A3(n19721), 
        .ZN(n19726) );
  NAND2_X1 U14460 ( .A1(n19714), .A2(n19726), .ZN(n12784) );
  INV_X1 U14461 ( .A(n12784), .ZN(n11926) );
  NAND3_X1 U14462 ( .A1(n12317), .A2(n11297), .A3(n11926), .ZN(n11621) );
  INV_X1 U14463 ( .A(n12317), .ZN(n11583) );
  AOI21_X1 U14464 ( .B1(n11581), .B2(n16408), .A(n11701), .ZN(n11582) );
  NAND2_X1 U14465 ( .A1(n11583), .A2(n11582), .ZN(n11620) );
  NOR2_X1 U14466 ( .A1(n11584), .A2(n11597), .ZN(n11585) );
  MUX2_X1 U14467 ( .A(n11736), .B(n11590), .S(n11646), .Z(n11644) );
  OAI21_X1 U14468 ( .B1(n11585), .B2(n11644), .A(n11591), .ZN(n11586) );
  NAND2_X1 U14469 ( .A1(n11586), .A2(n11594), .ZN(n19840) );
  INV_X1 U14470 ( .A(n16407), .ZN(n11690) );
  AND2_X1 U14471 ( .A1(n11280), .A2(n16421), .ZN(n11609) );
  NAND2_X1 U14472 ( .A1(n11690), .A2(n11609), .ZN(n11623) );
  AND2_X1 U14473 ( .A1(n11588), .A2(n11587), .ZN(n15472) );
  INV_X1 U14474 ( .A(n15472), .ZN(n16403) );
  INV_X1 U14475 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11589) );
  OAI21_X1 U14476 ( .B1(n12592), .B2(n16403), .A(n11589), .ZN(n19828) );
  NAND2_X1 U14477 ( .A1(n19828), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11601) );
  NAND2_X1 U14478 ( .A1(n11591), .A2(n11590), .ZN(n11596) );
  INV_X1 U14479 ( .A(n11596), .ZN(n11592) );
  NAND2_X1 U14480 ( .A1(n11593), .A2(n11592), .ZN(n11595) );
  OAI21_X1 U14481 ( .B1(n11597), .B2(n11596), .A(n13505), .ZN(n11598) );
  INV_X1 U14482 ( .A(n11598), .ZN(n11599) );
  NAND2_X1 U14483 ( .A1(n16395), .A2(n11599), .ZN(n11600) );
  NAND2_X1 U14484 ( .A1(n11601), .A2(n11600), .ZN(n19843) );
  NAND3_X1 U14485 ( .A1(n11690), .A2(n15526), .A3(n19843), .ZN(n11602) );
  NAND2_X1 U14486 ( .A1(n11603), .A2(n11602), .ZN(n11929) );
  MUX2_X1 U14487 ( .A(n11604), .B(n12046), .S(n16421), .Z(n11606) );
  NAND2_X1 U14488 ( .A1(n16395), .A2(n19714), .ZN(n11605) );
  NOR2_X1 U14489 ( .A1(n11606), .A2(n11605), .ZN(n11618) );
  INV_X1 U14490 ( .A(n11607), .ZN(n11608) );
  NAND2_X1 U14491 ( .A1(n11608), .A2(n16408), .ZN(n15473) );
  OAI21_X1 U14492 ( .B1(n11697), .B2(n11297), .A(n15473), .ZN(n11615) );
  INV_X1 U14493 ( .A(n9603), .ZN(n12103) );
  OAI21_X1 U14494 ( .B1(n11610), .B2(n12103), .A(n11609), .ZN(n11698) );
  NAND2_X1 U14495 ( .A1(n16421), .A2(n15543), .ZN(n11692) );
  NAND2_X1 U14496 ( .A1(n11692), .A2(n16408), .ZN(n11611) );
  NAND2_X1 U14497 ( .A1(n11611), .A2(n11307), .ZN(n11612) );
  NAND2_X1 U14498 ( .A1(n11612), .A2(n12046), .ZN(n11613) );
  AND2_X1 U14499 ( .A1(n11698), .A2(n11613), .ZN(n11614) );
  NAND3_X1 U14500 ( .A1(n11616), .A2(n16395), .A3(n11926), .ZN(n11617) );
  NAND2_X1 U14501 ( .A1(n11694), .A2(n11617), .ZN(n12318) );
  NOR3_X1 U14502 ( .A1(n11929), .A2(n11618), .A3(n12318), .ZN(n11619) );
  NAND3_X1 U14503 ( .A1(n11621), .A2(n11620), .A3(n11619), .ZN(n11622) );
  NOR2_X1 U14504 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16435), .ZN(n19713) );
  NAND2_X1 U14505 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19713), .ZN(n19146) );
  INV_X1 U14506 ( .A(n11623), .ZN(n19839) );
  NOR2_X1 U14507 ( .A1(n16288), .A2(n16383), .ZN(n11801) );
  NAND2_X1 U14508 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14509 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14510 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U14511 ( .A1(n13222), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11624) );
  INV_X1 U14512 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20845) );
  NAND2_X1 U14513 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14514 ( .A1(n13235), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11630) );
  NAND2_X1 U14515 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11629) );
  NAND2_X1 U14516 ( .A1(n12594), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U14517 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14518 ( .A1(n12598), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14519 ( .A1(n12600), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14520 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U14521 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14522 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11637) );
  AOI22_X1 U14523 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13229), .ZN(n11636) );
  AND3_X1 U14524 ( .A1(n11638), .A2(n11637), .A3(n11636), .ZN(n11639) );
  NAND4_X1 U14525 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n14343) );
  INV_X1 U14526 ( .A(n14343), .ZN(n11643) );
  INV_X2 U14527 ( .A(n11643), .ZN(n14896) );
  MUX2_X1 U14528 ( .A(n11644), .B(n11333), .S(n14828), .Z(n11654) );
  INV_X1 U14529 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14557) );
  NOR2_X1 U14530 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n11645) );
  MUX2_X1 U14531 ( .A(n11729), .B(n11645), .S(n14828), .Z(n11657) );
  AND2_X1 U14532 ( .A1(n11646), .A2(n11720), .ZN(n11670) );
  NAND2_X1 U14533 ( .A1(n11670), .A2(n11647), .ZN(n11648) );
  NAND2_X1 U14534 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  INV_X1 U14535 ( .A(n11679), .ZN(n11652) );
  NAND2_X1 U14536 ( .A1(n11656), .A2(n11650), .ZN(n11651) );
  NAND2_X1 U14537 ( .A1(n11652), .A2(n11651), .ZN(n14543) );
  OR2_X1 U14538 ( .A1(n11654), .A2(n11657), .ZN(n11655) );
  NAND2_X1 U14539 ( .A1(n11656), .A2(n11655), .ZN(n12837) );
  XNOR2_X1 U14540 ( .A(n12837), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12026) );
  INV_X1 U14541 ( .A(n11657), .ZN(n11660) );
  AND2_X1 U14542 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11658) );
  NAND2_X1 U14543 ( .A1(n14828), .A2(n11658), .ZN(n11659) );
  NAND2_X1 U14544 ( .A1(n11660), .A2(n11659), .ZN(n14553) );
  MUX2_X1 U14545 ( .A(n11721), .B(P2_EBX_REG_0__SCAN_IN), .S(n14828), .Z(
        n14566) );
  NAND2_X1 U14546 ( .A1(n14566), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12086) );
  OAI21_X1 U14547 ( .B1(n14553), .B2(n12786), .A(n12086), .ZN(n11662) );
  NAND2_X1 U14548 ( .A1(n14553), .A2(n12786), .ZN(n11661) );
  AND2_X1 U14549 ( .A1(n11662), .A2(n11661), .ZN(n12025) );
  NAND2_X1 U14550 ( .A1(n12026), .A2(n12025), .ZN(n12024) );
  INV_X1 U14551 ( .A(n12837), .ZN(n11663) );
  NAND2_X1 U14552 ( .A1(n11663), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11664) );
  AND2_X1 U14553 ( .A1(n12024), .A2(n11664), .ZN(n12765) );
  NAND2_X1 U14554 ( .A1(n12792), .A2(n11668), .ZN(n11669) );
  INV_X1 U14555 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19108) );
  MUX2_X1 U14556 ( .A(n11669), .B(n19108), .S(n14828), .Z(n11673) );
  NAND2_X1 U14557 ( .A1(n11671), .A2(n11670), .ZN(n11672) );
  XNOR2_X1 U14558 ( .A(n11679), .B(n11678), .ZN(n11674) );
  XNOR2_X1 U14559 ( .A(n11674), .B(n15118), .ZN(n15113) );
  INV_X1 U14560 ( .A(n11674), .ZN(n19105) );
  NAND2_X1 U14561 ( .A1(n19105), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11675) );
  MUX2_X1 U14562 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n11752), .S(n9590), .Z(n11680) );
  OAI21_X1 U14563 ( .B1(n11682), .B2(n11681), .A(n11687), .ZN(n14532) );
  INV_X1 U14564 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U14565 ( .A1(n11683), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11684) );
  NAND2_X1 U14566 ( .A1(n11685), .A2(n11643), .ZN(n11689) );
  MUX2_X1 U14567 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11758), .S(n11720), .Z(
        n11686) );
  NAND2_X1 U14568 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  NAND2_X1 U14569 ( .A1(n9930), .A2(n11688), .ZN(n12806) );
  XNOR2_X1 U14570 ( .A(n14783), .B(n14782), .ZN(n16286) );
  INV_X1 U14571 ( .A(n11771), .ZN(n11691) );
  NAND2_X1 U14572 ( .A1(n11690), .A2(n12792), .ZN(n19844) );
  NOR2_X1 U14573 ( .A1(n16286), .A2(n16373), .ZN(n11800) );
  NAND2_X1 U14574 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16362) );
  INV_X1 U14575 ( .A(n11692), .ZN(n11693) );
  NAND2_X1 U14576 ( .A1(n11771), .A2(n16398), .ZN(n15319) );
  NOR2_X1 U14577 ( .A1(n12786), .A2(n12087), .ZN(n11695) );
  INV_X1 U14578 ( .A(n11695), .ZN(n15435) );
  NOR2_X1 U14579 ( .A1(n12027), .A2(n15435), .ZN(n12037) );
  INV_X1 U14580 ( .A(n12037), .ZN(n11696) );
  NOR2_X1 U14581 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11695), .ZN(
        n12038) );
  AOI21_X1 U14582 ( .B1(n15319), .B2(n11696), .A(n12038), .ZN(n12773) );
  OAI21_X1 U14583 ( .B1(n11697), .B2(n12103), .A(n15526), .ZN(n15440) );
  NAND2_X1 U14584 ( .A1(n15440), .A2(n11698), .ZN(n11699) );
  NAND2_X1 U14585 ( .A1(n11699), .A2(n15537), .ZN(n11705) );
  NOR2_X1 U14586 ( .A1(n11700), .A2(n11701), .ZN(n11702) );
  NOR2_X1 U14587 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  NAND2_X1 U14588 ( .A1(n11705), .A2(n11704), .ZN(n11711) );
  MUX2_X1 U14589 ( .A(n12044), .B(n11707), .S(n11706), .Z(n11708) );
  AOI21_X1 U14590 ( .B1(n11708), .B2(n11700), .A(n15537), .ZN(n11709) );
  MUX2_X1 U14591 ( .A(n11709), .B(n11280), .S(n11297), .Z(n11710) );
  NOR2_X1 U14592 ( .A1(n11711), .A2(n11710), .ZN(n12302) );
  NAND2_X1 U14593 ( .A1(n12302), .A2(n11321), .ZN(n11712) );
  NAND2_X1 U14594 ( .A1(n11771), .A2(n11712), .ZN(n15316) );
  NAND3_X1 U14595 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12773), .A3(
        n16376), .ZN(n15421) );
  NOR2_X1 U14596 ( .A1(n16362), .A2(n15421), .ZN(n11718) );
  NAND2_X1 U14597 ( .A1(n13505), .A2(n12070), .ZN(n19801) );
  NOR2_X1 U14598 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19801), .ZN(n11713) );
  NAND2_X1 U14599 ( .A1(n11713), .A2(n16435), .ZN(n11795) );
  OR2_X1 U14600 ( .A1(n11771), .A2(n19111), .ZN(n16374) );
  INV_X1 U14601 ( .A(n12038), .ZN(n11714) );
  OR2_X1 U14602 ( .A1(n15319), .A2(n11714), .ZN(n11715) );
  OAI211_X1 U14603 ( .C1(n15316), .C2(n12037), .A(n16374), .B(n11715), .ZN(
        n12768) );
  AND2_X1 U14604 ( .A1(n16376), .A2(n11666), .ZN(n12772) );
  AOI21_X1 U14605 ( .B1(n16376), .B2(n16362), .A(n16355), .ZN(n11716) );
  INV_X1 U14606 ( .A(n11716), .ZN(n11717) );
  MUX2_X1 U14607 ( .A(n11718), .B(n11717), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n11799) );
  NOR2_X2 U14608 ( .A1(n16421), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11739) );
  INV_X1 U14609 ( .A(n11303), .ZN(n12065) );
  NAND2_X1 U14610 ( .A1(n11739), .A2(n12065), .ZN(n11734) );
  NAND2_X1 U14611 ( .A1(n12903), .A2(n11721), .ZN(n11723) );
  NAND2_X1 U14612 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14613 ( .A1(n11734), .A2(n11751), .A3(n11723), .A4(n11722), .ZN(
        n12055) );
  INV_X1 U14614 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12092) );
  NAND2_X1 U14615 ( .A1(n12103), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11724) );
  OAI211_X1 U14616 ( .C1(n16421), .C2(n12087), .A(n11724), .B(n12070), .ZN(
        n11725) );
  INV_X1 U14617 ( .A(n11725), .ZN(n11726) );
  OAI21_X1 U14618 ( .B1(n14361), .B2(n12092), .A(n11726), .ZN(n12054) );
  NAND2_X1 U14619 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  AOI22_X1 U14620 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n11719), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n11728) );
  XNOR2_X1 U14621 ( .A(n12056), .B(n11732), .ZN(n12123) );
  NAND2_X1 U14622 ( .A1(n11303), .A2(n9603), .ZN(n12052) );
  MUX2_X1 U14623 ( .A(n12052), .B(n19827), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11731) );
  NAND2_X1 U14624 ( .A1(n12903), .A2(n11729), .ZN(n11730) );
  NAND2_X1 U14625 ( .A1(n11731), .A2(n11730), .ZN(n12122) );
  NAND2_X1 U14626 ( .A1(n11732), .A2(n12056), .ZN(n11733) );
  OAI21_X1 U14627 ( .B1(n19817), .B2(n12070), .A(n11734), .ZN(n11735) );
  AOI21_X1 U14628 ( .B1(n12903), .B2(n11736), .A(n11735), .ZN(n11741) );
  AOI222_X1 U14629 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n11738), .B1(n11739), 
        .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n14358), .C2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U14630 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  NAND2_X1 U14631 ( .A1(n11738), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14632 ( .A1(n11719), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n11746) );
  NAND2_X1 U14633 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14634 ( .A1(n12903), .A2(n11743), .ZN(n11744) );
  AOI22_X1 U14635 ( .A1(n11738), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n14358), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14636 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12903), .B2(n11748), .ZN(n11749) );
  NAND2_X1 U14637 ( .A1(n11750), .A2(n11749), .ZN(n12563) );
  NAND2_X1 U14638 ( .A1(n11738), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14639 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U14640 ( .A1(n14358), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n11755) );
  INV_X1 U14641 ( .A(n11752), .ZN(n11753) );
  NAND2_X1 U14642 ( .A1(n12903), .A2(n11753), .ZN(n11754) );
  NAND4_X1 U14643 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n12561) );
  INV_X1 U14644 ( .A(n11758), .ZN(n11759) );
  NAND2_X1 U14645 ( .A1(n12903), .A2(n11759), .ZN(n11760) );
  NAND2_X1 U14646 ( .A1(n12560), .A2(n11760), .ZN(n11764) );
  INV_X1 U14647 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U14648 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U14649 ( .A1(n14358), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n11761) );
  OAI211_X1 U14650 ( .C1(n14361), .C2(n11792), .A(n11762), .B(n11761), .ZN(
        n11763) );
  NAND2_X1 U14651 ( .A1(n11764), .A2(n11763), .ZN(n12280) );
  OR2_X1 U14652 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NAND2_X1 U14653 ( .A1(n12280), .A2(n11765), .ZN(n12811) );
  AND2_X1 U14654 ( .A1(n11766), .A2(n9636), .ZN(n12303) );
  INV_X1 U14655 ( .A(n12303), .ZN(n16400) );
  NAND2_X1 U14656 ( .A1(n11287), .A2(n15473), .ZN(n16397) );
  NAND2_X1 U14657 ( .A1(n16397), .A2(n15526), .ZN(n11768) );
  NAND2_X1 U14658 ( .A1(n16400), .A2(n11768), .ZN(n11769) );
  NAND2_X1 U14659 ( .A1(n11771), .A2(n11769), .ZN(n16319) );
  AND2_X1 U14660 ( .A1(n11770), .A2(n11771), .ZN(n16369) );
  INV_X1 U14661 ( .A(n11774), .ZN(n11776) );
  NAND2_X1 U14662 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  OR2_X1 U14663 ( .A1(n11329), .A2(n15118), .ZN(n11782) );
  NAND2_X1 U14664 ( .A1(n14307), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U14665 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11778) );
  OAI211_X1 U14666 ( .C1(n13534), .C2(n19108), .A(n11779), .B(n11778), .ZN(
        n11780) );
  INV_X1 U14667 ( .A(n11780), .ZN(n11781) );
  OR2_X1 U14668 ( .A1(n11329), .A2(n11783), .ZN(n11789) );
  INV_X1 U14669 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11786) );
  NAND2_X1 U14670 ( .A1(n14307), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U14671 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11784) );
  OAI211_X1 U14672 ( .C1(n11786), .C2(n13534), .A(n11785), .B(n11784), .ZN(
        n11787) );
  INV_X1 U14673 ( .A(n11787), .ZN(n11788) );
  NAND2_X1 U14674 ( .A1(n11789), .A2(n11788), .ZN(n13084) );
  OR2_X1 U14675 ( .A1(n11329), .A2(n9772), .ZN(n11791) );
  AOI22_X1 U14676 ( .A1(n14308), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11790) );
  OAI211_X1 U14677 ( .C1(n13540), .C2(n11792), .A(n11791), .B(n11790), .ZN(
        n11793) );
  NOR2_X1 U14678 ( .A1(n13086), .A2(n11793), .ZN(n11794) );
  NOR2_X1 U14679 ( .A1(n12472), .A2(n11794), .ZN(n16290) );
  INV_X2 U14680 ( .A(n11795), .ZN(n19111) );
  NOR2_X1 U14681 ( .A1(n19089), .A2(n11792), .ZN(n11796) );
  AOI21_X1 U14682 ( .B1(n16369), .B2(n16290), .A(n11796), .ZN(n11797) );
  OAI21_X1 U14683 ( .B1(n12811), .B2(n16319), .A(n11797), .ZN(n11798) );
  OR4_X1 U14684 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        P2_U3040) );
  NOR2_X1 U14685 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n11802), .ZN(n16593)
         );
  INV_X2 U14686 ( .A(n20772), .ZN(U215) );
  INV_X1 U14687 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17685) );
  NAND2_X1 U14688 ( .A1(n17831), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16867) );
  INV_X1 U14689 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17785) );
  NOR2_X1 U14690 ( .A1(n17785), .A2(n16844), .ZN(n11803) );
  INV_X1 U14691 ( .A(n11803), .ZN(n17778) );
  NAND2_X1 U14692 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17734) );
  NAND2_X1 U14693 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17701) );
  INV_X1 U14694 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17927) );
  NOR2_X1 U14695 ( .A1(n17686), .A2(n17927), .ZN(n11804) );
  INV_X1 U14696 ( .A(n11804), .ZN(n17653) );
  NOR2_X1 U14697 ( .A1(n17655), .A2(n17927), .ZN(n16644) );
  AOI21_X1 U14698 ( .B1(n17685), .B2(n17653), .A(n16644), .ZN(n17688) );
  NOR2_X1 U14699 ( .A1(n17776), .A2(n17927), .ZN(n17770) );
  NAND2_X1 U14700 ( .A1(n11803), .A2(n17770), .ZN(n16820) );
  NOR2_X1 U14701 ( .A1(n10043), .A2(n16820), .ZN(n17732) );
  NAND2_X1 U14702 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17732), .ZN(
        n16805) );
  NOR2_X1 U14703 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16805), .ZN(
        n16800) );
  INV_X1 U14704 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16654) );
  INV_X1 U14705 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16667) );
  NAND2_X1 U14706 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17656) );
  INV_X1 U14707 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U14708 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17615) );
  NOR2_X1 U14709 ( .A1(n16729), .A2(n17615), .ZN(n17599) );
  NAND3_X1 U14710 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17610), .A3(
        n17599), .ZN(n17571) );
  INV_X1 U14711 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17592) );
  INV_X1 U14712 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17572) );
  AOI21_X1 U14713 ( .B1(n11804), .B2(n16800), .A(n9694), .ZN(n11805) );
  NOR2_X1 U14714 ( .A1(n17688), .A2(n11805), .ZN(n16645) );
  INV_X1 U14715 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18928) );
  INV_X1 U14716 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18938) );
  INV_X1 U14717 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16612) );
  NAND3_X1 U14718 ( .A1(n18928), .A2(n18938), .A3(n16612), .ZN(n18783) );
  NOR2_X1 U14719 ( .A1(n18885), .A2(n18783), .ZN(n16951) );
  AOI211_X1 U14720 ( .C1(n17688), .C2(n11805), .A(n16645), .B(n18781), .ZN(
        n11923) );
  NOR3_X1 U14721 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16968) );
  INV_X1 U14722 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17294) );
  NAND2_X1 U14723 ( .A1(n16968), .A2(n17294), .ZN(n16964) );
  NOR2_X1 U14724 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16964), .ZN(n16946) );
  INV_X1 U14725 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17281) );
  NAND2_X1 U14726 ( .A1(n16946), .A2(n17281), .ZN(n16936) );
  INV_X1 U14727 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20874) );
  NAND2_X1 U14728 ( .A1(n16915), .A2(n20874), .ZN(n16907) );
  INV_X1 U14729 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U14730 ( .A1(n16886), .A2(n17233), .ZN(n16872) );
  INV_X1 U14731 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16863) );
  NAND2_X1 U14732 ( .A1(n16871), .A2(n16863), .ZN(n16862) );
  INV_X1 U14733 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16841) );
  NAND2_X1 U14734 ( .A1(n16845), .A2(n16841), .ZN(n16840) );
  INV_X1 U14735 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U14736 ( .A1(n16817), .A2(n16811), .ZN(n16810) );
  INV_X1 U14737 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16791) );
  NAND2_X1 U14738 ( .A1(n16795), .A2(n16791), .ZN(n16790) );
  INV_X1 U14739 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16766) );
  NAND2_X1 U14740 ( .A1(n16772), .A2(n16766), .ZN(n16764) );
  NAND2_X1 U14741 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18919) );
  AOI22_X1 U14742 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11810) );
  INV_X4 U14743 ( .A(n9642), .ZN(n17270) );
  OR2_X2 U14744 ( .A1(n11806), .A2(n18740), .ZN(n17178) );
  INV_X4 U14745 ( .A(n17178), .ZN(n17237) );
  AOI22_X1 U14746 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11809) );
  INV_X4 U14747 ( .A(n17241), .ZN(n17185) );
  AOI22_X1 U14748 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11808) );
  BUF_X4 U14749 ( .A(n15740), .Z(n17244) );
  AOI22_X1 U14750 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11807) );
  NAND4_X1 U14751 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11821) );
  AOI22_X1 U14752 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11819) );
  BUF_X4 U14753 ( .A(n15736), .Z(n17269) );
  AOI22_X1 U14754 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11818) );
  BUF_X4 U14755 ( .A(n15729), .Z(n17271) );
  AOI22_X1 U14756 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11817) );
  BUF_X4 U14757 ( .A(n15737), .Z(n17238) );
  AOI22_X1 U14758 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11816) );
  NAND4_X1 U14759 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11820) );
  AOI22_X1 U14760 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14761 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17244), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17242), .ZN(n11824) );
  AOI22_X1 U14762 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14763 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17238), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17237), .ZN(n11822) );
  NAND4_X1 U14764 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11831) );
  AOI22_X1 U14765 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14766 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n15780), .ZN(n11828) );
  AOI22_X1 U14767 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17262), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14768 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17271), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17270), .ZN(n11826) );
  NAND4_X1 U14769 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11830) );
  AOI22_X1 U14770 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11835) );
  BUF_X4 U14771 ( .A(n15753), .Z(n17262) );
  AOI22_X1 U14772 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14773 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14774 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U14775 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11841) );
  AOI22_X1 U14776 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14777 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14778 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14779 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11836) );
  NAND4_X1 U14780 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11840) );
  AOI22_X1 U14781 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14782 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14783 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14784 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11842) );
  NAND4_X1 U14785 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11851) );
  AOI22_X1 U14786 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14787 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14788 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14789 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11846) );
  NAND4_X1 U14790 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11850) );
  AOI22_X1 U14791 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14792 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14793 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11852) );
  OAI21_X1 U14794 ( .B1(n10232), .B2(n18284), .A(n11852), .ZN(n11858) );
  AOI22_X1 U14795 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14796 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14797 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14798 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U14799 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  AOI211_X1 U14800 ( .C1(n17260), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11858), .B(n11857), .ZN(n11859) );
  NAND3_X1 U14801 ( .A1(n11861), .A2(n11860), .A3(n11859), .ZN(n15682) );
  AOI22_X1 U14802 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14803 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14804 ( .A1(n17239), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11862) );
  OAI21_X1 U14805 ( .B1(n15605), .B2(n20811), .A(n11862), .ZN(n11868) );
  INV_X2 U14806 ( .A(n10232), .ZN(n17261) );
  AOI22_X1 U14807 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14808 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14809 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14810 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U14811 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11867) );
  INV_X1 U14812 ( .A(n15683), .ZN(n18308) );
  AOI22_X1 U14813 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14814 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14815 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14816 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11871) );
  NAND4_X1 U14817 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n11880) );
  AOI22_X1 U14818 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14819 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14820 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14821 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U14822 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11879) );
  NOR2_X1 U14823 ( .A1(n18316), .A2(n17462), .ZN(n11900) );
  NAND4_X1 U14824 ( .A1(n18287), .A2(n18293), .A3(n11900), .A4(n11881), .ZN(
        n11892) );
  AOI22_X1 U14825 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14826 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14827 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11882) );
  OAI21_X1 U14828 ( .B1(n17207), .B2(n20791), .A(n11882), .ZN(n11888) );
  AOI22_X1 U14829 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14830 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14831 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14832 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U14833 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  INV_X1 U14834 ( .A(n11892), .ZN(n11902) );
  INV_X1 U14835 ( .A(n18287), .ZN(n11903) );
  NOR2_X1 U14836 ( .A1(n18300), .A2(n15682), .ZN(n15691) );
  NOR2_X1 U14837 ( .A1(n18300), .A2(n15683), .ZN(n18744) );
  NAND2_X1 U14838 ( .A1(n18274), .A2(n17462), .ZN(n15672) );
  INV_X1 U14839 ( .A(n15672), .ZN(n11893) );
  OAI21_X1 U14840 ( .B1(n18316), .B2(n18744), .A(n11893), .ZN(n13078) );
  OAI21_X1 U14841 ( .B1(n15691), .B2(n11894), .A(n13078), .ZN(n11901) );
  NAND2_X1 U14842 ( .A1(n18281), .A2(n15673), .ZN(n13074) );
  AOI21_X1 U14843 ( .B1(n17424), .B2(n11896), .A(n18293), .ZN(n11895) );
  AOI21_X1 U14844 ( .B1(n11896), .B2(n13074), .A(n11895), .ZN(n11899) );
  NOR2_X1 U14845 ( .A1(n18293), .A2(n15683), .ZN(n18722) );
  AOI21_X1 U14846 ( .B1(n18281), .B2(n18925), .A(n18744), .ZN(n11897) );
  OR3_X1 U14847 ( .A1(n18722), .A2(n11897), .A3(n13075), .ZN(n11898) );
  OAI211_X1 U14848 ( .C1(n11900), .C2(n11903), .A(n11899), .B(n11898), .ZN(
        n13077) );
  AOI21_X1 U14849 ( .B1(n11903), .B2(n11901), .A(n13077), .ZN(n15681) );
  NAND2_X1 U14850 ( .A1(n11902), .A2(n15681), .ZN(n15675) );
  NOR2_X1 U14851 ( .A1(n11903), .A2(n15682), .ZN(n18721) );
  NOR2_X1 U14852 ( .A1(n16445), .A2(n17462), .ZN(n15913) );
  AND2_X1 U14853 ( .A1(n17424), .A2(n15913), .ZN(n11904) );
  NAND2_X1 U14854 ( .A1(n18748), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13062) );
  INV_X1 U14855 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18755) );
  OAI22_X1 U14856 ( .A1(n18892), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18755), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11910) );
  OAI22_X1 U14857 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18759), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11907), .ZN(n11913) );
  NOR2_X1 U14858 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18759), .ZN(
        n11908) );
  NAND2_X1 U14859 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11907), .ZN(
        n11912) );
  AOI22_X1 U14860 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11913), .B1(
        n11908), .B2(n11912), .ZN(n13066) );
  OAI21_X1 U14861 ( .B1(n11911), .B2(n11910), .A(n13066), .ZN(n11909) );
  XOR2_X1 U14862 ( .A(n13062), .B(n13063), .Z(n11915) );
  INV_X1 U14863 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18716) );
  OAI22_X1 U14864 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18716), .B1(
        n11914), .B2(n11913), .ZN(n13064) );
  NOR2_X1 U14865 ( .A1(n18928), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18778) );
  NAND2_X1 U14866 ( .A1(n18778), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18773) );
  INV_X1 U14867 ( .A(n17501), .ZN(n16607) );
  NAND2_X1 U14868 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16445), .ZN(n11916) );
  AOI211_X4 U14869 ( .C1(n16612), .C2(n18919), .A(n11918), .B(n11916), .ZN(
        n16965) );
  AOI211_X1 U14870 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16764), .A(n16751), .B(
        n16995), .ZN(n11922) );
  NAND2_X1 U14871 ( .A1(n18885), .A2(n18872), .ZN(n18884) );
  INV_X1 U14872 ( .A(n18941), .ZN(n16947) );
  NAND2_X1 U14873 ( .A1(n18938), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18776) );
  INV_X1 U14874 ( .A(n18776), .ZN(n18647) );
  NAND2_X1 U14875 ( .A1(n18778), .A2(n18647), .ZN(n18772) );
  INV_X2 U14876 ( .A(n18936), .ZN(n18935) );
  OAI211_X1 U14877 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18799), .B(n18861), .ZN(n18792) );
  INV_X1 U14878 ( .A(n18792), .ZN(n18924) );
  OAI211_X1 U14879 ( .C1(n18924), .C2(n16445), .A(n18919), .B(n16612), .ZN(
        n18767) );
  INV_X1 U14880 ( .A(n18767), .ZN(n11917) );
  AOI211_X4 U14881 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16445), .A(n11917), .B(
        n11918), .ZN(n16976) );
  INV_X1 U14882 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n15572) );
  OAI22_X1 U14883 ( .A1(n17685), .A2(n16987), .B1(n16996), .B2(n15572), .ZN(
        n11921) );
  INV_X1 U14884 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18836) );
  INV_X1 U14885 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18833) );
  INV_X1 U14886 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18830) );
  INV_X1 U14887 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18828) );
  NOR3_X1 U14888 ( .A1(n18833), .A2(n18830), .A3(n18828), .ZN(n16760) );
  INV_X1 U14889 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18827) );
  INV_X1 U14890 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18823) );
  INV_X1 U14891 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18816) );
  INV_X1 U14892 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18811) );
  INV_X1 U14893 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18807) );
  NAND3_X1 U14894 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16954) );
  NOR2_X1 U14895 ( .A1(n18807), .A2(n16954), .ZN(n16931) );
  NAND2_X1 U14896 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16931), .ZN(n16916) );
  NOR2_X1 U14897 ( .A1(n18811), .A2(n16916), .ZN(n16912) );
  NAND2_X1 U14898 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16912), .ZN(n16894) );
  NOR2_X1 U14899 ( .A1(n18816), .A2(n16894), .ZN(n16829) );
  NAND4_X1 U14900 ( .A1(n16829), .A2(P3_REIP_REG_11__SCAN_IN), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16850) );
  NOR2_X1 U14901 ( .A1(n18823), .A2(n16850), .ZN(n16833) );
  NAND2_X1 U14902 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16833), .ZN(n16821) );
  NOR3_X1 U14903 ( .A1(n16989), .A2(n18827), .A3(n16821), .ZN(n16786) );
  AND2_X1 U14904 ( .A1(n16760), .A2(n16786), .ZN(n16778) );
  NAND2_X1 U14905 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16778), .ZN(n16771) );
  NOR2_X1 U14906 ( .A1(n18836), .A2(n16771), .ZN(n11919) );
  INV_X1 U14907 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18838) );
  INV_X1 U14908 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18834) );
  NOR3_X1 U14909 ( .A1(n18838), .A2(n18836), .A3(n18834), .ZN(n16740) );
  AND2_X1 U14910 ( .A1(n16760), .A2(n16740), .ZN(n16634) );
  NOR2_X1 U14911 ( .A1(n18827), .A2(n16821), .ZN(n16635) );
  NAND2_X1 U14912 ( .A1(n16635), .A2(n16999), .ZN(n16822) );
  INV_X1 U14913 ( .A(n16822), .ZN(n16759) );
  NAND2_X1 U14914 ( .A1(n16989), .A2(n16999), .ZN(n16997) );
  INV_X1 U14915 ( .A(n16997), .ZN(n16758) );
  AOI21_X1 U14916 ( .B1(n16634), .B2(n16759), .A(n16758), .ZN(n16747) );
  MUX2_X1 U14917 ( .A(n11919), .B(n16747), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n11920) );
  OR4_X1 U14918 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        P3_U2651) );
  AOI21_X1 U14919 ( .B1(n19799), .B2(n13505), .A(P2_READREQUEST_REG_SCAN_IN), 
        .ZN(n11925) );
  NAND2_X1 U14920 ( .A1(n18951), .A2(n11700), .ZN(n11924) );
  OAI21_X1 U14921 ( .B1(n18951), .B2(n11925), .A(n11924), .ZN(P2_U3612) );
  INV_X1 U14922 ( .A(n12320), .ZN(n11927) );
  AND2_X1 U14923 ( .A1(n11700), .A2(n19714), .ZN(n12319) );
  NOR3_X1 U14924 ( .A1(n11927), .A2(n12319), .A3(n11926), .ZN(n16402) );
  NOR2_X1 U14925 ( .A1(n16402), .A2(n19146), .ZN(n19845) );
  NOR2_X1 U14926 ( .A1(n16408), .A2(n19146), .ZN(n11928) );
  NAND2_X1 U14927 ( .A1(n11929), .A2(n11928), .ZN(n12079) );
  OAI21_X1 U14928 ( .B1(n19845), .B2(n11589), .A(n12079), .ZN(P2_U2819) );
  NAND2_X1 U14929 ( .A1(n16395), .A2(n12098), .ZN(n12834) );
  OAI21_X1 U14930 ( .B1(n16421), .B2(n19714), .A(n18946), .ZN(n11942) );
  AOI22_X1 U14931 ( .A1(n12795), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11942), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n11930) );
  NAND3_X1 U14932 ( .A1(n18946), .A2(n19714), .A3(n15526), .ZN(n11980) );
  AOI22_X1 U14933 ( .A1(n13482), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n13481), .ZN(n12753) );
  INV_X1 U14934 ( .A(n12753), .ZN(n13479) );
  NAND2_X1 U14935 ( .A1(n11988), .A2(n13479), .ZN(n11969) );
  NAND2_X1 U14936 ( .A1(n11930), .A2(n11969), .ZN(P2_U2981) );
  AOI22_X1 U14937 ( .A1(n12795), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11942), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14938 ( .A1(n13482), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13481), .ZN(n12620) );
  INV_X1 U14939 ( .A(n12620), .ZN(n14691) );
  NAND2_X1 U14940 ( .A1(n11988), .A2(n14691), .ZN(n11977) );
  NAND2_X1 U14941 ( .A1(n11931), .A2(n11977), .ZN(P2_U2979) );
  AOI22_X1 U14942 ( .A1(n12795), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11942), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n11935) );
  INV_X1 U14943 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n11932) );
  OR2_X1 U14944 ( .A1(n13481), .A2(n11932), .ZN(n11934) );
  NAND2_X1 U14945 ( .A1(n13481), .A2(BUF2_REG_10__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U14946 ( .A1(n11934), .A2(n11933), .ZN(n14704) );
  NAND2_X1 U14947 ( .A1(n11988), .A2(n14704), .ZN(n11973) );
  NAND2_X1 U14948 ( .A1(n11935), .A2(n11973), .ZN(P2_U2977) );
  AOI22_X1 U14949 ( .A1(n12795), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11942), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n11936) );
  OAI22_X1 U14950 ( .A1(n13481), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13482), .ZN(n12333) );
  INV_X1 U14951 ( .A(n12333), .ZN(n16229) );
  NAND2_X1 U14952 ( .A1(n11988), .A2(n16229), .ZN(n11965) );
  NAND2_X1 U14953 ( .A1(n11936), .A2(n11965), .ZN(P2_U2974) );
  AOI22_X1 U14954 ( .A1(n12795), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11942), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U14955 ( .A1(n13482), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13481), .ZN(n12818) );
  INV_X1 U14956 ( .A(n12818), .ZN(n14773) );
  NAND2_X1 U14957 ( .A1(n11988), .A2(n14773), .ZN(n11951) );
  NAND2_X1 U14958 ( .A1(n11937), .A2(n11951), .ZN(P2_U2952) );
  AOI22_X1 U14959 ( .A1(n12795), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11942), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n11941) );
  INV_X1 U14960 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n11938) );
  OR2_X1 U14961 ( .A1(n13481), .A2(n11938), .ZN(n11940) );
  NAND2_X1 U14962 ( .A1(n13481), .A2(BUF2_REG_9__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U14963 ( .A1(n11940), .A2(n11939), .ZN(n14709) );
  NAND2_X1 U14964 ( .A1(n11988), .A2(n14709), .ZN(n11961) );
  NAND2_X1 U14965 ( .A1(n11941), .A2(n11961), .ZN(P2_U2976) );
  AOI22_X1 U14966 ( .A1(n12795), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14967 ( .A1(n13482), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13481), .ZN(n15531) );
  INV_X1 U14968 ( .A(n15531), .ZN(n14752) );
  NAND2_X1 U14969 ( .A1(n11988), .A2(n14752), .ZN(n11955) );
  NAND2_X1 U14970 ( .A1(n11943), .A2(n11955), .ZN(P2_U2969) );
  AOI22_X1 U14971 ( .A1(n12795), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U14972 ( .A1(n13482), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13481), .ZN(n15548) );
  INV_X1 U14973 ( .A(n15548), .ZN(n14728) );
  NAND2_X1 U14974 ( .A1(n11988), .A2(n14728), .ZN(n11975) );
  NAND2_X1 U14975 ( .A1(n11944), .A2(n11975), .ZN(P2_U2972) );
  AOI22_X1 U14976 ( .A1(n12795), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11990), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U14977 ( .A1(n13482), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13481), .ZN(n15492) );
  INV_X1 U14978 ( .A(n15492), .ZN(n14721) );
  NAND2_X1 U14979 ( .A1(n11988), .A2(n14721), .ZN(n11957) );
  NAND2_X1 U14980 ( .A1(n11945), .A2(n11957), .ZN(P2_U2958) );
  AOI22_X1 U14981 ( .A1(n12795), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U14982 ( .A1(n13482), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13481), .ZN(n15542) );
  INV_X1 U14983 ( .A(n15542), .ZN(n14734) );
  NAND2_X1 U14984 ( .A1(n11988), .A2(n14734), .ZN(n11959) );
  NAND2_X1 U14985 ( .A1(n11946), .A2(n11959), .ZN(P2_U2971) );
  AOI22_X1 U14986 ( .A1(n12795), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n11950) );
  INV_X1 U14987 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n11947) );
  OR2_X1 U14988 ( .A1(n13481), .A2(n11947), .ZN(n11949) );
  NAND2_X1 U14989 ( .A1(n13481), .A2(BUF2_REG_8__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14990 ( .A1(n11949), .A2(n11948), .ZN(n14714) );
  NAND2_X1 U14991 ( .A1(n11988), .A2(n14714), .ZN(n11967) );
  NAND2_X1 U14992 ( .A1(n11950), .A2(n11967), .ZN(P2_U2975) );
  AOI22_X1 U14993 ( .A1(n12795), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14994 ( .A1(n11952), .A2(n11951), .ZN(P2_U2967) );
  AOI22_X1 U14995 ( .A1(n12795), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14996 ( .A1(n13482), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13481), .ZN(n15525) );
  INV_X1 U14997 ( .A(n15525), .ZN(n14761) );
  NAND2_X1 U14998 ( .A1(n11988), .A2(n14761), .ZN(n11971) );
  NAND2_X1 U14999 ( .A1(n11953), .A2(n11971), .ZN(P2_U2968) );
  AOI22_X1 U15000 ( .A1(n12795), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15001 ( .A1(n13482), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13481), .ZN(n15536) );
  INV_X1 U15002 ( .A(n15536), .ZN(n14742) );
  NAND2_X1 U15003 ( .A1(n11988), .A2(n14742), .ZN(n11963) );
  NAND2_X1 U15004 ( .A1(n11954), .A2(n11963), .ZN(P2_U2970) );
  AOI22_X1 U15005 ( .A1(n12795), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11990), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U15006 ( .A1(n11956), .A2(n11955), .ZN(P2_U2954) );
  AOI22_X1 U15007 ( .A1(n12795), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11990), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U15008 ( .A1(n11958), .A2(n11957), .ZN(P2_U2973) );
  AOI22_X1 U15009 ( .A1(n12795), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11990), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15010 ( .A1(n11960), .A2(n11959), .ZN(P2_U2956) );
  AOI22_X1 U15011 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U15012 ( .A1(n11962), .A2(n11961), .ZN(P2_U2961) );
  AOI22_X1 U15013 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U15014 ( .A1(n11964), .A2(n11963), .ZN(P2_U2955) );
  AOI22_X1 U15015 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U15016 ( .A1(n11966), .A2(n11965), .ZN(P2_U2959) );
  AOI22_X1 U15017 ( .A1(P2_EAX_REG_24__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n11968) );
  NAND2_X1 U15018 ( .A1(n11968), .A2(n11967), .ZN(P2_U2960) );
  AOI22_X1 U15019 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n11970) );
  NAND2_X1 U15020 ( .A1(n11970), .A2(n11969), .ZN(P2_U2966) );
  AOI22_X1 U15021 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U15022 ( .A1(n11972), .A2(n11971), .ZN(P2_U2953) );
  AOI22_X1 U15023 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U15024 ( .A1(n11974), .A2(n11973), .ZN(P2_U2962) );
  AOI22_X1 U15025 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15026 ( .A1(n11976), .A2(n11975), .ZN(P2_U2957) );
  AOI22_X1 U15027 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U15028 ( .A1(n11978), .A2(n11977), .ZN(P2_U2964) );
  AOI22_X1 U15029 ( .A1(n13482), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13481), .ZN(n12908) );
  AOI22_X1 U15030 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n12795), .B1(n11990), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n11979) );
  OAI21_X1 U15031 ( .B1(n12908), .B2(n11980), .A(n11979), .ZN(P2_U2982) );
  INV_X1 U15032 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19157) );
  INV_X1 U15033 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16551) );
  OR2_X1 U15034 ( .A1(n13481), .A2(n16551), .ZN(n11982) );
  NAND2_X1 U15035 ( .A1(n13481), .A2(BUF2_REG_11__SCAN_IN), .ZN(n11981) );
  AND2_X1 U15036 ( .A1(n11982), .A2(n11981), .ZN(n14697) );
  INV_X1 U15037 ( .A(n14697), .ZN(n19139) );
  NAND2_X1 U15038 ( .A1(n11988), .A2(n19139), .ZN(n11985) );
  NAND2_X1 U15039 ( .A1(n11990), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n11983) );
  OAI211_X1 U15040 ( .C1(n19145), .C2(n19157), .A(n11985), .B(n11983), .ZN(
        P2_U2963) );
  INV_X1 U15041 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19189) );
  NAND2_X1 U15042 ( .A1(n11990), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n11984) );
  OAI211_X1 U15043 ( .C1(n19145), .C2(n19189), .A(n11985), .B(n11984), .ZN(
        P2_U2978) );
  INV_X1 U15044 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19153) );
  INV_X1 U15045 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16548) );
  OR2_X1 U15046 ( .A1(n13481), .A2(n16548), .ZN(n11987) );
  NAND2_X1 U15047 ( .A1(n13481), .A2(BUF2_REG_13__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U15048 ( .A1(n11987), .A2(n11986), .ZN(n19136) );
  NAND2_X1 U15049 ( .A1(n11988), .A2(n19136), .ZN(n11992) );
  NAND2_X1 U15050 ( .A1(n11990), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n11989) );
  OAI211_X1 U15051 ( .C1(n19145), .C2(n19153), .A(n11992), .B(n11989), .ZN(
        P2_U2965) );
  INV_X1 U15052 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20783) );
  NAND2_X1 U15053 ( .A1(n11990), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n11991) );
  OAI211_X1 U15054 ( .C1(n19145), .C2(n20783), .A(n11992), .B(n11991), .ZN(
        P2_U2980) );
  NAND2_X1 U15055 ( .A1(n13000), .A2(n12976), .ZN(n11994) );
  NOR3_X1 U15056 ( .A1(n11997), .A2(n11996), .A3(n11995), .ZN(n11999) );
  OAI21_X1 U15057 ( .B1(n12000), .B2(n11999), .A(n11998), .ZN(n12961) );
  NAND2_X1 U15058 ( .A1(n12135), .A2(n12976), .ZN(n12002) );
  NAND2_X1 U15059 ( .A1(n20510), .A2(n20649), .ZN(n19852) );
  INV_X1 U15060 ( .A(n19852), .ZN(n12003) );
  AOI21_X1 U15061 ( .B1(n12002), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12003), 
        .ZN(n12001) );
  NAND2_X1 U15062 ( .A1(n12231), .A2(n12001), .ZN(P1_U2801) );
  NOR2_X1 U15063 ( .A1(n12003), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12006)
         );
  NAND2_X1 U15064 ( .A1(n20739), .A2(n12004), .ZN(n12005) );
  OAI21_X1 U15065 ( .B1(n20739), .B2(n12006), .A(n12005), .ZN(P1_U3487) );
  INV_X1 U15066 ( .A(n12973), .ZN(n12014) );
  OAI22_X1 U15067 ( .A1(n12014), .A2(n12131), .B1(n13000), .B2(n12135), .ZN(
        n19850) );
  NAND2_X1 U15068 ( .A1(n12007), .A2(n20668), .ZN(n15907) );
  INV_X1 U15069 ( .A(n15907), .ZN(n12629) );
  NOR3_X1 U15070 ( .A1(n12131), .A2(n13585), .A3(n12629), .ZN(n12008) );
  NAND2_X1 U15071 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20741) );
  INV_X1 U15072 ( .A(n20741), .ZN(n15905) );
  NOR2_X1 U15073 ( .A1(n12008), .A2(n15905), .ZN(n20743) );
  NOR2_X1 U15074 ( .A1(n19850), .A2(n20743), .ZN(n15876) );
  OR2_X1 U15075 ( .A1(n15876), .A2(n19849), .ZN(n19856) );
  INV_X1 U15076 ( .A(n19856), .ZN(n12023) );
  INV_X1 U15077 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12022) );
  INV_X1 U15078 ( .A(n12009), .ZN(n12142) );
  NAND2_X1 U15079 ( .A1(n12628), .A2(n12015), .ZN(n12010) );
  NAND2_X1 U15080 ( .A1(n12142), .A2(n12010), .ZN(n12991) );
  INV_X1 U15081 ( .A(n12991), .ZN(n12011) );
  AOI21_X1 U15082 ( .B1(n12012), .B2(n12978), .A(n12011), .ZN(n12013) );
  OAI22_X1 U15083 ( .A1(n12014), .A2(n12013), .B1(n12961), .B2(n12144), .ZN(
        n12020) );
  INV_X1 U15084 ( .A(n12634), .ZN(n12016) );
  AND2_X1 U15085 ( .A1(n12016), .A2(n12015), .ZN(n12017) );
  OR2_X1 U15086 ( .A1(n12018), .A2(n12017), .ZN(n12155) );
  NAND2_X1 U15087 ( .A1(n12166), .A2(n12959), .ZN(n12970) );
  NOR2_X1 U15088 ( .A1(n12155), .A2(n12970), .ZN(n12139) );
  INV_X1 U15089 ( .A(n12139), .ZN(n12986) );
  NOR2_X1 U15090 ( .A1(n12973), .A2(n12986), .ZN(n12019) );
  OAI21_X1 U15091 ( .B1(n12020), .B2(n12019), .A(n12500), .ZN(n15877) );
  OR2_X1 U15092 ( .A1(n19856), .A2(n15877), .ZN(n12021) );
  OAI21_X1 U15093 ( .B1(n12023), .B2(n12022), .A(n12021), .ZN(P1_U3484) );
  NOR3_X1 U15094 ( .A1(n15316), .A2(n12037), .A3(n12038), .ZN(n12030) );
  INV_X1 U15095 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19743) );
  NOR2_X1 U15096 ( .A1(n11795), .A2(n19743), .ZN(n19221) );
  INV_X1 U15097 ( .A(n12024), .ZN(n19219) );
  NOR2_X1 U15098 ( .A1(n12026), .A2(n12025), .ZN(n19220) );
  NOR3_X1 U15099 ( .A1(n16373), .A2(n19219), .A3(n19220), .ZN(n12029) );
  NOR2_X1 U15100 ( .A1(n16374), .A2(n12027), .ZN(n12028) );
  NOR4_X1 U15101 ( .A1(n12030), .A2(n19221), .A3(n12029), .A4(n12028), .ZN(
        n12042) );
  OAI21_X1 U15102 ( .B1(n12033), .B2(n12032), .A(n12031), .ZN(n19815) );
  OAI21_X1 U15103 ( .B1(n12036), .B2(n12035), .A(n12034), .ZN(n19214) );
  NOR2_X1 U15104 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  OAI22_X1 U15105 ( .A1(n16383), .A2(n19214), .B1(n12039), .B2(n15319), .ZN(
        n12040) );
  AOI21_X1 U15106 ( .B1(n16371), .B2(n19815), .A(n12040), .ZN(n12041) );
  OAI211_X1 U15107 ( .C1(n12200), .C2(n16309), .A(n12042), .B(n12041), .ZN(
        P2_U3044) );
  INV_X1 U15108 ( .A(n16401), .ZN(n12043) );
  NAND2_X1 U15109 ( .A1(n12043), .A2(n16398), .ZN(n12324) );
  INV_X1 U15110 ( .A(n12044), .ZN(n12045) );
  NAND3_X1 U15111 ( .A1(n12047), .A2(n12046), .A3(n12045), .ZN(n12048) );
  NAND2_X1 U15112 ( .A1(n12324), .A2(n12048), .ZN(n12049) );
  NAND2_X1 U15113 ( .A1(n12049), .A2(n12098), .ZN(n12051) );
  NAND2_X1 U15114 ( .A1(n18951), .A2(n12319), .ZN(n12050) );
  INV_X1 U15115 ( .A(n12052), .ZN(n12053) );
  NAND2_X1 U15116 ( .A1(n19144), .A2(n12053), .ZN(n13092) );
  INV_X1 U15117 ( .A(n13092), .ZN(n19140) );
  OR2_X1 U15118 ( .A1(n12055), .A2(n12054), .ZN(n12057) );
  AND2_X1 U15119 ( .A1(n12057), .A2(n12056), .ZN(n16370) );
  INV_X1 U15120 ( .A(n16370), .ZN(n12066) );
  INV_X1 U15121 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19213) );
  OAI22_X1 U15122 ( .A1(n14776), .A2(n12066), .B1(n19213), .B2(n19144), .ZN(
        n12068) );
  NAND2_X1 U15123 ( .A1(n15494), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15124 ( .A1(n12287), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19799), .B2(n19836), .ZN(n12059) );
  INV_X1 U15125 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15489) );
  NAND2_X1 U15126 ( .A1(n12070), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12061) );
  NOR2_X1 U15127 ( .A1(n15494), .A2(n12061), .ZN(n12062) );
  OAI21_X1 U15128 ( .B1(n16421), .B2(n15489), .A(n12062), .ZN(n12063) );
  INV_X1 U15129 ( .A(n12063), .ZN(n12064) );
  NOR2_X1 U15130 ( .A1(n19831), .A2(n12066), .ZN(n12127) );
  AOI211_X1 U15131 ( .C1(n19831), .C2(n12066), .A(n12127), .B(n14779), .ZN(
        n12067) );
  AOI211_X1 U15132 ( .C1(n19140), .C2(n14773), .A(n12068), .B(n12067), .ZN(
        n12069) );
  INV_X1 U15133 ( .A(n12069), .ZN(P2_U2919) );
  INV_X1 U15134 ( .A(n15448), .ZN(n15429) );
  NAND2_X1 U15135 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n14298) );
  OAI21_X1 U15136 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n16435), .ZN(n16427) );
  INV_X1 U15137 ( .A(n16427), .ZN(n12071) );
  AOI22_X4 U15138 ( .A1(n16435), .A2(n16428), .B1(n14298), .B2(n12071), .ZN(
        n19463) );
  AOI21_X1 U15139 ( .B1(n12786), .B2(n12073), .A(n12072), .ZN(n15433) );
  INV_X1 U15140 ( .A(n12079), .ZN(n12074) );
  XNOR2_X1 U15141 ( .A(n12086), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12075) );
  XNOR2_X1 U15142 ( .A(n12075), .B(n14553), .ZN(n15434) );
  INV_X1 U15143 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12076) );
  NOR2_X1 U15144 ( .A1(n19089), .A2(n12076), .ZN(n15431) );
  AOI21_X1 U15145 ( .B1(n16302), .B2(n15434), .A(n15431), .ZN(n12077) );
  INV_X1 U15146 ( .A(n12077), .ZN(n12083) );
  INV_X1 U15147 ( .A(n19801), .ZN(n18952) );
  OR2_X1 U15148 ( .A1(n19799), .A2(n18952), .ZN(n19818) );
  NAND2_X1 U15149 ( .A1(n19818), .A2(n16435), .ZN(n12078) );
  INV_X1 U15150 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n18957) );
  NAND2_X1 U15151 ( .A1(n18957), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U15152 ( .A1(n9864), .A2(n12080), .ZN(n12095) );
  INV_X1 U15153 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12081) );
  MUX2_X1 U15154 ( .A(n19215), .B(n16295), .S(n12081), .Z(n12082) );
  AOI211_X1 U15155 ( .C1(n15433), .C2(n19216), .A(n12083), .B(n12082), .ZN(
        n12084) );
  OAI21_X1 U15156 ( .B1(n15429), .B2(n15115), .A(n12084), .ZN(P2_U3013) );
  INV_X1 U15157 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n12085) );
  OAI222_X1 U15158 ( .A1(n12085), .A2(n19144), .B1(n13092), .B2(n15492), .C1(
        n12811), .C2(n19135), .ZN(P2_U2913) );
  OAI21_X1 U15159 ( .B1(n14566), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12086), .ZN(n16372) );
  NAND2_X1 U15160 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  NAND2_X1 U15161 ( .A1(n12090), .A2(n12089), .ZN(n16382) );
  INV_X1 U15162 ( .A(n16382), .ZN(n12091) );
  NAND2_X1 U15163 ( .A1(n19216), .A2(n12091), .ZN(n12093) );
  OR2_X1 U15164 ( .A1(n19089), .A2(n12092), .ZN(n16380) );
  OAI211_X1 U15165 ( .C1(n16372), .C2(n19218), .A(n12093), .B(n16380), .ZN(
        n12094) );
  INV_X1 U15166 ( .A(n12094), .ZN(n12097) );
  OAI21_X1 U15167 ( .B1(n19215), .B2(n12095), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12096) );
  OAI211_X1 U15168 ( .C1(n12120), .C2(n15115), .A(n12097), .B(n12096), .ZN(
        P2_U3014) );
  NAND2_X1 U15169 ( .A1(n16401), .A2(n12303), .ZN(n12322) );
  NAND2_X1 U15170 ( .A1(n12322), .A2(n11321), .ZN(n12099) );
  AND2_X2 U15171 ( .A1(n12099), .A2(n12098), .ZN(n14652) );
  INV_X1 U15172 ( .A(n13363), .ZN(n13309) );
  NAND2_X1 U15173 ( .A1(n13309), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12196) );
  NAND2_X1 U15174 ( .A1(n12287), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12101) );
  NAND2_X1 U15175 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19827), .ZN(
        n19461) );
  NAND2_X1 U15176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19836), .ZN(
        n19494) );
  NAND2_X1 U15177 ( .A1(n19461), .A2(n19494), .ZN(n19371) );
  NAND2_X1 U15178 ( .A1(n19799), .A2(n19371), .ZN(n19497) );
  NAND2_X1 U15179 ( .A1(n12101), .A2(n19497), .ZN(n12102) );
  NAND2_X1 U15180 ( .A1(n19823), .A2(n14658), .ZN(n12105) );
  NAND2_X1 U15181 ( .A1(n14652), .A2(n15448), .ZN(n12104) );
  OAI211_X1 U15182 ( .C1(n14652), .C2(n14557), .A(n12105), .B(n12104), .ZN(
        P2_U2886) );
  INV_X1 U15183 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12109) );
  INV_X1 U15184 ( .A(n12985), .ZN(n12176) );
  NAND2_X1 U15185 ( .A1(n12176), .A2(n12976), .ZN(n12106) );
  OAI22_X1 U15186 ( .A1(n12231), .A2(n12959), .B1(n12973), .B2(n12106), .ZN(
        n12107) );
  NAND2_X1 U15187 ( .A1(n19959), .A2(n12978), .ZN(n12372) );
  NAND2_X1 U15188 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16180) );
  NOR2_X1 U15189 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16180), .ZN(n19987) );
  NOR2_X4 U15190 ( .A1(n19959), .A2(n20742), .ZN(n19986) );
  AOI22_X1 U15191 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12108) );
  OAI21_X1 U15192 ( .B1(n12109), .B2(n12372), .A(n12108), .ZN(P1_U2907) );
  INV_X1 U15193 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15194 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12110) );
  OAI21_X1 U15195 ( .B1(n12111), .B2(n12372), .A(n12110), .ZN(P1_U2909) );
  AOI22_X1 U15196 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12112) );
  OAI21_X1 U15197 ( .B1(n13858), .B2(n12372), .A(n12112), .ZN(P1_U2908) );
  AOI22_X1 U15198 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12113) );
  OAI21_X1 U15199 ( .B1(n13867), .B2(n12372), .A(n12113), .ZN(P1_U2910) );
  INV_X1 U15200 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15201 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12114) );
  OAI21_X1 U15202 ( .B1(n12115), .B2(n12372), .A(n12114), .ZN(P1_U2911) );
  INV_X1 U15203 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15204 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12116) );
  OAI21_X1 U15205 ( .B1(n12117), .B2(n12372), .A(n12116), .ZN(P1_U2912) );
  INV_X1 U15206 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15207 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12118) );
  OAI21_X1 U15208 ( .B1(n12119), .B2(n12372), .A(n12118), .ZN(P1_U2906) );
  MUX2_X1 U15209 ( .A(n11317), .B(n12120), .S(n14652), .Z(n12121) );
  OAI21_X1 U15210 ( .B1(n14677), .B2(n19831), .A(n12121), .ZN(P2_U2887) );
  NAND2_X1 U15211 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  NAND2_X1 U15212 ( .A1(n12125), .A2(n12124), .ZN(n19825) );
  INV_X1 U15213 ( .A(n19825), .ZN(n15428) );
  NAND2_X1 U15214 ( .A1(n19820), .A2(n15428), .ZN(n12413) );
  OAI21_X1 U15215 ( .B1(n19820), .B2(n15428), .A(n12413), .ZN(n12126) );
  NOR2_X1 U15216 ( .A1(n12126), .A2(n12127), .ZN(n12415) );
  AOI21_X1 U15217 ( .B1(n12127), .B2(n12126), .A(n12415), .ZN(n12130) );
  AOI22_X1 U15218 ( .A1(n19129), .A2(n19825), .B1(n19131), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15219 ( .A1(n19140), .A2(n14761), .ZN(n12128) );
  OAI211_X1 U15220 ( .C1(n12130), .C2(n14779), .A(n12129), .B(n12128), .ZN(
        P2_U2918) );
  NAND2_X1 U15221 ( .A1(n12142), .A2(n12131), .ZN(n12172) );
  OR2_X1 U15222 ( .A1(n12132), .A2(n15905), .ZN(n12133) );
  NAND3_X1 U15223 ( .A1(n12135), .A2(n10345), .A3(n20741), .ZN(n12136) );
  INV_X1 U15224 ( .A(n12207), .ZN(n12151) );
  NAND2_X1 U15225 ( .A1(n12985), .A2(n12162), .ZN(n12138) );
  NAND3_X1 U15226 ( .A1(n12138), .A2(n12629), .A3(n20741), .ZN(n12148) );
  NAND2_X1 U15227 ( .A1(n12973), .A2(n12139), .ZN(n12496) );
  AOI21_X1 U15228 ( .B1(n10338), .B2(n12959), .A(n20101), .ZN(n12140) );
  NAND2_X1 U15229 ( .A1(n12141), .A2(n12140), .ZN(n12156) );
  NAND2_X1 U15230 ( .A1(n12142), .A2(n12156), .ZN(n12143) );
  NOR2_X1 U15231 ( .A1(n12634), .A2(n12145), .ZN(n12146) );
  NOR2_X1 U15232 ( .A1(n12971), .A2(n12146), .ZN(n12147) );
  OAI211_X1 U15233 ( .C1(n12973), .C2(n12148), .A(n12496), .B(n12147), .ZN(
        n12149) );
  INV_X1 U15234 ( .A(n12149), .ZN(n12150) );
  INV_X1 U15235 ( .A(n12442), .ZN(n15864) );
  NOR2_X1 U15236 ( .A1(n20650), .A2(n16180), .ZN(n16184) );
  AOI22_X1 U15237 ( .A1(n12976), .A2(n15864), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n16184), .ZN(n16175) );
  OAI21_X1 U15238 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20355), .A(n16175), 
        .ZN(n16172) );
  INV_X1 U15239 ( .A(n12152), .ZN(n12154) );
  OAI211_X1 U15240 ( .C1(n10344), .C2(n12208), .A(n12173), .B(n12500), .ZN(
        n12153) );
  AOI22_X1 U15241 ( .A1(n12154), .A2(n13646), .B1(n12959), .B2(n12153), .ZN(
        n12159) );
  INV_X1 U15242 ( .A(n12155), .ZN(n12158) );
  NAND4_X1 U15243 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12983) );
  NAND3_X1 U15244 ( .A1(n12162), .A2(n12161), .A3(n12160), .ZN(n12163) );
  NOR2_X1 U15245 ( .A1(n12983), .A2(n12163), .ZN(n12165) );
  NAND2_X1 U15246 ( .A1(n12165), .A2(n12164), .ZN(n14284) );
  AOI22_X1 U15247 ( .A1(n20207), .A2(n14284), .B1(n12166), .B2(n12170), .ZN(
        n15859) );
  INV_X1 U15248 ( .A(n16170), .ZN(n20724) );
  INV_X1 U15249 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U15250 ( .A1(n12170), .A2(n14285), .B1(n20051), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n12167) );
  OAI21_X1 U15251 ( .B1(n15859), .B2(n20724), .A(n12167), .ZN(n12168) );
  NOR2_X1 U15252 ( .A1(n12985), .A2(n12170), .ZN(n15860) );
  AOI22_X1 U15253 ( .A1(n16172), .A2(n12168), .B1(n16170), .B2(n15860), .ZN(
        n12169) );
  OAI21_X1 U15254 ( .B1(n16172), .B2(n12170), .A(n12169), .ZN(P1_U3474) );
  INV_X1 U15255 ( .A(n16172), .ZN(n20726) );
  INV_X1 U15256 ( .A(n14284), .ZN(n12181) );
  NAND2_X1 U15257 ( .A1(n12986), .A2(n12172), .ZN(n12426) );
  INV_X1 U15258 ( .A(n12426), .ZN(n12175) );
  OR2_X1 U15259 ( .A1(n14284), .A2(n12173), .ZN(n12434) );
  XNOR2_X1 U15260 ( .A(n14286), .B(n12174), .ZN(n12182) );
  MUX2_X1 U15261 ( .A(n12175), .B(n12434), .S(n12182), .Z(n12180) );
  NAND2_X1 U15262 ( .A1(n12176), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12178) );
  NOR2_X1 U15263 ( .A1(n12985), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14283) );
  INV_X1 U15264 ( .A(n14283), .ZN(n12177) );
  MUX2_X1 U15265 ( .A(n12178), .B(n12177), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12179) );
  OAI211_X1 U15266 ( .C1(n20479), .C2(n12181), .A(n12180), .B(n12179), .ZN(
        n12422) );
  NOR2_X1 U15267 ( .A1(n20649), .A2(n20051), .ZN(n14289) );
  INV_X1 U15268 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14075) );
  INV_X1 U15269 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20078) );
  OAI22_X1 U15270 ( .A1(n14075), .A2(n20078), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14290) );
  INV_X1 U15271 ( .A(n14290), .ZN(n12183) );
  AOI222_X1 U15272 ( .A1(n12422), .A2(n16170), .B1(n14289), .B2(n12183), .C1(
        n14285), .C2(n12182), .ZN(n12185) );
  NAND2_X1 U15273 ( .A1(n20726), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12184) );
  OAI21_X1 U15274 ( .B1(n20726), .B2(n12185), .A(n12184), .ZN(P1_U3472) );
  NAND2_X1 U15275 ( .A1(n15511), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15479) );
  INV_X1 U15276 ( .A(n15511), .ZN(n12187) );
  NAND2_X1 U15277 ( .A1(n12187), .A2(n19817), .ZN(n12188) );
  NAND2_X1 U15278 ( .A1(n15479), .A2(n12188), .ZN(n19304) );
  NOR2_X1 U15279 ( .A1(n19552), .A2(n19304), .ZN(n12189) );
  AOI21_X1 U15280 ( .B1(n12287), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12189), .ZN(n12190) );
  INV_X1 U15281 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12191) );
  NOR2_X1 U15282 ( .A1(n13363), .A2(n12191), .ZN(n12192) );
  NAND2_X1 U15283 ( .A1(n12194), .A2(n12193), .ZN(n12198) );
  INV_X1 U15284 ( .A(n12195), .ZN(n15443) );
  NAND2_X1 U15285 ( .A1(n15443), .A2(n12196), .ZN(n12197) );
  MUX2_X1 U15286 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n9592), .S(n14652), .Z(n12201) );
  AOI21_X1 U15287 ( .B1(n19812), .B2(n14658), .A(n12201), .ZN(n12202) );
  INV_X1 U15288 ( .A(n12202), .ZN(P2_U2885) );
  NAND2_X1 U15289 ( .A1(n12204), .A2(n12203), .ZN(n12205) );
  NAND2_X1 U15290 ( .A1(n12206), .A2(n12205), .ZN(n13770) );
  AND3_X1 U15291 ( .A1(n20124), .A2(n12976), .A3(n12208), .ZN(n12210) );
  NOR2_X1 U15292 ( .A1(n12500), .A2(n13848), .ZN(n12209) );
  NAND3_X1 U15293 ( .A1(n12211), .A2(n12210), .A3(n12209), .ZN(n12497) );
  NAND2_X1 U15294 ( .A1(n12214), .A2(n12500), .ZN(n12215) );
  NAND2_X2 U15295 ( .A1(n13917), .A2(n12215), .ZN(n13915) );
  INV_X1 U15296 ( .A(n20095), .ZN(n20097) );
  NAND2_X1 U15297 ( .A1(n20097), .A2(DATAI_0_), .ZN(n12217) );
  NAND2_X1 U15298 ( .A1(n20095), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12216) );
  AND2_X1 U15299 ( .A1(n12217), .A2(n12216), .ZN(n20107) );
  INV_X1 U15300 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20848) );
  OAI222_X1 U15301 ( .A1(n13770), .A2(n13915), .B1(n13920), .B2(n20107), .C1(
        n13917), .C2(n20848), .ZN(P1_U2904) );
  OAI21_X1 U15302 ( .B1(n12219), .B2(n12218), .A(n12335), .ZN(n12647) );
  NAND2_X1 U15303 ( .A1(n20097), .A2(DATAI_1_), .ZN(n12221) );
  NAND2_X1 U15304 ( .A1(n20095), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12220) );
  AND2_X1 U15305 ( .A1(n12221), .A2(n12220), .ZN(n20114) );
  INV_X1 U15306 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19985) );
  OAI222_X1 U15307 ( .A1(n12647), .A2(n13915), .B1(n13920), .B2(n20114), .C1(
        n13917), .C2(n19985), .ZN(P1_U2903) );
  INV_X1 U15308 ( .A(n12222), .ZN(n12223) );
  OAI21_X1 U15309 ( .B1(n20022), .B2(n12223), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12229) );
  OR2_X1 U15310 ( .A1(n12224), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U15311 ( .A1(n12226), .A2(n12225), .ZN(n20084) );
  NAND2_X1 U15312 ( .A1(n20021), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20091) );
  OAI21_X1 U15313 ( .B1(n16067), .B2(n20084), .A(n20091), .ZN(n12227) );
  INV_X1 U15314 ( .A(n12227), .ZN(n12228) );
  OAI211_X1 U15315 ( .C1(n13770), .C2(n20098), .A(n12229), .B(n12228), .ZN(
        P1_U2999) );
  AND2_X1 U15316 ( .A1(n20744), .A2(n15905), .ZN(n12230) );
  AND2_X2 U15317 ( .A1(n12259), .A2(n10345), .ZN(n20018) );
  INV_X2 U15318 ( .A(n12259), .ZN(n20017) );
  AOI22_X1 U15319 ( .A1(n20018), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n12232) );
  NAND2_X1 U15320 ( .A1(n12259), .A2(n12959), .ZN(n12261) );
  INV_X1 U15321 ( .A(n20114), .ZN(n13903) );
  NAND2_X1 U15322 ( .A1(n20003), .A2(n13903), .ZN(n12247) );
  NAND2_X1 U15323 ( .A1(n12232), .A2(n12247), .ZN(P1_U2953) );
  AOI22_X1 U15324 ( .A1(n20018), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n12233) );
  INV_X1 U15325 ( .A(n20107), .ZN(n13909) );
  NAND2_X1 U15326 ( .A1(n20003), .A2(n13909), .ZN(n12249) );
  NAND2_X1 U15327 ( .A1(n12233), .A2(n12249), .ZN(P1_U2952) );
  AOI22_X1 U15328 ( .A1(n20018), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U15329 ( .A1(n20097), .A2(DATAI_6_), .ZN(n12235) );
  NAND2_X1 U15330 ( .A1(n20095), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12234) );
  AND2_X1 U15331 ( .A1(n12235), .A2(n12234), .ZN(n20133) );
  INV_X1 U15332 ( .A(n20133), .ZN(n13880) );
  NAND2_X1 U15333 ( .A1(n20003), .A2(n13880), .ZN(n12407) );
  NAND2_X1 U15334 ( .A1(n12236), .A2(n12407), .ZN(P1_U2943) );
  AOI22_X1 U15335 ( .A1(n20018), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n12239) );
  NAND2_X1 U15336 ( .A1(n20097), .A2(DATAI_5_), .ZN(n12238) );
  NAND2_X1 U15337 ( .A1(n20095), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12237) );
  AND2_X1 U15338 ( .A1(n12238), .A2(n12237), .ZN(n20129) );
  INV_X1 U15339 ( .A(n20129), .ZN(n13884) );
  NAND2_X1 U15340 ( .A1(n20003), .A2(n13884), .ZN(n12403) );
  NAND2_X1 U15341 ( .A1(n12239), .A2(n12403), .ZN(P1_U2942) );
  AOI22_X1 U15342 ( .A1(n20018), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U15343 ( .A1(n20097), .A2(DATAI_4_), .ZN(n12241) );
  NAND2_X1 U15344 ( .A1(n20095), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12240) );
  AND2_X1 U15345 ( .A1(n12241), .A2(n12240), .ZN(n20125) );
  INV_X1 U15346 ( .A(n20125), .ZN(n12242) );
  NAND2_X1 U15347 ( .A1(n20003), .A2(n12242), .ZN(n12409) );
  NAND2_X1 U15348 ( .A1(n12243), .A2(n12409), .ZN(P1_U2941) );
  AOI22_X1 U15349 ( .A1(n20018), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U15350 ( .A1(n20097), .A2(DATAI_2_), .ZN(n12245) );
  NAND2_X1 U15351 ( .A1(n20095), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12244) );
  AND2_X1 U15352 ( .A1(n12245), .A2(n12244), .ZN(n20117) );
  INV_X1 U15353 ( .A(n20117), .ZN(n13899) );
  NAND2_X1 U15354 ( .A1(n20003), .A2(n13899), .ZN(n12405) );
  NAND2_X1 U15355 ( .A1(n12246), .A2(n12405), .ZN(P1_U2939) );
  AOI22_X1 U15356 ( .A1(n20018), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n12248) );
  NAND2_X1 U15357 ( .A1(n12248), .A2(n12247), .ZN(P1_U2938) );
  AOI22_X1 U15358 ( .A1(n20018), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U15359 ( .A1(n12250), .A2(n12249), .ZN(P1_U2937) );
  AOI22_X1 U15360 ( .A1(n20018), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n12253) );
  NAND2_X1 U15361 ( .A1(n20097), .A2(DATAI_3_), .ZN(n12252) );
  NAND2_X1 U15362 ( .A1(n20095), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12251) );
  AND2_X1 U15363 ( .A1(n12252), .A2(n12251), .ZN(n20121) );
  INV_X1 U15364 ( .A(n20121), .ZN(n13895) );
  NAND2_X1 U15365 ( .A1(n20003), .A2(n13895), .ZN(n12401) );
  NAND2_X1 U15366 ( .A1(n12253), .A2(n12401), .ZN(P1_U2940) );
  AOI22_X1 U15367 ( .A1(n20018), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U15368 ( .A1(n20097), .A2(DATAI_7_), .ZN(n12255) );
  NAND2_X1 U15369 ( .A1(n20095), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12254) );
  AND2_X1 U15370 ( .A1(n12255), .A2(n12254), .ZN(n20141) );
  INV_X1 U15371 ( .A(n20141), .ZN(n13877) );
  NAND2_X1 U15372 ( .A1(n20003), .A2(n13877), .ZN(n12411) );
  NAND2_X1 U15373 ( .A1(n12256), .A2(n12411), .ZN(P1_U2944) );
  INV_X1 U15374 ( .A(n20018), .ZN(n12400) );
  INV_X1 U15375 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12262) );
  INV_X1 U15376 ( .A(DATAI_15_), .ZN(n12258) );
  INV_X1 U15377 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12257) );
  MUX2_X1 U15378 ( .A(n12258), .B(n12257), .S(n20095), .Z(n13914) );
  INV_X1 U15379 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12260) );
  OAI222_X1 U15380 ( .A1(n12400), .A2(n12262), .B1(n12261), .B2(n13914), .C1(
        n12260), .C2(n12259), .ZN(P1_U2967) );
  INV_X1 U15381 ( .A(n14714), .ZN(n12283) );
  NAND2_X1 U15382 ( .A1(n11738), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15383 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12278) );
  NAND2_X1 U15384 ( .A1(n14358), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15385 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11415), .B1(
        n11402), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15386 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13236), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15387 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n13235), .ZN(n12264) );
  AOI22_X1 U15388 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12600), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U15389 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12275) );
  AOI22_X1 U15390 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15391 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12272) );
  INV_X1 U15392 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U15393 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13229), .ZN(
        n12267) );
  OAI21_X1 U15394 ( .B1(n12722), .B2(n12268), .A(n12267), .ZN(n12269) );
  AOI21_X1 U15395 ( .B1(n13222), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n12269), .ZN(n12271) );
  NAND2_X1 U15396 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12270) );
  NAND4_X1 U15397 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  NAND2_X1 U15398 ( .A1(n12903), .A2(n9633), .ZN(n12276) );
  NAND4_X1 U15399 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12282) );
  AOI222_X1 U15400 ( .A1(n11738), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n11739), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n14358), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n12331) );
  INV_X1 U15401 ( .A(n12280), .ZN(n12281) );
  AOI21_X1 U15402 ( .B1(n12903), .B2(n14343), .A(n12281), .ZN(n12332) );
  OAI21_X1 U15403 ( .B1(n12282), .B2(n9685), .A(n12355), .ZN(n19102) );
  INV_X1 U15404 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20780) );
  OAI222_X1 U15405 ( .A1(n13092), .A2(n12283), .B1(n19102), .B2(n19135), .C1(
        n19144), .C2(n20780), .ZN(P2_U2911) );
  NAND2_X1 U15406 ( .A1(n15479), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12285) );
  NAND2_X1 U15407 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19809), .ZN(
        n19367) );
  INV_X1 U15408 ( .A(n19367), .ZN(n19370) );
  NAND2_X1 U15409 ( .A1(n15511), .A2(n19370), .ZN(n19431) );
  NAND2_X1 U15410 ( .A1(n12285), .A2(n19431), .ZN(n12286) );
  AND2_X1 U15411 ( .A1(n12286), .A2(n19799), .ZN(n19544) );
  AOI21_X1 U15412 ( .B1(n12287), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19544), .ZN(n12288) );
  NOR2_X1 U15413 ( .A1(n13363), .A2(n20842), .ZN(n12290) );
  NAND2_X1 U15414 ( .A1(n12465), .A2(n12290), .ZN(n12568) );
  INV_X1 U15415 ( .A(n12464), .ZN(n12295) );
  NAND2_X1 U15416 ( .A1(n12461), .A2(n12459), .ZN(n12296) );
  INV_X1 U15417 ( .A(n12296), .ZN(n12294) );
  NAND2_X1 U15418 ( .A1(n12295), .A2(n12294), .ZN(n12298) );
  NAND2_X1 U15419 ( .A1(n12464), .A2(n12296), .ZN(n12297) );
  MUX2_X1 U15420 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n14546), .S(n14652), .Z(
        n12300) );
  AOI21_X1 U15421 ( .B1(n19803), .B2(n14658), .A(n12300), .ZN(n12301) );
  INV_X1 U15422 ( .A(n12301), .ZN(P2_U2884) );
  INV_X1 U15423 ( .A(n12302), .ZN(n15467) );
  NAND2_X1 U15424 ( .A1(n14546), .A2(n15467), .ZN(n12316) );
  NOR2_X1 U15425 ( .A1(n16398), .A2(n12303), .ZN(n15458) );
  INV_X1 U15426 ( .A(n12304), .ZN(n12305) );
  NAND2_X1 U15427 ( .A1(n12305), .A2(n11550), .ZN(n15459) );
  INV_X1 U15428 ( .A(n15459), .ZN(n15463) );
  INV_X1 U15429 ( .A(n12308), .ZN(n12309) );
  AOI21_X1 U15430 ( .B1(n12307), .B2(n12309), .A(n13426), .ZN(n12310) );
  OAI21_X1 U15431 ( .B1(n15458), .B2(n15463), .A(n12310), .ZN(n12313) );
  NAND2_X1 U15432 ( .A1(n12307), .A2(n12308), .ZN(n15462) );
  INV_X1 U15433 ( .A(n13426), .ZN(n15460) );
  NAND2_X1 U15434 ( .A1(n12311), .A2(n15460), .ZN(n15464) );
  OAI211_X1 U15435 ( .C1(n15458), .C2(n15459), .A(n15462), .B(n15464), .ZN(
        n12312) );
  MUX2_X1 U15436 ( .A(n12313), .B(n12312), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12314) );
  INV_X1 U15437 ( .A(n12314), .ZN(n12315) );
  NAND2_X1 U15438 ( .A1(n12316), .A2(n12315), .ZN(n16390) );
  AOI22_X1 U15439 ( .A1(n19803), .A2(n16428), .B1(n18952), .B2(n16390), .ZN(
        n12330) );
  NOR2_X1 U15440 ( .A1(n16435), .A2(n14298), .ZN(n16434) );
  NOR2_X1 U15441 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12070), .ZN(n12328) );
  INV_X1 U15442 ( .A(n15473), .ZN(n16404) );
  NAND2_X1 U15443 ( .A1(n12317), .A2(n16404), .ZN(n19147) );
  OR2_X1 U15444 ( .A1(n19147), .A2(n12784), .ZN(n12326) );
  INV_X1 U15445 ( .A(n12318), .ZN(n12323) );
  NAND2_X1 U15446 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  AND4_X1 U15447 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .ZN(
        n12325) );
  NOR2_X1 U15448 ( .A1(n16413), .A2(n19146), .ZN(n12327) );
  AOI211_X2 U15449 ( .C1(n16434), .C2(P2_FLUSH_REG_SCAN_IN), .A(n12328), .B(
        n12327), .ZN(n15474) );
  NAND2_X1 U15450 ( .A1(n15474), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12329) );
  OAI21_X1 U15451 ( .B1(n12330), .B2(n15474), .A(n12329), .ZN(P2_U3596) );
  INV_X1 U15452 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n12334) );
  AOI21_X1 U15453 ( .B1(n12332), .B2(n12331), .A(n9685), .ZN(n16348) );
  INV_X1 U15454 ( .A(n16348), .ZN(n14526) );
  OAI222_X1 U15455 ( .A1(n12334), .A2(n19144), .B1(n14526), .B2(n19135), .C1(
        n13092), .C2(n12333), .ZN(P2_U2912) );
  OAI21_X1 U15456 ( .B1(n10234), .B2(n10695), .A(n12336), .ZN(n12692) );
  INV_X1 U15457 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19983) );
  OAI222_X1 U15458 ( .A1(n12692), .A2(n13915), .B1(n13920), .B2(n20117), .C1(
        n13917), .C2(n19983), .ZN(P1_U2902) );
  AOI22_X1 U15459 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15460 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15461 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15462 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U15463 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12350) );
  AOI22_X1 U15464 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12604), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12348) );
  OR2_X1 U15465 ( .A1(n13211), .A2(n13270), .ZN(n12342) );
  AOI22_X1 U15466 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13122), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12341) );
  OAI211_X1 U15467 ( .C1(n13214), .C2(n12343), .A(n12342), .B(n12341), .ZN(
        n12344) );
  INV_X1 U15468 ( .A(n12344), .ZN(n12347) );
  NAND2_X1 U15469 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15470 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12345) );
  NAND4_X1 U15471 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12349) );
  NOR2_X1 U15472 ( .A1(n12350), .A2(n12349), .ZN(n12671) );
  INV_X1 U15473 ( .A(n12671), .ZN(n12351) );
  AOI22_X1 U15474 ( .A1(n11738), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12903), 
        .B2(n12351), .ZN(n12353) );
  AOI22_X1 U15475 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14358), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U15476 ( .A1(n12354), .A2(n12355), .ZN(n12356) );
  NAND2_X1 U15477 ( .A1(n12356), .A2(n10189), .ZN(n15390) );
  AOI22_X1 U15478 ( .A1(n19140), .A2(n14709), .B1(n19131), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n12357) );
  OAI21_X1 U15479 ( .B1(n19135), .B2(n15390), .A(n12357), .ZN(P2_U2910) );
  AOI22_X1 U15480 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12358) );
  OAI21_X1 U15481 ( .B1(n13889), .B2(n12372), .A(n12358), .ZN(P1_U2916) );
  INV_X1 U15482 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15483 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12359) );
  OAI21_X1 U15484 ( .B1(n12360), .B2(n12372), .A(n12359), .ZN(P1_U2913) );
  INV_X1 U15485 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15486 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12361) );
  OAI21_X1 U15487 ( .B1(n12362), .B2(n12372), .A(n12361), .ZN(P1_U2915) );
  INV_X1 U15488 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15489 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12363) );
  OAI21_X1 U15490 ( .B1(n12364), .B2(n12372), .A(n12363), .ZN(P1_U2919) );
  INV_X1 U15491 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15492 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12365) );
  OAI21_X1 U15493 ( .B1(n12366), .B2(n12372), .A(n12365), .ZN(P1_U2918) );
  INV_X1 U15494 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15495 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12367) );
  OAI21_X1 U15496 ( .B1(n12368), .B2(n12372), .A(n12367), .ZN(P1_U2917) );
  INV_X1 U15497 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15498 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12369) );
  OAI21_X1 U15499 ( .B1(n12370), .B2(n12372), .A(n12369), .ZN(P1_U2914) );
  INV_X1 U15500 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15501 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12371) );
  OAI21_X1 U15502 ( .B1(n12373), .B2(n12372), .A(n12371), .ZN(P1_U2920) );
  INV_X1 U15503 ( .A(n14704), .ZN(n12392) );
  INV_X1 U15504 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15505 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n14358), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15506 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15507 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15508 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15509 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12374) );
  NAND4_X1 U15510 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12386) );
  AOI22_X1 U15511 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13223), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15512 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13236), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12383) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12379) );
  NAND2_X1 U15514 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13229), .ZN(
        n12378) );
  OAI21_X1 U15515 ( .B1(n12722), .B2(n12379), .A(n12378), .ZN(n12380) );
  AOI21_X1 U15516 ( .B1(n13222), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n12380), .ZN(n12382) );
  NAND2_X1 U15517 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12381) );
  NAND4_X1 U15518 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12385) );
  NAND2_X1 U15519 ( .A1(n12903), .A2(n12694), .ZN(n12387) );
  OAI211_X1 U15520 ( .C1(n12675), .C2(n14361), .A(n12388), .B(n12387), .ZN(
        n12389) );
  OR2_X1 U15521 ( .A1(n12389), .A2(n12390), .ZN(n12391) );
  NAND2_X1 U15522 ( .A1(n12391), .A2(n16329), .ZN(n19086) );
  INV_X1 U15523 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19192) );
  OAI222_X1 U15524 ( .A1(n13092), .A2(n12392), .B1(n19086), .B2(n19135), .C1(
        n19144), .C2(n19192), .ZN(P2_U2909) );
  OAI21_X1 U15525 ( .B1(n12394), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12393), .ZN(n12395) );
  INV_X1 U15526 ( .A(n12395), .ZN(n20074) );
  INV_X1 U15527 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n12396) );
  NOR2_X1 U15528 ( .A1(n20068), .A2(n12396), .ZN(n20069) );
  AOI21_X1 U15529 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n20069), .ZN(n12397) );
  OAI21_X1 U15530 ( .B1(n20033), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12397), .ZN(n12398) );
  AOI21_X1 U15531 ( .B1(n20029), .B2(n20074), .A(n12398), .ZN(n12399) );
  OAI21_X1 U15532 ( .B1(n20098), .B2(n12647), .A(n12399), .ZN(P1_U2998) );
  AOI22_X1 U15533 ( .A1(n20018), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15534 ( .A1(n12402), .A2(n12401), .ZN(P1_U2955) );
  AOI22_X1 U15535 ( .A1(n20018), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U15536 ( .A1(n12404), .A2(n12403), .ZN(P1_U2957) );
  AOI22_X1 U15537 ( .A1(n20018), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15538 ( .A1(n12406), .A2(n12405), .ZN(P1_U2954) );
  AOI22_X1 U15539 ( .A1(n20018), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U15540 ( .A1(n12408), .A2(n12407), .ZN(P1_U2958) );
  AOI22_X1 U15541 ( .A1(n20018), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U15542 ( .A1(n12410), .A2(n12409), .ZN(P1_U2956) );
  AOI22_X1 U15543 ( .A1(n20018), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15544 ( .A1(n12412), .A2(n12411), .ZN(P1_U2959) );
  INV_X1 U15545 ( .A(n12413), .ZN(n12414) );
  NOR2_X1 U15546 ( .A1(n12415), .A2(n12414), .ZN(n12418) );
  INV_X1 U15547 ( .A(n19815), .ZN(n12416) );
  NAND2_X1 U15548 ( .A1(n15476), .A2(n12416), .ZN(n12528) );
  OAI21_X1 U15549 ( .B1(n15476), .B2(n12416), .A(n12528), .ZN(n12417) );
  NOR2_X1 U15550 ( .A1(n12417), .A2(n12418), .ZN(n12530) );
  AOI21_X1 U15551 ( .B1(n12418), .B2(n12417), .A(n12530), .ZN(n12421) );
  AOI22_X1 U15552 ( .A1(n19140), .A2(n14752), .B1(n19131), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n12420) );
  NAND2_X1 U15553 ( .A1(n19815), .A2(n19129), .ZN(n12419) );
  OAI211_X1 U15554 ( .C1(n12421), .C2(n14779), .A(n12420), .B(n12419), .ZN(
        P2_U2917) );
  NOR2_X1 U15555 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20649), .ZN(n12444) );
  MUX2_X1 U15556 ( .A(n12422), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n12442), .Z(n15869) );
  AOI22_X1 U15557 ( .A1(n12444), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15869), .B2(n20649), .ZN(n12439) );
  AOI21_X1 U15558 ( .B1(n14286), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12424), .ZN(n12423) );
  NOR2_X1 U15559 ( .A1(n10420), .A2(n12423), .ZN(n20723) );
  AOI21_X1 U15560 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12428), .A(
        n12425), .ZN(n12431) );
  NAND2_X1 U15561 ( .A1(n14283), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12430) );
  MUX2_X1 U15562 ( .A(n12425), .B(n12424), .S(n14286), .Z(n12427) );
  OAI21_X1 U15563 ( .B1(n12428), .B2(n12427), .A(n12426), .ZN(n12429) );
  OAI211_X1 U15564 ( .C1(n12431), .C2(n12985), .A(n12430), .B(n12429), .ZN(
        n12432) );
  INV_X1 U15565 ( .A(n12432), .ZN(n12433) );
  OAI21_X1 U15566 ( .B1(n12434), .B2(n20723), .A(n12433), .ZN(n12435) );
  AOI21_X1 U15567 ( .B1(n20103), .B2(n14284), .A(n12435), .ZN(n20725) );
  OR2_X1 U15568 ( .A1(n12442), .A2(n20725), .ZN(n12437) );
  NAND2_X1 U15569 ( .A1(n12442), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12436) );
  NAND2_X1 U15570 ( .A1(n12437), .A2(n12436), .ZN(n15870) );
  AOI22_X1 U15571 ( .A1(n15870), .A2(n20649), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12444), .ZN(n12438) );
  OR2_X1 U15572 ( .A1(n12439), .A2(n12438), .ZN(n15874) );
  INV_X1 U15573 ( .A(n12164), .ZN(n16171) );
  INV_X1 U15574 ( .A(n20234), .ZN(n20478) );
  XNOR2_X1 U15575 ( .A(n12440), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19935) );
  AOI21_X1 U15576 ( .B1(n16171), .B2(n19935), .A(n12442), .ZN(n12441) );
  AOI211_X1 U15577 ( .C1(n12442), .C2(n16173), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n12441), .ZN(n12443) );
  AOI21_X1 U15578 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n12444), .A(
        n12443), .ZN(n15880) );
  OAI21_X1 U15579 ( .B1(n15874), .B2(n14287), .A(n15880), .ZN(n12478) );
  OAI21_X1 U15580 ( .B1(n12478), .B2(P1_FLUSH_REG_SCAN_IN), .A(n16184), .ZN(
        n12445) );
  NOR2_X1 U15581 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20745) );
  INV_X1 U15582 ( .A(n20745), .ZN(n16176) );
  NAND2_X1 U15583 ( .A1(n12445), .A2(n20148), .ZN(n20093) );
  AND2_X1 U15584 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20355), .ZN(n14279) );
  OR2_X1 U15585 ( .A1(n9587), .A2(n20587), .ZN(n12447) );
  NAND2_X1 U15586 ( .A1(n20510), .A2(n20542), .ZN(n20476) );
  NAND2_X1 U15587 ( .A1(n12447), .A2(n20476), .ZN(n20446) );
  OAI21_X1 U15588 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9587), .A(n20446), 
        .ZN(n12448) );
  OAI21_X1 U15589 ( .B1(n14279), .B2(n20540), .A(n12448), .ZN(n12449) );
  NAND2_X1 U15590 ( .A1(n20093), .A2(n12449), .ZN(n12450) );
  OAI21_X1 U15591 ( .B1(n20093), .B2(n10622), .A(n12450), .ZN(P1_U3477) );
  OAI21_X1 U15592 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12762) );
  INV_X1 U15593 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19981) );
  OAI222_X1 U15594 ( .A1(n12762), .A2(n13915), .B1(n13920), .B2(n20121), .C1(
        n13917), .C2(n19981), .ZN(P1_U2901) );
  NOR2_X1 U15595 ( .A1(n20479), .A2(n14279), .ZN(n12456) );
  INV_X1 U15596 ( .A(n9587), .ZN(n14274) );
  NAND2_X1 U15597 ( .A1(n20510), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20514) );
  NOR2_X1 U15598 ( .A1(n14274), .A2(n20514), .ZN(n20593) );
  MUX2_X1 U15599 ( .A(n20593), .B(n20446), .S(n12454), .Z(n12455) );
  OAI21_X1 U15600 ( .B1(n12456), .B2(n12455), .A(n20093), .ZN(n12457) );
  OAI21_X1 U15601 ( .B1(n10625), .B2(n20093), .A(n12457), .ZN(P1_U3476) );
  NAND2_X1 U15602 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15494), .ZN(
        n12458) );
  INV_X1 U15603 ( .A(n12458), .ZN(n12463) );
  AND2_X1 U15604 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  NAND2_X1 U15605 ( .A1(n12461), .A2(n12460), .ZN(n12462) );
  INV_X1 U15606 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12466) );
  NOR2_X1 U15607 ( .A1(n13363), .A2(n12466), .ZN(n12569) );
  XNOR2_X1 U15608 ( .A(n12546), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12477) );
  INV_X1 U15609 ( .A(n12472), .ZN(n12470) );
  INV_X1 U15610 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n14518) );
  INV_X1 U15611 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16345) );
  OR2_X1 U15612 ( .A1(n11329), .A2(n16345), .ZN(n12468) );
  AOI22_X1 U15613 ( .A1(n14308), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12467) );
  OAI211_X1 U15614 ( .C1(n13540), .C2(n14518), .A(n12468), .B(n12467), .ZN(
        n12471) );
  INV_X1 U15615 ( .A(n12471), .ZN(n12469) );
  NAND2_X1 U15616 ( .A1(n12470), .A2(n12469), .ZN(n12473) );
  AND2_X1 U15617 ( .A1(n12473), .A2(n12544), .ZN(n16349) );
  INV_X1 U15618 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12474) );
  NOR2_X1 U15619 ( .A1(n14652), .A2(n12474), .ZN(n12475) );
  AOI21_X1 U15620 ( .B1(n16349), .B2(n14652), .A(n12475), .ZN(n12476) );
  OAI21_X1 U15621 ( .B1(n12477), .B2(n14677), .A(n12476), .ZN(P2_U2880) );
  NOR2_X1 U15622 ( .A1(n12478), .A2(n16180), .ZN(n15890) );
  OAI22_X1 U15623 ( .A1(n10688), .A2(n20587), .B1(n13768), .B2(n14279), .ZN(
        n12479) );
  OAI21_X1 U15624 ( .B1(n15890), .B2(n12479), .A(n20093), .ZN(n12480) );
  OAI21_X1 U15625 ( .B1(n20093), .B2(n20509), .A(n12480), .ZN(P1_U3478) );
  INV_X1 U15626 ( .A(n12481), .ZN(n12685) );
  INV_X1 U15627 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12482) );
  OAI22_X1 U15628 ( .A1(n14062), .A2(n12482), .B1(n20068), .B2(n20067), .ZN(
        n12483) );
  AOI21_X1 U15629 ( .B1(n12685), .B2(n16064), .A(n12483), .ZN(n12488) );
  OR2_X1 U15630 ( .A1(n12485), .A2(n12484), .ZN(n20062) );
  NAND3_X1 U15631 ( .A1(n20062), .A2(n12486), .A3(n20029), .ZN(n12487) );
  OAI211_X1 U15632 ( .C1(n12692), .C2(n20098), .A(n12488), .B(n12487), .ZN(
        P1_U2997) );
  INV_X1 U15633 ( .A(n16290), .ZN(n12495) );
  NOR2_X1 U15634 ( .A1(n12489), .A2(n12490), .ZN(n12492) );
  INV_X1 U15635 ( .A(n12546), .ZN(n12491) );
  OAI211_X1 U15636 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12492), .A(
        n12491), .B(n14658), .ZN(n12494) );
  NAND2_X1 U15637 ( .A1(n14659), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12493) );
  OAI211_X1 U15638 ( .C1(n12495), .C2(n14659), .A(n12494), .B(n12493), .ZN(
        P2_U2881) );
  OR2_X1 U15639 ( .A1(n12497), .A2(n13544), .ZN(n12498) );
  MUX2_X1 U15640 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12503) );
  OR2_X1 U15641 ( .A1(n13593), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12502) );
  NAND2_X1 U15642 ( .A1(n12503), .A2(n12502), .ZN(n12507) );
  INV_X1 U15644 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12504) );
  OR2_X1 U15645 ( .A1(n13579), .A2(n12504), .ZN(n12506) );
  NAND2_X1 U15646 ( .A1(n13646), .A2(n12504), .ZN(n12505) );
  NAND2_X1 U15647 ( .A1(n12506), .A2(n12505), .ZN(n12518) );
  XNOR2_X1 U15648 ( .A(n12507), .B(n12518), .ZN(n12645) );
  AOI21_X1 U15649 ( .B1(n12645), .B2(n13585), .A(n12507), .ZN(n12522) );
  INV_X1 U15650 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U15651 ( .A1(n13044), .A2(n12524), .ZN(n12512) );
  NAND2_X1 U15652 ( .A1(n13585), .A2(n12524), .ZN(n12510) );
  NAND2_X1 U15653 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12509) );
  NAND3_X1 U15654 ( .A1(n12510), .A2(n13579), .A3(n12509), .ZN(n12511) );
  AND2_X1 U15655 ( .A1(n12512), .A2(n12511), .ZN(n12521) );
  NAND2_X1 U15656 ( .A1(n12522), .A2(n12521), .ZN(n19931) );
  NAND2_X1 U15657 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12513) );
  NAND2_X1 U15658 ( .A1(n13579), .A2(n12513), .ZN(n12515) );
  INV_X1 U15659 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U15660 ( .A1(n13585), .A2(n12517), .ZN(n12514) );
  NAND2_X1 U15661 ( .A1(n12515), .A2(n12514), .ZN(n12516) );
  OAI21_X1 U15662 ( .B1(n13596), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12516), .ZN(
        n12663) );
  INV_X1 U15663 ( .A(n12663), .ZN(n19930) );
  XNOR2_X1 U15664 ( .A(n19931), .B(n19930), .ZN(n12648) );
  OAI222_X1 U15665 ( .A1(n12762), .A2(n16020), .B1(n19954), .B2(n12648), .C1(
        n13839), .C2(n12517), .ZN(P1_U2869) );
  INV_X1 U15666 ( .A(n12518), .ZN(n12520) );
  OR2_X1 U15667 ( .A1(n13593), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12519) );
  NAND2_X1 U15668 ( .A1(n12520), .A2(n12519), .ZN(n20082) );
  OAI222_X1 U15669 ( .A1(n13770), .A2(n16020), .B1(n13839), .B2(n12504), .C1(
        n20082), .C2(n19954), .ZN(P1_U2872) );
  OR2_X1 U15670 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  AND2_X1 U15671 ( .A1(n12523), .A2(n19931), .ZN(n20053) );
  INV_X1 U15672 ( .A(n20053), .ZN(n12525) );
  OAI22_X1 U15673 ( .A1(n19954), .A2(n12525), .B1(n12524), .B2(n13839), .ZN(
        n12526) );
  INV_X1 U15674 ( .A(n12526), .ZN(n12527) );
  OAI21_X1 U15675 ( .B1(n12692), .B2(n16020), .A(n12527), .ZN(P1_U2870) );
  INV_X1 U15676 ( .A(n12528), .ZN(n12529) );
  NOR2_X1 U15677 ( .A1(n12530), .A2(n12529), .ZN(n12533) );
  XNOR2_X1 U15678 ( .A(n12531), .B(n9708), .ZN(n19797) );
  XNOR2_X1 U15679 ( .A(n19803), .B(n19797), .ZN(n12532) );
  NOR2_X1 U15680 ( .A1(n12533), .A2(n12532), .ZN(n12566) );
  AOI21_X1 U15681 ( .B1(n12533), .B2(n12532), .A(n12566), .ZN(n12536) );
  AOI22_X1 U15682 ( .A1(n19140), .A2(n14742), .B1(n19131), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15683 ( .A1(n19797), .A2(n19129), .ZN(n12534) );
  OAI211_X1 U15684 ( .C1(n12536), .C2(n14779), .A(n12535), .B(n12534), .ZN(
        P2_U2916) );
  INV_X1 U15685 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15416) );
  OR2_X1 U15686 ( .A1(n11329), .A2(n15416), .ZN(n12542) );
  INV_X1 U15687 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12539) );
  NAND2_X1 U15688 ( .A1(n14307), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15689 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12537) );
  OAI211_X1 U15690 ( .C1(n12539), .C2(n13534), .A(n12538), .B(n12537), .ZN(
        n12540) );
  INV_X1 U15691 ( .A(n12540), .ZN(n12541) );
  AND2_X1 U15692 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  OR2_X1 U15693 ( .A1(n12545), .A2(n12553), .ZN(n15412) );
  OAI211_X1 U15694 ( .C1(n9710), .C2(n9633), .A(n14658), .B(n12672), .ZN(
        n12548) );
  NAND2_X1 U15695 ( .A1(n14659), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12547) );
  OAI211_X1 U15696 ( .C1(n15412), .C2(n14659), .A(n12548), .B(n12547), .ZN(
        P2_U2879) );
  XNOR2_X1 U15697 ( .A(n12672), .B(n12671), .ZN(n12556) );
  INV_X1 U15698 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12551) );
  INV_X1 U15699 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15397) );
  OR2_X1 U15700 ( .A1(n11329), .A2(n15397), .ZN(n12550) );
  AOI22_X1 U15701 ( .A1(n14308), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12549) );
  OAI211_X1 U15702 ( .C1(n13540), .C2(n12551), .A(n12550), .B(n12549), .ZN(
        n12552) );
  NOR2_X1 U15703 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  OR2_X1 U15704 ( .A1(n12697), .A2(n12554), .ZN(n15387) );
  INV_X1 U15705 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14509) );
  MUX2_X1 U15706 ( .A(n15387), .B(n14509), .S(n14659), .Z(n12555) );
  OAI21_X1 U15707 ( .B1(n12556), .B2(n14677), .A(n12555), .ZN(P2_U2878) );
  INV_X1 U15708 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19979) );
  XNOR2_X1 U15709 ( .A(n12451), .B(n10715), .ZN(n20027) );
  INV_X1 U15710 ( .A(n20027), .ZN(n12558) );
  OAI222_X1 U15711 ( .A1(n13917), .A2(n19979), .B1(n13920), .B2(n20125), .C1(
        n13915), .C2(n12558), .ZN(P1_U2900) );
  OAI21_X1 U15712 ( .B1(n12559), .B2(n12561), .A(n12560), .ZN(n16354) );
  NOR2_X1 U15713 ( .A1(n19803), .A2(n19797), .ZN(n12565) );
  INV_X1 U15714 ( .A(n12559), .ZN(n12562) );
  OAI21_X1 U15715 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n19106) );
  OAI21_X1 U15716 ( .B1(n12566), .B2(n12565), .A(n19106), .ZN(n13091) );
  INV_X1 U15717 ( .A(n14779), .ZN(n16233) );
  INV_X1 U15718 ( .A(n12567), .ZN(n12572) );
  INV_X1 U15719 ( .A(n12569), .ZN(n12570) );
  NAND2_X1 U15720 ( .A1(n12568), .A2(n12570), .ZN(n12571) );
  OAI21_X1 U15721 ( .B1(n12572), .B2(n12571), .A(n12489), .ZN(n13102) );
  INV_X1 U15722 ( .A(n13102), .ZN(n19117) );
  NAND3_X1 U15723 ( .A1(n13091), .A2(n16233), .A3(n19117), .ZN(n12574) );
  AOI22_X1 U15724 ( .A1(n19140), .A2(n14728), .B1(n19131), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12573) );
  OAI211_X1 U15725 ( .C1(n19135), .C2(n16354), .A(n12574), .B(n12573), .ZN(
        P2_U2914) );
  NAND2_X1 U15726 ( .A1(n11738), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U15727 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12590) );
  NAND2_X1 U15728 ( .A1(n14358), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15729 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13209), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15730 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15731 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15732 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12575) );
  NAND4_X1 U15733 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12587) );
  AOI22_X1 U15734 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12585) );
  INV_X1 U15735 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15736 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13229), .ZN(
        n12579) );
  OAI21_X1 U15737 ( .B1(n12722), .B2(n12580), .A(n12579), .ZN(n12581) );
  AOI21_X1 U15738 ( .B1(n11415), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n12581), .ZN(n12584) );
  AOI22_X1 U15739 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12583) );
  NAND2_X1 U15740 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12582) );
  NAND4_X1 U15741 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12586) );
  NAND2_X1 U15742 ( .A1(n12903), .A2(n12705), .ZN(n12588) );
  NAND4_X1 U15743 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n12619) );
  INV_X1 U15744 ( .A(n12592), .ZN(n13160) );
  INV_X1 U15745 ( .A(n13235), .ZN(n13159) );
  OAI22_X1 U15746 ( .A1(n13160), .A2(n13326), .B1(n13159), .B2(n12593), .ZN(
        n12596) );
  INV_X1 U15747 ( .A(n13223), .ZN(n13162) );
  INV_X1 U15748 ( .A(n12594), .ZN(n13161) );
  OAI22_X1 U15749 ( .A1(n13162), .A2(n15541), .B1(n13161), .B2(n13327), .ZN(
        n12595) );
  NOR2_X1 U15750 ( .A1(n12596), .A2(n12595), .ZN(n12616) );
  INV_X1 U15751 ( .A(n12597), .ZN(n13180) );
  INV_X1 U15752 ( .A(n12598), .ZN(n13179) );
  OAI22_X1 U15753 ( .A1(n13180), .A2(n13328), .B1(n13179), .B2(n13329), .ZN(
        n12603) );
  INV_X1 U15754 ( .A(n12599), .ZN(n13182) );
  INV_X1 U15755 ( .A(n12600), .ZN(n13181) );
  OAI22_X1 U15756 ( .A1(n13182), .A2(n12601), .B1(n13181), .B2(n13149), .ZN(
        n12602) );
  NOR2_X1 U15757 ( .A1(n12603), .A2(n12602), .ZN(n12615) );
  NAND2_X1 U15758 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U15759 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12608) );
  NAND2_X1 U15760 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12607) );
  INV_X1 U15761 ( .A(n12604), .ZN(n12605) );
  INV_X1 U15762 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20842) );
  OR2_X1 U15763 ( .A1(n12605), .A2(n20842), .ZN(n12606) );
  AND4_X1 U15764 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12614) );
  OR2_X1 U15765 ( .A1(n13211), .A2(n13320), .ZN(n12611) );
  AOI22_X1 U15766 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13122), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12610) );
  OAI211_X1 U15767 ( .C1(n13214), .C2(n13158), .A(n12611), .B(n12610), .ZN(
        n12612) );
  INV_X1 U15768 ( .A(n12612), .ZN(n12613) );
  NAND4_X1 U15769 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12702) );
  AOI22_X1 U15770 ( .A1(n11738), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n12903), 
        .B2(n12702), .ZN(n12618) );
  AOI22_X1 U15771 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n14358), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12617) );
  OAI21_X1 U15772 ( .B1(n12619), .B2(n16328), .A(n14493), .ZN(n19061) );
  INV_X1 U15773 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19187) );
  OAI222_X1 U15774 ( .A1(n13092), .A2(n12620), .B1(n19061), .B2(n19135), .C1(
        n19144), .C2(n19187), .ZN(P2_U2907) );
  NAND3_X1 U15775 ( .A1(n20650), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n13622), 
        .ZN(n12621) );
  NAND3_X1 U15776 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_3__SCAN_IN), .A3(n20745), .ZN(n15895) );
  NAND3_X1 U15777 ( .A1(n20068), .A2(n12621), .A3(n15895), .ZN(n12622) );
  INV_X1 U15778 ( .A(n12623), .ZN(n12624) );
  NAND2_X1 U15779 ( .A1(n12624), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13599) );
  INV_X1 U15780 ( .A(n13599), .ZN(n12625) );
  NAND2_X1 U15781 ( .A1(n12625), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12626) );
  INV_X1 U15782 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13638) );
  XNOR2_X1 U15783 ( .A(n12626), .B(n13638), .ZN(n13925) );
  NOR2_X1 U15784 ( .A1(n13925), .A2(n20649), .ZN(n12627) );
  OAI21_X1 U15785 ( .B1(n12635), .B2(n12628), .A(n15943), .ZN(n19942) );
  INV_X1 U15786 ( .A(n19942), .ZN(n13771) );
  NOR2_X1 U15787 ( .A1(n12635), .A2(n20101), .ZN(n12637) );
  OAI21_X1 U15788 ( .B1(n12959), .B2(n12629), .A(n20741), .ZN(n12962) );
  NOR2_X1 U15789 ( .A1(n12962), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12636) );
  AND2_X1 U15790 ( .A1(n13585), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12631) );
  NOR2_X1 U15791 ( .A1(n12636), .A2(n12631), .ZN(n12630) );
  NAND2_X1 U15792 ( .A1(n20741), .A2(n20542), .ZN(n15884) );
  NAND2_X1 U15793 ( .A1(n12631), .A2(n15884), .ZN(n12632) );
  NOR2_X2 U15794 ( .A1(n12635), .A2(n12632), .ZN(n19914) );
  AND2_X1 U15795 ( .A1(n19914), .A2(n12645), .ZN(n12643) );
  AND2_X1 U15796 ( .A1(n13925), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12633) );
  NOR2_X1 U15797 ( .A1(n12635), .A2(n12634), .ZN(n19936) );
  INV_X1 U15798 ( .A(n20540), .ZN(n20544) );
  NAND2_X1 U15799 ( .A1(n19936), .A2(n20544), .ZN(n12641) );
  INV_X1 U15800 ( .A(n19889), .ZN(n12952) );
  INV_X1 U15801 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12638) );
  OAI22_X1 U15802 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n19890), .B1(n12638), 
        .B2(n19926), .ZN(n12639) );
  AOI21_X1 U15803 ( .B1(n12952), .B2(P1_REIP_REG_1__SCAN_IN), .A(n12639), .ZN(
        n12640) );
  OAI211_X1 U15804 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19948), .A(
        n12641), .B(n12640), .ZN(n12642) );
  AOI211_X1 U15805 ( .C1(P1_EBX_REG_1__SCAN_IN), .C2(n19934), .A(n12643), .B(
        n12642), .ZN(n12644) );
  OAI21_X1 U15806 ( .B1(n13771), .B2(n12647), .A(n12644), .ZN(P1_U2839) );
  XNOR2_X1 U15807 ( .A(n12645), .B(n13585), .ZN(n20070) );
  AOI22_X1 U15808 ( .A1(n19950), .A2(n20070), .B1(n13828), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n12646) );
  OAI21_X1 U15809 ( .B1(n16020), .B2(n12647), .A(n12646), .ZN(P1_U2871) );
  INV_X1 U15810 ( .A(n12648), .ZN(n20044) );
  AOI22_X1 U15811 ( .A1(n19914), .A2(n20044), .B1(n19936), .B2(n20103), .ZN(
        n12651) );
  OAI221_X1 U15812 ( .B1(n19890), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19890), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n19889), .ZN(n12649) );
  AOI22_X1 U15813 ( .A1(n19901), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n12649), .ZN(n12650) );
  OAI211_X1 U15814 ( .C1(n12758), .C2(n19948), .A(n12651), .B(n12650), .ZN(
        n12653) );
  INV_X1 U15815 ( .A(n19890), .ZN(n19923) );
  INV_X1 U15816 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20675) );
  AND4_X1 U15817 ( .A1(n19923), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n20675), .A4(
        P1_REIP_REG_1__SCAN_IN), .ZN(n12652) );
  AOI211_X1 U15818 ( .C1(P1_EBX_REG_3__SCAN_IN), .C2(n19934), .A(n12653), .B(
        n12652), .ZN(n12654) );
  OAI21_X1 U15819 ( .B1(n13771), .B2(n12762), .A(n12654), .ZN(P1_U2837) );
  NAND2_X1 U15820 ( .A1(n12656), .A2(n12655), .ZN(n12657) );
  INV_X1 U15821 ( .A(n19918), .ZN(n12670) );
  OAI222_X1 U15822 ( .A1(n12670), .A2(n13915), .B1(n13920), .B2(n20129), .C1(
        n13917), .C2(n10720), .ZN(P1_U2899) );
  INV_X1 U15823 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U15824 ( .A1(n13044), .A2(n19958), .ZN(n12662) );
  NAND2_X1 U15825 ( .A1(n13585), .A2(n19958), .ZN(n12660) );
  NAND2_X1 U15826 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12659) );
  NAND3_X1 U15827 ( .A1(n12660), .A2(n13579), .A3(n12659), .ZN(n12661) );
  AND2_X1 U15828 ( .A1(n12662), .A2(n12661), .ZN(n19928) );
  NAND2_X1 U15829 ( .A1(n12663), .A2(n19928), .ZN(n12664) );
  NAND2_X1 U15830 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12665) );
  NAND2_X1 U15831 ( .A1(n13579), .A2(n12665), .ZN(n12667) );
  INV_X1 U15832 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n12669) );
  NAND2_X1 U15833 ( .A1(n13585), .A2(n12669), .ZN(n12666) );
  NAND2_X1 U15834 ( .A1(n12667), .A2(n12666), .ZN(n12668) );
  OAI21_X1 U15835 ( .B1(n13596), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12668), .ZN(
        n16149) );
  XNOR2_X1 U15836 ( .A(n19932), .B(n16149), .ZN(n19913) );
  INV_X1 U15837 ( .A(n19913), .ZN(n16162) );
  OAI222_X1 U15838 ( .A1(n12670), .A2(n16020), .B1(n19954), .B2(n16162), .C1(
        n12669), .C2(n13839), .ZN(P1_U2867) );
  XNOR2_X1 U15839 ( .A(n12704), .B(n12702), .ZN(n12683) );
  INV_X1 U15840 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15374) );
  OR2_X1 U15841 ( .A1(n11329), .A2(n15374), .ZN(n12674) );
  AOI22_X1 U15842 ( .A1(n14308), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12673) );
  OAI211_X1 U15843 ( .C1(n13540), .C2(n12675), .A(n12674), .B(n12673), .ZN(
        n12696) );
  INV_X1 U15844 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12678) );
  INV_X1 U15845 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16336) );
  OR2_X1 U15846 ( .A1(n11329), .A2(n16336), .ZN(n12677) );
  AOI22_X1 U15847 ( .A1(n14308), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12676) );
  OAI211_X1 U15848 ( .C1(n13540), .C2(n12678), .A(n12677), .B(n12676), .ZN(
        n12679) );
  OR2_X1 U15849 ( .A1(n12699), .A2(n12679), .ZN(n12680) );
  AND2_X1 U15850 ( .A1(n12680), .A2(n12709), .ZN(n19071) );
  INV_X1 U15851 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19068) );
  NOR2_X1 U15852 ( .A1(n14652), .A2(n19068), .ZN(n12681) );
  AOI21_X1 U15853 ( .B1(n19071), .B2(n14652), .A(n12681), .ZN(n12682) );
  OAI21_X1 U15854 ( .B1(n12683), .B2(n14677), .A(n12682), .ZN(P2_U2876) );
  INV_X1 U15855 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20067) );
  NAND3_X1 U15856 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n19923), .A3(n20067), 
        .ZN(n12691) );
  INV_X1 U15857 ( .A(n20479), .ZN(n20348) );
  AOI22_X1 U15858 ( .A1(n19914), .A2(n20053), .B1(n19936), .B2(n20348), .ZN(
        n12689) );
  NAND2_X1 U15859 ( .A1(n19934), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12688) );
  OAI21_X1 U15860 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19890), .A(n19889), .ZN(
        n12684) );
  AOI22_X1 U15861 ( .A1(n19901), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n12684), .ZN(n12687) );
  NAND2_X1 U15862 ( .A1(n19879), .A2(n12685), .ZN(n12686) );
  AND4_X1 U15863 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12690) );
  OAI211_X1 U15864 ( .C1(n13771), .C2(n12692), .A(n12691), .B(n12690), .ZN(
        P1_U2838) );
  INV_X1 U15865 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n20801) );
  INV_X1 U15866 ( .A(n12704), .ZN(n12693) );
  OAI211_X1 U15867 ( .C1(n12695), .C2(n12694), .A(n12693), .B(n14658), .ZN(
        n12701) );
  NOR2_X1 U15868 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  OR2_X1 U15869 ( .A1(n12699), .A2(n12698), .ZN(n15109) );
  INV_X1 U15870 ( .A(n15109), .ZN(n19082) );
  NAND2_X1 U15871 ( .A1(n19082), .A2(n14652), .ZN(n12700) );
  OAI211_X1 U15872 ( .C1(n14652), .C2(n20801), .A(n12701), .B(n12700), .ZN(
        P2_U2877) );
  INV_X1 U15873 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12713) );
  AND2_X1 U15874 ( .A1(n12704), .A2(n12702), .ZN(n12706) );
  AND2_X1 U15875 ( .A1(n12702), .A2(n12705), .ZN(n12703) );
  OAI211_X1 U15876 ( .C1(n12706), .C2(n12705), .A(n14658), .B(n12909), .ZN(
        n12712) );
  INV_X1 U15877 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15097) );
  OAI22_X1 U15878 ( .A1(n13534), .A2(n12713), .B1(n13505), .B2(n15097), .ZN(
        n12708) );
  INV_X1 U15879 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16322) );
  NOR2_X1 U15880 ( .A1(n11329), .A2(n16322), .ZN(n12707) );
  AOI211_X1 U15881 ( .C1(n14307), .C2(P2_REIP_REG_12__SCAN_IN), .A(n12708), 
        .B(n12707), .ZN(n12710) );
  AOI21_X1 U15882 ( .B1(n12710), .B2(n12709), .A(n14489), .ZN(n19057) );
  NAND2_X1 U15883 ( .A1(n19057), .A2(n14652), .ZN(n12711) );
  OAI211_X1 U15884 ( .C1(n14652), .C2(n12713), .A(n12712), .B(n12711), .ZN(
        P2_U2875) );
  INV_X1 U15885 ( .A(n19951), .ZN(n12715) );
  OAI222_X1 U15886 ( .A1(n13915), .A2(n12715), .B1(n13920), .B2(n20133), .C1(
        n13917), .C2(n10730), .ZN(P1_U2898) );
  INV_X1 U15887 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U15888 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n14358), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15889 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13209), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15890 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15891 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12600), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15892 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13236), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12716) );
  NAND4_X1 U15893 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n12729) );
  AOI22_X1 U15894 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15895 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13229), .ZN(
        n12720) );
  OAI21_X1 U15896 ( .B1(n12722), .B2(n12721), .A(n12720), .ZN(n12723) );
  AOI21_X1 U15897 ( .B1(n11415), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n12723), .ZN(n12726) );
  AOI22_X1 U15898 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12604), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U15899 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12724) );
  NAND4_X1 U15900 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12728) );
  NOR2_X1 U15901 ( .A1(n12729), .A2(n12728), .ZN(n12910) );
  INV_X1 U15902 ( .A(n12910), .ZN(n12730) );
  NAND2_X1 U15903 ( .A1(n12903), .A2(n12730), .ZN(n12731) );
  OAI211_X1 U15904 ( .C1(n14361), .C2(n12920), .A(n12732), .B(n12731), .ZN(
        n12750) );
  INV_X1 U15905 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16244) );
  NOR2_X1 U15906 ( .A1(n12888), .A2(n16244), .ZN(n12749) );
  INV_X1 U15907 ( .A(n12903), .ZN(n12747) );
  AOI22_X1 U15908 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15909 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15910 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15911 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12733) );
  NAND4_X1 U15912 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12746) );
  AOI22_X1 U15913 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12744) );
  OR2_X1 U15914 ( .A1(n13211), .A2(n13369), .ZN(n12738) );
  AOI22_X1 U15915 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13122), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12737) );
  OAI211_X1 U15916 ( .C1(n13214), .C2(n12739), .A(n12738), .B(n12737), .ZN(
        n12740) );
  INV_X1 U15917 ( .A(n12740), .ZN(n12743) );
  NAND2_X1 U15918 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12742) );
  NAND2_X1 U15919 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12741) );
  NAND4_X1 U15920 ( .A1(n12744), .A2(n12743), .A3(n12742), .A4(n12741), .ZN(
        n12745) );
  NOR2_X1 U15921 ( .A1(n12746), .A2(n12745), .ZN(n14675) );
  INV_X1 U15922 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n14499) );
  OAI22_X1 U15923 ( .A1(n12747), .A2(n14675), .B1(n14361), .B2(n14499), .ZN(
        n12748) );
  AOI211_X1 U15924 ( .C1(P2_EAX_REG_13__SCAN_IN), .C2(n11719), .A(n12749), .B(
        n12748), .ZN(n14494) );
  OR2_X1 U15925 ( .A1(n12750), .A2(n9688), .ZN(n12752) );
  NAND2_X1 U15926 ( .A1(n12752), .A2(n12751), .ZN(n19049) );
  INV_X1 U15927 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19184) );
  OAI222_X1 U15928 ( .A1(n13092), .A2(n12753), .B1(n19049), .B2(n19135), .C1(
        n19144), .C2(n19184), .ZN(P2_U2905) );
  OAI21_X1 U15929 ( .B1(n12756), .B2(n12755), .A(n12754), .ZN(n12757) );
  INV_X1 U15930 ( .A(n12757), .ZN(n20045) );
  NAND2_X1 U15931 ( .A1(n20045), .A2(n20029), .ZN(n12761) );
  AND2_X1 U15932 ( .A1(n20021), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20043) );
  NOR2_X1 U15933 ( .A1(n20033), .A2(n12758), .ZN(n12759) );
  AOI211_X1 U15934 ( .C1(n20022), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20043), .B(n12759), .ZN(n12760) );
  OAI211_X1 U15935 ( .C1(n20098), .C2(n12762), .A(n12761), .B(n12760), .ZN(
        P1_U2996) );
  NAND2_X1 U15936 ( .A1(n12764), .A2(n12763), .ZN(n12766) );
  XNOR2_X1 U15937 ( .A(n12766), .B(n12765), .ZN(n12783) );
  INV_X1 U15938 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19745) );
  NOR2_X1 U15939 ( .A1(n19745), .A2(n11795), .ZN(n12767) );
  AOI21_X1 U15940 ( .B1(n12768), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12767), .ZN(n12770) );
  NAND2_X1 U15941 ( .A1(n19797), .A2(n16371), .ZN(n12769) );
  OAI211_X1 U15942 ( .C1(n16309), .C2(n11363), .A(n12770), .B(n12769), .ZN(
        n12771) );
  AOI21_X1 U15943 ( .B1(n12773), .B2(n12772), .A(n12771), .ZN(n12776) );
  NAND2_X1 U15944 ( .A1(n11653), .A2(n12774), .ZN(n12779) );
  NAND3_X1 U15945 ( .A1(n12780), .A2(n12779), .A3(n16358), .ZN(n12775) );
  OAI211_X1 U15946 ( .C1(n12783), .C2(n16373), .A(n12776), .B(n12775), .ZN(
        P2_U3043) );
  AOI21_X1 U15947 ( .B1(n14541), .B2(n12787), .A(n12789), .ZN(n14539) );
  OAI22_X1 U15948 ( .A1(n14541), .A2(n16305), .B1(n19745), .B2(n11795), .ZN(
        n12778) );
  NOR2_X1 U15949 ( .A1(n11363), .A2(n15115), .ZN(n12777) );
  AOI211_X1 U15950 ( .C1(n16295), .C2(n14539), .A(n12778), .B(n12777), .ZN(
        n12782) );
  NAND3_X1 U15951 ( .A1(n12780), .A2(n12779), .A3(n19216), .ZN(n12781) );
  OAI211_X1 U15952 ( .C1(n12783), .C2(n19218), .A(n12782), .B(n12781), .ZN(
        P2_U3011) );
  NOR2_X1 U15953 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12784), .ZN(n16420) );
  INV_X1 U15954 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20790) );
  INV_X1 U15955 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16252) );
  INV_X1 U15956 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20861) );
  NAND2_X1 U15957 ( .A1(n14338), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14337) );
  INV_X1 U15958 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15054) );
  INV_X1 U15959 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14325) );
  INV_X1 U15960 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15005) );
  INV_X1 U15961 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14986) );
  INV_X1 U15962 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U15963 ( .A1(n14317), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14315) );
  INV_X1 U15964 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14928) );
  NAND2_X1 U15965 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14305) );
  AOI21_X1 U15966 ( .B1(n16306), .B2(n12788), .A(n9629), .ZN(n16294) );
  INV_X1 U15967 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U15968 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12087), .B1(n14562), 
        .B2(n16435), .ZN(n15439) );
  AOI22_X1 U15969 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12786), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16435), .ZN(n14552) );
  NOR2_X1 U15970 ( .A1(n15439), .A2(n14552), .ZN(n14551) );
  OAI21_X1 U15971 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12787), .ZN(n19223) );
  NAND2_X1 U15972 ( .A1(n14551), .A2(n19223), .ZN(n14537) );
  NOR2_X1 U15973 ( .A1(n14539), .A2(n14537), .ZN(n19119) );
  OAI21_X1 U15974 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12789), .A(
        n12788), .ZN(n19118) );
  NAND2_X1 U15975 ( .A1(n19119), .A2(n19118), .ZN(n14527) );
  NOR2_X1 U15976 ( .A1(n16294), .A2(n14527), .ZN(n14328) );
  NOR2_X1 U15977 ( .A1(n19094), .A2(n14328), .ZN(n12790) );
  OAI21_X1 U15978 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9629), .A(
        n14327), .ZN(n16293) );
  XNOR2_X1 U15979 ( .A(n12790), .B(n16293), .ZN(n12791) );
  NAND4_X1 U15980 ( .A1(n16425), .A2(n16435), .A3(n18957), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19717) );
  INV_X1 U15981 ( .A(n19717), .ZN(n19098) );
  NAND2_X1 U15982 ( .A1(n12791), .A2(n19098), .ZN(n12810) );
  AND2_X1 U15983 ( .A1(n18951), .A2(n12792), .ZN(n12805) );
  INV_X1 U15984 ( .A(n12805), .ZN(n12793) );
  NAND2_X1 U15985 ( .A1(n19714), .A2(n18957), .ZN(n12802) );
  INV_X1 U15986 ( .A(n16420), .ZN(n12794) );
  AND2_X1 U15987 ( .A1(n12795), .A2(n12794), .ZN(n14364) );
  INV_X1 U15988 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14574) );
  AND3_X1 U15989 ( .A1(n18946), .A2(n12802), .A3(n14574), .ZN(n12796) );
  INV_X1 U15990 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12801) );
  AND3_X1 U15991 ( .A1(n16425), .A2(n19713), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16417) );
  INV_X1 U15992 ( .A(n16417), .ZN(n12797) );
  NAND3_X1 U15993 ( .A1(n19717), .A2(n19089), .A3(n12797), .ZN(n12798) );
  NAND2_X1 U15994 ( .A1(n19091), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16207) );
  INV_X2 U15995 ( .A(n16207), .ZN(n19103) );
  OAI21_X1 U15996 ( .B1(n11792), .B2(n19091), .A(n19089), .ZN(n12799) );
  AOI21_X1 U15997 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19103), .A(
        n12799), .ZN(n12800) );
  OAI21_X1 U15998 ( .B1(n19109), .B2(n12801), .A(n12800), .ZN(n12808) );
  INV_X1 U15999 ( .A(n12802), .ZN(n12803) );
  NOR2_X1 U16000 ( .A1(n12803), .A2(n14574), .ZN(n12804) );
  NOR2_X1 U16001 ( .A1(n12806), .A2(n19075), .ZN(n12807) );
  AOI211_X1 U16002 ( .C1(n16290), .C2(n19115), .A(n12808), .B(n12807), .ZN(
        n12809) );
  OAI211_X1 U16003 ( .C1(n12811), .C2(n19107), .A(n12810), .B(n12809), .ZN(
        P2_U2849) );
  NAND2_X1 U16004 ( .A1(n19803), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19658) );
  NAND3_X1 U16005 ( .A1(n19827), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19545) );
  OAI21_X1 U16006 ( .B1(n19658), .B2(n19338), .A(n19545), .ZN(n12815) );
  NOR2_X1 U16007 ( .A1(n19836), .A2(n19545), .ZN(n19591) );
  INV_X1 U16008 ( .A(n19591), .ZN(n19606) );
  AND2_X1 U16009 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19606), .ZN(n12812) );
  NAND2_X1 U16010 ( .A1(n12813), .A2(n12812), .ZN(n12817) );
  NAND2_X1 U16011 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19606), .ZN(n12814) );
  INV_X1 U16012 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12821) );
  INV_X1 U16013 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16544) );
  INV_X1 U16014 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18263) );
  OAI22_X2 U16015 ( .A1(n16544), .A2(n15564), .B1(n18263), .B2(n15563), .ZN(
        n19662) );
  NOR2_X2 U16016 ( .A1(n19598), .A2(n19338), .ZN(n19593) );
  INV_X1 U16017 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18265) );
  INV_X1 U16018 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U16019 ( .A1(n19642), .A2(n19662), .B1(n19593), .B2(n19605), .ZN(
        n12820) );
  OAI21_X1 U16020 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19545), .A(n16425), 
        .ZN(n12816) );
  NOR2_X2 U16021 ( .A1(n12818), .A2(n19463), .ZN(n19653) );
  NAND2_X1 U16022 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19655), .ZN(n15493) );
  NOR2_X2 U16023 ( .A1(n16408), .A2(n15493), .ZN(n19652) );
  AOI22_X1 U16024 ( .A1(n19592), .A2(n19653), .B1(n19652), .B2(n19591), .ZN(
        n12819) );
  OAI211_X1 U16025 ( .C1(n19597), .C2(n12821), .A(n12820), .B(n12819), .ZN(
        P2_U3152) );
  INV_X1 U16026 ( .A(n19658), .ZN(n19459) );
  INV_X1 U16027 ( .A(n19800), .ZN(n12822) );
  NAND2_X1 U16028 ( .A1(n19459), .A2(n12822), .ZN(n12827) );
  NAND2_X1 U16029 ( .A1(n19817), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19498) );
  INV_X1 U16030 ( .A(n19498), .ZN(n19427) );
  NAND2_X1 U16031 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19427), .ZN(
        n12828) );
  NAND2_X1 U16032 ( .A1(n15511), .A2(n19427), .ZN(n12823) );
  INV_X1 U16033 ( .A(n12823), .ZN(n19537) );
  AND2_X1 U16034 ( .A1(n12823), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U16035 ( .A1(n12825), .A2(n12824), .ZN(n12830) );
  OAI211_X1 U16036 ( .C1(n19537), .C2(n12070), .A(n12830), .B(n19655), .ZN(
        n12826) );
  INV_X1 U16037 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16038 ( .A1(n19549), .A2(n19662), .B1(n19539), .B2(n19605), .ZN(
        n12832) );
  OAI21_X1 U16039 ( .B1(n12828), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16425), 
        .ZN(n12829) );
  AND2_X1 U16040 ( .A1(n12830), .A2(n12829), .ZN(n19538) );
  AOI22_X1 U16041 ( .A1(n19538), .A2(n19653), .B1(n19652), .B2(n19537), .ZN(
        n12831) );
  OAI211_X1 U16042 ( .C1(n19543), .C2(n12833), .A(n12832), .B(n12831), .ZN(
        P2_U3136) );
  NOR2_X1 U16043 ( .A1(n15473), .A2(n12834), .ZN(n19116) );
  INV_X1 U16044 ( .A(n19116), .ZN(n18947) );
  NOR2_X1 U16045 ( .A1(n19094), .A2(n14551), .ZN(n12835) );
  XNOR2_X1 U16046 ( .A(n12835), .B(n19223), .ZN(n12836) );
  NAND2_X1 U16047 ( .A1(n12836), .A2(n19098), .ZN(n12843) );
  NOR2_X1 U16048 ( .A1(n19075), .A2(n12837), .ZN(n12841) );
  AOI22_X1 U16049 ( .A1(n19087), .A2(P2_EBX_REG_2__SCAN_IN), .B1(n19815), .B2(
        n19070), .ZN(n12839) );
  NAND2_X1 U16050 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19103), .ZN(
        n12838) );
  OAI211_X1 U16051 ( .C1(n19091), .C2(n19743), .A(n12839), .B(n12838), .ZN(
        n12840) );
  OAI211_X1 U16052 ( .C1(n15476), .C2(n18947), .A(n12843), .B(n12842), .ZN(
        P2_U2853) );
  OR2_X1 U16053 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  AND2_X1 U16054 ( .A1(n12844), .A2(n12847), .ZN(n19888) );
  INV_X1 U16055 ( .A(n19888), .ZN(n12861) );
  INV_X1 U16056 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n12860) );
  INV_X1 U16057 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19953) );
  NAND2_X1 U16058 ( .A1(n13044), .A2(n19953), .ZN(n12852) );
  NAND2_X1 U16059 ( .A1(n13585), .A2(n19953), .ZN(n12850) );
  NAND2_X1 U16060 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12849) );
  NAND3_X1 U16061 ( .A1(n12850), .A2(n13579), .A3(n12849), .ZN(n12851) );
  AND2_X1 U16062 ( .A1(n12852), .A2(n12851), .ZN(n16148) );
  NAND2_X1 U16063 ( .A1(n16149), .A2(n16148), .ZN(n12853) );
  NAND2_X1 U16064 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12854) );
  NAND2_X1 U16065 ( .A1(n13579), .A2(n12854), .ZN(n12856) );
  NAND2_X1 U16066 ( .A1(n13585), .A2(n12860), .ZN(n12855) );
  NAND2_X1 U16067 ( .A1(n12856), .A2(n12855), .ZN(n12857) );
  OAI21_X1 U16068 ( .B1(n13596), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12857), .ZN(
        n12859) );
  INV_X1 U16069 ( .A(n12869), .ZN(n12858) );
  OAI21_X1 U16070 ( .B1(n16150), .B2(n12859), .A(n12858), .ZN(n19900) );
  OAI222_X1 U16071 ( .A1(n12861), .A2(n16020), .B1(n13839), .B2(n12860), .C1(
        n19954), .C2(n19900), .ZN(P1_U2865) );
  OAI222_X1 U16072 ( .A1(n12861), .A2(n13915), .B1(n13920), .B2(n20141), .C1(
        n19975), .C2(n13917), .ZN(P1_U2897) );
  INV_X1 U16073 ( .A(n12844), .ZN(n12863) );
  OAI21_X1 U16074 ( .B1(n12863), .B2(n10224), .A(n12862), .ZN(n13032) );
  INV_X1 U16075 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U16076 ( .A1(n13044), .A2(n12883), .ZN(n12867) );
  NAND2_X1 U16077 ( .A1(n13585), .A2(n12883), .ZN(n12865) );
  NAND2_X1 U16078 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12864) );
  NAND3_X1 U16079 ( .A1(n12865), .A2(n13579), .A3(n12864), .ZN(n12866) );
  AND2_X1 U16080 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  OR2_X1 U16081 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  AND2_X1 U16082 ( .A1(n12937), .A2(n12870), .ZN(n16139) );
  INV_X1 U16083 ( .A(n16139), .ZN(n12871) );
  OAI22_X1 U16084 ( .A1(n19954), .A2(n12871), .B1(n12883), .B2(n13839), .ZN(
        n12872) );
  INV_X1 U16085 ( .A(n12872), .ZN(n12873) );
  OAI21_X1 U16086 ( .B1(n13032), .B2(n16020), .A(n12873), .ZN(P1_U2864) );
  INV_X1 U16087 ( .A(DATAI_8_), .ZN(n12875) );
  NAND2_X1 U16088 ( .A1(n20095), .A2(BUF1_REG_8__SCAN_IN), .ZN(n12874) );
  OAI21_X1 U16089 ( .B1(n20095), .B2(n12875), .A(n12874), .ZN(n19990) );
  AOI22_X1 U16090 ( .A1(n13059), .A2(n19990), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n13906), .ZN(n12876) );
  OAI21_X1 U16091 ( .B1(n13032), .B2(n13915), .A(n12876), .ZN(P1_U2896) );
  INV_X1 U16092 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20673) );
  NAND3_X1 U16093 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19925) );
  NOR2_X1 U16094 ( .A1(n20673), .A2(n19925), .ZN(n19891) );
  INV_X1 U16095 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n12877) );
  NAND3_X1 U16096 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n12880) );
  NOR2_X1 U16097 ( .A1(n12877), .A2(n12880), .ZN(n13756) );
  NAND2_X1 U16098 ( .A1(n19891), .A2(n13756), .ZN(n13633) );
  NOR2_X1 U16099 ( .A1(n12952), .A2(n13633), .ZN(n12878) );
  NOR2_X1 U16100 ( .A1(n15982), .A2(n12878), .ZN(n12886) );
  AOI21_X1 U16101 ( .B1(n19901), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20021), .ZN(n12879) );
  OAI21_X1 U16102 ( .B1(n13028), .B2(n19948), .A(n12879), .ZN(n12885) );
  INV_X1 U16103 ( .A(n19891), .ZN(n19922) );
  NOR2_X1 U16104 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n12880), .ZN(n12881) );
  AOI22_X1 U16105 ( .A1(n19914), .A2(n16139), .B1(n19917), .B2(n12881), .ZN(
        n12882) );
  OAI21_X1 U16106 ( .B1(n12883), .B2(n16011), .A(n12882), .ZN(n12884) );
  AOI211_X1 U16107 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n12886), .A(n12885), .B(
        n12884), .ZN(n12887) );
  OAI21_X1 U16108 ( .B1(n15943), .B2(n13032), .A(n12887), .ZN(P1_U2832) );
  NAND2_X1 U16109 ( .A1(n11738), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U16110 ( .A1(n14358), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16111 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12905) );
  AOI22_X1 U16112 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U16113 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n13235), .ZN(n12891) );
  AOI22_X1 U16114 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16115 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12600), .B1(
        n12599), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12889) );
  NAND4_X1 U16116 ( .A1(n12892), .A2(n12891), .A3(n12890), .A4(n12889), .ZN(
        n12901) );
  AOI22_X1 U16117 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12899) );
  INV_X1 U16118 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n19492) );
  INV_X1 U16119 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n19333) );
  OR2_X1 U16120 ( .A1(n13211), .A2(n19333), .ZN(n12894) );
  AOI22_X1 U16121 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13229), .ZN(n12893) );
  OAI211_X1 U16122 ( .C1(n13214), .C2(n19492), .A(n12894), .B(n12893), .ZN(
        n12895) );
  INV_X1 U16123 ( .A(n12895), .ZN(n12898) );
  NAND2_X1 U16124 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U16125 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12896) );
  NAND4_X1 U16126 ( .A1(n12899), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n12900) );
  NOR2_X1 U16127 ( .A1(n12901), .A2(n12900), .ZN(n14670) );
  INV_X1 U16128 ( .A(n14670), .ZN(n12902) );
  NAND2_X1 U16129 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  NAND4_X1 U16130 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n14770) );
  XNOR2_X1 U16131 ( .A(n14770), .B(n14769), .ZN(n19037) );
  INV_X1 U16132 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19182) );
  OAI222_X1 U16133 ( .A1(n19037), .A2(n19135), .B1(n13092), .B2(n12908), .C1(
        n19144), .C2(n19182), .ZN(P2_U2904) );
  INV_X1 U16134 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12927) );
  OAI21_X1 U16135 ( .B1(n12909), .B2(n14675), .A(n12910), .ZN(n12912) );
  NAND3_X1 U16136 ( .A1(n12912), .A2(n14658), .A3(n13103), .ZN(n12926) );
  OR2_X1 U16137 ( .A1(n11329), .A2(n16244), .ZN(n12917) );
  INV_X1 U16138 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U16139 ( .A1(n14307), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U16140 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12913) );
  OAI211_X1 U16141 ( .C1(n13534), .C2(n14345), .A(n12914), .B(n12913), .ZN(
        n12915) );
  INV_X1 U16142 ( .A(n12915), .ZN(n12916) );
  NAND2_X1 U16143 ( .A1(n12917), .A2(n12916), .ZN(n14490) );
  INV_X1 U16144 ( .A(n14492), .ZN(n12922) );
  INV_X1 U16145 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15365) );
  OR2_X1 U16146 ( .A1(n11329), .A2(n15365), .ZN(n12919) );
  AOI22_X1 U16147 ( .A1(n14308), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12918) );
  OAI211_X1 U16148 ( .C1(n13540), .C2(n12920), .A(n12919), .B(n12918), .ZN(
        n12923) );
  INV_X1 U16149 ( .A(n12923), .ZN(n12921) );
  NAND2_X1 U16150 ( .A1(n12922), .A2(n12921), .ZN(n12924) );
  AND2_X1 U16151 ( .A1(n12924), .A2(n14672), .ZN(n19045) );
  NAND2_X1 U16152 ( .A1(n14652), .A2(n19045), .ZN(n12925) );
  OAI211_X1 U16153 ( .C1(n14652), .C2(n12927), .A(n12926), .B(n12925), .ZN(
        P2_U2873) );
  AOI21_X1 U16154 ( .B1(n12929), .B2(n12862), .A(n12928), .ZN(n19880) );
  INV_X1 U16155 ( .A(n19880), .ZN(n12940) );
  INV_X1 U16156 ( .A(DATAI_9_), .ZN(n12931) );
  NAND2_X1 U16157 ( .A1(n20095), .A2(BUF1_REG_9__SCAN_IN), .ZN(n12930) );
  OAI21_X1 U16158 ( .B1(n20095), .B2(n12931), .A(n12930), .ZN(n19992) );
  AOI22_X1 U16159 ( .A1(n13059), .A2(n19992), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n13906), .ZN(n12932) );
  OAI21_X1 U16160 ( .B1(n12940), .B2(n13915), .A(n12932), .ZN(P1_U2895) );
  INV_X1 U16161 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U16162 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12933) );
  NAND2_X1 U16163 ( .A1(n13579), .A2(n12933), .ZN(n12935) );
  NAND2_X1 U16164 ( .A1(n13585), .A2(n12939), .ZN(n12934) );
  AOI22_X1 U16165 ( .A1(n13584), .A2(n12939), .B1(n12935), .B2(n12934), .ZN(
        n12936) );
  NAND2_X1 U16166 ( .A1(n12937), .A2(n12936), .ZN(n12938) );
  NAND2_X1 U16167 ( .A1(n12948), .A2(n12938), .ZN(n19875) );
  OAI222_X1 U16168 ( .A1(n12940), .A2(n16020), .B1(n13839), .B2(n12939), .C1(
        n19875), .C2(n19954), .ZN(P1_U2863) );
  NOR2_X1 U16169 ( .A1(n12928), .A2(n12942), .ZN(n12943) );
  OR2_X1 U16170 ( .A1(n12941), .A2(n12943), .ZN(n14056) );
  INV_X1 U16171 ( .A(DATAI_10_), .ZN(n12945) );
  NAND2_X1 U16172 ( .A1(n20095), .A2(BUF1_REG_10__SCAN_IN), .ZN(n12944) );
  OAI21_X1 U16173 ( .B1(n20095), .B2(n12945), .A(n12944), .ZN(n19994) );
  AOI22_X1 U16174 ( .A1(n13059), .A2(n19994), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n13906), .ZN(n12946) );
  OAI21_X1 U16175 ( .B1(n14056), .B2(n13915), .A(n12946), .ZN(P1_U2894) );
  MUX2_X1 U16176 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12947) );
  NAND2_X1 U16177 ( .A1(n10231), .A2(n12947), .ZN(n12949) );
  AOI21_X1 U16178 ( .B1(n12949), .B2(n12948), .A(n13017), .ZN(n16130) );
  AOI22_X1 U16179 ( .A1(n19950), .A2(n16130), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n13828), .ZN(n12950) );
  OAI21_X1 U16180 ( .B1(n14056), .B2(n16020), .A(n12950), .ZN(P1_U2862) );
  INV_X1 U16181 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19874) );
  AOI211_X1 U16182 ( .C1(n19923), .C2(n13633), .A(n12952), .B(n19874), .ZN(
        n19884) );
  NAND2_X1 U16183 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n12951) );
  NOR3_X1 U16184 ( .A1(n12952), .A2(n13633), .A3(n12951), .ZN(n15955) );
  NOR2_X1 U16185 ( .A1(n15982), .A2(n15955), .ZN(n16015) );
  OAI21_X1 U16186 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n19884), .A(n16015), 
        .ZN(n12958) );
  INV_X1 U16187 ( .A(n12953), .ZN(n14053) );
  INV_X1 U16188 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16189 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n19934), .B1(n19914), 
        .B2(n16130), .ZN(n12954) );
  OAI211_X1 U16190 ( .C1(n19926), .C2(n12955), .A(n12954), .B(n20068), .ZN(
        n12956) );
  AOI21_X1 U16191 ( .B1(n19879), .B2(n14053), .A(n12956), .ZN(n12957) );
  OAI211_X1 U16192 ( .C1(n14056), .C2(n15943), .A(n12958), .B(n12957), .ZN(
        P1_U2830) );
  INV_X1 U16193 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16158) );
  NAND2_X1 U16194 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20038) );
  INV_X1 U16195 ( .A(n20038), .ZN(n12998) );
  NAND2_X1 U16196 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12998), .ZN(
        n14066) );
  AOI21_X1 U16197 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12996) );
  INV_X1 U16198 ( .A(n12996), .ZN(n20050) );
  NAND2_X1 U16199 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20052) );
  AOI21_X1 U16200 ( .B1(n12959), .B2(n15907), .A(n15905), .ZN(n12960) );
  AND2_X1 U16201 ( .A1(n12961), .A2(n12960), .ZN(n12968) );
  INV_X1 U16202 ( .A(n12962), .ZN(n12964) );
  NAND2_X1 U16203 ( .A1(n13844), .A2(n12978), .ZN(n12963) );
  AOI21_X1 U16204 ( .B1(n12965), .B2(n12964), .A(n12963), .ZN(n12966) );
  NOR2_X1 U16205 ( .A1(n12973), .A2(n12966), .ZN(n12967) );
  MUX2_X1 U16206 ( .A(n12968), .B(n12967), .S(n10344), .Z(n12969) );
  INV_X1 U16207 ( .A(n12969), .ZN(n12975) );
  INV_X1 U16208 ( .A(n12970), .ZN(n12972) );
  AOI21_X1 U16209 ( .B1(n12973), .B2(n12972), .A(n12971), .ZN(n12974) );
  NAND2_X1 U16210 ( .A1(n12975), .A2(n12974), .ZN(n12977) );
  MUX2_X1 U16211 ( .A(n12979), .B(n10344), .S(n12978), .Z(n12981) );
  NAND2_X1 U16212 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  NOR2_X1 U16213 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  OR2_X2 U16214 ( .A1(n13005), .A2(n12985), .ZN(n14232) );
  NAND2_X1 U16215 ( .A1(n20051), .A2(n14232), .ZN(n20076) );
  NAND2_X1 U16216 ( .A1(n20050), .A2(n16120), .ZN(n20049) );
  NOR2_X1 U16217 ( .A1(n14066), .A2(n20049), .ZN(n16154) );
  INV_X1 U16218 ( .A(n16154), .ZN(n14260) );
  NOR2_X1 U16219 ( .A1(n16158), .A2(n14260), .ZN(n16142) );
  INV_X1 U16220 ( .A(n16142), .ZN(n13009) );
  NAND2_X1 U16221 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  XNOR2_X1 U16222 ( .A(n12990), .B(n12989), .ZN(n16079) );
  OAI21_X1 U16223 ( .B1(n20124), .B2(n13001), .A(n12991), .ZN(n12992) );
  NOR2_X1 U16224 ( .A1(n10357), .A2(n12992), .ZN(n12993) );
  NAND2_X1 U16225 ( .A1(n16079), .A2(n20075), .ZN(n13008) );
  NAND2_X1 U16226 ( .A1(n14263), .A2(n20073), .ZN(n20077) );
  INV_X1 U16227 ( .A(n20077), .ZN(n14217) );
  INV_X1 U16228 ( .A(n20056), .ZN(n12999) );
  NOR2_X1 U16229 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20038), .ZN(
        n16164) );
  INV_X1 U16230 ( .A(n14085), .ZN(n14234) );
  NAND2_X1 U16231 ( .A1(n14234), .A2(n20051), .ZN(n12995) );
  NAND2_X1 U16232 ( .A1(n13005), .A2(n20068), .ZN(n12994) );
  INV_X1 U16233 ( .A(n20072), .ZN(n20057) );
  AOI21_X1 U16234 ( .B1(n20058), .B2(n20052), .A(n20057), .ZN(n20036) );
  NOR2_X1 U16235 ( .A1(n14066), .A2(n12996), .ZN(n14262) );
  OR2_X1 U16236 ( .A1(n20073), .A2(n14262), .ZN(n12997) );
  OAI211_X1 U16237 ( .C1(n14263), .C2(n12998), .A(n20036), .B(n12997), .ZN(
        n16160) );
  AOI21_X1 U16238 ( .B1(n12999), .B2(n16164), .A(n16160), .ZN(n16159) );
  OAI21_X1 U16239 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14217), .A(
        n16159), .ZN(n16140) );
  NAND2_X1 U16240 ( .A1(n13000), .A2(n10345), .ZN(n15885) );
  INV_X1 U16241 ( .A(n13001), .ZN(n13002) );
  NAND2_X1 U16242 ( .A1(n13002), .A2(n20124), .ZN(n13003) );
  AND2_X1 U16243 ( .A1(n15885), .A2(n13003), .ZN(n13004) );
  INV_X1 U16244 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19893) );
  OAI22_X1 U16245 ( .A1(n20083), .A2(n19900), .B1(n19893), .B2(n20068), .ZN(
        n13006) );
  AOI21_X1 U16246 ( .B1(n16140), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13006), .ZN(n13007) );
  OAI211_X1 U16247 ( .C1(n13009), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13008), .B(n13007), .ZN(P1_U3024) );
  OR2_X1 U16248 ( .A1(n12941), .A2(n13011), .ZN(n13012) );
  NAND2_X1 U16249 ( .A1(n13010), .A2(n13012), .ZN(n13035) );
  XNOR2_X1 U16250 ( .A(n13035), .B(n13033), .ZN(n16075) );
  INV_X1 U16251 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16073) );
  NAND2_X1 U16252 ( .A1(n13579), .A2(n16073), .ZN(n13014) );
  INV_X1 U16253 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U16254 ( .A1(n13585), .A2(n16012), .ZN(n13013) );
  NAND3_X1 U16255 ( .A1(n13014), .A2(n12501), .A3(n13013), .ZN(n13015) );
  OAI21_X1 U16256 ( .B1(n13596), .B2(P1_EBX_REG_11__SCAN_IN), .A(n13015), .ZN(
        n13016) );
  NOR2_X1 U16257 ( .A1(n13017), .A2(n13016), .ZN(n13018) );
  OR2_X1 U16258 ( .A1(n14251), .A2(n13018), .ZN(n16123) );
  OAI22_X1 U16259 ( .A1(n19954), .A2(n16123), .B1(n16012), .B2(n13839), .ZN(
        n13019) );
  AOI21_X1 U16260 ( .B1(n16075), .B2(n19956), .A(n13019), .ZN(n13020) );
  INV_X1 U16261 ( .A(n13020), .ZN(P1_U2861) );
  INV_X1 U16262 ( .A(n16075), .ZN(n13024) );
  INV_X1 U16263 ( .A(DATAI_11_), .ZN(n13022) );
  NAND2_X1 U16264 ( .A1(n20095), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13021) );
  OAI21_X1 U16265 ( .B1(n20095), .B2(n13022), .A(n13021), .ZN(n19996) );
  AOI22_X1 U16266 ( .A1(n13059), .A2(n19996), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n13906), .ZN(n13023) );
  OAI21_X1 U16267 ( .B1(n13024), .B2(n13915), .A(n13023), .ZN(P1_U2893) );
  XNOR2_X1 U16268 ( .A(n13026), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13027) );
  XNOR2_X1 U16269 ( .A(n13025), .B(n13027), .ZN(n16141) );
  NAND2_X1 U16270 ( .A1(n16141), .A2(n20029), .ZN(n13031) );
  AND2_X1 U16271 ( .A1(n20021), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n16138) );
  NOR2_X1 U16272 ( .A1(n20033), .A2(n13028), .ZN(n13029) );
  AOI211_X1 U16273 ( .C1(n20022), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16138), .B(n13029), .ZN(n13030) );
  OAI211_X1 U16274 ( .C1(n20098), .C2(n13032), .A(n13031), .B(n13030), .ZN(
        P1_U2991) );
  INV_X1 U16275 ( .A(n13033), .ZN(n13034) );
  OAI21_X1 U16276 ( .B1(n13035), .B2(n13034), .A(n13010), .ZN(n13037) );
  NAND2_X1 U16277 ( .A1(n13037), .A2(n13036), .ZN(n13755) );
  OAI21_X1 U16278 ( .B1(n13037), .B2(n13036), .A(n13755), .ZN(n16005) );
  INV_X1 U16279 ( .A(DATAI_12_), .ZN(n13039) );
  NAND2_X1 U16280 ( .A1(n20095), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16281 ( .B1(n20095), .B2(n13039), .A(n13038), .ZN(n19998) );
  AOI22_X1 U16282 ( .A1(n13059), .A2(n19998), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n13906), .ZN(n13040) );
  OAI21_X1 U16283 ( .B1(n16005), .B2(n13915), .A(n13040), .ZN(P1_U2892) );
  AOI21_X1 U16284 ( .B1(n13043), .B2(n13041), .A(n13042), .ZN(n16059) );
  INV_X1 U16285 ( .A(n16059), .ZN(n13061) );
  INV_X1 U16286 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16026) );
  NAND2_X1 U16287 ( .A1(n13044), .A2(n16026), .ZN(n13048) );
  NAND2_X1 U16288 ( .A1(n13585), .A2(n16026), .ZN(n13046) );
  NAND2_X1 U16289 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13045) );
  NAND3_X1 U16290 ( .A1(n13046), .A2(n13579), .A3(n13045), .ZN(n13047) );
  AND2_X1 U16291 ( .A1(n13048), .A2(n13047), .ZN(n14250) );
  INV_X1 U16292 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13840) );
  NAND2_X1 U16293 ( .A1(n13584), .A2(n13840), .ZN(n13052) );
  NAND2_X1 U16294 ( .A1(n13579), .A2(n14077), .ZN(n13050) );
  NAND2_X1 U16295 ( .A1(n13585), .A2(n13840), .ZN(n13049) );
  NAND3_X1 U16296 ( .A1(n13050), .A2(n12501), .A3(n13049), .ZN(n13051) );
  AND2_X1 U16297 ( .A1(n13052), .A2(n13051), .ZN(n13757) );
  MUX2_X1 U16298 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13053) );
  NAND2_X1 U16299 ( .A1(n10229), .A2(n13053), .ZN(n13054) );
  AND2_X1 U16300 ( .A1(n13759), .A2(n13054), .ZN(n13055) );
  NOR2_X1 U16301 ( .A1(n9706), .A2(n13055), .ZN(n16109) );
  AOI22_X1 U16302 ( .A1(n16109), .A2(n19950), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n13828), .ZN(n13056) );
  OAI21_X1 U16303 ( .B1(n13061), .B2(n16020), .A(n13056), .ZN(P1_U2858) );
  INV_X1 U16304 ( .A(DATAI_14_), .ZN(n13058) );
  NAND2_X1 U16305 ( .A1(n20095), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13057) );
  OAI21_X1 U16306 ( .B1(n20095), .B2(n13058), .A(n13057), .ZN(n20002) );
  AOI22_X1 U16307 ( .A1(n13059), .A2(n20002), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n13906), .ZN(n13060) );
  OAI21_X1 U16308 ( .B1(n13061), .B2(n13915), .A(n13060), .ZN(P1_U2890) );
  NAND3_X1 U16309 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17293) );
  NAND3_X1 U16310 ( .A1(n15676), .A2(n15691), .A3(n18722), .ZN(n15674) );
  OAI21_X1 U16311 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18748), .A(
        n13062), .ZN(n15685) );
  NOR2_X1 U16312 ( .A1(n13063), .A2(n15685), .ZN(n13065) );
  AOI211_X1 U16313 ( .C1(n13066), .C2(n13065), .A(n15684), .B(n13064), .ZN(
        n18707) );
  INV_X1 U16314 ( .A(n18707), .ZN(n16439) );
  NAND3_X1 U16315 ( .A1(n18316), .A2(n18293), .A3(n13067), .ZN(n13068) );
  OAI21_X1 U16316 ( .B1(n15674), .B2(n16439), .A(n13068), .ZN(n15912) );
  NOR2_X1 U16317 ( .A1(n18773), .A2(n18274), .ZN(n16440) );
  NAND2_X1 U16318 ( .A1(n18316), .A2(n17305), .ZN(n17307) );
  NOR2_X1 U16319 ( .A1(n17293), .A2(n17307), .ZN(n17297) );
  INV_X1 U16320 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17306) );
  INV_X1 U16321 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17301) );
  NOR2_X1 U16322 ( .A1(n17306), .A2(n17301), .ZN(n13069) );
  AOI21_X1 U16323 ( .B1(n17305), .B2(n13069), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n13070) );
  NOR2_X1 U16324 ( .A1(n17297), .A2(n13070), .ZN(n13071) );
  MUX2_X1 U16325 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B(n13071), .S(n17300), 
        .Z(P3_U2701) );
  INV_X1 U16326 ( .A(n18719), .ZN(n18734) );
  OAI21_X1 U16327 ( .B1(n18734), .B2(n18880), .A(n18716), .ZN(n15662) );
  NAND2_X1 U16328 ( .A1(n18735), .A2(n15662), .ZN(n18714) );
  NOR2_X1 U16329 ( .A1(n18884), .A2(n18714), .ZN(n13083) );
  INV_X1 U16330 ( .A(n18919), .ZN(n18926) );
  NOR2_X1 U16331 ( .A1(n18926), .A2(n16614), .ZN(n13081) );
  NAND2_X1 U16332 ( .A1(n18274), .A2(n17502), .ZN(n18768) );
  INV_X1 U16333 ( .A(n18768), .ZN(n17500) );
  NOR2_X1 U16334 ( .A1(n15677), .A2(n17500), .ZN(n13072) );
  NOR2_X1 U16335 ( .A1(n13075), .A2(n13074), .ZN(n13076) );
  OAI211_X1 U16336 ( .C1(n18293), .C2(n18744), .A(n15676), .B(n13076), .ZN(
        n15814) );
  NOR2_X1 U16337 ( .A1(n15814), .A2(n13077), .ZN(n13080) );
  OAI21_X1 U16338 ( .B1(n13080), .B2(n13079), .A(n13078), .ZN(n15689) );
  AOI211_X1 U16339 ( .C1(n13081), .C2(n17461), .A(n15914), .B(n15689), .ZN(
        n13082) );
  OAI21_X1 U16340 ( .B1(n16439), .B2(n15674), .A(n13082), .ZN(n18742) );
  NOR2_X1 U16341 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18872), .ZN(n18267) );
  INV_X1 U16342 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16618) );
  NAND3_X1 U16343 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18871)
         );
  NOR2_X1 U16344 ( .A1(n16618), .A2(n18871), .ZN(n15664) );
  AOI211_X1 U16345 ( .C1(n18923), .C2(n18742), .A(n18267), .B(n15664), .ZN(
        n18906) );
  MUX2_X1 U16346 ( .A(n13083), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18906), .Z(P3_U3284) );
  XOR2_X1 U16347 ( .A(n12489), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13090)
         );
  INV_X1 U16348 ( .A(n13084), .ZN(n13087) );
  INV_X1 U16349 ( .A(n13085), .ZN(n13099) );
  AOI21_X1 U16350 ( .B1(n13087), .B2(n13099), .A(n13086), .ZN(n16357) );
  NOR2_X1 U16351 ( .A1(n14652), .A2(n11786), .ZN(n13088) );
  AOI21_X1 U16352 ( .B1(n16357), .B2(n14652), .A(n13088), .ZN(n13089) );
  OAI21_X1 U16353 ( .B1(n13090), .B2(n14677), .A(n13089), .ZN(P2_U2882) );
  XOR2_X1 U16354 ( .A(n13102), .B(n13091), .Z(n13096) );
  INV_X1 U16355 ( .A(n19106), .ZN(n13094) );
  INV_X1 U16356 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19202) );
  OAI22_X1 U16357 ( .A1(n13092), .A2(n15542), .B1(n19202), .B2(n19144), .ZN(
        n13093) );
  AOI21_X1 U16358 ( .B1(n13094), .B2(n19129), .A(n13093), .ZN(n13095) );
  OAI21_X1 U16359 ( .B1(n13096), .B2(n14779), .A(n13095), .ZN(P2_U2915) );
  NAND2_X1 U16360 ( .A1(n13098), .A2(n13097), .ZN(n13100) );
  NAND2_X1 U16361 ( .A1(n13100), .A2(n13099), .ZN(n19113) );
  MUX2_X1 U16362 ( .A(n19108), .B(n19113), .S(n14652), .Z(n13101) );
  OAI21_X1 U16363 ( .B1(n13102), .B2(n14677), .A(n13101), .ZN(P2_U2883) );
  AOI22_X1 U16364 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16365 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n13235), .ZN(n13106) );
  AOI22_X1 U16366 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16367 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12600), .B1(
        n12599), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13104) );
  NAND4_X1 U16368 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13116) );
  INV_X1 U16369 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U16370 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13109) );
  AOI22_X1 U16371 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n13229), .ZN(n13108) );
  OAI211_X1 U16372 ( .C1(n13214), .C2(n13250), .A(n13109), .B(n13108), .ZN(
        n13110) );
  INV_X1 U16373 ( .A(n13110), .ZN(n13114) );
  AOI22_X1 U16374 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U16375 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13112) );
  NAND2_X1 U16376 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13111) );
  NAND4_X1 U16377 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n13115) );
  NAND2_X1 U16378 ( .A1(n14662), .A2(n14663), .ZN(n14654) );
  INV_X1 U16379 ( .A(n14654), .ZN(n13133) );
  AOI22_X1 U16380 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16381 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16382 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16383 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13117) );
  NAND4_X1 U16384 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13117), .ZN(
        n13131) );
  AOI22_X1 U16385 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13129) );
  OR2_X1 U16386 ( .A1(n13211), .A2(n13121), .ZN(n13124) );
  AOI22_X1 U16387 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13122), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13123) );
  OAI211_X1 U16388 ( .C1(n13214), .C2(n11360), .A(n13124), .B(n13123), .ZN(
        n13125) );
  INV_X1 U16389 ( .A(n13125), .ZN(n13128) );
  NAND2_X1 U16390 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13127) );
  NAND2_X1 U16391 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13126) );
  NAND4_X1 U16392 ( .A1(n13129), .A2(n13128), .A3(n13127), .A4(n13126), .ZN(
        n13130) );
  NOR2_X1 U16393 ( .A1(n13131), .A2(n13130), .ZN(n14657) );
  AOI22_X1 U16394 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16395 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16396 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16397 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U16398 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13148) );
  AOI22_X1 U16399 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13146) );
  INV_X1 U16400 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13141) );
  INV_X1 U16401 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13138) );
  OR2_X1 U16402 ( .A1(n13211), .A2(n13138), .ZN(n13140) );
  AOI22_X1 U16403 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13139) );
  OAI211_X1 U16404 ( .C1(n13214), .C2(n13141), .A(n13140), .B(n13139), .ZN(
        n13142) );
  INV_X1 U16405 ( .A(n13142), .ZN(n13145) );
  NAND2_X1 U16406 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13144) );
  NAND2_X1 U16407 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13143) );
  NAND4_X1 U16408 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n13147) );
  NOR2_X1 U16409 ( .A1(n13148), .A2(n13147), .ZN(n14645) );
  AOI22_X1 U16410 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13157) );
  OR2_X1 U16411 ( .A1(n13211), .A2(n13149), .ZN(n13151) );
  AOI22_X1 U16412 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13150) );
  OAI211_X1 U16413 ( .C1(n13214), .C2(n13152), .A(n13151), .B(n13150), .ZN(
        n13153) );
  INV_X1 U16414 ( .A(n13153), .ZN(n13156) );
  NAND2_X1 U16415 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13155) );
  NAND2_X1 U16416 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13154) );
  AND4_X1 U16417 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13168) );
  OAI22_X1 U16418 ( .A1(n13160), .A2(n20842), .B1(n13159), .B2(n13158), .ZN(
        n13164) );
  OAI22_X1 U16419 ( .A1(n13162), .A2(n13320), .B1(n13161), .B2(n13329), .ZN(
        n13163) );
  NOR2_X1 U16420 ( .A1(n13164), .A2(n13163), .ZN(n13167) );
  AOI22_X1 U16421 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13166) );
  AOI22_X1 U16422 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13165) );
  NAND4_X1 U16423 ( .A1(n13168), .A2(n13167), .A3(n13166), .A4(n13165), .ZN(
        n14637) );
  AOI22_X1 U16424 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13177) );
  INV_X1 U16425 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13172) );
  INV_X1 U16426 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13169) );
  OR2_X1 U16427 ( .A1(n13211), .A2(n13169), .ZN(n13171) );
  AOI22_X1 U16428 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13170) );
  OAI211_X1 U16429 ( .C1(n13214), .C2(n13172), .A(n13171), .B(n13170), .ZN(
        n13173) );
  INV_X1 U16430 ( .A(n13173), .ZN(n13176) );
  NAND2_X1 U16431 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13175) );
  NAND2_X1 U16432 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13174) );
  AND4_X1 U16433 ( .A1(n13177), .A2(n13176), .A3(n13175), .A4(n13174), .ZN(
        n13188) );
  AOI22_X1 U16434 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U16435 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13186) );
  INV_X1 U16436 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13352) );
  INV_X1 U16437 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13178) );
  OAI22_X1 U16438 ( .A1(n13180), .A2(n13352), .B1(n13179), .B2(n13178), .ZN(
        n13184) );
  INV_X1 U16439 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13354) );
  INV_X1 U16440 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13345) );
  OAI22_X1 U16441 ( .A1(n13182), .A2(n13354), .B1(n13181), .B2(n13345), .ZN(
        n13183) );
  NOR2_X1 U16442 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  NAND4_X1 U16443 ( .A1(n13188), .A2(n13187), .A3(n13186), .A4(n13185), .ZN(
        n14632) );
  AOI22_X1 U16444 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16445 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16446 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16447 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12600), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13189) );
  NAND4_X1 U16448 ( .A1(n13192), .A2(n13191), .A3(n13190), .A4(n13189), .ZN(
        n13203) );
  AOI22_X1 U16449 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13201) );
  OR2_X1 U16450 ( .A1(n13211), .A2(n13193), .ZN(n13195) );
  AOI22_X1 U16451 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13229), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13194) );
  OAI211_X1 U16452 ( .C1(n13214), .C2(n13196), .A(n13195), .B(n13194), .ZN(
        n13197) );
  INV_X1 U16453 ( .A(n13197), .ZN(n13200) );
  NAND2_X1 U16454 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13199) );
  NAND2_X1 U16455 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13198) );
  NAND4_X1 U16456 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        n13202) );
  NOR2_X1 U16457 ( .A1(n13203), .A2(n13202), .ZN(n14628) );
  INV_X1 U16458 ( .A(n14628), .ZN(n13204) );
  AOI22_X1 U16459 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13223), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16460 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n13235), .ZN(n13207) );
  AOI22_X1 U16461 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U16462 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12600), .B1(
        n12599), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13205) );
  NAND4_X1 U16463 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        n13221) );
  AOI22_X1 U16464 ( .A1(n13209), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13219) );
  OR2_X1 U16465 ( .A1(n13211), .A2(n13210), .ZN(n13213) );
  AOI22_X1 U16466 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n13229), .ZN(n13212) );
  OAI211_X1 U16467 ( .C1(n13214), .C2(n13395), .A(n13213), .B(n13212), .ZN(
        n13215) );
  INV_X1 U16468 ( .A(n13215), .ZN(n13218) );
  NAND2_X1 U16469 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13217) );
  NAND2_X1 U16470 ( .A1(n11415), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13216) );
  NAND4_X1 U16471 ( .A1(n13219), .A2(n13218), .A3(n13217), .A4(n13216), .ZN(
        n13220) );
  NOR2_X1 U16472 ( .A1(n13221), .A2(n13220), .ZN(n14619) );
  AOI22_X1 U16473 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12592), .B1(
        n11415), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13228) );
  AOI22_X1 U16474 ( .A1(n13223), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13222), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16475 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12594), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U16476 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12600), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13225) );
  NAND4_X1 U16477 ( .A1(n13228), .A2(n13227), .A3(n13226), .A4(n13225), .ZN(
        n13241) );
  AOI22_X1 U16478 ( .A1(n11402), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12598), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13239) );
  INV_X1 U16479 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19542) );
  NAND2_X1 U16480 ( .A1(n12599), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13232) );
  AOI22_X1 U16481 ( .A1(n13230), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n13229), .ZN(n13231) );
  OAI211_X1 U16482 ( .C1(n19542), .C2(n13233), .A(n13232), .B(n13231), .ZN(
        n13234) );
  INV_X1 U16483 ( .A(n13234), .ZN(n13238) );
  AOI22_X1 U16484 ( .A1(n13236), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13235), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13237) );
  NAND3_X1 U16485 ( .A1(n13239), .A2(n13238), .A3(n13237), .ZN(n13240) );
  NOR2_X1 U16486 ( .A1(n13241), .A2(n13240), .ZN(n13262) );
  INV_X1 U16487 ( .A(n13262), .ZN(n13261) );
  INV_X1 U16488 ( .A(n11388), .ZN(n13416) );
  INV_X1 U16489 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19315) );
  OAI22_X1 U16490 ( .A1(n13242), .A2(n15489), .B1(n13416), .B2(n19315), .ZN(
        n13245) );
  INV_X1 U16491 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15524) );
  INV_X1 U16492 ( .A(n13425), .ZN(n13398) );
  INV_X1 U16493 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13243) );
  OAI22_X1 U16494 ( .A1(n15460), .A2(n15524), .B1(n13398), .B2(n13243), .ZN(
        n13244) );
  NOR2_X1 U16495 ( .A1(n13245), .A2(n13244), .ZN(n13248) );
  AOI22_X1 U16496 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16497 ( .A1(n11383), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13246) );
  XNOR2_X1 U16498 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13418) );
  NAND4_X1 U16499 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13418), .ZN(
        n13260) );
  INV_X1 U16500 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13251) );
  OAI22_X1 U16501 ( .A1(n13242), .A2(n13251), .B1(n9597), .B2(n13250), .ZN(
        n13255) );
  INV_X1 U16502 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13253) );
  INV_X1 U16503 ( .A(n11383), .ZN(n13378) );
  INV_X1 U16504 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13252) );
  OAI22_X1 U16505 ( .A1(n13416), .A2(n13253), .B1(n13378), .B2(n13252), .ZN(
        n13254) );
  NOR2_X1 U16506 ( .A1(n13255), .A2(n13254), .ZN(n13258) );
  INV_X1 U16507 ( .A(n13418), .ZN(n13423) );
  AOI22_X1 U16508 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U16509 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13256) );
  NAND4_X1 U16510 ( .A1(n13258), .A2(n13423), .A3(n13257), .A4(n13256), .ZN(
        n13259) );
  NAND2_X1 U16511 ( .A1(n13260), .A2(n13259), .ZN(n13288) );
  INV_X1 U16512 ( .A(n13288), .ZN(n13264) );
  NAND2_X1 U16513 ( .A1(n13261), .A2(n13264), .ZN(n13267) );
  OAI21_X1 U16514 ( .B1(n16421), .B2(n13288), .A(n13262), .ZN(n13263) );
  OAI21_X1 U16515 ( .B1(n13267), .B2(n16421), .A(n13263), .ZN(n13289) );
  NAND2_X1 U16516 ( .A1(n16421), .A2(n13264), .ZN(n14615) );
  INV_X1 U16517 ( .A(n13267), .ZN(n13286) );
  OAI22_X1 U16518 ( .A1(n15460), .A2(n15530), .B1(n13398), .B2(n13268), .ZN(
        n13272) );
  OAI22_X1 U16519 ( .A1(n13416), .A2(n13270), .B1(n13378), .B2(n13269), .ZN(
        n13271) );
  NOR2_X1 U16520 ( .A1(n13272), .A2(n13271), .ZN(n13275) );
  AOI22_X1 U16521 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16522 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13273) );
  NAND4_X1 U16523 ( .A1(n13275), .A2(n13274), .A3(n13273), .A4(n13418), .ZN(
        n13285) );
  OAI22_X1 U16524 ( .A1(n15460), .A2(n19526), .B1(n13398), .B2(n13276), .ZN(
        n13280) );
  OAI22_X1 U16525 ( .A1(n13416), .A2(n13278), .B1(n13378), .B2(n13277), .ZN(
        n13279) );
  NOR2_X1 U16526 ( .A1(n13280), .A2(n13279), .ZN(n13283) );
  AOI22_X1 U16527 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16528 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13281) );
  NAND4_X1 U16529 ( .A1(n13283), .A2(n13423), .A3(n13282), .A4(n13281), .ZN(
        n13284) );
  AND2_X1 U16530 ( .A1(n13285), .A2(n13284), .ZN(n13287) );
  NAND2_X1 U16531 ( .A1(n13286), .A2(n13287), .ZN(n13290) );
  OAI211_X1 U16532 ( .C1(n13286), .C2(n13287), .A(n13309), .B(n13290), .ZN(
        n14608) );
  NAND2_X1 U16533 ( .A1(n16421), .A2(n13287), .ZN(n14610) );
  INV_X1 U16534 ( .A(n13290), .ZN(n13310) );
  INV_X1 U16535 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15535) );
  INV_X1 U16536 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13291) );
  OAI22_X1 U16537 ( .A1(n15460), .A2(n15535), .B1(n13398), .B2(n13291), .ZN(
        n13295) );
  INV_X1 U16538 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13293) );
  INV_X1 U16539 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13292) );
  OAI22_X1 U16540 ( .A1(n13416), .A2(n13293), .B1(n13378), .B2(n13292), .ZN(
        n13294) );
  NOR2_X1 U16541 ( .A1(n13295), .A2(n13294), .ZN(n13298) );
  AOI22_X1 U16542 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16543 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13296) );
  NAND4_X1 U16544 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13418), .ZN(
        n13308) );
  INV_X1 U16545 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20775) );
  OAI22_X1 U16546 ( .A1(n13299), .A2(n13398), .B1(n15460), .B2(n20775), .ZN(
        n13303) );
  INV_X1 U16547 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13301) );
  INV_X1 U16548 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13300) );
  OAI22_X1 U16549 ( .A1(n13416), .A2(n13301), .B1(n13378), .B2(n13300), .ZN(
        n13302) );
  NOR2_X1 U16550 ( .A1(n13303), .A2(n13302), .ZN(n13306) );
  AOI22_X1 U16551 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16552 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13304) );
  NAND4_X1 U16553 ( .A1(n13306), .A2(n13423), .A3(n13305), .A4(n13304), .ZN(
        n13307) );
  AND2_X1 U16554 ( .A1(n13308), .A2(n13307), .ZN(n13312) );
  NAND2_X1 U16555 ( .A1(n13310), .A2(n13312), .ZN(n13338) );
  OAI211_X1 U16556 ( .C1(n13310), .C2(n13312), .A(n13309), .B(n13338), .ZN(
        n13315) );
  INV_X1 U16557 ( .A(n13315), .ZN(n13311) );
  INV_X1 U16558 ( .A(n13312), .ZN(n13313) );
  NOR2_X1 U16559 ( .A1(n15526), .A2(n13313), .ZN(n14603) );
  OR2_X2 U16560 ( .A1(n13316), .A2(n13315), .ZN(n13317) );
  OAI22_X1 U16561 ( .A1(n15460), .A2(n15541), .B1(n13398), .B2(n13318), .ZN(
        n13322) );
  OAI22_X1 U16562 ( .A1(n13416), .A2(n13320), .B1(n13378), .B2(n13319), .ZN(
        n13321) );
  NOR2_X1 U16563 ( .A1(n13322), .A2(n13321), .ZN(n13325) );
  AOI22_X1 U16564 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16565 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13323) );
  NAND4_X1 U16566 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13418), .ZN(
        n13337) );
  OAI22_X1 U16567 ( .A1(n15460), .A2(n13327), .B1(n13398), .B2(n13326), .ZN(
        n13331) );
  OAI22_X1 U16568 ( .A1(n13416), .A2(n13329), .B1(n13378), .B2(n13328), .ZN(
        n13330) );
  NOR2_X1 U16569 ( .A1(n13331), .A2(n13330), .ZN(n13335) );
  AOI22_X1 U16570 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13334) );
  AOI22_X1 U16571 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13333) );
  NAND4_X1 U16572 ( .A1(n13335), .A2(n13423), .A3(n13334), .A4(n13333), .ZN(
        n13336) );
  NAND2_X1 U16573 ( .A1(n13337), .A2(n13336), .ZN(n13340) );
  AOI21_X1 U16574 ( .B1(n13338), .B2(n13340), .A(n13363), .ZN(n13339) );
  OR2_X1 U16575 ( .A1(n13338), .A2(n13340), .ZN(n13364) );
  NAND2_X1 U16576 ( .A1(n13339), .A2(n13364), .ZN(n13342) );
  NOR2_X1 U16577 ( .A1(n15526), .A2(n13340), .ZN(n14598) );
  INV_X1 U16578 ( .A(n13341), .ZN(n13343) );
  INV_X1 U16579 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15547) );
  INV_X1 U16580 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13344) );
  OAI22_X1 U16581 ( .A1(n15460), .A2(n15547), .B1(n13398), .B2(n13344), .ZN(
        n13348) );
  INV_X1 U16582 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13346) );
  OAI22_X1 U16583 ( .A1(n13416), .A2(n13346), .B1(n13378), .B2(n13345), .ZN(
        n13347) );
  NOR2_X1 U16584 ( .A1(n13348), .A2(n13347), .ZN(n13351) );
  AOI22_X1 U16585 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16586 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13349) );
  NAND4_X1 U16587 ( .A1(n13351), .A2(n13350), .A3(n13349), .A4(n13418), .ZN(
        n13362) );
  INV_X1 U16588 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13353) );
  OAI22_X1 U16589 ( .A1(n15460), .A2(n13353), .B1(n13398), .B2(n13352), .ZN(
        n13357) );
  INV_X1 U16590 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13355) );
  OAI22_X1 U16591 ( .A1(n13416), .A2(n13355), .B1(n13378), .B2(n13354), .ZN(
        n13356) );
  NOR2_X1 U16592 ( .A1(n13357), .A2(n13356), .ZN(n13360) );
  AOI22_X1 U16593 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U16594 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13358) );
  NAND4_X1 U16595 ( .A1(n13360), .A2(n13423), .A3(n13359), .A4(n13358), .ZN(
        n13361) );
  NAND2_X1 U16596 ( .A1(n13362), .A2(n13361), .ZN(n13366) );
  NOR2_X1 U16597 ( .A1(n13364), .A2(n13366), .ZN(n13407) );
  NOR2_X1 U16598 ( .A1(n15526), .A2(n13366), .ZN(n14594) );
  NAND2_X1 U16599 ( .A1(n14592), .A2(n14594), .ZN(n14593) );
  OAI22_X1 U16600 ( .A1(n15460), .A2(n15552), .B1(n13398), .B2(n13367), .ZN(
        n13371) );
  OAI22_X1 U16601 ( .A1(n13416), .A2(n13369), .B1(n13378), .B2(n13368), .ZN(
        n13370) );
  NOR2_X1 U16602 ( .A1(n13371), .A2(n13370), .ZN(n13374) );
  AOI22_X1 U16603 ( .A1(n9599), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16604 ( .A1(n9600), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13372) );
  NAND4_X1 U16605 ( .A1(n13374), .A2(n13373), .A3(n13372), .A4(n13418), .ZN(
        n13388) );
  OAI22_X1 U16606 ( .A1(n15460), .A2(n13376), .B1(n13398), .B2(n13375), .ZN(
        n13381) );
  OAI22_X1 U16607 ( .A1(n13416), .A2(n13379), .B1(n13378), .B2(n13377), .ZN(
        n13380) );
  NOR2_X1 U16608 ( .A1(n13381), .A2(n13380), .ZN(n13386) );
  AOI22_X1 U16609 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U16610 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13384) );
  NAND4_X1 U16611 ( .A1(n13386), .A2(n13423), .A3(n13385), .A4(n13384), .ZN(
        n13387) );
  NAND2_X1 U16612 ( .A1(n13388), .A2(n13387), .ZN(n14588) );
  AOI21_X1 U16613 ( .B1(n14593), .B2(n14587), .A(n14588), .ZN(n14578) );
  OAI22_X1 U16614 ( .A1(n13242), .A2(n15497), .B1(n11522), .B2(n9597), .ZN(
        n13391) );
  OAI22_X1 U16615 ( .A1(n15460), .A2(n15557), .B1(n13398), .B2(n13389), .ZN(
        n13390) );
  NOR2_X1 U16616 ( .A1(n13391), .A2(n13390), .ZN(n13394) );
  AOI22_X1 U16617 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U16618 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13392) );
  NAND4_X1 U16619 ( .A1(n13394), .A2(n13393), .A3(n13392), .A4(n13418), .ZN(
        n13406) );
  OAI22_X1 U16620 ( .A1(n13242), .A2(n13396), .B1(n9597), .B2(n13395), .ZN(
        n13401) );
  OAI22_X1 U16621 ( .A1(n15460), .A2(n13399), .B1(n13398), .B2(n13397), .ZN(
        n13400) );
  NOR2_X1 U16622 ( .A1(n13401), .A2(n13400), .ZN(n13404) );
  AOI22_X1 U16623 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11383), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16624 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13402) );
  NAND4_X1 U16625 ( .A1(n13404), .A2(n13423), .A3(n13403), .A4(n13402), .ZN(
        n13405) );
  NAND2_X1 U16626 ( .A1(n13406), .A2(n13405), .ZN(n13411) );
  INV_X1 U16627 ( .A(n13407), .ZN(n14586) );
  INV_X1 U16628 ( .A(n14588), .ZN(n13408) );
  NAND2_X1 U16629 ( .A1(n15526), .A2(n13408), .ZN(n13409) );
  OR2_X1 U16630 ( .A1(n14586), .A2(n13409), .ZN(n13410) );
  NOR2_X1 U16631 ( .A1(n13410), .A2(n13411), .ZN(n13412) );
  AOI21_X1 U16632 ( .B1(n13411), .B2(n13410), .A(n13412), .ZN(n14577) );
  NAND2_X1 U16633 ( .A1(n14578), .A2(n14577), .ZN(n14579) );
  INV_X1 U16634 ( .A(n13412), .ZN(n13413) );
  NAND2_X1 U16635 ( .A1(n14579), .A2(n13413), .ZN(n13436) );
  AOI22_X1 U16636 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U16637 ( .A1(n13421), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13414) );
  OAI211_X1 U16638 ( .C1(n19333), .C2(n13416), .A(n13415), .B(n13414), .ZN(
        n13433) );
  AOI22_X1 U16639 ( .A1(n9608), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13420) );
  AOI22_X1 U16640 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13419) );
  NAND3_X1 U16641 ( .A1(n13420), .A2(n13419), .A3(n13418), .ZN(n13432) );
  AOI22_X1 U16642 ( .A1(n11260), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13382), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U16643 ( .A1(n11388), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13383), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13422) );
  NAND3_X1 U16644 ( .A1(n13424), .A2(n13423), .A3(n13422), .ZN(n13431) );
  AOI22_X1 U16645 ( .A1(n13426), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13425), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U16646 ( .A1(n11383), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13427) );
  OAI211_X1 U16647 ( .C1(n13429), .C2(n19492), .A(n13428), .B(n13427), .ZN(
        n13430) );
  OAI22_X1 U16648 ( .A1(n13433), .A2(n13432), .B1(n13431), .B2(n13430), .ZN(
        n13434) );
  INV_X1 U16649 ( .A(n13434), .ZN(n13435) );
  XNOR2_X1 U16650 ( .A(n13436), .B(n13435), .ZN(n13543) );
  AND2_X1 U16651 ( .A1(n14828), .A2(n9603), .ZN(n13437) );
  INV_X1 U16652 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19768) );
  NAND2_X1 U16653 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13439) );
  NAND2_X1 U16654 ( .A1(n11719), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n13438) );
  OAI211_X1 U16655 ( .C1(n14361), .C2(n19768), .A(n13439), .B(n13438), .ZN(
        n14481) );
  INV_X1 U16656 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19761) );
  NAND2_X1 U16657 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13441) );
  NAND2_X1 U16658 ( .A1(n14358), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U16659 ( .C1(n14361), .C2(n19761), .A(n13441), .B(n13440), .ZN(
        n14768) );
  INV_X1 U16660 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n13444) );
  NAND2_X1 U16661 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13443) );
  NAND2_X1 U16662 ( .A1(n14358), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U16663 ( .C1(n14361), .C2(n13444), .A(n13443), .B(n13442), .ZN(
        n14758) );
  INV_X1 U16664 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19764) );
  NAND2_X1 U16665 ( .A1(n14358), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U16666 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13445) );
  OAI211_X1 U16667 ( .C1(n14361), .C2(n19764), .A(n13446), .B(n13445), .ZN(
        n14749) );
  AOI22_X1 U16668 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n14358), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U16669 ( .A1(n11738), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13447) );
  NOR2_X2 U16670 ( .A1(n14750), .A2(n14741), .ZN(n14480) );
  NAND2_X1 U16671 ( .A1(n14481), .A2(n14480), .ZN(n14465) );
  INV_X2 U16672 ( .A(n14465), .ZN(n13452) );
  INV_X1 U16673 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19770) );
  NAND2_X1 U16674 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13450) );
  NAND2_X1 U16675 ( .A1(n14358), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n13449) );
  OAI211_X1 U16676 ( .C1(n14361), .C2(n19770), .A(n13450), .B(n13449), .ZN(
        n13451) );
  INV_X1 U16677 ( .A(n13451), .ZN(n14466) );
  INV_X1 U16678 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19772) );
  NAND2_X1 U16679 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13454) );
  NAND2_X1 U16680 ( .A1(n11719), .A2(P2_EAX_REG_22__SCAN_IN), .ZN(n13453) );
  OAI211_X1 U16681 ( .C1(n14361), .C2(n19772), .A(n13454), .B(n13453), .ZN(
        n13455) );
  INV_X1 U16682 ( .A(n13455), .ZN(n14718) );
  INV_X1 U16683 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19773) );
  NAND2_X1 U16684 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13457) );
  NAND2_X1 U16685 ( .A1(n11719), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n13456) );
  OAI211_X1 U16686 ( .C1(n14361), .C2(n19773), .A(n13457), .B(n13456), .ZN(
        n14445) );
  INV_X1 U16687 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19775) );
  NAND2_X1 U16688 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13459) );
  NAND2_X1 U16689 ( .A1(n11719), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n13458) );
  OAI211_X1 U16690 ( .C1(n14361), .C2(n19775), .A(n13459), .B(n13458), .ZN(
        n14429) );
  INV_X1 U16691 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19777) );
  NAND2_X1 U16692 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13461) );
  NAND2_X1 U16693 ( .A1(n11719), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n13460) );
  OAI211_X1 U16694 ( .C1(n14361), .C2(n19777), .A(n13461), .B(n13460), .ZN(
        n13462) );
  INV_X1 U16695 ( .A(n13462), .ZN(n14406) );
  INV_X1 U16696 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19779) );
  NAND2_X1 U16697 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13464) );
  NAND2_X1 U16698 ( .A1(n11719), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n13463) );
  OAI211_X1 U16699 ( .C1(n14361), .C2(n19779), .A(n13464), .B(n13463), .ZN(
        n14398) );
  INV_X1 U16700 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U16701 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13467) );
  NAND2_X1 U16702 ( .A1(n11719), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n13466) );
  OAI211_X1 U16703 ( .C1(n14361), .C2(n14961), .A(n13467), .B(n13466), .ZN(
        n14374) );
  NAND2_X1 U16704 ( .A1(n14397), .A2(n14374), .ZN(n14687) );
  INV_X1 U16705 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19782) );
  NAND2_X1 U16706 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13469) );
  NAND2_X1 U16707 ( .A1(n14358), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n13468) );
  OAI211_X1 U16708 ( .C1(n14361), .C2(n19782), .A(n13469), .B(n13468), .ZN(
        n14689) );
  INV_X1 U16709 ( .A(n14689), .ZN(n13470) );
  OR2_X2 U16710 ( .A1(n14687), .A2(n13470), .ZN(n14688) );
  NAND2_X1 U16711 ( .A1(n11738), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U16712 ( .A1(n14358), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16713 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13472) );
  AND3_X1 U16714 ( .A1(n13474), .A2(n13473), .A3(n13472), .ZN(n14680) );
  OR2_X2 U16715 ( .A1(n14688), .A2(n14680), .ZN(n14682) );
  INV_X1 U16716 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16717 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13476) );
  NAND2_X1 U16718 ( .A1(n14358), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n13475) );
  OAI211_X1 U16719 ( .C1(n14361), .C2(n13539), .A(n13476), .B(n13475), .ZN(
        n13477) );
  INV_X1 U16720 ( .A(n13477), .ZN(n14357) );
  XNOR2_X1 U16721 ( .A(n14682), .B(n14357), .ZN(n16187) );
  INV_X1 U16722 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19151) );
  OAI22_X1 U16723 ( .A1(n14776), .A2(n16187), .B1(n19144), .B2(n19151), .ZN(
        n13478) );
  AOI21_X1 U16724 ( .B1(n16230), .B2(n13479), .A(n13478), .ZN(n13485) );
  OR2_X1 U16725 ( .A1(n19131), .A2(n13480), .ZN(n13483) );
  NOR2_X2 U16726 ( .A1(n13483), .A2(n13481), .ZN(n19132) );
  NOR2_X2 U16727 ( .A1(n13483), .A2(n13482), .ZN(n19130) );
  AOI22_X1 U16728 ( .A1(n19132), .A2(BUF1_REG_30__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13484) );
  OAI211_X1 U16729 ( .C1(n13543), .C2(n14779), .A(n13485), .B(n13484), .ZN(
        P2_U2889) );
  INV_X1 U16730 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U16731 ( .A1(n14307), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U16732 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13486) );
  OAI211_X1 U16733 ( .C1(n13534), .C2(n14832), .A(n13487), .B(n13486), .ZN(
        n13488) );
  AOI21_X1 U16734 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n13488), .ZN(n14671) );
  INV_X1 U16735 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15341) );
  OR2_X1 U16736 ( .A1(n11329), .A2(n15341), .ZN(n13490) );
  AOI22_X1 U16737 ( .A1(n14308), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n13489) );
  OAI211_X1 U16738 ( .C1(n13540), .C2(n19761), .A(n13490), .B(n13489), .ZN(
        n14665) );
  INV_X1 U16739 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U16740 ( .A1(n14307), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16741 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13491) );
  OAI211_X1 U16742 ( .C1(n13534), .C2(n13493), .A(n13492), .B(n13491), .ZN(
        n13494) );
  AOI21_X1 U16743 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13494), .ZN(n14653) );
  INV_X1 U16744 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U16745 ( .A1(n14307), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U16746 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13495) );
  OAI211_X1 U16747 ( .C1(n13534), .C2(n13497), .A(n13496), .B(n13495), .ZN(
        n13498) );
  AOI21_X1 U16748 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n13498), .ZN(n14646) );
  INV_X1 U16749 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15298) );
  OR2_X1 U16750 ( .A1(n11329), .A2(n15298), .ZN(n13502) );
  INV_X1 U16751 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n14351) );
  OAI22_X1 U16752 ( .A1(n13534), .A2(n14351), .B1(n13505), .B2(n15054), .ZN(
        n13500) );
  INV_X1 U16753 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19766) );
  NOR2_X1 U16754 ( .A1(n13540), .A2(n19766), .ZN(n13499) );
  NOR2_X1 U16755 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  INV_X1 U16756 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15281) );
  OR2_X1 U16757 ( .A1(n11329), .A2(n15281), .ZN(n13504) );
  AOI22_X1 U16758 ( .A1(n14308), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n13503) );
  OAI211_X1 U16759 ( .C1(n13540), .C2(n19768), .A(n13504), .B(n13503), .ZN(
        n14478) );
  INV_X1 U16760 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15270) );
  OR2_X1 U16761 ( .A1(n11329), .A2(n15270), .ZN(n13509) );
  INV_X1 U16762 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14454) );
  INV_X1 U16763 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13505) );
  OAI22_X1 U16764 ( .A1(n13534), .A2(n14454), .B1(n13505), .B2(n14325), .ZN(
        n13507) );
  NOR2_X1 U16765 ( .A1(n13540), .A2(n19770), .ZN(n13506) );
  NOR2_X1 U16766 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  INV_X1 U16767 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n13512) );
  NAND2_X1 U16768 ( .A1(n14307), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13511) );
  NAND2_X1 U16769 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13510) );
  OAI211_X1 U16770 ( .C1(n13534), .C2(n13512), .A(n13511), .B(n13510), .ZN(
        n13513) );
  AOI21_X1 U16771 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n13513), .ZN(n14620) );
  INV_X1 U16772 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15245) );
  OR2_X1 U16773 ( .A1(n11329), .A2(n15245), .ZN(n13515) );
  AOI22_X1 U16774 ( .A1(n14308), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n13514) );
  OAI211_X1 U16775 ( .C1(n13540), .C2(n19773), .A(n13515), .B(n13514), .ZN(
        n14442) );
  INV_X1 U16776 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15225) );
  OR2_X1 U16777 ( .A1(n11329), .A2(n15225), .ZN(n13517) );
  AOI22_X1 U16778 ( .A1(n14308), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n13516) );
  OAI211_X1 U16779 ( .C1(n13540), .C2(n19775), .A(n13517), .B(n13516), .ZN(
        n14426) );
  INV_X1 U16780 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20824) );
  OR2_X1 U16781 ( .A1(n11329), .A2(n20824), .ZN(n13521) );
  INV_X1 U16782 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14604) );
  OAI22_X1 U16783 ( .A1(n13534), .A2(n14604), .B1(n13505), .B2(n14986), .ZN(
        n13519) );
  NOR2_X1 U16784 ( .A1(n13540), .A2(n19777), .ZN(n13518) );
  NOR2_X1 U16785 ( .A1(n13519), .A2(n13518), .ZN(n13520) );
  AND2_X1 U16786 ( .A1(n13521), .A2(n13520), .ZN(n14404) );
  NAND2_X1 U16787 ( .A1(n14307), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13523) );
  NAND2_X1 U16788 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13522) );
  OAI211_X1 U16789 ( .C1(n13534), .C2(n9922), .A(n13523), .B(n13522), .ZN(
        n13524) );
  AOI21_X1 U16790 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13524), .ZN(n14386) );
  INV_X1 U16791 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16792 ( .A1(n14307), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13526) );
  NAND2_X1 U16793 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13525) );
  OAI211_X1 U16794 ( .C1(n13534), .C2(n13527), .A(n13526), .B(n13525), .ZN(
        n13528) );
  AOI21_X1 U16795 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13528), .ZN(n14370) );
  INV_X1 U16796 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14937) );
  OR2_X1 U16797 ( .A1(n11329), .A2(n14937), .ZN(n13530) );
  AOI22_X1 U16798 ( .A1(n14308), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n13529) );
  OAI211_X1 U16799 ( .C1(n13540), .C2(n19782), .A(n13530), .B(n13529), .ZN(
        n14582) );
  INV_X1 U16800 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U16801 ( .A1(n14307), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U16802 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13531) );
  OAI211_X1 U16803 ( .C1(n13534), .C2(n13533), .A(n13532), .B(n13531), .ZN(
        n13535) );
  AOI21_X1 U16804 ( .B1(n13536), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13535), .ZN(n14575) );
  INV_X1 U16805 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15125) );
  OR2_X1 U16806 ( .A1(n11329), .A2(n15125), .ZN(n13538) );
  AOI22_X1 U16807 ( .A1(n14308), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13537) );
  OAI211_X1 U16808 ( .C1(n13540), .C2(n13539), .A(n13538), .B(n13537), .ZN(
        n14303) );
  NAND2_X1 U16809 ( .A1(n16189), .A2(n14652), .ZN(n13542) );
  NAND2_X1 U16810 ( .A1(n14659), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13541) );
  OAI211_X1 U16811 ( .C1(n13543), .C2(n14677), .A(n13542), .B(n13541), .ZN(
        P2_U2857) );
  AOI22_X1 U16812 ( .A1(n13593), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13544), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13598) );
  NAND2_X1 U16813 ( .A1(n13593), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U16814 ( .A1(n13544), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13545) );
  NAND2_X1 U16815 ( .A1(n13546), .A2(n13545), .ZN(n13649) );
  NAND2_X1 U16816 ( .A1(n13579), .A2(n13547), .ZN(n13549) );
  INV_X1 U16817 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U16818 ( .A1(n13585), .A2(n13836), .ZN(n13548) );
  NAND3_X1 U16819 ( .A1(n13549), .A2(n12501), .A3(n13548), .ZN(n13550) );
  OAI21_X1 U16820 ( .B1(n13596), .B2(P1_EBX_REG_15__SCAN_IN), .A(n13550), .ZN(
        n13833) );
  MUX2_X1 U16821 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13551) );
  OAI21_X1 U16822 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n13593), .A(
        n13551), .ZN(n13552) );
  INV_X1 U16823 ( .A(n13552), .ZN(n13825) );
  INV_X1 U16824 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U16825 ( .A1(n13584), .A2(n15970), .ZN(n13557) );
  INV_X1 U16826 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U16827 ( .A1(n13579), .A2(n13553), .ZN(n13555) );
  NAND2_X1 U16828 ( .A1(n13585), .A2(n15970), .ZN(n13554) );
  NAND3_X1 U16829 ( .A1(n13555), .A2(n12501), .A3(n13554), .ZN(n13556) );
  AND2_X1 U16830 ( .A1(n13557), .A2(n13556), .ZN(n13818) );
  MUX2_X1 U16831 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13558) );
  OAI21_X1 U16832 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n13593), .A(
        n13558), .ZN(n13812) );
  INV_X1 U16833 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14191) );
  NAND2_X1 U16834 ( .A1(n13579), .A2(n14191), .ZN(n13560) );
  INV_X1 U16835 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U16836 ( .A1(n13585), .A2(n13806), .ZN(n13559) );
  NAND3_X1 U16837 ( .A1(n13560), .A2(n12501), .A3(n13559), .ZN(n13561) );
  OAI21_X1 U16838 ( .B1(n13596), .B2(P1_EBX_REG_19__SCAN_IN), .A(n13561), .ZN(
        n13804) );
  INV_X1 U16839 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n20792) );
  NAND2_X1 U16840 ( .A1(n13585), .A2(n20792), .ZN(n13563) );
  NAND2_X1 U16841 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13562) );
  NAND3_X1 U16842 ( .A1(n13563), .A2(n13579), .A3(n13562), .ZN(n13564) );
  OAI21_X1 U16843 ( .B1(n13590), .B2(P1_EBX_REG_20__SCAN_IN), .A(n13564), .ZN(
        n14187) );
  INV_X1 U16844 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U16845 ( .A1(n13584), .A2(n13797), .ZN(n13568) );
  NAND2_X1 U16846 ( .A1(n13579), .A2(n14182), .ZN(n13566) );
  NAND2_X1 U16847 ( .A1(n13585), .A2(n13797), .ZN(n13565) );
  NAND3_X1 U16848 ( .A1(n13566), .A2(n12501), .A3(n13565), .ZN(n13567) );
  AND2_X1 U16849 ( .A1(n13568), .A2(n13567), .ZN(n13794) );
  INV_X1 U16850 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n20887) );
  NAND2_X1 U16851 ( .A1(n13585), .A2(n20887), .ZN(n13570) );
  NAND2_X1 U16852 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13569) );
  NAND3_X1 U16853 ( .A1(n13570), .A2(n13579), .A3(n13569), .ZN(n13571) );
  OAI21_X1 U16854 ( .B1(n13590), .B2(P1_EBX_REG_22__SCAN_IN), .A(n13571), .ZN(
        n13748) );
  INV_X1 U16855 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U16856 ( .A1(n13584), .A2(n13788), .ZN(n13576) );
  NAND2_X1 U16857 ( .A1(n12501), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13572) );
  NAND2_X1 U16858 ( .A1(n13579), .A2(n13572), .ZN(n13574) );
  NAND2_X1 U16859 ( .A1(n13585), .A2(n13788), .ZN(n13573) );
  NAND2_X1 U16860 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  AND2_X1 U16861 ( .A1(n13576), .A2(n13575), .ZN(n13786) );
  MUX2_X1 U16862 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13577) );
  OAI21_X1 U16863 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n13593), .A(
        n13577), .ZN(n13727) );
  NOR2_X1 U16864 ( .A1(n13786), .A2(n13727), .ZN(n13578) );
  NAND2_X1 U16865 ( .A1(n13579), .A2(n14146), .ZN(n13581) );
  INV_X1 U16866 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n13783) );
  NAND2_X1 U16867 ( .A1(n13585), .A2(n13783), .ZN(n13580) );
  NAND3_X1 U16868 ( .A1(n13581), .A2(n12508), .A3(n13580), .ZN(n13582) );
  OAI21_X1 U16869 ( .B1(n13596), .B2(P1_EBX_REG_25__SCAN_IN), .A(n13582), .ZN(
        n13714) );
  MUX2_X1 U16870 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13583) );
  OAI21_X1 U16871 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n13593), .A(
        n13583), .ZN(n13696) );
  INV_X1 U16872 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13781) );
  NAND2_X1 U16873 ( .A1(n13584), .A2(n13781), .ZN(n13589) );
  NAND2_X1 U16874 ( .A1(n13579), .A2(n10619), .ZN(n13587) );
  NAND2_X1 U16875 ( .A1(n13585), .A2(n13781), .ZN(n13586) );
  NAND3_X1 U16876 ( .A1(n13587), .A2(n12501), .A3(n13586), .ZN(n13588) );
  AND2_X1 U16877 ( .A1(n13589), .A2(n13588), .ZN(n13681) );
  MUX2_X1 U16878 ( .A(n13590), .B(n12501), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13591) );
  OAI21_X1 U16879 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13593), .A(
        n13591), .ZN(n13673) );
  INV_X1 U16880 ( .A(n13673), .ZN(n13592) );
  OR2_X1 U16881 ( .A1(n13593), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13595) );
  INV_X1 U16882 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U16883 ( .A1(n13585), .A2(n13778), .ZN(n13594) );
  NAND2_X1 U16884 ( .A1(n13595), .A2(n13594), .ZN(n13644) );
  OAI22_X1 U16885 ( .A1(n13644), .A2(n13646), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13596), .ZN(n13662) );
  MUX2_X1 U16886 ( .A(n13649), .B(n13646), .S(n9643), .Z(n13597) );
  INV_X1 U16887 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13654) );
  XNOR2_X1 U16888 ( .A(n13599), .B(n13654), .ZN(n13934) );
  AOI22_X1 U16889 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10420), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13606) );
  AOI22_X1 U16890 ( .A1(n10314), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13600), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U16891 ( .A1(n13602), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U16892 ( .A1(n10407), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10994), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13603) );
  NAND4_X1 U16893 ( .A1(n13606), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        n13617) );
  AOI22_X1 U16894 ( .A1(n10993), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13607), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U16895 ( .A1(n10441), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13608), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U16896 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13609), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U16897 ( .A1(n13611), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13610), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13612) );
  NAND4_X1 U16898 ( .A1(n13615), .A2(n13614), .A3(n13613), .A4(n13612), .ZN(
        n13616) );
  NOR2_X1 U16899 ( .A1(n13617), .A2(n13616), .ZN(n13621) );
  NOR2_X1 U16900 ( .A1(n13619), .A2(n13618), .ZN(n13620) );
  XOR2_X1 U16901 ( .A(n13621), .B(n13620), .Z(n13626) );
  AOI21_X1 U16902 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n10675), .A(
        n13622), .ZN(n13624) );
  NAND2_X1 U16903 ( .A1(n10690), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13623) );
  OAI211_X1 U16904 ( .C1(n13626), .C2(n13625), .A(n13624), .B(n13623), .ZN(
        n13627) );
  OAI21_X1 U16905 ( .B1(n10823), .B2(n13934), .A(n13627), .ZN(n13653) );
  AOI22_X1 U16906 ( .A1(n10690), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13629), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U16907 ( .A1(n13927), .A2(n19904), .ZN(n13643) );
  INV_X1 U16908 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20703) );
  INV_X1 U16909 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20701) );
  INV_X1 U16910 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20691) );
  INV_X1 U16911 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14256) );
  INV_X1 U16912 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16122) );
  INV_X1 U16913 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20685) );
  INV_X1 U16914 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20686) );
  NOR4_X1 U16915 ( .A1(n14256), .A2(n16122), .A3(n20685), .A4(n20686), .ZN(
        n15991) );
  NAND3_X1 U16916 ( .A1(n15991), .A2(P1_REIP_REG_16__SCAN_IN), .A3(
        P1_REIP_REG_15__SCAN_IN), .ZN(n15975) );
  NOR2_X1 U16917 ( .A1(n20691), .A2(n15975), .ZN(n15956) );
  NAND4_X1 U16918 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n15956), .ZN(n15948) );
  INV_X1 U16919 ( .A(n15948), .ZN(n13631) );
  NAND2_X1 U16920 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n13631), .ZN(n13632) );
  NOR2_X1 U16921 ( .A1(n13633), .A2(n13632), .ZN(n15938) );
  NAND2_X1 U16922 ( .A1(n15938), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15928) );
  NAND3_X1 U16923 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n13634) );
  OR2_X1 U16924 ( .A1(n15928), .A2(n13634), .ZN(n13730) );
  NOR2_X1 U16925 ( .A1(n20701), .A2(n13730), .ZN(n13711) );
  NAND2_X1 U16926 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n13711), .ZN(n13639) );
  NOR2_X1 U16927 ( .A1(n20703), .A2(n13639), .ZN(n13635) );
  AND2_X1 U16928 ( .A1(n19889), .A2(n13635), .ZN(n13636) );
  OR2_X1 U16929 ( .A1(n15982), .A2(n13636), .ZN(n13687) );
  INV_X1 U16930 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20821) );
  INV_X1 U16931 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U16932 ( .B1(n20821), .B2(n13940), .A(n19923), .ZN(n13637) );
  NAND2_X1 U16933 ( .A1(n13687), .A2(n13637), .ZN(n13674) );
  INV_X1 U16934 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20710) );
  NOR2_X1 U16935 ( .A1(n13674), .A2(n20710), .ZN(n13666) );
  AOI21_X1 U16936 ( .B1(n13666), .B2(P1_REIP_REG_30__SCAN_IN), .A(n15982), 
        .ZN(n13655) );
  INV_X1 U16937 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n13775) );
  OAI22_X1 U16938 ( .A1(n16011), .A2(n13775), .B1(n13638), .B2(n19926), .ZN(
        n13641) );
  OR2_X1 U16939 ( .A1(n19890), .A2(n13639), .ZN(n13700) );
  NOR3_X1 U16940 ( .A1(n13700), .A2(n20821), .A3(n20703), .ZN(n13675) );
  NAND3_X1 U16941 ( .A1(n13675), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n13657) );
  INV_X1 U16942 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13932) );
  NOR3_X1 U16943 ( .A1(n13657), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13932), 
        .ZN(n13640) );
  AOI211_X1 U16944 ( .C1(n13655), .C2(P1_REIP_REG_31__SCAN_IN), .A(n13641), 
        .B(n13640), .ZN(n13642) );
  OAI211_X1 U16945 ( .C1(n14065), .C2(n19939), .A(n13643), .B(n13642), .ZN(
        P1_U2809) );
  NAND2_X1 U16946 ( .A1(n9643), .A2(n13646), .ZN(n13645) );
  NAND2_X1 U16947 ( .A1(n13645), .A2(n13644), .ZN(n13648) );
  OR2_X1 U16948 ( .A1(n13671), .A2(n13646), .ZN(n13647) );
  NAND2_X1 U16949 ( .A1(n13648), .A2(n13647), .ZN(n13651) );
  INV_X1 U16950 ( .A(n13649), .ZN(n13650) );
  NAND2_X1 U16951 ( .A1(n13936), .A2(n19904), .ZN(n13661) );
  OAI22_X1 U16952 ( .A1(n13654), .A2(n19926), .B1(n19948), .B2(n13934), .ZN(
        n13659) );
  INV_X1 U16953 ( .A(n13655), .ZN(n13656) );
  AOI21_X1 U16954 ( .B1(n13932), .B2(n13657), .A(n13656), .ZN(n13658) );
  AOI211_X1 U16955 ( .C1(n19934), .C2(P1_EBX_REG_30__SCAN_IN), .A(n13659), .B(
        n13658), .ZN(n13660) );
  OAI211_X1 U16956 ( .C1(n14104), .C2(n19939), .A(n13661), .B(n13660), .ZN(
        P1_U2810) );
  OAI21_X1 U16957 ( .B1(n13671), .B2(n13662), .A(n9643), .ZN(n13777) );
  INV_X1 U16958 ( .A(n13777), .ZN(n14113) );
  AOI21_X1 U16959 ( .B1(n13675), .B2(P1_REIP_REG_28__SCAN_IN), .A(
        P1_REIP_REG_29__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U16960 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19901), .B1(
        n19879), .B2(n13663), .ZN(n13665) );
  NAND2_X1 U16961 ( .A1(n19934), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13664) );
  OAI211_X1 U16962 ( .C1(n13667), .C2(n13666), .A(n13665), .B(n13664), .ZN(
        n13668) );
  AOI21_X1 U16963 ( .B1(n14113), .B2(n19914), .A(n13668), .ZN(n13669) );
  OAI21_X1 U16964 ( .B1(n13857), .B2(n15943), .A(n13669), .ZN(P1_U2811) );
  AOI21_X1 U16965 ( .B1(n13670), .B2(n9614), .A(n11151), .ZN(n13944) );
  INV_X1 U16966 ( .A(n13944), .ZN(n13863) );
  INV_X1 U16967 ( .A(n13682), .ZN(n13672) );
  AOI21_X1 U16968 ( .B1(n13673), .B2(n13672), .A(n13671), .ZN(n14120) );
  INV_X1 U16969 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13780) );
  OAI21_X1 U16970 ( .B1(n13675), .B2(P1_REIP_REG_28__SCAN_IN), .A(n13674), 
        .ZN(n13678) );
  INV_X1 U16971 ( .A(n13942), .ZN(n13676) );
  AOI22_X1 U16972 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19901), .B1(
        n19879), .B2(n13676), .ZN(n13677) );
  OAI211_X1 U16973 ( .C1(n16011), .C2(n13780), .A(n13678), .B(n13677), .ZN(
        n13679) );
  AOI21_X1 U16974 ( .B1(n14120), .B2(n19914), .A(n13679), .ZN(n13680) );
  OAI21_X1 U16975 ( .B1(n13863), .B2(n15943), .A(n13680), .ZN(P1_U2812) );
  AND2_X1 U16976 ( .A1(n9665), .A2(n13681), .ZN(n13683) );
  OR2_X1 U16977 ( .A1(n13683), .A2(n13682), .ZN(n14126) );
  INV_X1 U16978 ( .A(n9614), .ZN(n13685) );
  AOI21_X1 U16979 ( .B1(n13686), .B2(n13684), .A(n13685), .ZN(n13954) );
  NAND2_X1 U16980 ( .A1(n13954), .A2(n19904), .ZN(n13692) );
  INV_X1 U16981 ( .A(n13687), .ZN(n13701) );
  AOI22_X1 U16982 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19901), .B1(
        n19879), .B2(n13950), .ZN(n13688) );
  OAI21_X1 U16983 ( .B1(n16011), .B2(n13781), .A(n13688), .ZN(n13690) );
  NOR3_X1 U16984 ( .A1(n13700), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n20703), 
        .ZN(n13689) );
  AOI211_X1 U16985 ( .C1(n13701), .C2(P1_REIP_REG_27__SCAN_IN), .A(n13690), 
        .B(n13689), .ZN(n13691) );
  OAI211_X1 U16986 ( .C1(n19939), .C2(n14126), .A(n13692), .B(n13691), .ZN(
        P1_U2813) );
  INV_X1 U16987 ( .A(n13684), .ZN(n13694) );
  AOI21_X1 U16988 ( .B1(n13695), .B2(n13693), .A(n13694), .ZN(n13962) );
  NAND2_X1 U16989 ( .A1(n13716), .A2(n13696), .ZN(n13697) );
  NAND2_X1 U16990 ( .A1(n9665), .A2(n13697), .ZN(n14132) );
  OAI22_X1 U16991 ( .A1(n13698), .A2(n19926), .B1(n19948), .B2(n13960), .ZN(
        n13699) );
  AOI21_X1 U16992 ( .B1(n19934), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13699), .ZN(
        n13704) );
  INV_X1 U16993 ( .A(n13700), .ZN(n13702) );
  OAI21_X1 U16994 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n13702), .A(n13701), 
        .ZN(n13703) );
  OAI211_X1 U16995 ( .C1(n14132), .C2(n19939), .A(n13704), .B(n13703), .ZN(
        n13705) );
  AOI21_X1 U16996 ( .B1(n13962), .B2(n19904), .A(n13705), .ZN(n13706) );
  INV_X1 U16997 ( .A(n13706), .ZN(P1_U2814) );
  OAI21_X1 U16998 ( .B1(n13707), .B2(n13708), .A(n13693), .ZN(n13974) );
  INV_X1 U16999 ( .A(n13730), .ZN(n13709) );
  AOI21_X1 U17000 ( .B1(n13709), .B2(n19889), .A(n15982), .ZN(n13728) );
  NAND2_X1 U17001 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n13710) );
  OAI211_X1 U17002 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n13711), .A(n19923), 
        .B(n13710), .ZN(n13713) );
  AOI22_X1 U17003 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19901), .B1(
        n19879), .B2(n13967), .ZN(n13712) );
  OAI211_X1 U17004 ( .C1(n16011), .C2(n13783), .A(n13713), .B(n13712), .ZN(
        n13718) );
  OR2_X1 U17005 ( .A1(n13725), .A2(n13714), .ZN(n13715) );
  NAND2_X1 U17006 ( .A1(n13716), .A2(n13715), .ZN(n14140) );
  NOR2_X1 U17007 ( .A1(n14140), .A2(n19939), .ZN(n13717) );
  AOI211_X1 U17008 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n13728), .A(n13718), 
        .B(n13717), .ZN(n13719) );
  OAI21_X1 U17009 ( .B1(n13974), .B2(n15943), .A(n13719), .ZN(P1_U2815) );
  INV_X1 U17010 ( .A(n13707), .ZN(n13722) );
  OAI21_X1 U17011 ( .B1(n13723), .B2(n13721), .A(n13722), .ZN(n13983) );
  INV_X1 U17012 ( .A(n13786), .ZN(n13724) );
  NAND2_X1 U17013 ( .A1(n13787), .A2(n13724), .ZN(n13726) );
  AOI21_X1 U17014 ( .B1(n13727), .B2(n13726), .A(n13725), .ZN(n14155) );
  INV_X1 U17015 ( .A(n13728), .ZN(n15919) );
  OAI22_X1 U17016 ( .A1(n13729), .A2(n19926), .B1(n19948), .B2(n13975), .ZN(
        n13732) );
  NOR3_X1 U17017 ( .A1(n19890), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n13730), 
        .ZN(n13731) );
  AOI211_X1 U17018 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n19934), .A(n13732), .B(
        n13731), .ZN(n13733) );
  OAI21_X1 U17019 ( .B1(n15919), .B2(n20701), .A(n13733), .ZN(n13734) );
  AOI21_X1 U17020 ( .B1(n14155), .B2(n19914), .A(n13734), .ZN(n13735) );
  OAI21_X1 U17021 ( .B1(n13983), .B2(n15943), .A(n13735), .ZN(P1_U2816) );
  INV_X1 U17022 ( .A(n13737), .ZN(n13738) );
  AOI21_X1 U17023 ( .B1(n13739), .B2(n13736), .A(n13738), .ZN(n13993) );
  INV_X1 U17024 ( .A(n13993), .ZN(n13883) );
  INV_X1 U17025 ( .A(n15928), .ZN(n13740) );
  OAI21_X1 U17026 ( .B1(n19890), .B2(n13740), .A(n19889), .ZN(n15942) );
  INV_X1 U17027 ( .A(n15942), .ZN(n13741) );
  OAI21_X1 U17028 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19890), .A(n13741), 
        .ZN(n13747) );
  INV_X1 U17029 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n13742) );
  NOR3_X1 U17030 ( .A1(n19890), .A2(n13742), .A3(n15928), .ZN(n15918) );
  INV_X1 U17031 ( .A(n15918), .ZN(n13745) );
  AOI22_X1 U17032 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19901), .B1(
        n19879), .B2(n13996), .ZN(n13744) );
  NAND2_X1 U17033 ( .A1(n19934), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13743) );
  OAI211_X1 U17034 ( .C1(n13745), .C2(P1_REIP_REG_22__SCAN_IN), .A(n13744), 
        .B(n13743), .ZN(n13746) );
  AOI21_X1 U17035 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n13747), .A(n13746), 
        .ZN(n13751) );
  AND2_X1 U17036 ( .A1(n13796), .A2(n13748), .ZN(n13749) );
  NOR2_X1 U17037 ( .A1(n13787), .A2(n13749), .ZN(n14171) );
  NAND2_X1 U17038 ( .A1(n14171), .A2(n19914), .ZN(n13750) );
  OAI211_X1 U17039 ( .C1(n13883), .C2(n15943), .A(n13751), .B(n13750), .ZN(
        P1_U2818) );
  INV_X1 U17040 ( .A(n13752), .ZN(n13754) );
  INV_X1 U17041 ( .A(n13041), .ZN(n13753) );
  AOI21_X1 U17042 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(n14050) );
  INV_X1 U17043 ( .A(n14050), .ZN(n13921) );
  INV_X1 U17044 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20877) );
  NAND2_X1 U17045 ( .A1(n13756), .A2(n19917), .ZN(n19873) );
  INV_X1 U17046 ( .A(n16016), .ZN(n15974) );
  NOR3_X1 U17047 ( .A1(n14256), .A2(n16122), .A3(n15974), .ZN(n15999) );
  NAND2_X1 U17048 ( .A1(n14253), .A2(n13757), .ZN(n13758) );
  NAND2_X1 U17049 ( .A1(n13759), .A2(n13758), .ZN(n14238) );
  AND3_X1 U17050 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15955), .ZN(n15983) );
  OR2_X1 U17051 ( .A1(n15982), .A2(n15983), .ZN(n16008) );
  OAI22_X1 U17052 ( .A1(n19939), .A2(n14238), .B1(n20686), .B2(n16008), .ZN(
        n13765) );
  INV_X1 U17053 ( .A(n14048), .ZN(n13762) );
  INV_X1 U17054 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U17055 ( .B1(n19926), .B2(n13760), .A(n20068), .ZN(n13761) );
  AOI21_X1 U17056 ( .B1(n19879), .B2(n13762), .A(n13761), .ZN(n13763) );
  OAI21_X1 U17057 ( .B1(n16011), .B2(n13840), .A(n13763), .ZN(n13764) );
  AOI211_X1 U17058 ( .C1(n15999), .C2(n20686), .A(n13765), .B(n13764), .ZN(
        n13766) );
  OAI21_X1 U17059 ( .B1(n13921), .B2(n15943), .A(n13766), .ZN(P1_U2827) );
  INV_X1 U17060 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20733) );
  INV_X1 U17061 ( .A(n19936), .ZN(n13769) );
  OAI21_X1 U17062 ( .B1(n19901), .B2(n19879), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13767) );
  OAI21_X1 U17063 ( .B1(n13769), .B2(n13768), .A(n13767), .ZN(n13773) );
  OAI22_X1 U17064 ( .A1(n19939), .A2(n20082), .B1(n13771), .B2(n13770), .ZN(
        n13772) );
  AOI211_X1 U17065 ( .C1(P1_EBX_REG_0__SCAN_IN), .C2(n19934), .A(n13773), .B(
        n13772), .ZN(n13774) );
  OAI21_X1 U17066 ( .B1(n15982), .B2(n20733), .A(n13774), .ZN(P1_U2840) );
  OAI22_X1 U17067 ( .A1(n14065), .A2(n19954), .B1(n13775), .B2(n13839), .ZN(
        P1_U2841) );
  INV_X1 U17068 ( .A(n13936), .ZN(n13852) );
  INV_X1 U17069 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13776) );
  OAI222_X1 U17070 ( .A1(n16020), .A2(n13852), .B1(n19954), .B2(n14104), .C1(
        n13776), .C2(n13839), .ZN(P1_U2842) );
  OAI222_X1 U17071 ( .A1(n13778), .A2(n13839), .B1(n19954), .B2(n13777), .C1(
        n13857), .C2(n16020), .ZN(P1_U2843) );
  INV_X1 U17072 ( .A(n14120), .ZN(n13779) );
  OAI222_X1 U17073 ( .A1(n13780), .A2(n13839), .B1(n19954), .B2(n13779), .C1(
        n13863), .C2(n16020), .ZN(P1_U2844) );
  INV_X1 U17074 ( .A(n13954), .ZN(n13866) );
  OAI222_X1 U17075 ( .A1(n13781), .A2(n13839), .B1(n19954), .B2(n14126), .C1(
        n13866), .C2(n16020), .ZN(P1_U2845) );
  INV_X1 U17076 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n13782) );
  INV_X1 U17077 ( .A(n13962), .ZN(n13872) );
  OAI222_X1 U17078 ( .A1(n13782), .A2(n13839), .B1(n19954), .B2(n14132), .C1(
        n13872), .C2(n16020), .ZN(P1_U2846) );
  OAI222_X1 U17079 ( .A1(n13783), .A2(n13839), .B1(n19954), .B2(n14140), .C1(
        n13974), .C2(n16020), .ZN(P1_U2847) );
  AOI22_X1 U17080 ( .A1(n14155), .A2(n19950), .B1(n13828), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n13784) );
  OAI21_X1 U17081 ( .B1(n13983), .B2(n16020), .A(n13784), .ZN(P1_U2848) );
  AOI21_X1 U17082 ( .B1(n13785), .B2(n13737), .A(n13721), .ZN(n13988) );
  INV_X1 U17083 ( .A(n13988), .ZN(n15921) );
  XNOR2_X1 U17084 ( .A(n13787), .B(n13786), .ZN(n15923) );
  INV_X1 U17085 ( .A(n15923), .ZN(n13789) );
  OAI222_X1 U17086 ( .A1(n15921), .A2(n16020), .B1(n19954), .B2(n13789), .C1(
        n13788), .C2(n13839), .ZN(P1_U2849) );
  NAND2_X1 U17087 ( .A1(n13993), .A2(n19956), .ZN(n13791) );
  NAND2_X1 U17088 ( .A1(n14171), .A2(n19950), .ZN(n13790) );
  OAI211_X1 U17089 ( .C1(n20887), .C2(n13839), .A(n13791), .B(n13790), .ZN(
        P1_U2850) );
  OAI21_X1 U17090 ( .B1(n13792), .B2(n13793), .A(n13736), .ZN(n15933) );
  NAND2_X1 U17091 ( .A1(n14190), .A2(n13794), .ZN(n13795) );
  NAND2_X1 U17092 ( .A1(n13796), .A2(n13795), .ZN(n15937) );
  OAI22_X1 U17093 ( .A1(n15937), .A2(n19954), .B1(n13797), .B2(n13839), .ZN(
        n13798) );
  INV_X1 U17094 ( .A(n13798), .ZN(n13799) );
  OAI21_X1 U17095 ( .B1(n15933), .B2(n16020), .A(n13799), .ZN(P1_U2851) );
  AND2_X1 U17096 ( .A1(n13801), .A2(n13802), .ZN(n13803) );
  NOR2_X1 U17097 ( .A1(n13800), .A2(n13803), .ZN(n15954) );
  OR2_X1 U17098 ( .A1(n13814), .A2(n13804), .ZN(n13805) );
  NAND2_X1 U17099 ( .A1(n14188), .A2(n13805), .ZN(n15960) );
  OAI22_X1 U17100 ( .A1(n15960), .A2(n19954), .B1(n13806), .B2(n13839), .ZN(
        n13807) );
  AOI21_X1 U17101 ( .B1(n15954), .B2(n19956), .A(n13807), .ZN(n13808) );
  INV_X1 U17102 ( .A(n13808), .ZN(P1_U2853) );
  NAND2_X1 U17103 ( .A1(n13809), .A2(n13810), .ZN(n13811) );
  AND2_X1 U17104 ( .A1(n13801), .A2(n13811), .ZN(n15965) );
  INV_X1 U17105 ( .A(n15965), .ZN(n13902) );
  INV_X1 U17106 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n13815) );
  AND2_X1 U17107 ( .A1(n13820), .A2(n13812), .ZN(n13813) );
  OR2_X1 U17108 ( .A1(n13814), .A2(n13813), .ZN(n15963) );
  OAI222_X1 U17109 ( .A1(n13902), .A2(n16020), .B1(n13839), .B2(n13815), .C1(
        n15963), .C2(n19954), .ZN(P1_U2854) );
  OAI21_X1 U17110 ( .B1(n13816), .B2(n13817), .A(n13809), .ZN(n14036) );
  INV_X1 U17111 ( .A(n14036), .ZN(n15978) );
  NAND2_X1 U17112 ( .A1(n13827), .A2(n13818), .ZN(n13819) );
  NAND2_X1 U17113 ( .A1(n13820), .A2(n13819), .ZN(n15981) );
  OAI22_X1 U17114 ( .A1(n15981), .A2(n19954), .B1(n15970), .B2(n13839), .ZN(
        n13821) );
  AOI21_X1 U17115 ( .B1(n15978), .B2(n19956), .A(n13821), .ZN(n13822) );
  INV_X1 U17116 ( .A(n13822), .ZN(P1_U2855) );
  AOI21_X1 U17117 ( .B1(n13824), .B2(n13823), .A(n13816), .ZN(n16035) );
  INV_X1 U17118 ( .A(n16035), .ZN(n13913) );
  OR2_X1 U17119 ( .A1(n13835), .A2(n13825), .ZN(n13826) );
  AND2_X1 U17120 ( .A1(n13827), .A2(n13826), .ZN(n16096) );
  AOI22_X1 U17121 ( .A1(n16096), .A2(n19950), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n13828), .ZN(n13829) );
  OAI21_X1 U17122 ( .B1(n13913), .B2(n16020), .A(n13829), .ZN(P1_U2856) );
  INV_X1 U17123 ( .A(n13823), .ZN(n13830) );
  AOI21_X1 U17124 ( .B1(n13832), .B2(n13831), .A(n13830), .ZN(n16047) );
  NOR2_X1 U17125 ( .A1(n9706), .A2(n13833), .ZN(n13834) );
  OR2_X1 U17126 ( .A1(n13835), .A2(n13834), .ZN(n16101) );
  OAI22_X1 U17127 ( .A1(n16101), .A2(n19954), .B1(n13836), .B2(n13839), .ZN(
        n13837) );
  AOI21_X1 U17128 ( .B1(n16047), .B2(n19956), .A(n13837), .ZN(n13838) );
  INV_X1 U17129 ( .A(n13838), .ZN(P1_U2857) );
  OAI22_X1 U17130 ( .A1(n19954), .A2(n14238), .B1(n13840), .B2(n13839), .ZN(
        n13841) );
  AOI21_X1 U17131 ( .B1(n14050), .B2(n19956), .A(n13841), .ZN(n13842) );
  INV_X1 U17132 ( .A(n13842), .ZN(P1_U2859) );
  NOR2_X1 U17133 ( .A1(n13844), .A2(n20097), .ZN(n13843) );
  NAND2_X1 U17134 ( .A1(n13917), .A2(n13843), .ZN(n13890) );
  INV_X1 U17135 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16517) );
  NAND3_X1 U17136 ( .A1(n13927), .A2(n20136), .A3(n13917), .ZN(n13847) );
  NOR3_X1 U17137 ( .A1(n13906), .A2(n20095), .A3(n13844), .ZN(n13845) );
  AOI22_X1 U17138 ( .A1(n13908), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n13906), .ZN(n13846) );
  OAI211_X1 U17139 ( .C1(n13890), .C2(n16517), .A(n13847), .B(n13846), .ZN(
        P1_U2873) );
  AOI22_X1 U17140 ( .A1(n13907), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n13906), .ZN(n13851) );
  NOR3_X1 U17141 ( .A1(n13906), .A2(n20136), .A3(n13848), .ZN(n13849) );
  AOI22_X1 U17142 ( .A1(n13910), .A2(n20002), .B1(n13908), .B2(DATAI_30_), 
        .ZN(n13850) );
  OAI211_X1 U17143 ( .C1(n13852), .C2(n13915), .A(n13851), .B(n13850), .ZN(
        P1_U2874) );
  AOI22_X1 U17144 ( .A1(n13907), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n13906), .ZN(n13856) );
  INV_X1 U17145 ( .A(DATAI_13_), .ZN(n13854) );
  NAND2_X1 U17146 ( .A1(n20095), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13853) );
  OAI21_X1 U17147 ( .B1(n20095), .B2(n13854), .A(n13853), .ZN(n20000) );
  AOI22_X1 U17148 ( .A1(n13910), .A2(n20000), .B1(n13908), .B2(DATAI_29_), 
        .ZN(n13855) );
  OAI211_X1 U17149 ( .C1(n13857), .C2(n13915), .A(n13856), .B(n13855), .ZN(
        P1_U2875) );
  INV_X1 U17150 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n13859) );
  OAI22_X1 U17151 ( .A1(n13890), .A2(n13859), .B1(n13858), .B2(n13917), .ZN(
        n13860) );
  INV_X1 U17152 ( .A(n13860), .ZN(n13862) );
  AOI22_X1 U17153 ( .A1(n13910), .A2(n19998), .B1(n13908), .B2(DATAI_28_), 
        .ZN(n13861) );
  OAI211_X1 U17154 ( .C1(n13863), .C2(n13915), .A(n13862), .B(n13861), .ZN(
        P1_U2876) );
  AOI22_X1 U17155 ( .A1(n13907), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n13906), .ZN(n13865) );
  AOI22_X1 U17156 ( .A1(n13910), .A2(n19996), .B1(n13908), .B2(DATAI_27_), 
        .ZN(n13864) );
  OAI211_X1 U17157 ( .C1(n13866), .C2(n13915), .A(n13865), .B(n13864), .ZN(
        P1_U2877) );
  INV_X1 U17158 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n13868) );
  OAI22_X1 U17159 ( .A1(n13890), .A2(n13868), .B1(n13867), .B2(n13917), .ZN(
        n13869) );
  INV_X1 U17160 ( .A(n13869), .ZN(n13871) );
  AOI22_X1 U17161 ( .A1(n13910), .A2(n19994), .B1(n13908), .B2(DATAI_26_), 
        .ZN(n13870) );
  OAI211_X1 U17162 ( .C1(n13872), .C2(n13915), .A(n13871), .B(n13870), .ZN(
        P1_U2878) );
  AOI22_X1 U17163 ( .A1(n13907), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n13906), .ZN(n13874) );
  AOI22_X1 U17164 ( .A1(n13910), .A2(n19992), .B1(n13908), .B2(DATAI_25_), 
        .ZN(n13873) );
  OAI211_X1 U17165 ( .C1(n13974), .C2(n13915), .A(n13874), .B(n13873), .ZN(
        P1_U2879) );
  AOI22_X1 U17166 ( .A1(n13907), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n13906), .ZN(n13876) );
  AOI22_X1 U17167 ( .A1(n13910), .A2(n19990), .B1(n13908), .B2(DATAI_24_), 
        .ZN(n13875) );
  OAI211_X1 U17168 ( .C1(n13983), .C2(n13915), .A(n13876), .B(n13875), .ZN(
        P1_U2880) );
  AOI22_X1 U17169 ( .A1(n13907), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n13906), .ZN(n13879) );
  AOI22_X1 U17170 ( .A1(n13910), .A2(n13877), .B1(n13908), .B2(DATAI_23_), 
        .ZN(n13878) );
  OAI211_X1 U17171 ( .C1(n15921), .C2(n13915), .A(n13879), .B(n13878), .ZN(
        P1_U2881) );
  AOI22_X1 U17172 ( .A1(n13907), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n13906), .ZN(n13882) );
  AOI22_X1 U17173 ( .A1(n13910), .A2(n13880), .B1(n13908), .B2(DATAI_22_), 
        .ZN(n13881) );
  OAI211_X1 U17174 ( .C1(n13883), .C2(n13915), .A(n13882), .B(n13881), .ZN(
        P1_U2882) );
  AOI22_X1 U17175 ( .A1(n13907), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n13906), .ZN(n13886) );
  AOI22_X1 U17176 ( .A1(n13910), .A2(n13884), .B1(n13908), .B2(DATAI_21_), 
        .ZN(n13885) );
  OAI211_X1 U17177 ( .C1(n15933), .C2(n13915), .A(n13886), .B(n13885), .ZN(
        P1_U2883) );
  NOR2_X1 U17178 ( .A1(n13800), .A2(n13887), .ZN(n13888) );
  OR2_X1 U17179 ( .A1(n13792), .A2(n13888), .ZN(n16021) );
  INV_X1 U17180 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16536) );
  INV_X1 U17181 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13889) );
  OAI22_X1 U17182 ( .A1(n13890), .A2(n16536), .B1(n13889), .B2(n13917), .ZN(
        n13893) );
  INV_X1 U17183 ( .A(n13910), .ZN(n13891) );
  NOR2_X1 U17184 ( .A1(n13891), .A2(n20125), .ZN(n13892) );
  AOI211_X1 U17185 ( .C1(n13908), .C2(DATAI_20_), .A(n13893), .B(n13892), .ZN(
        n13894) );
  OAI21_X1 U17186 ( .B1(n16021), .B2(n13915), .A(n13894), .ZN(P1_U2884) );
  INV_X1 U17187 ( .A(n15954), .ZN(n13898) );
  AOI22_X1 U17188 ( .A1(n13907), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n13906), .ZN(n13897) );
  AOI22_X1 U17189 ( .A1(n13910), .A2(n13895), .B1(n13908), .B2(DATAI_19_), 
        .ZN(n13896) );
  OAI211_X1 U17190 ( .C1(n13898), .C2(n13915), .A(n13897), .B(n13896), .ZN(
        P1_U2885) );
  AOI22_X1 U17191 ( .A1(n13907), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n13906), .ZN(n13901) );
  AOI22_X1 U17192 ( .A1(n13910), .A2(n13899), .B1(n13908), .B2(DATAI_18_), 
        .ZN(n13900) );
  OAI211_X1 U17193 ( .C1(n13902), .C2(n13915), .A(n13901), .B(n13900), .ZN(
        P1_U2886) );
  AOI22_X1 U17194 ( .A1(n13907), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n13906), .ZN(n13905) );
  AOI22_X1 U17195 ( .A1(n13910), .A2(n13903), .B1(n13908), .B2(DATAI_17_), 
        .ZN(n13904) );
  OAI211_X1 U17196 ( .C1(n14036), .C2(n13915), .A(n13905), .B(n13904), .ZN(
        P1_U2887) );
  AOI22_X1 U17197 ( .A1(n13907), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n13906), .ZN(n13912) );
  AOI22_X1 U17198 ( .A1(n13910), .A2(n13909), .B1(n13908), .B2(DATAI_16_), 
        .ZN(n13911) );
  OAI211_X1 U17199 ( .C1(n13913), .C2(n13915), .A(n13912), .B(n13911), .ZN(
        P1_U2888) );
  INV_X1 U17200 ( .A(n16047), .ZN(n13916) );
  OAI222_X1 U17201 ( .A1(n13916), .A2(n13915), .B1(n13920), .B2(n13914), .C1(
        n13917), .C2(n12262), .ZN(P1_U2889) );
  INV_X1 U17202 ( .A(n20000), .ZN(n13919) );
  OAI222_X1 U17203 ( .A1(n13921), .A2(n13915), .B1(n13920), .B2(n13919), .C1(
        n13918), .C2(n13917), .ZN(P1_U2891) );
  INV_X1 U17204 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14115) );
  NAND2_X1 U17205 ( .A1(n20021), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U17206 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13924) );
  OAI211_X1 U17207 ( .C1(n20033), .C2(n13925), .A(n14096), .B(n13924), .ZN(
        n13926) );
  AOI21_X1 U17208 ( .B1(n13927), .B2(n20028), .A(n13926), .ZN(n13928) );
  OAI21_X1 U17209 ( .B1(n14102), .B2(n16067), .A(n13928), .ZN(P1_U2968) );
  XNOR2_X1 U17210 ( .A(n13931), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14108) );
  NOR2_X1 U17211 ( .A1(n20068), .A2(n13932), .ZN(n14105) );
  AOI21_X1 U17212 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14105), .ZN(n13933) );
  OAI21_X1 U17213 ( .B1(n20033), .B2(n13934), .A(n13933), .ZN(n13935) );
  AOI21_X1 U17214 ( .B1(n13936), .B2(n20028), .A(n13935), .ZN(n13937) );
  OAI21_X1 U17215 ( .B1(n14108), .B2(n16067), .A(n13937), .ZN(P1_U2969) );
  XOR2_X1 U17216 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n13939), .Z(
        n14123) );
  NOR2_X1 U17217 ( .A1(n20068), .A2(n13940), .ZN(n14119) );
  AOI21_X1 U17218 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14119), .ZN(n13941) );
  OAI21_X1 U17219 ( .B1(n20033), .B2(n13942), .A(n13941), .ZN(n13943) );
  AOI21_X1 U17220 ( .B1(n13944), .B2(n20028), .A(n13943), .ZN(n13945) );
  OAI21_X1 U17221 ( .B1(n16067), .B2(n14123), .A(n13945), .ZN(P1_U2971) );
  NAND2_X1 U17222 ( .A1(n13946), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13948) );
  MUX2_X1 U17223 ( .A(n13948), .B(n13947), .S(n14000), .Z(n13949) );
  XNOR2_X1 U17224 ( .A(n13949), .B(n10619), .ZN(n14131) );
  NAND2_X1 U17225 ( .A1(n16064), .A2(n13950), .ZN(n13951) );
  NAND2_X1 U17226 ( .A1(n20021), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U17227 ( .C1(n14062), .C2(n13952), .A(n13951), .B(n14125), .ZN(
        n13953) );
  AOI21_X1 U17228 ( .B1(n13954), .B2(n20028), .A(n13953), .ZN(n13955) );
  OAI21_X1 U17229 ( .B1(n16067), .B2(n14131), .A(n13955), .ZN(P1_U2972) );
  OR2_X1 U17230 ( .A1(n13956), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13957) );
  NAND2_X1 U17231 ( .A1(n13958), .A2(n13957), .ZN(n14139) );
  NOR2_X1 U17232 ( .A1(n20068), .A2(n20703), .ZN(n14134) );
  AOI21_X1 U17233 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14134), .ZN(n13959) );
  OAI21_X1 U17234 ( .B1(n20033), .B2(n13960), .A(n13959), .ZN(n13961) );
  AOI21_X1 U17235 ( .B1(n13962), .B2(n20028), .A(n13961), .ZN(n13963) );
  OAI21_X1 U17236 ( .B1(n16067), .B2(n14139), .A(n13963), .ZN(P1_U2973) );
  INV_X1 U17237 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n13964) );
  NOR2_X1 U17238 ( .A1(n20068), .A2(n13964), .ZN(n14141) );
  INV_X1 U17239 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13965) );
  NOR2_X1 U17240 ( .A1(n14062), .A2(n13965), .ZN(n13966) );
  AOI211_X1 U17241 ( .C1(n16064), .C2(n13967), .A(n14141), .B(n13966), .ZN(
        n13973) );
  AOI21_X1 U17242 ( .B1(n13968), .B2(n16055), .A(n14165), .ZN(n13977) );
  NOR2_X1 U17243 ( .A1(n13985), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13969) );
  MUX2_X1 U17244 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n13969), .S(
        n14000), .Z(n13970) );
  OAI21_X1 U17245 ( .B1(n13977), .B2(n14086), .A(n13970), .ZN(n13971) );
  XNOR2_X1 U17246 ( .A(n13971), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14149) );
  NAND2_X1 U17247 ( .A1(n14149), .A2(n20029), .ZN(n13972) );
  OAI211_X1 U17248 ( .C1(n13974), .C2(n20098), .A(n13973), .B(n13972), .ZN(
        P1_U2974) );
  NOR2_X1 U17249 ( .A1(n20068), .A2(n20701), .ZN(n14154) );
  NOR2_X1 U17250 ( .A1(n20033), .A2(n13975), .ZN(n13976) );
  AOI211_X1 U17251 ( .C1(n20022), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14154), .B(n13976), .ZN(n13982) );
  NOR2_X1 U17252 ( .A1(n13985), .A2(n16055), .ZN(n13979) );
  MUX2_X1 U17253 ( .A(n13979), .B(n13978), .S(n13977), .Z(n13980) );
  XNOR2_X1 U17254 ( .A(n13980), .B(n14086), .ZN(n14151) );
  NAND2_X1 U17255 ( .A1(n14151), .A2(n20029), .ZN(n13981) );
  OAI211_X1 U17256 ( .C1(n13983), .C2(n20098), .A(n13982), .B(n13981), .ZN(
        P1_U2975) );
  XNOR2_X1 U17257 ( .A(n16055), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13984) );
  XNOR2_X1 U17258 ( .A(n13985), .B(n13984), .ZN(n14169) );
  NAND2_X1 U17259 ( .A1(n16064), .A2(n15917), .ZN(n13986) );
  NAND2_X1 U17260 ( .A1(n20021), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14163) );
  OAI211_X1 U17261 ( .C1(n14062), .C2(n15926), .A(n13986), .B(n14163), .ZN(
        n13987) );
  AOI21_X1 U17262 ( .B1(n13988), .B2(n20028), .A(n13987), .ZN(n13989) );
  OAI21_X1 U17263 ( .B1(n14169), .B2(n16067), .A(n13989), .ZN(P1_U2976) );
  NAND2_X1 U17264 ( .A1(n13991), .A2(n13990), .ZN(n13992) );
  XOR2_X1 U17265 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n13992), .Z(
        n14177) );
  NAND2_X1 U17266 ( .A1(n13993), .A2(n20028), .ZN(n13998) );
  INV_X1 U17267 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20698) );
  NOR2_X1 U17268 ( .A1(n20068), .A2(n20698), .ZN(n14170) );
  INV_X1 U17269 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13994) );
  NOR2_X1 U17270 ( .A1(n14062), .A2(n13994), .ZN(n13995) );
  AOI211_X1 U17271 ( .C1(n16064), .C2(n13996), .A(n14170), .B(n13995), .ZN(
        n13997) );
  OAI211_X1 U17272 ( .C1(n14177), .C2(n16067), .A(n13998), .B(n13997), .ZN(
        P1_U2977) );
  INV_X1 U17273 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14210) );
  OAI21_X1 U17274 ( .B1(n16070), .B2(n14210), .A(n13999), .ZN(n14017) );
  NAND2_X1 U17275 ( .A1(n14000), .A2(n14191), .ZN(n14015) );
  NAND2_X1 U17276 ( .A1(n16070), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14014) );
  OAI22_X1 U17277 ( .A1(n14017), .A2(n14015), .B1(n13999), .B2(n14014), .ZN(
        n14009) );
  NAND2_X1 U17278 ( .A1(n14009), .A2(n14008), .ZN(n14007) );
  INV_X1 U17279 ( .A(n14014), .ZN(n14001) );
  NAND2_X1 U17280 ( .A1(n14001), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14002) );
  OAI22_X1 U17281 ( .A1(n14007), .A2(n16055), .B1(n13999), .B2(n14002), .ZN(
        n14003) );
  XNOR2_X1 U17282 ( .A(n14003), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14185) );
  NAND2_X1 U17283 ( .A1(n20021), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17284 ( .B1(n14062), .B2(n15927), .A(n14178), .ZN(n14005) );
  NOR2_X1 U17285 ( .A1(n15933), .A2(n20098), .ZN(n14004) );
  AOI211_X1 U17286 ( .C1(n16064), .C2(n15935), .A(n14005), .B(n14004), .ZN(
        n14006) );
  OAI21_X1 U17287 ( .B1(n14185), .B2(n16067), .A(n14006), .ZN(P1_U2978) );
  OAI21_X1 U17288 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14186) );
  NAND2_X1 U17289 ( .A1(n14186), .A2(n20029), .ZN(n14013) );
  INV_X1 U17290 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14010) );
  NOR2_X1 U17291 ( .A1(n20068), .A2(n14010), .ZN(n14193) );
  NOR2_X1 U17292 ( .A1(n20033), .A2(n15947), .ZN(n14011) );
  AOI211_X1 U17293 ( .C1(n20022), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14193), .B(n14011), .ZN(n14012) );
  OAI211_X1 U17294 ( .C1(n16021), .C2(n20098), .A(n14013), .B(n14012), .ZN(
        P1_U2979) );
  NAND2_X1 U17295 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  XNOR2_X1 U17296 ( .A(n14017), .B(n14016), .ZN(n14207) );
  NAND2_X1 U17297 ( .A1(n15954), .A2(n20028), .ZN(n14020) );
  INV_X1 U17298 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20693) );
  NOR2_X1 U17299 ( .A1(n20068), .A2(n20693), .ZN(n14200) );
  INV_X1 U17300 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15951) );
  NOR2_X1 U17301 ( .A1(n14062), .A2(n15951), .ZN(n14018) );
  AOI211_X1 U17302 ( .C1(n16064), .C2(n15949), .A(n14200), .B(n14018), .ZN(
        n14019) );
  OAI211_X1 U17303 ( .C1(n14207), .C2(n16067), .A(n14020), .B(n14019), .ZN(
        P1_U2980) );
  OAI21_X1 U17304 ( .B1(n14022), .B2(n14021), .A(n13999), .ZN(n14220) );
  NAND2_X1 U17305 ( .A1(n16064), .A2(n15962), .ZN(n14023) );
  NAND2_X1 U17306 ( .A1(n20021), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14208) );
  OAI211_X1 U17307 ( .C1(n14062), .C2(n14024), .A(n14023), .B(n14208), .ZN(
        n14025) );
  AOI21_X1 U17308 ( .B1(n15965), .B2(n20028), .A(n14025), .ZN(n14026) );
  OAI21_X1 U17309 ( .B1(n16067), .B2(n14220), .A(n14026), .ZN(P1_U2981) );
  NAND2_X1 U17310 ( .A1(n14027), .A2(n14028), .ZN(n16052) );
  INV_X1 U17311 ( .A(n14029), .ZN(n14031) );
  OAI21_X1 U17312 ( .B1(n16052), .B2(n14031), .A(n14030), .ZN(n14032) );
  MUX2_X1 U17313 ( .A(n14034), .B(n14033), .S(n14032), .Z(n14035) );
  XNOR2_X1 U17314 ( .A(n14035), .B(n13553), .ZN(n14226) );
  NAND2_X1 U17315 ( .A1(n20021), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14221) );
  OAI21_X1 U17316 ( .B1(n14062), .B2(n15971), .A(n14221), .ZN(n14038) );
  NOR2_X1 U17317 ( .A1(n14036), .A2(n20098), .ZN(n14037) );
  AOI211_X1 U17318 ( .C1(n16064), .C2(n15973), .A(n14038), .B(n14037), .ZN(
        n14039) );
  OAI21_X1 U17319 ( .B1(n14226), .B2(n16067), .A(n14039), .ZN(P1_U2982) );
  NAND2_X1 U17320 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14040) );
  NAND2_X1 U17321 ( .A1(n16055), .A2(n14040), .ZN(n16050) );
  INV_X1 U17322 ( .A(n16050), .ZN(n14042) );
  OAI22_X1 U17323 ( .A1(n14027), .A2(n14042), .B1(n14041), .B2(n16055), .ZN(
        n14245) );
  INV_X1 U17324 ( .A(n14044), .ZN(n14043) );
  OAI21_X1 U17325 ( .B1(n16070), .B2(n14248), .A(n14043), .ZN(n14244) );
  NOR2_X1 U17326 ( .A1(n14245), .A2(n14244), .ZN(n14243) );
  NOR2_X1 U17327 ( .A1(n14243), .A2(n14044), .ZN(n14045) );
  XOR2_X1 U17328 ( .A(n14046), .B(n14045), .Z(n14242) );
  AOI22_X1 U17329 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U17330 ( .B1(n20033), .B2(n14048), .A(n14047), .ZN(n14049) );
  AOI21_X1 U17331 ( .B1(n14050), .B2(n20028), .A(n14049), .ZN(n14051) );
  OAI21_X1 U17332 ( .B1(n14242), .B2(n16067), .A(n14051), .ZN(P1_U2986) );
  MUX2_X1 U17333 ( .A(n16069), .B(n14027), .S(n16070), .Z(n14052) );
  XNOR2_X1 U17334 ( .A(n14052), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16133) );
  NOR2_X1 U17335 ( .A1(n20068), .A2(n20877), .ZN(n16129) );
  AOI21_X1 U17336 ( .B1(n20022), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16129), .ZN(n14055) );
  NAND2_X1 U17337 ( .A1(n16064), .A2(n14053), .ZN(n14054) );
  OAI211_X1 U17338 ( .C1(n14056), .C2(n20098), .A(n14055), .B(n14054), .ZN(
        n14057) );
  AOI21_X1 U17339 ( .B1(n16133), .B2(n20029), .A(n14057), .ZN(n14058) );
  INV_X1 U17340 ( .A(n14058), .ZN(P1_U2989) );
  MUX2_X1 U17341 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n10604), .S(
        n16070), .Z(n14060) );
  XOR2_X1 U17342 ( .A(n14060), .B(n14059), .Z(n14271) );
  NAND2_X1 U17343 ( .A1(n16064), .A2(n19878), .ZN(n14061) );
  NAND2_X1 U17344 ( .A1(n20021), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14267) );
  OAI211_X1 U17345 ( .C1(n14062), .C2(n19876), .A(n14061), .B(n14267), .ZN(
        n14063) );
  AOI21_X1 U17346 ( .B1(n19880), .B2(n20028), .A(n14063), .ZN(n14064) );
  OAI21_X1 U17347 ( .B1(n14271), .B2(n16067), .A(n14064), .ZN(P1_U2990) );
  INV_X1 U17348 ( .A(n14065), .ZN(n14100) );
  NOR2_X1 U17349 ( .A1(n20052), .A2(n14066), .ZN(n14261) );
  INV_X1 U17350 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16136) );
  NAND3_X1 U17351 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14264) );
  NOR3_X1 U17352 ( .A1(n16136), .A2(n10604), .A3(n14264), .ZN(n14068) );
  NAND2_X1 U17353 ( .A1(n14261), .A2(n14068), .ZN(n14247) );
  NOR3_X1 U17354 ( .A1(n14248), .A2(n16073), .A3(n14247), .ZN(n14231) );
  INV_X1 U17355 ( .A(n14231), .ZN(n14233) );
  NOR2_X1 U17356 ( .A1(n14085), .A2(n14233), .ZN(n14067) );
  NAND2_X1 U17357 ( .A1(n14067), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14070) );
  INV_X1 U17358 ( .A(n20073), .ZN(n20055) );
  AND2_X1 U17359 ( .A1(n14068), .A2(n14262), .ZN(n16121) );
  AND2_X1 U17360 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16121), .ZN(
        n14249) );
  NAND2_X1 U17361 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14249), .ZN(
        n14076) );
  INV_X1 U17362 ( .A(n14076), .ZN(n14237) );
  NAND2_X1 U17363 ( .A1(n20055), .A2(n14237), .ZN(n14069) );
  NOR2_X1 U17364 ( .A1(n14077), .A2(n14233), .ZN(n14227) );
  INV_X1 U17365 ( .A(n14227), .ZN(n14235) );
  INV_X1 U17366 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16100) );
  NOR3_X1 U17367 ( .A1(n13547), .A2(n16100), .A3(n13553), .ZN(n14216) );
  NAND3_X1 U17368 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n14216), .ZN(n14202) );
  INV_X1 U17369 ( .A(n14202), .ZN(n14071) );
  NAND2_X1 U17370 ( .A1(n14071), .A2(n9723), .ZN(n14080) );
  NOR2_X1 U17371 ( .A1(n14209), .A2(n14080), .ZN(n14183) );
  NAND2_X1 U17372 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14082) );
  INV_X1 U17373 ( .A(n14082), .ZN(n14072) );
  AND2_X1 U17374 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U17375 ( .A1(n14143), .A2(n14093), .ZN(n14124) );
  INV_X1 U17376 ( .A(n14074), .ZN(n14094) );
  OR2_X1 U17377 ( .A1(n14124), .A2(n14094), .ZN(n14111) );
  NAND3_X1 U17378 ( .A1(n14075), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14098) );
  NOR2_X1 U17379 ( .A1(n14077), .A2(n14076), .ZN(n16115) );
  NOR2_X1 U17380 ( .A1(n20073), .A2(n16115), .ZN(n14215) );
  OAI21_X1 U17381 ( .B1(n14215), .B2(n14202), .A(n20077), .ZN(n14078) );
  INV_X1 U17382 ( .A(n14078), .ZN(n14079) );
  OAI21_X1 U17383 ( .B1(n14263), .B2(n14227), .A(n20072), .ZN(n14214) );
  OR2_X1 U17384 ( .A1(n14079), .A2(n14214), .ZN(n14205) );
  AND2_X1 U17385 ( .A1(n20077), .A2(n14080), .ZN(n14081) );
  NOR2_X1 U17386 ( .A1(n14205), .A2(n14081), .ZN(n14179) );
  NAND2_X1 U17387 ( .A1(n20077), .A2(n14082), .ZN(n14083) );
  AND2_X1 U17388 ( .A1(n14179), .A2(n14083), .ZN(n14166) );
  NAND2_X1 U17389 ( .A1(n20055), .A2(n14165), .ZN(n14084) );
  AND2_X1 U17390 ( .A1(n14166), .A2(n14084), .ZN(n14156) );
  NAND2_X1 U17391 ( .A1(n20073), .A2(n14085), .ZN(n20087) );
  NAND2_X1 U17392 ( .A1(n20087), .A2(n14086), .ZN(n14087) );
  NAND2_X1 U17393 ( .A1(n14156), .A2(n14087), .ZN(n14088) );
  NOR2_X1 U17394 ( .A1(n14088), .A2(n20077), .ZN(n14092) );
  INV_X1 U17395 ( .A(n14092), .ZN(n14095) );
  INV_X1 U17396 ( .A(n14088), .ZN(n14091) );
  NAND2_X1 U17397 ( .A1(n20058), .A2(n14089), .ZN(n14090) );
  AOI21_X1 U17398 ( .B1(n14093), .B2(n14147), .A(n14092), .ZN(n14129) );
  AOI21_X1 U17399 ( .B1(n14094), .B2(n14095), .A(n14129), .ZN(n14116) );
  OAI211_X1 U17400 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14217), .A(
        n14116), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14107) );
  NAND3_X1 U17401 ( .A1(n14107), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14095), .ZN(n14097) );
  OAI211_X1 U17402 ( .C1(n14111), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        n14099) );
  AOI21_X1 U17403 ( .B1(n20071), .B2(n14100), .A(n14099), .ZN(n14101) );
  OAI21_X1 U17404 ( .B1(n14102), .B2(n20085), .A(n14101), .ZN(P1_U3000) );
  INV_X1 U17405 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14103) );
  OAI21_X1 U17406 ( .B1(n14111), .B2(n14115), .A(n14103), .ZN(n14106) );
  OAI21_X1 U17407 ( .B1(n14111), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14110), .ZN(n14112) );
  AOI21_X1 U17408 ( .B1(n14113), .B2(n20071), .A(n14112), .ZN(n14114) );
  XNOR2_X1 U17409 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14117) );
  NOR2_X1 U17410 ( .A1(n14124), .A2(n14117), .ZN(n14118) );
  AOI211_X1 U17411 ( .C1(n14120), .C2(n20071), .A(n14119), .B(n14118), .ZN(
        n14122) );
  NAND2_X1 U17412 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14121) );
  OAI211_X1 U17413 ( .C1(n14123), .C2(n20085), .A(n14122), .B(n14121), .ZN(
        P1_U3003) );
  NOR2_X1 U17414 ( .A1(n14124), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14128) );
  OAI21_X1 U17415 ( .B1(n14126), .B2(n20083), .A(n14125), .ZN(n14127) );
  AOI211_X1 U17416 ( .C1(n14129), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14128), .B(n14127), .ZN(n14130) );
  OAI21_X1 U17417 ( .B1(n14131), .B2(n20085), .A(n14130), .ZN(P1_U3004) );
  XNOR2_X1 U17418 ( .A(n14146), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14135) );
  NOR2_X1 U17419 ( .A1(n14132), .A2(n20083), .ZN(n14133) );
  AOI211_X1 U17420 ( .C1(n14135), .C2(n14143), .A(n14134), .B(n14133), .ZN(
        n14138) );
  INV_X1 U17421 ( .A(n14147), .ZN(n14136) );
  NAND2_X1 U17422 ( .A1(n14136), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14137) );
  OAI211_X1 U17423 ( .C1(n14139), .C2(n20085), .A(n14138), .B(n14137), .ZN(
        P1_U3005) );
  INV_X1 U17424 ( .A(n14140), .ZN(n14142) );
  AOI21_X1 U17425 ( .B1(n14142), .B2(n20071), .A(n14141), .ZN(n14145) );
  NAND2_X1 U17426 ( .A1(n14143), .A2(n14146), .ZN(n14144) );
  OAI211_X1 U17427 ( .C1(n14147), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14148) );
  AOI21_X1 U17428 ( .B1(n14149), .B2(n20075), .A(n14148), .ZN(n14150) );
  INV_X1 U17429 ( .A(n14150), .ZN(P1_U3006) );
  INV_X1 U17430 ( .A(n14151), .ZN(n14161) );
  INV_X1 U17431 ( .A(n14162), .ZN(n14152) );
  NOR3_X1 U17432 ( .A1(n14152), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14165), .ZN(n14153) );
  AOI211_X1 U17433 ( .C1(n20071), .C2(n14155), .A(n14154), .B(n14153), .ZN(
        n14160) );
  OAI21_X1 U17434 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14157), .A(
        n14156), .ZN(n14158) );
  NAND2_X1 U17435 ( .A1(n14158), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14159) );
  OAI211_X1 U17436 ( .C1(n14161), .C2(n20085), .A(n14160), .B(n14159), .ZN(
        P1_U3007) );
  NAND2_X1 U17437 ( .A1(n14162), .A2(n14165), .ZN(n14164) );
  OAI211_X1 U17438 ( .C1(n14166), .C2(n14165), .A(n14164), .B(n14163), .ZN(
        n14167) );
  AOI21_X1 U17439 ( .B1(n20071), .B2(n15923), .A(n14167), .ZN(n14168) );
  OAI21_X1 U17440 ( .B1(n14169), .B2(n20085), .A(n14168), .ZN(P1_U3008) );
  XNOR2_X1 U17441 ( .A(n14182), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14175) );
  INV_X1 U17442 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14173) );
  AOI21_X1 U17443 ( .B1(n14171), .B2(n20071), .A(n14170), .ZN(n14172) );
  OAI21_X1 U17444 ( .B1(n14179), .B2(n14173), .A(n14172), .ZN(n14174) );
  AOI21_X1 U17445 ( .B1(n14183), .B2(n14175), .A(n14174), .ZN(n14176) );
  OAI21_X1 U17446 ( .B1(n14177), .B2(n20085), .A(n14176), .ZN(P1_U3009) );
  OAI21_X1 U17447 ( .B1(n15937), .B2(n20083), .A(n14178), .ZN(n14181) );
  NOR2_X1 U17448 ( .A1(n14179), .A2(n14182), .ZN(n14180) );
  AOI211_X1 U17449 ( .C1(n14183), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14184) );
  OAI21_X1 U17450 ( .B1(n14185), .B2(n20085), .A(n14184), .ZN(P1_U3010) );
  INV_X1 U17451 ( .A(n14186), .ZN(n14199) );
  NAND2_X1 U17452 ( .A1(n14188), .A2(n14187), .ZN(n14189) );
  NAND2_X1 U17453 ( .A1(n14190), .A2(n14189), .ZN(n16019) );
  INV_X1 U17454 ( .A(n16019), .ZN(n14194) );
  NOR4_X1 U17455 ( .A1(n14209), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14191), .A4(n14202), .ZN(n14192) );
  AOI211_X1 U17456 ( .C1(n20071), .C2(n14194), .A(n14193), .B(n14192), .ZN(
        n14198) );
  AOI21_X1 U17457 ( .B1(n14195), .B2(n14232), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14196) );
  OAI21_X1 U17458 ( .B1(n14196), .B2(n14205), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14197) );
  OAI211_X1 U17459 ( .C1(n14199), .C2(n20085), .A(n14198), .B(n14197), .ZN(
        P1_U3011) );
  INV_X1 U17460 ( .A(n14200), .ZN(n14201) );
  OAI21_X1 U17461 ( .B1(n15960), .B2(n20083), .A(n14201), .ZN(n14204) );
  NOR3_X1 U17462 ( .A1(n14209), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14202), .ZN(n14203) );
  AOI211_X1 U17463 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14205), .A(
        n14204), .B(n14203), .ZN(n14206) );
  OAI21_X1 U17464 ( .B1(n14207), .B2(n20085), .A(n14206), .ZN(P1_U3012) );
  INV_X1 U17465 ( .A(n15963), .ZN(n14213) );
  INV_X1 U17466 ( .A(n14208), .ZN(n14212) );
  NOR2_X1 U17467 ( .A1(n16114), .A2(n14209), .ZN(n16104) );
  AND3_X1 U17468 ( .A1(n14210), .A2(n14216), .A3(n16104), .ZN(n14211) );
  AOI211_X1 U17469 ( .C1(n14213), .C2(n20071), .A(n14212), .B(n14211), .ZN(
        n14219) );
  AOI211_X1 U17470 ( .C1(n16114), .C2(n20077), .A(n14215), .B(n14214), .ZN(
        n16107) );
  OAI21_X1 U17471 ( .B1(n14217), .B2(n14216), .A(n16107), .ZN(n14223) );
  NAND2_X1 U17472 ( .A1(n14223), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14218) );
  OAI211_X1 U17473 ( .C1(n14220), .C2(n20085), .A(n14219), .B(n14218), .ZN(
        P1_U3013) );
  NAND2_X1 U17474 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16094) );
  INV_X1 U17475 ( .A(n16104), .ZN(n16093) );
  OAI21_X1 U17476 ( .B1(n16094), .B2(n16093), .A(n13553), .ZN(n14224) );
  OAI21_X1 U17477 ( .B1(n15981), .B2(n20083), .A(n14221), .ZN(n14222) );
  AOI21_X1 U17478 ( .B1(n14224), .B2(n14223), .A(n14222), .ZN(n14225) );
  OAI21_X1 U17479 ( .B1(n14226), .B2(n20085), .A(n14225), .ZN(P1_U3014) );
  NOR2_X1 U17480 ( .A1(n14227), .A2(n14232), .ZN(n14230) );
  NOR2_X1 U17481 ( .A1(n20068), .A2(n20686), .ZN(n14229) );
  NOR2_X1 U17482 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14228), .ZN(
        n16113) );
  AOI211_X1 U17483 ( .C1(n14231), .C2(n14230), .A(n14229), .B(n16113), .ZN(
        n14241) );
  INV_X1 U17484 ( .A(n14232), .ZN(n20089) );
  AOI22_X1 U17485 ( .A1(n20089), .A2(n14235), .B1(n14234), .B2(n14233), .ZN(
        n14236) );
  OAI211_X1 U17486 ( .C1(n14237), .C2(n20073), .A(n20072), .B(n14236), .ZN(
        n16112) );
  INV_X1 U17487 ( .A(n14238), .ZN(n14239) );
  AOI22_X1 U17488 ( .A1(n16112), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20071), .B2(n14239), .ZN(n14240) );
  OAI211_X1 U17489 ( .C1(n14242), .C2(n20085), .A(n14241), .B(n14240), .ZN(
        P1_U3018) );
  AOI21_X1 U17490 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n16068) );
  NOR2_X1 U17491 ( .A1(n16068), .A2(n20085), .ZN(n14259) );
  OAI21_X1 U17492 ( .B1(n14249), .B2(n20073), .A(n20072), .ZN(n14246) );
  AOI21_X1 U17493 ( .B1(n20058), .B2(n14247), .A(n14246), .ZN(n16127) );
  AOI221_X1 U17494 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16127), 
        .C1(n20056), .C2(n16127), .A(n14248), .ZN(n14258) );
  NAND3_X1 U17495 ( .A1(n14249), .A2(n14248), .A3(n16120), .ZN(n14255) );
  OR2_X1 U17496 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  AND2_X1 U17497 ( .A1(n14253), .A2(n14252), .ZN(n16024) );
  NAND2_X1 U17498 ( .A1(n20071), .A2(n16024), .ZN(n14254) );
  OAI211_X1 U17499 ( .C1(n14256), .C2(n20068), .A(n14255), .B(n14254), .ZN(
        n14257) );
  OR3_X1 U17500 ( .A1(n14259), .A2(n14258), .A3(n14257), .ZN(P1_U3019) );
  NOR2_X1 U17501 ( .A1(n14264), .A2(n14260), .ZN(n16131) );
  AOI21_X1 U17502 ( .B1(n14263), .B2(n14262), .A(n14261), .ZN(n14265) );
  OAI21_X1 U17503 ( .B1(n14265), .B2(n14264), .A(n20077), .ZN(n14266) );
  AND2_X1 U17504 ( .A1(n14266), .A2(n20072), .ZN(n16137) );
  NOR2_X1 U17505 ( .A1(n16137), .A2(n10604), .ZN(n14269) );
  OAI21_X1 U17506 ( .B1(n20083), .B2(n19875), .A(n14267), .ZN(n14268) );
  AOI211_X1 U17507 ( .C1(n16131), .C2(n10604), .A(n14269), .B(n14268), .ZN(
        n14270) );
  OAI21_X1 U17508 ( .B1(n14271), .B2(n20085), .A(n14270), .ZN(P1_U3022) );
  INV_X1 U17509 ( .A(n20103), .ZN(n20349) );
  INV_X1 U17510 ( .A(n14273), .ZN(n14272) );
  NAND2_X1 U17511 ( .A1(n12454), .A2(n14273), .ZN(n20595) );
  MUX2_X1 U17512 ( .A(n20325), .B(n20595), .S(n14274), .Z(n14276) );
  INV_X1 U17513 ( .A(n12454), .ZN(n14275) );
  NAND3_X1 U17514 ( .A1(n14276), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20451), 
        .ZN(n14277) );
  OAI211_X1 U17515 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20099), .A(n14277), 
        .B(n20510), .ZN(n14278) );
  OAI21_X1 U17516 ( .B1(n20349), .B2(n14279), .A(n14278), .ZN(n14280) );
  MUX2_X1 U17517 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14280), .S(
        n20093), .Z(P1_U3475) );
  NOR3_X1 U17518 ( .A1(n14281), .A2(n14286), .A3(n14287), .ZN(n14282) );
  AOI211_X1 U17519 ( .C1(n20544), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n15862) );
  INV_X1 U17520 ( .A(n14285), .ZN(n20722) );
  NOR3_X1 U17521 ( .A1(n14287), .A2(n14286), .A3(n20722), .ZN(n14288) );
  AOI21_X1 U17522 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14291) );
  OAI21_X1 U17523 ( .B1(n15862), .B2(n20724), .A(n14291), .ZN(n14292) );
  MUX2_X1 U17524 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14292), .S(
        n16172), .Z(P1_U3473) );
  INV_X1 U17525 ( .A(n19726), .ZN(n14293) );
  NAND2_X1 U17526 ( .A1(n15526), .A2(n14293), .ZN(n14295) );
  OAI21_X1 U17527 ( .B1(n14293), .B2(n18957), .A(n16421), .ZN(n14294) );
  MUX2_X1 U17528 ( .A(n14295), .B(n14294), .S(n11280), .Z(n14297) );
  INV_X1 U17529 ( .A(n19714), .ZN(n19733) );
  OAI21_X1 U17530 ( .B1(n19733), .B2(n16425), .A(n16427), .ZN(n14296) );
  OAI21_X1 U17531 ( .B1(n14297), .B2(n16435), .A(n14296), .ZN(n14302) );
  NOR2_X1 U17532 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14298), .ZN(n19210) );
  AOI21_X1 U17533 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n14299), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14300) );
  AOI211_X1 U17534 ( .C1(n19190), .C2(n19714), .A(n14300), .B(n18951), .ZN(
        n14301) );
  MUX2_X1 U17535 ( .A(n14302), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14301), 
        .Z(P2_U3610) );
  INV_X1 U17536 ( .A(n14303), .ZN(n14304) );
  INV_X1 U17537 ( .A(n14305), .ZN(n14306) );
  NAND2_X1 U17538 ( .A1(n11770), .A2(n14306), .ZN(n14312) );
  NAND2_X1 U17539 ( .A1(n14307), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14311) );
  NAND2_X1 U17540 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U17541 ( .A1(n14308), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14309) );
  NAND4_X1 U17542 ( .A1(n14312), .A2(n14311), .A3(n14310), .A4(n14309), .ZN(
        n14313) );
  XNOR2_X1 U17543 ( .A(n14315), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16190) );
  OAI21_X1 U17544 ( .B1(n14317), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14315), .ZN(n14941) );
  INV_X1 U17545 ( .A(n14941), .ZN(n16205) );
  AND2_X1 U17546 ( .A1(n9714), .A2(n14316), .ZN(n14318) );
  OR2_X1 U17547 ( .A1(n14318), .A2(n14317), .ZN(n14955) );
  INV_X1 U17548 ( .A(n14955), .ZN(n16223) );
  OAI21_X1 U17549 ( .B1(n14320), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n9714), .ZN(n14963) );
  INV_X1 U17550 ( .A(n14963), .ZN(n14382) );
  INV_X1 U17551 ( .A(n14322), .ZN(n14321) );
  AOI21_X1 U17552 ( .B1(n10122), .B2(n14321), .A(n14320), .ZN(n14975) );
  AOI21_X1 U17553 ( .B1(n14323), .B2(n14986), .A(n14322), .ZN(n14988) );
  OAI21_X1 U17554 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14324), .A(
        n14323), .ZN(n14996) );
  INV_X1 U17555 ( .A(n14996), .ZN(n14424) );
  AOI21_X1 U17556 ( .B1(n15005), .B2(n14341), .A(n14324), .ZN(n15007) );
  NAND2_X1 U17557 ( .A1(n14325), .A2(n14339), .ZN(n14326) );
  AND2_X1 U17558 ( .A1(n14326), .A2(n10116), .ZN(n14459) );
  AOI21_X1 U17559 ( .B1(n15054), .B2(n14337), .A(n14340), .ZN(n18980) );
  AOI21_X1 U17560 ( .B1(n20790), .B2(n14336), .A(n14338), .ZN(n19003) );
  AOI21_X1 U17561 ( .B1(n14334), .B2(n20861), .A(n9687), .ZN(n19031) );
  AOI21_X1 U17562 ( .B1(n16252), .B2(n14332), .A(n14335), .ZN(n16241) );
  AOI21_X1 U17563 ( .B1(n16262), .B2(n14331), .A(n14333), .ZN(n19064) );
  AOI21_X1 U17564 ( .B1(n16269), .B2(n14329), .A(n9686), .ZN(n16263) );
  AOI21_X1 U17565 ( .B1(n16285), .B2(n14327), .A(n14330), .ZN(n16275) );
  NAND2_X1 U17566 ( .A1(n14328), .A2(n16293), .ZN(n14515) );
  NOR2_X1 U17567 ( .A1(n16275), .A2(n14515), .ZN(n19093) );
  OAI21_X1 U17568 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14330), .A(
        n14329), .ZN(n19095) );
  NAND2_X1 U17569 ( .A1(n19093), .A2(n19095), .ZN(n14503) );
  NOR2_X1 U17570 ( .A1(n16263), .A2(n14503), .ZN(n19079) );
  OAI21_X1 U17571 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9686), .A(
        n14331), .ZN(n19080) );
  NAND2_X1 U17572 ( .A1(n19079), .A2(n19080), .ZN(n19062) );
  NOR2_X1 U17573 ( .A1(n19064), .A2(n19062), .ZN(n19054) );
  OAI21_X1 U17574 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14333), .A(
        n14332), .ZN(n19055) );
  NAND2_X1 U17575 ( .A1(n19054), .A2(n19055), .ZN(n14487) );
  NOR2_X1 U17576 ( .A1(n16241), .A2(n14487), .ZN(n19042) );
  OAI21_X1 U17577 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14335), .A(
        n14334), .ZN(n19043) );
  NAND2_X1 U17578 ( .A1(n19042), .A2(n19043), .ZN(n19030) );
  NOR2_X1 U17579 ( .A1(n19031), .A2(n19030), .ZN(n19014) );
  OAI21_X1 U17580 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9687), .A(
        n14336), .ZN(n19016) );
  NAND2_X1 U17581 ( .A1(n19014), .A2(n19016), .ZN(n19001) );
  NOR2_X1 U17582 ( .A1(n19003), .A2(n19001), .ZN(n18993) );
  OAI21_X1 U17583 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14338), .A(
        n14337), .ZN(n18994) );
  NAND2_X1 U17584 ( .A1(n18993), .A2(n18994), .ZN(n18978) );
  NOR2_X1 U17585 ( .A1(n18980), .A2(n18978), .ZN(n14474) );
  OAI21_X1 U17586 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14340), .A(
        n14339), .ZN(n15042) );
  OAI21_X1 U17587 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14342), .A(
        n14341), .ZN(n15850) );
  NOR2_X1 U17588 ( .A1(n19094), .A2(n14439), .ZN(n14423) );
  NOR2_X1 U17589 ( .A1(n14424), .A2(n14423), .ZN(n14422) );
  NOR2_X1 U17590 ( .A1(n19094), .A2(n14422), .ZN(n14415) );
  NOR2_X1 U17591 ( .A1(n14988), .A2(n14415), .ZN(n14414) );
  NOR2_X1 U17592 ( .A1(n19094), .A2(n14414), .ZN(n14390) );
  NOR2_X1 U17593 ( .A1(n14975), .A2(n14390), .ZN(n14389) );
  NOR2_X1 U17594 ( .A1(n19094), .A2(n14389), .ZN(n14381) );
  NOR2_X1 U17595 ( .A1(n14382), .A2(n14381), .ZN(n14380) );
  NOR2_X1 U17596 ( .A1(n19094), .A2(n14380), .ZN(n16222) );
  NOR2_X1 U17597 ( .A1(n16223), .A2(n16222), .ZN(n16221) );
  NOR2_X1 U17598 ( .A1(n19094), .A2(n16221), .ZN(n16204) );
  NOR2_X1 U17599 ( .A1(n16205), .A2(n16204), .ZN(n16203) );
  NOR2_X1 U17600 ( .A1(n19094), .A2(n16203), .ZN(n16191) );
  NOR2_X1 U17601 ( .A1(n16190), .A2(n16191), .ZN(n16192) );
  NOR2_X1 U17602 ( .A1(n19094), .A2(n19717), .ZN(n14565) );
  NAND2_X1 U17603 ( .A1(n16192), .A2(n14565), .ZN(n14369) );
  MUX2_X1 U17604 ( .A(n12474), .B(n14343), .S(n11720), .Z(n14519) );
  NAND2_X1 U17605 ( .A1(n14828), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14785) );
  NAND2_X1 U17606 ( .A1(n14828), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14344) );
  NOR2_X1 U17607 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n14346) );
  NOR2_X1 U17608 ( .A1(n9590), .A2(n14346), .ZN(n14347) );
  INV_X1 U17609 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U17610 ( .A1(n14664), .A2(n13493), .ZN(n14348) );
  NAND2_X1 U17611 ( .A1(n14828), .A2(n14348), .ZN(n14349) );
  NAND2_X1 U17612 ( .A1(n14828), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14842) );
  NOR2_X1 U17613 ( .A1(n11720), .A2(n14351), .ZN(n14825) );
  INV_X1 U17614 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14633) );
  NAND2_X1 U17615 ( .A1(n14828), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14868) );
  INV_X1 U17616 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14352) );
  NOR2_X1 U17617 ( .A1(n9590), .A2(n14352), .ZN(n14436) );
  INV_X1 U17618 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14611) );
  INV_X1 U17619 ( .A(n14371), .ZN(n14353) );
  INV_X1 U17620 ( .A(n14395), .ZN(n14356) );
  NAND2_X1 U17621 ( .A1(n14828), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14372) );
  INV_X1 U17622 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14354) );
  NOR2_X1 U17623 ( .A1(n9590), .A2(n14354), .ZN(n14879) );
  NAND2_X1 U17624 ( .A1(n14828), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14889) );
  NOR2_X1 U17625 ( .A1(n14893), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14355) );
  MUX2_X1 U17626 ( .A(n14356), .B(n14355), .S(n14828), .Z(n14897) );
  NOR2_X2 U17627 ( .A1(n14682), .A2(n14357), .ZN(n14363) );
  INV_X1 U17628 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U17629 ( .A1(n13471), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14360) );
  NAND2_X1 U17630 ( .A1(n14358), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n14359) );
  OAI211_X1 U17631 ( .C1(n14917), .C2(n14361), .A(n14360), .B(n14359), .ZN(
        n14362) );
  AOI22_X1 U17632 ( .A1(n14364), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19103), .ZN(n14366) );
  NAND2_X1 U17633 ( .A1(n19112), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14365) );
  OAI211_X1 U17634 ( .C1(n19127), .C2(n19107), .A(n14366), .B(n14365), .ZN(
        n14367) );
  AOI21_X1 U17635 ( .B1(n14897), .B2(n19104), .A(n14367), .ZN(n14368) );
  OAI211_X1 U17636 ( .C1(n15140), .C2(n19021), .A(n14369), .B(n14368), .ZN(
        P2_U2824) );
  AOI21_X1 U17637 ( .B1(n14370), .B2(n14388), .A(n14583), .ZN(n15180) );
  OR2_X1 U17638 ( .A1(n14372), .A2(n14371), .ZN(n14373) );
  NAND2_X1 U17639 ( .A1(n14881), .A2(n14373), .ZN(n14781) );
  OR2_X1 U17640 ( .A1(n14397), .A2(n14374), .ZN(n14375) );
  AND2_X1 U17641 ( .A1(n14687), .A2(n14375), .ZN(n15184) );
  NAND2_X1 U17642 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19087), .ZN(n14377) );
  AOI22_X1 U17643 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19112), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19103), .ZN(n14376) );
  NAND2_X1 U17644 ( .A1(n14377), .A2(n14376), .ZN(n14378) );
  AOI21_X1 U17645 ( .B1(n15184), .B2(n19070), .A(n14378), .ZN(n14379) );
  OAI21_X1 U17646 ( .B1(n14781), .B2(n19075), .A(n14379), .ZN(n14384) );
  AOI211_X1 U17647 ( .C1(n14382), .C2(n14381), .A(n14380), .B(n19717), .ZN(
        n14383) );
  AOI211_X1 U17648 ( .C1(n19115), .C2(n15180), .A(n14384), .B(n14383), .ZN(
        n14385) );
  INV_X1 U17649 ( .A(n14385), .ZN(P2_U2828) );
  NAND2_X1 U17650 ( .A1(n9644), .A2(n14386), .ZN(n14387) );
  NAND2_X1 U17651 ( .A1(n14388), .A2(n14387), .ZN(n15202) );
  AOI211_X1 U17652 ( .C1(n14975), .C2(n14390), .A(n14389), .B(n19717), .ZN(
        n14391) );
  INV_X1 U17653 ( .A(n14391), .ZN(n14403) );
  NAND2_X1 U17654 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n14392), .ZN(n14393) );
  NOR2_X1 U17655 ( .A1(n11720), .A2(n14393), .ZN(n14394) );
  NOR2_X1 U17656 ( .A1(n14395), .A2(n14394), .ZN(n14885) );
  OAI21_X1 U17657 ( .B1(n14396), .B2(n14398), .A(n13465), .ZN(n15206) );
  AOI22_X1 U17658 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19112), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19087), .ZN(n14400) );
  NAND2_X1 U17659 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19103), .ZN(
        n14399) );
  OAI211_X1 U17660 ( .C1(n15206), .C2(n19107), .A(n14400), .B(n14399), .ZN(
        n14401) );
  AOI21_X1 U17661 ( .B1(n14885), .B2(n19104), .A(n14401), .ZN(n14402) );
  OAI211_X1 U17662 ( .C1(n19021), .C2(n15202), .A(n14403), .B(n14402), .ZN(
        P2_U2829) );
  NAND2_X1 U17663 ( .A1(n9661), .A2(n14404), .ZN(n14405) );
  NAND2_X1 U17664 ( .A1(n9644), .A2(n14405), .ZN(n15212) );
  NAND2_X1 U17665 ( .A1(n14428), .A2(n14406), .ZN(n14407) );
  NAND2_X1 U17666 ( .A1(n14408), .A2(n14407), .ZN(n15217) );
  NAND2_X1 U17667 ( .A1(n14828), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14409) );
  MUX2_X1 U17668 ( .A(n14409), .B(P2_EBX_REG_25__SCAN_IN), .S(n14419), .Z(
        n14410) );
  NAND2_X1 U17669 ( .A1(n14410), .A2(n14819), .ZN(n14884) );
  OAI22_X1 U17670 ( .A1(n14884), .A2(n19075), .B1(n16207), .B2(n14986), .ZN(
        n14411) );
  INV_X1 U17671 ( .A(n14411), .ZN(n14413) );
  AOI22_X1 U17672 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19112), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19087), .ZN(n14412) );
  OAI211_X1 U17673 ( .C1(n15217), .C2(n19107), .A(n14413), .B(n14412), .ZN(
        n14417) );
  AOI211_X1 U17674 ( .C1(n14988), .C2(n14415), .A(n14414), .B(n19717), .ZN(
        n14416) );
  NOR2_X1 U17675 ( .A1(n14417), .A2(n14416), .ZN(n14418) );
  OAI21_X1 U17676 ( .B1(n15212), .B2(n19021), .A(n14418), .ZN(P2_U2830) );
  NAND2_X1 U17677 ( .A1(n14828), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14421) );
  INV_X1 U17678 ( .A(n14419), .ZN(n14420) );
  OAI211_X1 U17679 ( .C1(n14438), .C2(n14421), .A(n14420), .B(n14819), .ZN(
        n14874) );
  AOI211_X1 U17680 ( .C1(n14424), .C2(n14423), .A(n14422), .B(n19717), .ZN(
        n14425) );
  INV_X1 U17681 ( .A(n14425), .ZN(n14435) );
  OR2_X1 U17682 ( .A1(n14444), .A2(n14426), .ZN(n14427) );
  NAND2_X1 U17683 ( .A1(n9661), .A2(n14427), .ZN(n15232) );
  INV_X1 U17684 ( .A(n15232), .ZN(n14433) );
  OAI21_X1 U17685 ( .B1(n14447), .B2(n14429), .A(n14428), .ZN(n15228) );
  AOI22_X1 U17686 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19112), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19087), .ZN(n14431) );
  NAND2_X1 U17687 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19103), .ZN(
        n14430) );
  OAI211_X1 U17688 ( .C1(n15228), .C2(n19107), .A(n14431), .B(n14430), .ZN(
        n14432) );
  AOI21_X1 U17689 ( .B1(n14433), .B2(n19115), .A(n14432), .ZN(n14434) );
  OAI211_X1 U17690 ( .C1(n19075), .C2(n14874), .A(n14435), .B(n14434), .ZN(
        P2_U2831) );
  AND2_X1 U17691 ( .A1(n14871), .A2(n14436), .ZN(n14437) );
  INV_X1 U17692 ( .A(n14873), .ZN(n14453) );
  AOI211_X1 U17693 ( .C1(n15007), .C2(n14440), .A(n14439), .B(n19717), .ZN(
        n14441) );
  INV_X1 U17694 ( .A(n14441), .ZN(n14452) );
  NOR2_X1 U17695 ( .A1(n14622), .A2(n14442), .ZN(n14443) );
  OR2_X1 U17696 ( .A1(n14444), .A2(n14443), .ZN(n15009) );
  INV_X1 U17697 ( .A(n15009), .ZN(n15242) );
  NOR2_X1 U17698 ( .A1(n9648), .A2(n14445), .ZN(n14446) );
  OR2_X1 U17699 ( .A1(n14447), .A2(n14446), .ZN(n16231) );
  NAND2_X1 U17700 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19087), .ZN(n14449) );
  AOI22_X1 U17701 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19112), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19103), .ZN(n14448) );
  OAI211_X1 U17702 ( .C1(n19107), .C2(n16231), .A(n14449), .B(n14448), .ZN(
        n14450) );
  AOI21_X1 U17703 ( .B1(n15242), .B2(n19115), .A(n14450), .ZN(n14451) );
  OAI211_X1 U17704 ( .C1(n19075), .C2(n14453), .A(n14452), .B(n14451), .ZN(
        P2_U2832) );
  NOR2_X1 U17705 ( .A1(n9590), .A2(n14454), .ZN(n14457) );
  AOI21_X1 U17706 ( .B1(n14457), .B2(n14456), .A(n14455), .ZN(n14814) );
  INV_X1 U17707 ( .A(n14814), .ZN(n14471) );
  INV_X1 U17708 ( .A(n14459), .ZN(n15031) );
  INV_X1 U17709 ( .A(n14473), .ZN(n14458) );
  AOI221_X1 U17710 ( .B1(n14459), .B2(n14473), .C1(n15031), .C2(n14458), .A(
        n19717), .ZN(n14461) );
  OAI22_X1 U17711 ( .A1(n19109), .A2(n14454), .B1(n19770), .B2(n19091), .ZN(
        n14460) );
  AOI211_X1 U17712 ( .C1(n19103), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14461), .B(n14460), .ZN(n14470) );
  NAND2_X1 U17713 ( .A1(n14462), .A2(n14463), .ZN(n14464) );
  AND2_X1 U17714 ( .A1(n14621), .A2(n14464), .ZN(n15268) );
  NAND2_X1 U17715 ( .A1(n14483), .A2(n14466), .ZN(n14467) );
  NAND2_X1 U17716 ( .A1(n14719), .A2(n14467), .ZN(n15265) );
  INV_X1 U17717 ( .A(n15265), .ZN(n14468) );
  AOI22_X1 U17718 ( .A1(n15268), .A2(n19115), .B1(n14468), .B2(n19070), .ZN(
        n14469) );
  OAI211_X1 U17719 ( .C1(n14471), .C2(n19075), .A(n14470), .B(n14469), .ZN(
        P2_U2834) );
  NAND3_X1 U17720 ( .A1(n14827), .A2(P2_EBX_REG_20__SCAN_IN), .A3(n14828), 
        .ZN(n14472) );
  OAI211_X1 U17721 ( .C1(n14827), .C2(P2_EBX_REG_20__SCAN_IN), .A(n14472), .B(
        n14819), .ZN(n14816) );
  NAND2_X1 U17722 ( .A1(n19094), .A2(n19098), .ZN(n14563) );
  AOI22_X1 U17723 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19112), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19103), .ZN(n14476) );
  OAI211_X1 U17724 ( .C1(n14474), .C2(n15042), .A(n19098), .B(n14473), .ZN(
        n14475) );
  OAI211_X1 U17725 ( .C1(n14563), .C2(n15042), .A(n14476), .B(n14475), .ZN(
        n14477) );
  INV_X1 U17726 ( .A(n14477), .ZN(n14486) );
  OR2_X1 U17727 ( .A1(n14640), .A2(n14478), .ZN(n14479) );
  NAND2_X1 U17728 ( .A1(n14462), .A2(n14479), .ZN(n15045) );
  INV_X1 U17729 ( .A(n15045), .ZN(n15283) );
  OR2_X1 U17730 ( .A1(n14481), .A2(n14480), .ZN(n14482) );
  NAND2_X1 U17731 ( .A1(n14483), .A2(n14482), .ZN(n15286) );
  OAI22_X1 U17732 ( .A1(n19109), .A2(n14633), .B1(n15286), .B2(n19107), .ZN(
        n14484) );
  AOI21_X1 U17733 ( .B1(n15283), .B2(n19115), .A(n14484), .ZN(n14485) );
  OAI211_X1 U17734 ( .C1(n19075), .C2(n14816), .A(n14486), .B(n14485), .ZN(
        P2_U2835) );
  NAND2_X1 U17735 ( .A1(n9591), .A2(n14487), .ZN(n14488) );
  XNOR2_X1 U17736 ( .A(n16241), .B(n14488), .ZN(n14501) );
  NOR2_X1 U17737 ( .A1(n14490), .A2(n14489), .ZN(n14491) );
  NOR2_X1 U17738 ( .A1(n14492), .A2(n14491), .ZN(n16249) );
  NAND2_X1 U17739 ( .A1(n16249), .A2(n19115), .ZN(n14498) );
  AOI21_X1 U17740 ( .B1(n14494), .B2(n14493), .A(n9688), .ZN(n19137) );
  XNOR2_X1 U17741 ( .A(n14812), .B(n9707), .ZN(n14858) );
  AOI22_X1 U17742 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19103), .B1(
        n19104), .B2(n14858), .ZN(n14495) );
  OAI21_X1 U17743 ( .B1(n19109), .B2(n14345), .A(n14495), .ZN(n14496) );
  AOI211_X1 U17744 ( .C1(n19137), .C2(n19070), .A(n19111), .B(n14496), .ZN(
        n14497) );
  OAI211_X1 U17745 ( .C1(n19091), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        n14500) );
  AOI21_X1 U17746 ( .B1(n14501), .B2(n19098), .A(n14500), .ZN(n14502) );
  INV_X1 U17747 ( .A(n14502), .ZN(P2_U2842) );
  NAND2_X1 U17748 ( .A1(n9591), .A2(n14503), .ZN(n14504) );
  XNOR2_X1 U17749 ( .A(n16263), .B(n14504), .ZN(n14505) );
  NAND2_X1 U17750 ( .A1(n14505), .A2(n19098), .ZN(n14514) );
  NAND2_X1 U17751 ( .A1(n14828), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14506) );
  XNOR2_X1 U17752 ( .A(n14507), .B(n14506), .ZN(n14800) );
  AOI22_X1 U17753 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19103), .B1(
        n19104), .B2(n14800), .ZN(n14508) );
  OAI21_X1 U17754 ( .B1(n19109), .B2(n14509), .A(n14508), .ZN(n14510) );
  NOR2_X1 U17755 ( .A1(n19111), .A2(n14510), .ZN(n14511) );
  OAI21_X1 U17756 ( .B1(n19107), .B2(n15390), .A(n14511), .ZN(n14512) );
  AOI21_X1 U17757 ( .B1(n19112), .B2(P2_REIP_REG_9__SCAN_IN), .A(n14512), .ZN(
        n14513) );
  OAI211_X1 U17758 ( .C1(n15387), .C2(n19021), .A(n14514), .B(n14513), .ZN(
        P2_U2846) );
  NAND2_X1 U17759 ( .A1(n9591), .A2(n14515), .ZN(n14516) );
  XNOR2_X1 U17760 ( .A(n16275), .B(n14516), .ZN(n14517) );
  NAND2_X1 U17761 ( .A1(n14517), .A2(n19098), .ZN(n14525) );
  OAI21_X1 U17762 ( .B1(n19091), .B2(n14518), .A(n19089), .ZN(n14523) );
  XNOR2_X1 U17763 ( .A(n14520), .B(n9929), .ZN(n14789) );
  AOI22_X1 U17764 ( .A1(n14789), .A2(n19104), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19087), .ZN(n14521) );
  OAI21_X1 U17765 ( .B1(n16285), .B2(n16207), .A(n14521), .ZN(n14522) );
  AOI211_X1 U17766 ( .C1(n16349), .C2(n19115), .A(n14523), .B(n14522), .ZN(
        n14524) );
  OAI211_X1 U17767 ( .C1(n19107), .C2(n14526), .A(n14525), .B(n14524), .ZN(
        P2_U2848) );
  NAND2_X1 U17768 ( .A1(n9591), .A2(n14527), .ZN(n14528) );
  XNOR2_X1 U17769 ( .A(n16294), .B(n14528), .ZN(n14529) );
  NAND2_X1 U17770 ( .A1(n14529), .A2(n19098), .ZN(n14536) );
  INV_X1 U17771 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14531) );
  AOI22_X1 U17772 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19103), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19087), .ZN(n14530) );
  OAI211_X1 U17773 ( .C1(n19091), .C2(n14531), .A(n14530), .B(n19089), .ZN(
        n14534) );
  NOR2_X1 U17774 ( .A1(n19075), .A2(n14532), .ZN(n14533) );
  AOI211_X1 U17775 ( .C1(n16357), .C2(n19115), .A(n14534), .B(n14533), .ZN(
        n14535) );
  OAI211_X1 U17776 ( .C1(n19107), .C2(n16354), .A(n14536), .B(n14535), .ZN(
        P2_U2850) );
  NAND2_X1 U17777 ( .A1(n9591), .A2(n14537), .ZN(n14538) );
  XNOR2_X1 U17778 ( .A(n14539), .B(n14538), .ZN(n14540) );
  NAND2_X1 U17779 ( .A1(n14540), .A2(n19098), .ZN(n14550) );
  OAI22_X1 U17780 ( .A1(n14541), .A2(n16207), .B1(n19745), .B2(n19091), .ZN(
        n14545) );
  OAI22_X1 U17781 ( .A1(n19075), .A2(n14543), .B1(n19109), .B2(n14542), .ZN(
        n14544) );
  AOI211_X1 U17782 ( .C1(n19797), .C2(n19070), .A(n14545), .B(n14544), .ZN(
        n14549) );
  NAND2_X1 U17783 ( .A1(n19803), .A2(n19116), .ZN(n14548) );
  NAND2_X1 U17784 ( .A1(n14546), .A2(n19115), .ZN(n14547) );
  NAND4_X1 U17785 ( .A1(n14550), .A2(n14549), .A3(n14548), .A4(n14547), .ZN(
        P2_U2852) );
  AOI211_X1 U17786 ( .C1(n15439), .C2(n14552), .A(n19094), .B(n14551), .ZN(
        n15447) );
  INV_X1 U17787 ( .A(n15447), .ZN(n14561) );
  OAI22_X1 U17788 ( .A1(n19075), .A2(n14553), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14563), .ZN(n14554) );
  AOI21_X1 U17789 ( .B1(n19070), .B2(n19825), .A(n14554), .ZN(n14555) );
  OAI21_X1 U17790 ( .B1(n15429), .B2(n19021), .A(n14555), .ZN(n14559) );
  AOI22_X1 U17791 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19103), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19112), .ZN(n14556) );
  OAI21_X1 U17792 ( .B1(n19109), .B2(n14557), .A(n14556), .ZN(n14558) );
  AOI211_X1 U17793 ( .C1(n19116), .C2(n19823), .A(n14559), .B(n14558), .ZN(
        n14560) );
  OAI21_X1 U17794 ( .B1(n14561), .B2(n19717), .A(n14560), .ZN(P2_U2854) );
  AOI21_X1 U17795 ( .B1(n16207), .B2(n14563), .A(n14562), .ZN(n14564) );
  AOI21_X1 U17796 ( .B1(n14565), .B2(n15439), .A(n14564), .ZN(n14571) );
  AOI22_X1 U17797 ( .A1(n19087), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n16370), .B2(
        n19070), .ZN(n14568) );
  NAND2_X1 U17798 ( .A1(n19104), .A2(n14566), .ZN(n14567) );
  OAI211_X1 U17799 ( .C1(n12092), .C2(n19091), .A(n14568), .B(n14567), .ZN(
        n14569) );
  AOI21_X1 U17800 ( .B1(n16368), .B2(n19115), .A(n14569), .ZN(n14570) );
  OAI211_X1 U17801 ( .C1(n18947), .C2(n19831), .A(n14571), .B(n14570), .ZN(
        P2_U2855) );
  INV_X1 U17802 ( .A(n15140), .ZN(n14572) );
  NAND2_X1 U17803 ( .A1(n14572), .A2(n14652), .ZN(n14573) );
  OAI21_X1 U17804 ( .B1(n14652), .B2(n14574), .A(n14573), .ZN(P2_U2856) );
  NAND2_X1 U17805 ( .A1(n14585), .A2(n14575), .ZN(n14576) );
  NAND2_X1 U17806 ( .A1(n9653), .A2(n14576), .ZN(n16212) );
  OR2_X1 U17807 ( .A1(n14578), .A2(n14577), .ZN(n14679) );
  NAND3_X1 U17808 ( .A1(n14679), .A2(n14579), .A3(n14658), .ZN(n14581) );
  NAND2_X1 U17809 ( .A1(n14659), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14580) );
  OAI211_X1 U17810 ( .C1(n14659), .C2(n16212), .A(n14581), .B(n14580), .ZN(
        P2_U2858) );
  OR2_X1 U17811 ( .A1(n14583), .A2(n14582), .ZN(n14584) );
  NAND2_X1 U17812 ( .A1(n14585), .A2(n14584), .ZN(n16218) );
  NAND2_X1 U17813 ( .A1(n14587), .A2(n14586), .ZN(n14589) );
  XNOR2_X1 U17814 ( .A(n14589), .B(n14588), .ZN(n14695) );
  NAND2_X1 U17815 ( .A1(n14695), .A2(n14658), .ZN(n14591) );
  NAND2_X1 U17816 ( .A1(n14659), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14590) );
  OAI211_X1 U17817 ( .C1(n16218), .C2(n14659), .A(n14591), .B(n14590), .ZN(
        P2_U2859) );
  OAI21_X1 U17818 ( .B1(n14592), .B2(n14594), .A(n14593), .ZN(n14702) );
  NAND2_X1 U17819 ( .A1(n14659), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17820 ( .A1(n15180), .A2(n14652), .ZN(n14595) );
  OAI211_X1 U17821 ( .C1(n14702), .C2(n14677), .A(n14596), .B(n14595), .ZN(
        P2_U2860) );
  OAI21_X1 U17822 ( .B1(n14599), .B2(n14598), .A(n14597), .ZN(n14707) );
  NOR2_X1 U17823 ( .A1(n15202), .A2(n14659), .ZN(n14600) );
  AOI21_X1 U17824 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14659), .A(n14600), .ZN(
        n14601) );
  OAI21_X1 U17825 ( .B1(n14707), .B2(n14677), .A(n14601), .ZN(P2_U2861) );
  MUX2_X1 U17826 ( .A(n15212), .B(n14604), .S(n14659), .Z(n14605) );
  OAI21_X1 U17827 ( .B1(n14712), .B2(n14677), .A(n14605), .ZN(P2_U2862) );
  AOI21_X1 U17828 ( .B1(n14606), .B2(n14608), .A(n14607), .ZN(n14609) );
  XOR2_X1 U17829 ( .A(n14610), .B(n14609), .Z(n14717) );
  MUX2_X1 U17830 ( .A(n15232), .B(n14611), .S(n14659), .Z(n14612) );
  OAI21_X1 U17831 ( .B1(n14717), .B2(n14677), .A(n14612), .ZN(P2_U2863) );
  AOI21_X1 U17832 ( .B1(n14613), .B2(n14615), .A(n14614), .ZN(n16234) );
  NAND2_X1 U17833 ( .A1(n16234), .A2(n14658), .ZN(n14617) );
  NAND2_X1 U17834 ( .A1(n14659), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14616) );
  OAI211_X1 U17835 ( .C1(n15009), .C2(n14659), .A(n14617), .B(n14616), .ZN(
        P2_U2864) );
  AOI21_X1 U17836 ( .B1(n14619), .B2(n14618), .A(n13265), .ZN(n14726) );
  NAND2_X1 U17837 ( .A1(n14726), .A2(n14658), .ZN(n14625) );
  AND2_X1 U17838 ( .A1(n14621), .A2(n14620), .ZN(n14623) );
  OR2_X1 U17839 ( .A1(n14623), .A2(n14622), .ZN(n15250) );
  INV_X1 U17840 ( .A(n15250), .ZN(n15855) );
  NAND2_X1 U17841 ( .A1(n15855), .A2(n14652), .ZN(n14624) );
  OAI211_X1 U17842 ( .C1(n14652), .C2(n13512), .A(n14625), .B(n14624), .ZN(
        P2_U2865) );
  INV_X1 U17843 ( .A(n14618), .ZN(n14627) );
  AOI21_X1 U17844 ( .B1(n14628), .B2(n14626), .A(n14627), .ZN(n14732) );
  NAND2_X1 U17845 ( .A1(n14732), .A2(n14658), .ZN(n14630) );
  NAND2_X1 U17846 ( .A1(n15268), .A2(n14652), .ZN(n14629) );
  OAI211_X1 U17847 ( .C1(n14652), .C2(n14454), .A(n14630), .B(n14629), .ZN(
        P2_U2866) );
  OAI21_X1 U17848 ( .B1(n14631), .B2(n14632), .A(n14626), .ZN(n14739) );
  MUX2_X1 U17849 ( .A(n15045), .B(n14633), .S(n14659), .Z(n14634) );
  OAI21_X1 U17850 ( .B1(n14739), .B2(n14677), .A(n14634), .ZN(P2_U2867) );
  INV_X1 U17851 ( .A(n14631), .ZN(n14636) );
  OAI21_X1 U17852 ( .B1(n14635), .B2(n14637), .A(n14636), .ZN(n14748) );
  AND2_X1 U17853 ( .A1(n14649), .A2(n14638), .ZN(n14639) );
  NOR2_X1 U17854 ( .A1(n14640), .A2(n14639), .ZN(n18986) );
  INV_X1 U17855 ( .A(n18986), .ZN(n15294) );
  NOR2_X1 U17856 ( .A1(n15294), .A2(n14659), .ZN(n14641) );
  AOI21_X1 U17857 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14659), .A(n14641), .ZN(
        n14642) );
  OAI21_X1 U17858 ( .B1(n14748), .B2(n14677), .A(n14642), .ZN(P2_U2868) );
  AOI21_X1 U17859 ( .B1(n14645), .B2(n14644), .A(n14635), .ZN(n14756) );
  NAND2_X1 U17860 ( .A1(n14756), .A2(n14658), .ZN(n14651) );
  NAND2_X1 U17861 ( .A1(n14647), .A2(n14646), .ZN(n14648) );
  AND2_X1 U17862 ( .A1(n14649), .A2(n14648), .ZN(n18996) );
  NAND2_X1 U17863 ( .A1(n18996), .A2(n14652), .ZN(n14650) );
  OAI211_X1 U17864 ( .C1(n14652), .C2(n13497), .A(n14651), .B(n14650), .ZN(
        P2_U2869) );
  XNOR2_X1 U17865 ( .A(n14667), .B(n14653), .ZN(n19008) );
  INV_X1 U17866 ( .A(n14644), .ZN(n14656) );
  AOI21_X1 U17867 ( .B1(n14657), .B2(n14655), .A(n14656), .ZN(n14766) );
  NAND2_X1 U17868 ( .A1(n14766), .A2(n14658), .ZN(n14661) );
  NAND2_X1 U17869 ( .A1(n14659), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14660) );
  OAI211_X1 U17870 ( .C1(n19008), .C2(n14659), .A(n14661), .B(n14660), .ZN(
        P2_U2870) );
  OAI21_X1 U17871 ( .B1(n14662), .B2(n14663), .A(n14655), .ZN(n14780) );
  OR2_X1 U17872 ( .A1(n14652), .A2(n14664), .ZN(n14669) );
  OR2_X1 U17873 ( .A1(n9696), .A2(n14665), .ZN(n14666) );
  AND2_X1 U17874 ( .A1(n14667), .A2(n14666), .ZN(n19019) );
  NAND2_X1 U17875 ( .A1(n14652), .A2(n19019), .ZN(n14668) );
  OAI211_X1 U17876 ( .C1(n14780), .C2(n14677), .A(n14669), .B(n14668), .ZN(
        P2_U2871) );
  XNOR2_X1 U17877 ( .A(n13103), .B(n14670), .ZN(n14674) );
  XNOR2_X1 U17878 ( .A(n14672), .B(n14671), .ZN(n15343) );
  MUX2_X1 U17879 ( .A(n14832), .B(n15343), .S(n14652), .Z(n14673) );
  OAI21_X1 U17880 ( .B1(n14674), .B2(n14677), .A(n14673), .ZN(P2_U2872) );
  XNOR2_X1 U17881 ( .A(n12909), .B(n14675), .ZN(n14678) );
  INV_X1 U17882 ( .A(n16249), .ZN(n16308) );
  MUX2_X1 U17883 ( .A(n14345), .B(n16308), .S(n14652), .Z(n14676) );
  OAI21_X1 U17884 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(P2_U2874) );
  NAND3_X1 U17885 ( .A1(n14679), .A2(n14579), .A3(n16233), .ZN(n14686) );
  NAND2_X1 U17886 ( .A1(n14688), .A2(n14680), .ZN(n14681) );
  AOI22_X1 U17887 ( .A1(n19129), .A2(n16215), .B1(n19131), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U17888 ( .A1(n19132), .A2(BUF1_REG_29__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U17889 ( .A1(n16230), .A2(n19136), .ZN(n14683) );
  NAND4_X1 U17890 ( .A1(n14686), .A2(n14685), .A3(n14684), .A4(n14683), .ZN(
        P2_U2890) );
  INV_X1 U17891 ( .A(n14687), .ZN(n14690) );
  OAI21_X1 U17892 ( .B1(n14690), .B2(n14689), .A(n14688), .ZN(n15169) );
  AOI22_X1 U17893 ( .A1(n19132), .A2(BUF1_REG_28__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U17894 ( .A1(n16230), .A2(n14691), .B1(n19131), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n14692) );
  OAI211_X1 U17895 ( .C1(n14776), .C2(n15169), .A(n14693), .B(n14692), .ZN(
        n14694) );
  AOI21_X1 U17896 ( .B1(n14695), .B2(n16233), .A(n14694), .ZN(n14696) );
  INV_X1 U17897 ( .A(n14696), .ZN(P2_U2891) );
  INV_X1 U17898 ( .A(n16230), .ZN(n14698) );
  OAI22_X1 U17899 ( .A1(n14698), .A2(n14697), .B1(n19144), .B2(n19157), .ZN(
        n14699) );
  AOI21_X1 U17900 ( .B1(n19129), .B2(n15184), .A(n14699), .ZN(n14701) );
  AOI22_X1 U17901 ( .A1(n19132), .A2(BUF1_REG_27__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14700) );
  OAI211_X1 U17902 ( .C1(n14702), .C2(n14779), .A(n14701), .B(n14700), .ZN(
        P2_U2892) );
  INV_X1 U17903 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20893) );
  OAI22_X1 U17904 ( .A1(n14776), .A2(n15206), .B1(n19144), .B2(n20893), .ZN(
        n14703) );
  AOI21_X1 U17905 ( .B1(n16230), .B2(n14704), .A(n14703), .ZN(n14706) );
  AOI22_X1 U17906 ( .A1(n19132), .A2(BUF1_REG_26__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14705) );
  OAI211_X1 U17907 ( .C1(n14707), .C2(n14779), .A(n14706), .B(n14705), .ZN(
        P2_U2893) );
  INV_X1 U17908 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19160) );
  OAI22_X1 U17909 ( .A1(n14776), .A2(n15217), .B1(n19144), .B2(n19160), .ZN(
        n14708) );
  AOI21_X1 U17910 ( .B1(n16230), .B2(n14709), .A(n14708), .ZN(n14711) );
  AOI22_X1 U17911 ( .A1(n19132), .A2(BUF1_REG_25__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14710) );
  OAI211_X1 U17912 ( .C1(n14712), .C2(n14779), .A(n14711), .B(n14710), .ZN(
        P2_U2894) );
  INV_X1 U17913 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19162) );
  OAI22_X1 U17914 ( .A1(n14776), .A2(n15228), .B1(n19144), .B2(n19162), .ZN(
        n14713) );
  AOI21_X1 U17915 ( .B1(n16230), .B2(n14714), .A(n14713), .ZN(n14716) );
  AOI22_X1 U17916 ( .A1(n19132), .A2(BUF1_REG_24__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14715) );
  OAI211_X1 U17917 ( .C1(n14717), .C2(n14779), .A(n14716), .B(n14715), .ZN(
        P2_U2895) );
  AND2_X1 U17918 ( .A1(n14719), .A2(n14718), .ZN(n14720) );
  NOR2_X1 U17919 ( .A1(n9648), .A2(n14720), .ZN(n15854) );
  INV_X1 U17920 ( .A(n15854), .ZN(n14724) );
  AOI22_X1 U17921 ( .A1(n19132), .A2(BUF1_REG_22__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U17922 ( .A1(n16230), .A2(n14721), .B1(n19131), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n14722) );
  OAI211_X1 U17923 ( .C1(n14776), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        n14725) );
  AOI21_X1 U17924 ( .B1(n14726), .B2(n16233), .A(n14725), .ZN(n14727) );
  INV_X1 U17925 ( .A(n14727), .ZN(P2_U2897) );
  AOI22_X1 U17926 ( .A1(n19132), .A2(BUF1_REG_21__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14730) );
  AOI22_X1 U17927 ( .A1(n16230), .A2(n14728), .B1(n19131), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14729) );
  OAI211_X1 U17928 ( .C1(n14776), .C2(n15265), .A(n14730), .B(n14729), .ZN(
        n14731) );
  AOI21_X1 U17929 ( .B1(n14732), .B2(n16233), .A(n14731), .ZN(n14733) );
  INV_X1 U17930 ( .A(n14733), .ZN(P2_U2898) );
  AOI22_X1 U17931 ( .A1(n19132), .A2(BUF1_REG_20__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U17932 ( .A1(n16230), .A2(n14734), .B1(n19131), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n14735) );
  OAI211_X1 U17933 ( .C1(n14776), .C2(n15286), .A(n14736), .B(n14735), .ZN(
        n14737) );
  INV_X1 U17934 ( .A(n14737), .ZN(n14738) );
  OAI21_X1 U17935 ( .B1(n14739), .B2(n14779), .A(n14738), .ZN(P2_U2899) );
  INV_X1 U17936 ( .A(n14750), .ZN(n14740) );
  XNOR2_X1 U17937 ( .A(n14741), .B(n14740), .ZN(n18985) );
  INV_X1 U17938 ( .A(n18985), .ZN(n14745) );
  AOI22_X1 U17939 ( .A1(n19132), .A2(BUF1_REG_19__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U17940 ( .A1(n16230), .A2(n14742), .B1(n19131), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14743) );
  OAI211_X1 U17941 ( .C1(n14776), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        n14746) );
  INV_X1 U17942 ( .A(n14746), .ZN(n14747) );
  OAI21_X1 U17943 ( .B1(n14748), .B2(n14779), .A(n14747), .ZN(P2_U2900) );
  OR2_X1 U17944 ( .A1(n14760), .A2(n14749), .ZN(n14751) );
  NAND2_X1 U17945 ( .A1(n14751), .A2(n14750), .ZN(n19000) );
  AOI22_X1 U17946 ( .A1(n19132), .A2(BUF1_REG_18__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U17947 ( .A1(n16230), .A2(n14752), .B1(n19131), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n14753) );
  OAI211_X1 U17948 ( .C1(n14776), .C2(n19000), .A(n14754), .B(n14753), .ZN(
        n14755) );
  AOI21_X1 U17949 ( .B1(n14756), .B2(n16233), .A(n14755), .ZN(n14757) );
  INV_X1 U17950 ( .A(n14757), .ZN(P2_U2901) );
  NOR2_X1 U17951 ( .A1(n14772), .A2(n14758), .ZN(n14759) );
  NOR2_X1 U17952 ( .A1(n14760), .A2(n14759), .ZN(n19009) );
  INV_X1 U17953 ( .A(n19009), .ZN(n14764) );
  AOI22_X1 U17954 ( .A1(n19132), .A2(BUF1_REG_17__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U17955 ( .A1(n16230), .A2(n14761), .B1(n19131), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14762) );
  OAI211_X1 U17956 ( .C1(n14776), .C2(n14764), .A(n14763), .B(n14762), .ZN(
        n14765) );
  AOI21_X1 U17957 ( .B1(n14766), .B2(n16233), .A(n14765), .ZN(n14767) );
  INV_X1 U17958 ( .A(n14767), .ZN(P2_U2902) );
  AOI21_X1 U17959 ( .B1(n14770), .B2(n14769), .A(n14768), .ZN(n14771) );
  OR2_X1 U17960 ( .A1(n14772), .A2(n14771), .ZN(n19020) );
  AOI22_X1 U17961 ( .A1(n19132), .A2(BUF1_REG_16__SCAN_IN), .B1(n19130), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n14775) );
  AOI22_X1 U17962 ( .A1(n16230), .A2(n14773), .B1(n19131), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U17963 ( .C1(n14776), .C2(n19020), .A(n14775), .B(n14774), .ZN(
        n14777) );
  INV_X1 U17964 ( .A(n14777), .ZN(n14778) );
  OAI21_X1 U17965 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(P2_U2903) );
  INV_X1 U17966 ( .A(n14785), .ZN(n14786) );
  XNOR2_X1 U17967 ( .A(n14787), .B(n14786), .ZN(n19088) );
  AND2_X1 U17968 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14911) );
  NAND2_X1 U17969 ( .A1(n19088), .A2(n14911), .ZN(n15407) );
  NAND2_X1 U17970 ( .A1(n14789), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16277) );
  NAND2_X1 U17971 ( .A1(n19088), .A2(n14896), .ZN(n14788) );
  NAND2_X1 U17972 ( .A1(n14788), .A2(n15416), .ZN(n15408) );
  INV_X1 U17973 ( .A(n14789), .ZN(n14790) );
  NAND2_X1 U17974 ( .A1(n14790), .A2(n16345), .ZN(n16276) );
  AND2_X1 U17975 ( .A1(n15408), .A2(n16276), .ZN(n14791) );
  AOI21_X1 U17976 ( .B1(n14800), .B2(n14896), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15395) );
  INV_X1 U17977 ( .A(n15395), .ZN(n14792) );
  NAND2_X1 U17978 ( .A1(n14796), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14793) );
  OAI21_X1 U17979 ( .B1(n14793), .B2(n11720), .A(n14819), .ZN(n14794) );
  INV_X1 U17980 ( .A(n14794), .ZN(n14795) );
  OAI21_X1 U17981 ( .B1(n14796), .B2(P2_EBX_REG_10__SCAN_IN), .A(n14795), .ZN(
        n19076) );
  OR2_X1 U17982 ( .A1(n19076), .A2(n11643), .ZN(n14797) );
  NAND2_X1 U17983 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14798) );
  OR2_X1 U17984 ( .A1(n19076), .A2(n14798), .ZN(n15105) );
  INV_X1 U17985 ( .A(n15105), .ZN(n14802) );
  AND2_X1 U17986 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14799) );
  NAND2_X1 U17987 ( .A1(n14800), .A2(n14799), .ZN(n15394) );
  INV_X1 U17988 ( .A(n14804), .ZN(n14805) );
  NAND2_X1 U17989 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n14805), .ZN(n14806) );
  NOR2_X1 U17990 ( .A1(n11720), .A2(n14806), .ZN(n14807) );
  OR2_X1 U17991 ( .A1(n14808), .A2(n14807), .ZN(n19065) );
  OAI21_X1 U17992 ( .B1(n19065), .B2(n11643), .A(n16336), .ZN(n16254) );
  NAND2_X1 U17993 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14809) );
  NAND3_X1 U17994 ( .A1(n14828), .A2(n14810), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n14811) );
  NAND2_X1 U17995 ( .A1(n14812), .A2(n14811), .ZN(n19050) );
  XOR2_X1 U17996 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n14813), .Z(
        n15095) );
  NAND2_X1 U17997 ( .A1(n14814), .A2(n14896), .ZN(n14866) );
  INV_X1 U17998 ( .A(n14866), .ZN(n14815) );
  NOR2_X1 U17999 ( .A1(n14815), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15020) );
  NOR2_X1 U18000 ( .A1(n14816), .A2(n11643), .ZN(n14852) );
  INV_X1 U18001 ( .A(n14852), .ZN(n14817) );
  NAND2_X1 U18002 ( .A1(n14817), .A2(n15281), .ZN(n15027) );
  INV_X1 U18003 ( .A(n15027), .ZN(n15037) );
  NOR2_X1 U18004 ( .A1(n11720), .A2(n14664), .ZN(n14818) );
  MUX2_X1 U18005 ( .A(n14664), .B(n14818), .S(n14834), .Z(n14821) );
  INV_X1 U18006 ( .A(n14819), .ZN(n14820) );
  AND2_X1 U18007 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14822) );
  NAND2_X1 U18008 ( .A1(n19017), .A2(n14822), .ZN(n15024) );
  INV_X1 U18009 ( .A(n19017), .ZN(n14823) );
  OAI21_X1 U18010 ( .B1(n14823), .B2(n11643), .A(n15341), .ZN(n14824) );
  NAND2_X1 U18011 ( .A1(n15024), .A2(n14824), .ZN(n15077) );
  NAND2_X1 U18012 ( .A1(n14846), .A2(n14825), .ZN(n14826) );
  AND2_X1 U18013 ( .A1(n14827), .A2(n14826), .ZN(n18981) );
  NAND2_X1 U18014 ( .A1(n18981), .A2(n14896), .ZN(n14853) );
  INV_X1 U18015 ( .A(n15049), .ZN(n14850) );
  OAI211_X1 U18016 ( .C1(n14834), .C2(P2_EBX_REG_16__SCAN_IN), .A(
        P2_EBX_REG_17__SCAN_IN), .B(n14828), .ZN(n14829) );
  AND2_X1 U18017 ( .A1(n14844), .A2(n14829), .ZN(n19004) );
  INV_X1 U18018 ( .A(n14856), .ZN(n14831) );
  INV_X1 U18019 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14830) );
  OR2_X1 U18020 ( .A1(n14838), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14840) );
  NOR2_X1 U18021 ( .A1(n9590), .A2(n14832), .ZN(n14833) );
  NAND2_X1 U18022 ( .A1(n14840), .A2(n14833), .ZN(n14835) );
  NAND2_X1 U18023 ( .A1(n14835), .A2(n14834), .ZN(n19027) );
  INV_X1 U18024 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15322) );
  OAI21_X1 U18025 ( .B1(n19027), .B2(n11643), .A(n15322), .ZN(n15084) );
  NAND2_X1 U18026 ( .A1(n14858), .A2(n14896), .ZN(n14836) );
  NAND2_X1 U18027 ( .A1(n14836), .A2(n16244), .ZN(n16246) );
  NAND2_X1 U18028 ( .A1(n15084), .A2(n16246), .ZN(n14837) );
  NOR2_X1 U18029 ( .A1(n15068), .A2(n14837), .ZN(n14849) );
  NAND2_X1 U18030 ( .A1(n14828), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14839) );
  MUX2_X1 U18031 ( .A(n14828), .B(n14839), .S(n14838), .Z(n14841) );
  NAND2_X1 U18032 ( .A1(n19038), .A2(n14896), .ZN(n14862) );
  NAND2_X1 U18033 ( .A1(n14862), .A2(n15365), .ZN(n15354) );
  INV_X1 U18034 ( .A(n14842), .ZN(n14843) );
  NAND2_X1 U18035 ( .A1(n14844), .A2(n14843), .ZN(n14845) );
  NAND2_X1 U18036 ( .A1(n14846), .A2(n14845), .ZN(n18990) );
  OR2_X1 U18037 ( .A1(n18990), .A2(n11643), .ZN(n14847) );
  INV_X1 U18038 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15310) );
  INV_X1 U18039 ( .A(n15060), .ZN(n14848) );
  NAND4_X1 U18040 ( .A1(n14850), .A2(n14849), .A3(n15354), .A4(n14848), .ZN(
        n14851) );
  AND2_X1 U18041 ( .A1(n14852), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15038) );
  INV_X1 U18042 ( .A(n15038), .ZN(n14865) );
  INV_X1 U18043 ( .A(n14853), .ZN(n14854) );
  NAND2_X1 U18044 ( .A1(n14854), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15026) );
  INV_X1 U18045 ( .A(n15026), .ZN(n15050) );
  NAND2_X1 U18046 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14855) );
  NOR2_X1 U18047 ( .A1(n18990), .A2(n14855), .ZN(n15059) );
  INV_X1 U18048 ( .A(n15059), .ZN(n14860) );
  NAND2_X1 U18049 ( .A1(n14856), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15069) );
  NAND2_X1 U18050 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14857) );
  NOR2_X1 U18051 ( .A1(n19027), .A2(n14857), .ZN(n15023) );
  INV_X1 U18052 ( .A(n15023), .ZN(n15085) );
  INV_X1 U18053 ( .A(n14858), .ZN(n14859) );
  NAND4_X1 U18054 ( .A1(n14860), .A2(n15069), .A3(n15085), .A4(n16245), .ZN(
        n14861) );
  NOR2_X1 U18055 ( .A1(n15050), .A2(n14861), .ZN(n14864) );
  INV_X1 U18056 ( .A(n14862), .ZN(n14863) );
  NAND2_X1 U18057 ( .A1(n14863), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15355) );
  NAND4_X1 U18058 ( .A1(n14865), .A2(n14864), .A3(n15024), .A4(n15355), .ZN(
        n14867) );
  NOR2_X1 U18059 ( .A1(n14866), .A2(n15270), .ZN(n15021) );
  INV_X1 U18060 ( .A(n14868), .ZN(n14869) );
  NAND2_X1 U18061 ( .A1(n9646), .A2(n14869), .ZN(n14870) );
  AND2_X1 U18062 ( .A1(n14871), .A2(n14870), .ZN(n15856) );
  AOI21_X1 U18063 ( .B1(n15856), .B2(n14896), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15012) );
  NAND3_X1 U18064 ( .A1(n15856), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14896), .ZN(n15013) );
  NOR2_X1 U18065 ( .A1(n11643), .A2(n15245), .ZN(n14872) );
  NOR2_X1 U18066 ( .A1(n14874), .A2(n11643), .ZN(n14992) );
  NAND2_X1 U18067 ( .A1(n14885), .A2(n14896), .ZN(n14875) );
  XOR2_X1 U18068 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14875), .Z(
        n14968) );
  INV_X1 U18069 ( .A(n14968), .ZN(n14878) );
  OR2_X1 U18070 ( .A1(n14884), .A2(n11643), .ZN(n14876) );
  AND2_X2 U18071 ( .A1(n14876), .A2(n20824), .ZN(n14981) );
  INV_X1 U18072 ( .A(n14879), .ZN(n14880) );
  XNOR2_X1 U18073 ( .A(n14881), .B(n14880), .ZN(n16217) );
  NAND2_X1 U18074 ( .A1(n16217), .A2(n14896), .ZN(n14882) );
  NAND2_X1 U18075 ( .A1(n14882), .A2(n14937), .ZN(n14951) );
  INV_X1 U18076 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U18077 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14883) );
  NAND3_X1 U18078 ( .A1(n14885), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14896), .ZN(n14886) );
  XNOR2_X1 U18079 ( .A(n14890), .B(n14889), .ZN(n14895) );
  INV_X1 U18080 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14936) );
  OAI21_X1 U18081 ( .B1(n14895), .B2(n11643), .A(n14936), .ZN(n14932) );
  NAND2_X1 U18082 ( .A1(n14828), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14892) );
  XNOR2_X1 U18083 ( .A(n14893), .B(n14892), .ZN(n14894) );
  AOI21_X1 U18084 ( .B1(n14894), .B2(n14896), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14924) );
  INV_X1 U18085 ( .A(n14894), .ZN(n16194) );
  INV_X1 U18086 ( .A(n14895), .ZN(n16210) );
  NAND3_X1 U18087 ( .A1(n16210), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14896), .ZN(n14933) );
  NAND2_X1 U18088 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  XNOR2_X1 U18089 ( .A(n14898), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14899) );
  NAND2_X1 U18090 ( .A1(n16279), .A2(n16345), .ZN(n14906) );
  INV_X1 U18091 ( .A(n16279), .ZN(n14907) );
  NAND2_X1 U18092 ( .A1(n14907), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14908) );
  NOR2_X1 U18093 ( .A1(n14910), .A2(n11643), .ZN(n14909) );
  XNOR2_X1 U18094 ( .A(n14909), .B(n15416), .ZN(n15403) );
  INV_X1 U18095 ( .A(n14910), .ZN(n14912) );
  NAND2_X1 U18096 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  AND2_X1 U18097 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15366) );
  AND2_X1 U18098 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16331) );
  AND2_X1 U18099 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14914) );
  AND3_X1 U18100 ( .A1(n15366), .A2(n16331), .A3(n14914), .ZN(n15318) );
  AND3_X1 U18101 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U18102 ( .A1(n15318), .A2(n14915), .ZN(n15304) );
  NOR2_X1 U18103 ( .A1(n15310), .A2(n15304), .ZN(n15278) );
  NAND3_X1 U18104 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n15278), .ZN(n15264) );
  NOR2_X1 U18105 ( .A1(n15264), .A2(n15270), .ZN(n15124) );
  INV_X1 U18106 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15256) );
  AND2_X2 U18107 ( .A1(n14995), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14984) );
  AND2_X2 U18108 ( .A1(n14984), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14972) );
  NAND2_X1 U18109 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U18110 ( .A1(n14938), .A2(n15125), .ZN(n14916) );
  XOR2_X1 U18111 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14916), .Z(
        n15142) );
  NOR2_X1 U18112 ( .A1(n19089), .A2(n14917), .ZN(n15122) );
  NOR2_X1 U18113 ( .A1(n19224), .A2(n14918), .ZN(n14919) );
  AOI211_X1 U18114 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19215), .A(
        n15122), .B(n14919), .ZN(n14920) );
  OAI21_X1 U18115 ( .B1(n15140), .B2(n15115), .A(n14920), .ZN(n14921) );
  AOI21_X1 U18116 ( .B1(n15142), .B2(n19216), .A(n14921), .ZN(n14922) );
  NAND2_X1 U18117 ( .A1(n14923), .A2(n14933), .ZN(n14926) );
  NOR2_X1 U18118 ( .A1(n14924), .A2(n9660), .ZN(n14925) );
  XNOR2_X1 U18119 ( .A(n14926), .B(n14925), .ZN(n15154) );
  INV_X1 U18120 ( .A(n15115), .ZN(n19227) );
  NAND2_X1 U18121 ( .A1(n16295), .A2(n16190), .ZN(n14927) );
  NAND2_X1 U18122 ( .A1(n19111), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15148) );
  OAI211_X1 U18123 ( .C1(n16305), .C2(n14928), .A(n14927), .B(n15148), .ZN(
        n14930) );
  OAI21_X1 U18124 ( .B1(n15154), .B2(n19218), .A(n14931), .ZN(P2_U2984) );
  NAND2_X1 U18125 ( .A1(n14933), .A2(n14932), .ZN(n14935) );
  XOR2_X1 U18126 ( .A(n14935), .B(n14934), .Z(n15167) );
  OAI21_X1 U18127 ( .B1(n14964), .B2(n14937), .A(n14936), .ZN(n14939) );
  AND2_X1 U18128 ( .A1(n14939), .A2(n14938), .ZN(n15165) );
  INV_X1 U18129 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n14940) );
  NOR2_X1 U18130 ( .A1(n19089), .A2(n14940), .ZN(n15155) );
  NOR2_X1 U18131 ( .A1(n19224), .A2(n14941), .ZN(n14942) );
  AOI211_X1 U18132 ( .C1(n19215), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15155), .B(n14942), .ZN(n14943) );
  OAI21_X1 U18133 ( .B1(n16212), .B2(n15115), .A(n14943), .ZN(n14944) );
  AOI21_X1 U18134 ( .B1(n15165), .B2(n19216), .A(n14944), .ZN(n14945) );
  OAI21_X1 U18135 ( .B1(n15167), .B2(n19218), .A(n14945), .ZN(P2_U2985) );
  NAND2_X1 U18136 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  XNOR2_X1 U18137 ( .A(n14954), .B(n14953), .ZN(n15178) );
  XNOR2_X1 U18138 ( .A(n14964), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15176) );
  NOR2_X1 U18139 ( .A1(n19089), .A2(n19782), .ZN(n15172) );
  NOR2_X1 U18140 ( .A1(n19224), .A2(n14955), .ZN(n14956) );
  AOI211_X1 U18141 ( .C1(n19215), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15172), .B(n14956), .ZN(n14957) );
  OAI21_X1 U18142 ( .B1(n16218), .B2(n15115), .A(n14957), .ZN(n14958) );
  AOI21_X1 U18143 ( .B1(n15176), .B2(n19216), .A(n14958), .ZN(n14959) );
  OAI21_X1 U18144 ( .B1(n15178), .B2(n19218), .A(n14959), .ZN(P2_U2986) );
  XNOR2_X1 U18145 ( .A(n14960), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15193) );
  NOR2_X1 U18146 ( .A1(n19089), .A2(n14961), .ZN(n15181) );
  AOI21_X1 U18147 ( .B1(n19215), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15181), .ZN(n14962) );
  OAI21_X1 U18148 ( .B1(n19224), .B2(n14963), .A(n14962), .ZN(n14966) );
  OAI21_X1 U18149 ( .B1(n14972), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14964), .ZN(n15188) );
  NOR2_X1 U18150 ( .A1(n15188), .A2(n16287), .ZN(n14965) );
  OAI21_X1 U18151 ( .B1(n15193), .B2(n19218), .A(n14967), .ZN(P2_U2987) );
  AOI21_X1 U18152 ( .B1(n14982), .B2(n14979), .A(n14981), .ZN(n14969) );
  MUX2_X1 U18153 ( .A(n14979), .B(n14969), .S(n14968), .Z(n14970) );
  NAND2_X1 U18154 ( .A1(n14971), .A2(n14970), .ZN(n15211) );
  INV_X1 U18155 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15200) );
  INV_X1 U18156 ( .A(n14984), .ZN(n14973) );
  AOI21_X1 U18157 ( .B1(n15200), .B2(n14973), .A(n14972), .ZN(n15209) );
  NAND2_X1 U18158 ( .A1(n19111), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15204) );
  OAI21_X1 U18159 ( .B1(n16305), .B2(n10122), .A(n15204), .ZN(n14974) );
  AOI21_X1 U18160 ( .B1(n16295), .B2(n14975), .A(n14974), .ZN(n14976) );
  OAI21_X1 U18161 ( .B1(n15202), .B2(n15115), .A(n14976), .ZN(n14977) );
  AOI21_X1 U18162 ( .B1(n15209), .B2(n19216), .A(n14977), .ZN(n14978) );
  OAI21_X1 U18163 ( .B1(n15211), .B2(n19218), .A(n14978), .ZN(P2_U2988) );
  INV_X1 U18164 ( .A(n14979), .ZN(n14980) );
  NOR2_X1 U18165 ( .A1(n14981), .A2(n14980), .ZN(n14983) );
  XOR2_X1 U18166 ( .A(n14983), .B(n14982), .Z(n15224) );
  INV_X1 U18167 ( .A(n14995), .ZN(n14985) );
  AOI21_X1 U18168 ( .B1(n20824), .B2(n14985), .A(n14984), .ZN(n15222) );
  NOR2_X1 U18169 ( .A1(n19089), .A2(n19777), .ZN(n15215) );
  NOR2_X1 U18170 ( .A1(n16305), .A2(n14986), .ZN(n14987) );
  AOI211_X1 U18171 ( .C1(n14988), .C2(n16295), .A(n15215), .B(n14987), .ZN(
        n14989) );
  OAI21_X1 U18172 ( .B1(n15212), .B2(n15115), .A(n14989), .ZN(n14990) );
  AOI21_X1 U18173 ( .B1(n15222), .B2(n19216), .A(n14990), .ZN(n14991) );
  OAI21_X1 U18174 ( .B1(n15224), .B2(n19218), .A(n14991), .ZN(P2_U2989) );
  XNOR2_X1 U18175 ( .A(n14992), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14993) );
  XNOR2_X1 U18176 ( .A(n14994), .B(n14993), .ZN(n15237) );
  AOI21_X1 U18177 ( .B1(n15225), .B2(n15003), .A(n14995), .ZN(n15235) );
  OAI22_X1 U18178 ( .A1(n19775), .A2(n11795), .B1(n19224), .B2(n14996), .ZN(
        n14997) );
  AOI21_X1 U18179 ( .B1(n19215), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14997), .ZN(n14998) );
  OAI21_X1 U18180 ( .B1(n15232), .B2(n15115), .A(n14998), .ZN(n14999) );
  AOI21_X1 U18181 ( .B1(n15235), .B2(n19216), .A(n14999), .ZN(n15000) );
  OAI21_X1 U18182 ( .B1(n15237), .B2(n19218), .A(n15000), .ZN(P2_U2990) );
  XNOR2_X1 U18183 ( .A(n15002), .B(n15001), .ZN(n15249) );
  INV_X1 U18184 ( .A(n15003), .ZN(n15004) );
  AOI21_X1 U18185 ( .B1(n15245), .B2(n15259), .A(n15004), .ZN(n15247) );
  NOR2_X1 U18186 ( .A1(n19089), .A2(n19773), .ZN(n15241) );
  NOR2_X1 U18187 ( .A1(n16305), .A2(n15005), .ZN(n15006) );
  AOI211_X1 U18188 ( .C1(n15007), .C2(n16295), .A(n15241), .B(n15006), .ZN(
        n15008) );
  OAI21_X1 U18189 ( .B1(n15009), .B2(n15115), .A(n15008), .ZN(n15010) );
  AOI21_X1 U18190 ( .B1(n15247), .B2(n19216), .A(n15010), .ZN(n15011) );
  OAI21_X1 U18191 ( .B1(n15249), .B2(n19218), .A(n15011), .ZN(P2_U2991) );
  NAND2_X1 U18192 ( .A1(n9795), .A2(n15013), .ZN(n15014) );
  XNOR2_X1 U18193 ( .A(n15015), .B(n15014), .ZN(n15262) );
  OAI22_X1 U18194 ( .A1(n19772), .A2(n19089), .B1(n19224), .B2(n15850), .ZN(
        n15017) );
  NOR2_X1 U18195 ( .A1(n15250), .A2(n15115), .ZN(n15016) );
  AOI211_X1 U18196 ( .C1(n19215), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15017), .B(n15016), .ZN(n15019) );
  NAND2_X1 U18197 ( .A1(n15033), .A2(n15256), .ZN(n15258) );
  NAND3_X1 U18198 ( .A1(n15259), .A2(n19216), .A3(n15258), .ZN(n15018) );
  OAI211_X1 U18199 ( .C1(n15262), .C2(n19218), .A(n15019), .B(n15018), .ZN(
        P2_U2992) );
  NOR2_X1 U18200 ( .A1(n15021), .A2(n15020), .ZN(n15029) );
  INV_X1 U18201 ( .A(n16246), .ZN(n15022) );
  NAND2_X1 U18202 ( .A1(n15357), .A2(n15354), .ZN(n15359) );
  INV_X1 U18203 ( .A(n15024), .ZN(n15025) );
  AOI211_X2 U18204 ( .C1(n15048), .C2(n15026), .A(n15049), .B(n15060), .ZN(
        n15040) );
  AOI21_X1 U18205 ( .B1(n15040), .B2(n15027), .A(n15038), .ZN(n15028) );
  XOR2_X1 U18206 ( .A(n15029), .B(n15028), .Z(n15276) );
  NOR2_X1 U18207 ( .A1(n19089), .A2(n19770), .ZN(n15267) );
  AOI21_X1 U18208 ( .B1(n19215), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15267), .ZN(n15030) );
  OAI21_X1 U18209 ( .B1(n19224), .B2(n15031), .A(n15030), .ZN(n15035) );
  NOR2_X1 U18210 ( .A1(n15386), .A2(n15264), .ZN(n15041) );
  OAI21_X1 U18211 ( .B1(n15041), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15033), .ZN(n15263) );
  NOR2_X1 U18212 ( .A1(n15263), .A2(n16287), .ZN(n15034) );
  AOI211_X1 U18213 ( .C1(n19227), .C2(n15268), .A(n15035), .B(n15034), .ZN(
        n15036) );
  OAI21_X1 U18214 ( .B1(n15276), .B2(n19218), .A(n15036), .ZN(P2_U2993) );
  NOR2_X1 U18215 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  XNOR2_X1 U18216 ( .A(n15040), .B(n15039), .ZN(n15291) );
  AND2_X1 U18217 ( .A1(n15032), .A2(n15278), .ZN(n15063) );
  NAND2_X1 U18218 ( .A1(n15063), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15055) );
  AOI21_X1 U18219 ( .B1(n15055), .B2(n15281), .A(n15041), .ZN(n15289) );
  NOR2_X1 U18220 ( .A1(n19089), .A2(n19768), .ZN(n15282) );
  NOR2_X1 U18221 ( .A1(n19224), .A2(n15042), .ZN(n15043) );
  AOI211_X1 U18222 ( .C1(n19215), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15282), .B(n15043), .ZN(n15044) );
  OAI21_X1 U18223 ( .B1(n15045), .B2(n15115), .A(n15044), .ZN(n15046) );
  AOI21_X1 U18224 ( .B1(n15289), .B2(n19216), .A(n15046), .ZN(n15047) );
  OAI21_X1 U18225 ( .B1(n15291), .B2(n19218), .A(n15047), .ZN(P2_U2994) );
  NOR2_X1 U18226 ( .A1(n15048), .A2(n15060), .ZN(n15052) );
  NOR2_X1 U18227 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  XNOR2_X1 U18228 ( .A(n15052), .B(n15051), .ZN(n15303) );
  NAND2_X1 U18229 ( .A1(n16295), .A2(n18980), .ZN(n15053) );
  NAND2_X1 U18230 ( .A1(n19111), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15293) );
  OAI211_X1 U18231 ( .C1(n16305), .C2(n15054), .A(n15053), .B(n15293), .ZN(
        n15057) );
  OAI21_X1 U18232 ( .B1(n15063), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15055), .ZN(n15292) );
  NOR2_X1 U18233 ( .A1(n15292), .A2(n16287), .ZN(n15056) );
  AOI211_X1 U18234 ( .C1(n19227), .C2(n18986), .A(n15057), .B(n15056), .ZN(
        n15058) );
  OAI21_X1 U18235 ( .B1(n15303), .B2(n19218), .A(n15058), .ZN(P2_U2995) );
  NOR2_X1 U18236 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  XNOR2_X1 U18237 ( .A(n9677), .B(n15061), .ZN(n15315) );
  INV_X1 U18238 ( .A(n15304), .ZN(n15062) );
  NAND2_X1 U18239 ( .A1(n15032), .A2(n15062), .ZN(n15074) );
  AOI21_X1 U18240 ( .B1(n15310), .B2(n15074), .A(n15063), .ZN(n15313) );
  NAND2_X1 U18241 ( .A1(n18996), .A2(n19227), .ZN(n15065) );
  NOR2_X1 U18242 ( .A1(n11795), .A2(n19764), .ZN(n15307) );
  AOI21_X1 U18243 ( .B1(n19215), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15307), .ZN(n15064) );
  OAI211_X1 U18244 ( .C1(n18994), .C2(n19224), .A(n15065), .B(n15064), .ZN(
        n15066) );
  AOI21_X1 U18245 ( .B1(n15313), .B2(n19216), .A(n15066), .ZN(n15067) );
  OAI21_X1 U18246 ( .B1(n15315), .B2(n19218), .A(n15067), .ZN(P2_U2996) );
  NAND2_X1 U18247 ( .A1(n10080), .A2(n15069), .ZN(n15070) );
  XNOR2_X1 U18248 ( .A(n15071), .B(n15070), .ZN(n15329) );
  NAND2_X1 U18249 ( .A1(n19111), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15324) );
  OAI21_X1 U18250 ( .B1(n16305), .B2(n20790), .A(n15324), .ZN(n15073) );
  NOR2_X1 U18251 ( .A1(n19008), .A2(n15115), .ZN(n15072) );
  AOI211_X1 U18252 ( .C1(n16295), .C2(n19003), .A(n15073), .B(n15072), .ZN(
        n15076) );
  OAI211_X1 U18253 ( .C1(n15323), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19216), .B(n15074), .ZN(n15075) );
  OAI211_X1 U18254 ( .C1(n15329), .C2(n19218), .A(n15076), .B(n15075), .ZN(
        P2_U2997) );
  NAND2_X1 U18255 ( .A1(n15078), .A2(n15077), .ZN(n15331) );
  NAND2_X1 U18256 ( .A1(n15331), .A2(n16302), .ZN(n15083) );
  NOR2_X1 U18257 ( .A1(n19089), .A2(n19761), .ZN(n15335) );
  AOI21_X1 U18258 ( .B1(n19215), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15335), .ZN(n15079) );
  OAI21_X1 U18259 ( .B1(n19224), .B2(n19016), .A(n15079), .ZN(n15081) );
  AOI211_X1 U18260 ( .C1(n15341), .C2(n15334), .A(n16287), .B(n15323), .ZN(
        n15080) );
  AOI211_X1 U18261 ( .C1(n19227), .C2(n19019), .A(n15081), .B(n15080), .ZN(
        n15082) );
  OAI21_X1 U18262 ( .B1(n15330), .B2(n15083), .A(n15082), .ZN(P2_U2998) );
  NAND2_X1 U18263 ( .A1(n15085), .A2(n15084), .ZN(n15087) );
  XOR2_X1 U18264 ( .A(n15087), .B(n15086), .Z(n15353) );
  INV_X1 U18265 ( .A(n15362), .ZN(n15089) );
  INV_X1 U18266 ( .A(n15334), .ZN(n15088) );
  AOI21_X1 U18267 ( .B1(n15322), .B2(n15089), .A(n15088), .ZN(n15351) );
  AOI22_X1 U18268 ( .A1(n19215), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19111), .ZN(n15091) );
  NAND2_X1 U18269 ( .A1(n16295), .A2(n19031), .ZN(n15090) );
  OAI211_X1 U18270 ( .C1(n15343), .C2(n15115), .A(n15091), .B(n15090), .ZN(
        n15092) );
  AOI21_X1 U18271 ( .B1(n15351), .B2(n19216), .A(n15092), .ZN(n15093) );
  OAI21_X1 U18272 ( .B1(n15353), .B2(n19218), .A(n15093), .ZN(P2_U2999) );
  NAND2_X1 U18273 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15360), .ZN(
        n16243) );
  OAI21_X1 U18274 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15360), .A(
        n16243), .ZN(n16327) );
  OAI21_X1 U18275 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n16324) );
  INV_X1 U18276 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19755) );
  OAI22_X1 U18277 ( .A1(n19755), .A2(n19089), .B1(n19224), .B2(n19055), .ZN(
        n15100) );
  INV_X1 U18278 ( .A(n19057), .ZN(n15098) );
  OAI22_X1 U18279 ( .A1(n15098), .A2(n15115), .B1(n16305), .B2(n15097), .ZN(
        n15099) );
  AOI211_X1 U18280 ( .C1(n16324), .C2(n16302), .A(n15100), .B(n15099), .ZN(
        n15101) );
  OAI21_X1 U18281 ( .B1(n16327), .B2(n16287), .A(n15101), .ZN(P2_U3002) );
  INV_X1 U18282 ( .A(n16256), .ZN(n15102) );
  OAI21_X1 U18283 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15385), .A(
        n15102), .ZN(n15384) );
  NAND2_X1 U18284 ( .A1(n15103), .A2(n15394), .ZN(n15108) );
  INV_X1 U18285 ( .A(n15104), .ZN(n15106) );
  NAND2_X1 U18286 ( .A1(n15106), .A2(n15105), .ZN(n15107) );
  XNOR2_X1 U18287 ( .A(n15108), .B(n15107), .ZN(n15382) );
  OAI22_X1 U18288 ( .A1(n12675), .A2(n19089), .B1(n19224), .B2(n19080), .ZN(
        n15111) );
  OAI22_X1 U18289 ( .A1(n15109), .A2(n15115), .B1(n16305), .B2(n10120), .ZN(
        n15110) );
  AOI211_X1 U18290 ( .C1(n15382), .C2(n16302), .A(n15111), .B(n15110), .ZN(
        n15112) );
  OAI21_X1 U18291 ( .B1(n15384), .B2(n16287), .A(n15112), .ZN(P2_U3004) );
  XNOR2_X1 U18292 ( .A(n15114), .B(n15113), .ZN(n15427) );
  INV_X1 U18293 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19746) );
  OAI22_X1 U18294 ( .A1(n19746), .A2(n19089), .B1(n19224), .B2(n19118), .ZN(
        n15117) );
  NOR2_X1 U18295 ( .A1(n19113), .A2(n15115), .ZN(n15116) );
  AOI211_X1 U18296 ( .C1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n19215), .A(
        n15117), .B(n15116), .ZN(n15121) );
  XNOR2_X1 U18297 ( .A(n15119), .B(n15118), .ZN(n15424) );
  NAND2_X1 U18298 ( .A1(n15424), .A2(n19216), .ZN(n15120) );
  OAI211_X1 U18299 ( .C1(n15427), .C2(n19218), .A(n15121), .B(n15120), .ZN(
        P2_U3010) );
  INV_X1 U18300 ( .A(n15122), .ZN(n15126) );
  NOR2_X1 U18301 ( .A1(n15123), .A2(n15182), .ZN(n15137) );
  INV_X1 U18302 ( .A(n15137), .ZN(n15145) );
  NAND3_X1 U18303 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15197) );
  NOR2_X1 U18304 ( .A1(n16345), .A2(n15416), .ZN(n15411) );
  INV_X1 U18305 ( .A(n15411), .ZN(n15131) );
  INV_X1 U18306 ( .A(n16362), .ZN(n15128) );
  INV_X1 U18307 ( .A(n15421), .ZN(n16363) );
  NAND3_X1 U18308 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15128), .A3(
        n16363), .ZN(n16346) );
  NOR2_X1 U18309 ( .A1(n15131), .A2(n16346), .ZN(n15398) );
  INV_X1 U18310 ( .A(n15398), .ZN(n15364) );
  INV_X1 U18311 ( .A(n15124), .ZN(n15133) );
  NOR2_X1 U18312 ( .A1(n15364), .A2(n15133), .ZN(n15257) );
  NAND3_X1 U18313 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n15257), .ZN(n15227) );
  NOR2_X1 U18314 ( .A1(n15197), .A2(n15227), .ZN(n15183) );
  INV_X1 U18315 ( .A(n15183), .ZN(n15170) );
  OAI211_X1 U18316 ( .C1(n19127), .C2(n16319), .A(n15126), .B(n10227), .ZN(
        n15127) );
  INV_X1 U18317 ( .A(n15127), .ZN(n15139) );
  INV_X1 U18318 ( .A(n16376), .ZN(n15363) );
  NAND2_X1 U18319 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15128), .ZN(
        n15129) );
  AND2_X1 U18320 ( .A1(n16376), .A2(n15129), .ZN(n15130) );
  NOR2_X1 U18321 ( .A1(n16355), .A2(n15130), .ZN(n16344) );
  NAND2_X1 U18322 ( .A1(n16376), .A2(n15131), .ZN(n15132) );
  NAND2_X1 U18323 ( .A1(n16344), .A2(n15132), .ZN(n15392) );
  AND2_X1 U18324 ( .A1(n16376), .A2(n15133), .ZN(n15134) );
  OR2_X1 U18325 ( .A1(n15392), .A2(n15134), .ZN(n15238) );
  NAND2_X1 U18326 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U18327 ( .A1(n15238), .A2(n15239), .ZN(n15196) );
  INV_X1 U18328 ( .A(n15197), .ZN(n15135) );
  NAND2_X1 U18329 ( .A1(n15196), .A2(n15135), .ZN(n15136) );
  NAND2_X1 U18330 ( .A1(n16344), .A2(n15363), .ZN(n15194) );
  NAND2_X1 U18331 ( .A1(n15136), .A2(n15194), .ZN(n15179) );
  OAI211_X1 U18332 ( .C1(n15363), .C2(n15137), .A(n15179), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15146) );
  NAND3_X1 U18333 ( .A1(n15146), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15194), .ZN(n15138) );
  OAI211_X1 U18334 ( .C1(n15140), .C2(n16309), .A(n15139), .B(n15138), .ZN(
        n15141) );
  AOI21_X1 U18335 ( .B1(n15142), .B2(n16358), .A(n15141), .ZN(n15143) );
  OAI21_X1 U18336 ( .B1(n15144), .B2(n16373), .A(n15143), .ZN(P2_U3015) );
  NOR2_X1 U18337 ( .A1(n15145), .A2(n15170), .ZN(n15147) );
  OAI21_X1 U18338 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15147), .A(
        n15146), .ZN(n15149) );
  OAI211_X1 U18339 ( .C1(n16187), .C2(n16319), .A(n15149), .B(n15148), .ZN(
        n15152) );
  NOR2_X1 U18340 ( .A1(n15150), .A2(n16383), .ZN(n15151) );
  OAI21_X1 U18341 ( .B1(n15154), .B2(n16373), .A(n15153), .ZN(P2_U3016) );
  INV_X1 U18342 ( .A(n16215), .ZN(n15159) );
  INV_X1 U18343 ( .A(n15155), .ZN(n15158) );
  OAI21_X1 U18344 ( .B1(n15182), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15156) );
  OAI211_X1 U18345 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15156), .B(n15183), .ZN(
        n15157) );
  OAI211_X1 U18346 ( .C1(n16319), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15160) );
  INV_X1 U18347 ( .A(n15160), .ZN(n15163) );
  NAND2_X1 U18348 ( .A1(n15182), .A2(n15183), .ZN(n15161) );
  NAND2_X1 U18349 ( .A1(n15179), .A2(n15161), .ZN(n15168) );
  NAND2_X1 U18350 ( .A1(n15168), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15162) );
  OAI211_X1 U18351 ( .C1(n16212), .C2(n16309), .A(n15163), .B(n15162), .ZN(
        n15164) );
  AOI21_X1 U18352 ( .B1(n15165), .B2(n16358), .A(n15164), .ZN(n15166) );
  OAI21_X1 U18353 ( .B1(n15167), .B2(n16373), .A(n15166), .ZN(P2_U3017) );
  NAND2_X1 U18354 ( .A1(n15168), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15174) );
  INV_X1 U18355 ( .A(n15169), .ZN(n16219) );
  NOR3_X1 U18356 ( .A1(n15182), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15170), .ZN(n15171) );
  AOI211_X1 U18357 ( .C1(n16371), .C2(n16219), .A(n15172), .B(n15171), .ZN(
        n15173) );
  OAI211_X1 U18358 ( .C1(n16218), .C2(n16309), .A(n15174), .B(n15173), .ZN(
        n15175) );
  AOI21_X1 U18359 ( .B1(n15176), .B2(n16358), .A(n15175), .ZN(n15177) );
  OAI21_X1 U18360 ( .B1(n15178), .B2(n16373), .A(n15177), .ZN(P2_U3018) );
  INV_X1 U18361 ( .A(n15179), .ZN(n15191) );
  INV_X1 U18362 ( .A(n15180), .ZN(n15187) );
  AOI21_X1 U18363 ( .B1(n15183), .B2(n15182), .A(n15181), .ZN(n15186) );
  NAND2_X1 U18364 ( .A1(n16371), .A2(n15184), .ZN(n15185) );
  OAI211_X1 U18365 ( .C1(n15187), .C2(n16309), .A(n15186), .B(n15185), .ZN(
        n15190) );
  NOR2_X1 U18366 ( .A1(n15188), .A2(n16383), .ZN(n15189) );
  OAI21_X1 U18367 ( .B1(n15193), .B2(n16373), .A(n15192), .ZN(P2_U3019) );
  INV_X1 U18368 ( .A(n15194), .ZN(n15195) );
  OR2_X1 U18369 ( .A1(n15196), .A2(n15195), .ZN(n15226) );
  INV_X1 U18370 ( .A(n15227), .ZN(n15198) );
  NAND2_X1 U18371 ( .A1(n15197), .A2(n15198), .ZN(n15201) );
  NAND3_X1 U18372 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n15198), .ZN(n15199) );
  AOI22_X1 U18373 ( .A1(n15226), .A2(n15201), .B1(n15200), .B2(n15199), .ZN(
        n15208) );
  INV_X1 U18374 ( .A(n15202), .ZN(n15203) );
  NAND2_X1 U18375 ( .A1(n15203), .A2(n16369), .ZN(n15205) );
  OAI211_X1 U18376 ( .C1(n16319), .C2(n15206), .A(n15205), .B(n15204), .ZN(
        n15207) );
  AOI211_X1 U18377 ( .C1(n15209), .C2(n16358), .A(n15208), .B(n15207), .ZN(
        n15210) );
  OAI21_X1 U18378 ( .B1(n15211), .B2(n16373), .A(n15210), .ZN(P2_U3020) );
  INV_X1 U18379 ( .A(n15212), .ZN(n15219) );
  XNOR2_X1 U18380 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15213) );
  NOR2_X1 U18381 ( .A1(n15213), .A2(n15227), .ZN(n15214) );
  NOR2_X1 U18382 ( .A1(n15215), .A2(n15214), .ZN(n15216) );
  OAI21_X1 U18383 ( .B1(n16319), .B2(n15217), .A(n15216), .ZN(n15218) );
  AOI21_X1 U18384 ( .B1(n15219), .B2(n16369), .A(n15218), .ZN(n15220) );
  OAI21_X1 U18385 ( .B1(n15226), .B2(n20824), .A(n15220), .ZN(n15221) );
  AOI21_X1 U18386 ( .B1(n15222), .B2(n16358), .A(n15221), .ZN(n15223) );
  OAI21_X1 U18387 ( .B1(n15224), .B2(n16373), .A(n15223), .ZN(P2_U3021) );
  NOR2_X1 U18388 ( .A1(n15226), .A2(n15225), .ZN(n15234) );
  NOR2_X1 U18389 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15227), .ZN(
        n15230) );
  NOR2_X1 U18390 ( .A1(n16319), .A2(n15228), .ZN(n15229) );
  AOI211_X1 U18391 ( .C1(n19111), .C2(P2_REIP_REG_24__SCAN_IN), .A(n15230), 
        .B(n15229), .ZN(n15231) );
  OAI21_X1 U18392 ( .B1(n15232), .B2(n16309), .A(n15231), .ZN(n15233) );
  AOI211_X1 U18393 ( .C1(n15235), .C2(n16358), .A(n15234), .B(n15233), .ZN(
        n15236) );
  OAI21_X1 U18394 ( .B1(n15237), .B2(n16373), .A(n15236), .ZN(P2_U3022) );
  INV_X1 U18395 ( .A(n15238), .ZN(n15254) );
  OAI211_X1 U18396 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15257), .B(n15239), .ZN(
        n15244) );
  NOR2_X1 U18397 ( .A1(n16319), .A2(n16231), .ZN(n15240) );
  AOI211_X1 U18398 ( .C1(n15242), .C2(n16369), .A(n15241), .B(n15240), .ZN(
        n15243) );
  OAI211_X1 U18399 ( .C1(n15254), .C2(n15245), .A(n15244), .B(n15243), .ZN(
        n15246) );
  AOI21_X1 U18400 ( .B1(n15247), .B2(n16358), .A(n15246), .ZN(n15248) );
  OAI21_X1 U18401 ( .B1(n15249), .B2(n16373), .A(n15248), .ZN(P2_U3023) );
  NOR2_X1 U18402 ( .A1(n19772), .A2(n11795), .ZN(n15252) );
  NOR2_X1 U18403 ( .A1(n15250), .A2(n16309), .ZN(n15251) );
  AOI211_X1 U18404 ( .C1(n16371), .C2(n15854), .A(n15252), .B(n15251), .ZN(
        n15253) );
  OAI21_X1 U18405 ( .B1(n15254), .B2(n15256), .A(n15253), .ZN(n15255) );
  AOI21_X1 U18406 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n15261) );
  NAND3_X1 U18407 ( .A1(n15259), .A2(n16358), .A3(n15258), .ZN(n15260) );
  OAI211_X1 U18408 ( .C1(n15262), .C2(n16373), .A(n15261), .B(n15260), .ZN(
        P2_U3024) );
  INV_X1 U18409 ( .A(n15263), .ZN(n15274) );
  NOR3_X1 U18410 ( .A1(n15364), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15264), .ZN(n15273) );
  AOI21_X1 U18411 ( .B1(n15264), .B2(n16376), .A(n15392), .ZN(n15271) );
  NOR2_X1 U18412 ( .A1(n16319), .A2(n15265), .ZN(n15266) );
  AOI211_X1 U18413 ( .C1(n15268), .C2(n16369), .A(n15267), .B(n15266), .ZN(
        n15269) );
  OAI21_X1 U18414 ( .B1(n15271), .B2(n15270), .A(n15269), .ZN(n15272) );
  AOI211_X1 U18415 ( .C1(n15274), .C2(n16358), .A(n15273), .B(n15272), .ZN(
        n15275) );
  OAI21_X1 U18416 ( .B1(n15276), .B2(n16373), .A(n15275), .ZN(P2_U3025) );
  NAND2_X1 U18417 ( .A1(n15398), .A2(n15318), .ZN(n15349) );
  NAND3_X1 U18418 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15277) );
  NOR2_X1 U18419 ( .A1(n15349), .A2(n15277), .ZN(n15305) );
  NAND3_X1 U18420 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15298), .ZN(n15297) );
  INV_X1 U18421 ( .A(n15278), .ZN(n15279) );
  AND2_X1 U18422 ( .A1(n16376), .A2(n15279), .ZN(n15280) );
  NOR2_X1 U18423 ( .A1(n15392), .A2(n15280), .ZN(n15299) );
  AOI21_X1 U18424 ( .B1(n15297), .B2(n15299), .A(n15281), .ZN(n15288) );
  NAND4_X1 U18425 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n15281), .ZN(n15285) );
  AOI21_X1 U18426 ( .B1(n15283), .B2(n16369), .A(n15282), .ZN(n15284) );
  OAI211_X1 U18427 ( .C1(n16319), .C2(n15286), .A(n15285), .B(n15284), .ZN(
        n15287) );
  AOI211_X1 U18428 ( .C1(n15289), .C2(n16358), .A(n15288), .B(n15287), .ZN(
        n15290) );
  OAI21_X1 U18429 ( .B1(n15291), .B2(n16373), .A(n15290), .ZN(P2_U3026) );
  INV_X1 U18430 ( .A(n15292), .ZN(n15301) );
  OAI21_X1 U18431 ( .B1(n15294), .B2(n16309), .A(n15293), .ZN(n15295) );
  AOI21_X1 U18432 ( .B1(n16371), .B2(n18985), .A(n15295), .ZN(n15296) );
  OAI211_X1 U18433 ( .C1(n15299), .C2(n15298), .A(n15297), .B(n15296), .ZN(
        n15300) );
  AOI21_X1 U18434 ( .B1(n15301), .B2(n16358), .A(n15300), .ZN(n15302) );
  OAI21_X1 U18435 ( .B1(n15303), .B2(n16373), .A(n15302), .ZN(P2_U3027) );
  AOI21_X1 U18436 ( .B1(n16376), .B2(n15304), .A(n15392), .ZN(n15311) );
  NAND2_X1 U18437 ( .A1(n15305), .A2(n15310), .ZN(n15309) );
  NOR2_X1 U18438 ( .A1(n16319), .A2(n19000), .ZN(n15306) );
  AOI211_X1 U18439 ( .C1(n18996), .C2(n16369), .A(n15307), .B(n15306), .ZN(
        n15308) );
  OAI211_X1 U18440 ( .C1(n15311), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15312) );
  AOI21_X1 U18441 ( .B1(n15313), .B2(n16358), .A(n15312), .ZN(n15314) );
  OAI21_X1 U18442 ( .B1(n15315), .B2(n16373), .A(n15314), .ZN(P2_U3028) );
  INV_X1 U18443 ( .A(n15316), .ZN(n15321) );
  INV_X1 U18444 ( .A(n15392), .ZN(n15317) );
  OAI21_X1 U18445 ( .B1(n15363), .B2(n15318), .A(n15317), .ZN(n15346) );
  AOI21_X1 U18446 ( .B1(n16383), .B2(n15319), .A(n15323), .ZN(n15320) );
  NOR2_X1 U18447 ( .A1(n15349), .A2(n15322), .ZN(n15332) );
  AOI22_X1 U18448 ( .A1(n15323), .A2(n16358), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15332), .ZN(n15327) );
  OAI21_X1 U18449 ( .B1(n16309), .B2(n19008), .A(n15324), .ZN(n15325) );
  AOI21_X1 U18450 ( .B1(n16371), .B2(n19009), .A(n15325), .ZN(n15326) );
  OAI21_X1 U18451 ( .B1(n15327), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15326), .ZN(n15328) );
  NAND3_X1 U18452 ( .A1(n10086), .A2(n16360), .A3(n15331), .ZN(n15340) );
  INV_X1 U18453 ( .A(n15332), .ZN(n15333) );
  OAI21_X1 U18454 ( .B1(n15334), .B2(n16383), .A(n15333), .ZN(n15338) );
  AOI21_X1 U18455 ( .B1(n16369), .B2(n19019), .A(n15335), .ZN(n15336) );
  OAI21_X1 U18456 ( .B1(n16319), .B2(n19020), .A(n15336), .ZN(n15337) );
  AOI21_X1 U18457 ( .B1(n15338), .B2(n15341), .A(n15337), .ZN(n15339) );
  OAI211_X1 U18458 ( .C1(n15342), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        P2_U3030) );
  INV_X1 U18459 ( .A(n15343), .ZN(n19033) );
  INV_X1 U18460 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19759) );
  NOR2_X1 U18461 ( .A1(n19759), .A2(n11795), .ZN(n15345) );
  NOR2_X1 U18462 ( .A1(n16319), .A2(n19037), .ZN(n15344) );
  AOI211_X1 U18463 ( .C1(n16369), .C2(n19033), .A(n15345), .B(n15344), .ZN(
        n15348) );
  NAND2_X1 U18464 ( .A1(n15346), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15347) );
  OAI211_X1 U18465 ( .C1(n15349), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15348), .B(n15347), .ZN(n15350) );
  AOI21_X1 U18466 ( .B1(n15351), .B2(n16358), .A(n15350), .ZN(n15352) );
  OAI21_X1 U18467 ( .B1(n15353), .B2(n16373), .A(n15352), .ZN(P2_U3031) );
  INV_X1 U18468 ( .A(n15355), .ZN(n15358) );
  AND2_X1 U18469 ( .A1(n15355), .A2(n15354), .ZN(n15356) );
  OAI22_X1 U18470 ( .A1(n15359), .A2(n15358), .B1(n15357), .B2(n15356), .ZN(
        n16239) );
  NOR2_X1 U18471 ( .A1(n16242), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15361) );
  AOI21_X1 U18472 ( .B1(n15397), .B2(n16376), .A(n15392), .ZN(n16337) );
  OAI21_X1 U18473 ( .B1(n15363), .B2(n16331), .A(n16337), .ZN(n16321) );
  NOR2_X1 U18474 ( .A1(n12920), .A2(n11795), .ZN(n15368) );
  INV_X1 U18475 ( .A(n15366), .ZN(n16314) );
  NOR2_X1 U18476 ( .A1(n15397), .A2(n15364), .ZN(n16333) );
  NAND2_X1 U18477 ( .A1(n16331), .A2(n16333), .ZN(n16313) );
  AOI221_X1 U18478 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15366), 
        .C1(n15365), .C2(n16314), .A(n16313), .ZN(n15367) );
  AOI211_X1 U18479 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16321), .A(
        n15368), .B(n15367), .ZN(n15371) );
  INV_X1 U18480 ( .A(n19049), .ZN(n15369) );
  AOI22_X1 U18481 ( .A1(n16371), .A2(n15369), .B1(n16369), .B2(n19045), .ZN(
        n15370) );
  OAI211_X1 U18482 ( .C1(n16238), .C2(n16383), .A(n15371), .B(n15370), .ZN(
        n15372) );
  INV_X1 U18483 ( .A(n15372), .ZN(n15373) );
  OAI21_X1 U18484 ( .B1(n16239), .B2(n16373), .A(n15373), .ZN(P2_U3032) );
  NOR2_X1 U18485 ( .A1(n16337), .A2(n15374), .ZN(n15381) );
  NAND2_X1 U18486 ( .A1(n19082), .A2(n16369), .ZN(n15379) );
  NOR2_X1 U18487 ( .A1(n12675), .A2(n11795), .ZN(n15377) );
  INV_X1 U18488 ( .A(n16333), .ZN(n15375) );
  NOR2_X1 U18489 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15375), .ZN(
        n15376) );
  NOR2_X1 U18490 ( .A1(n15377), .A2(n15376), .ZN(n15378) );
  OAI211_X1 U18491 ( .C1(n16319), .C2(n19086), .A(n15379), .B(n15378), .ZN(
        n15380) );
  AOI211_X1 U18492 ( .C1(n15382), .C2(n16360), .A(n15381), .B(n15380), .ZN(
        n15383) );
  OAI21_X1 U18493 ( .B1(n15384), .B2(n16383), .A(n15383), .ZN(P2_U3036) );
  AOI21_X1 U18494 ( .B1(n15386), .B2(n15397), .A(n15385), .ZN(n16266) );
  NAND2_X1 U18495 ( .A1(n16266), .A2(n16358), .ZN(n15402) );
  INV_X1 U18496 ( .A(n15387), .ZN(n16264) );
  NAND2_X1 U18497 ( .A1(n16369), .A2(n16264), .ZN(n15389) );
  NAND2_X1 U18498 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19111), .ZN(n15388) );
  OAI211_X1 U18499 ( .C1(n15390), .C2(n16319), .A(n15389), .B(n15388), .ZN(
        n15391) );
  AOI21_X1 U18500 ( .B1(n15392), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15391), .ZN(n15401) );
  NOR2_X1 U18501 ( .A1(n15395), .A2(n14801), .ZN(n15396) );
  XNOR2_X1 U18502 ( .A(n15393), .B(n15396), .ZN(n16265) );
  NAND2_X1 U18503 ( .A1(n16265), .A2(n16360), .ZN(n15400) );
  NAND2_X1 U18504 ( .A1(n15398), .A2(n15397), .ZN(n15399) );
  NAND4_X1 U18505 ( .A1(n15402), .A2(n15401), .A3(n15400), .A4(n15399), .ZN(
        P2_U3037) );
  XNOR2_X1 U18506 ( .A(n15404), .B(n15403), .ZN(n16271) );
  NAND2_X1 U18507 ( .A1(n15405), .A2(n16276), .ZN(n15406) );
  NAND2_X1 U18508 ( .A1(n15406), .A2(n16277), .ZN(n15410) );
  AND2_X1 U18509 ( .A1(n15408), .A2(n15407), .ZN(n15409) );
  XNOR2_X1 U18510 ( .A(n15410), .B(n15409), .ZN(n16270) );
  INV_X1 U18511 ( .A(n16270), .ZN(n15419) );
  AOI211_X1 U18512 ( .C1(n16345), .C2(n15416), .A(n15411), .B(n16346), .ZN(
        n15418) );
  INV_X1 U18513 ( .A(n15412), .ZN(n19097) );
  INV_X1 U18514 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n15413) );
  OAI22_X1 U18515 ( .A1(n16319), .A2(n19102), .B1(n19089), .B2(n15413), .ZN(
        n15414) );
  AOI21_X1 U18516 ( .B1(n16369), .B2(n19097), .A(n15414), .ZN(n15415) );
  OAI21_X1 U18517 ( .B1(n16344), .B2(n15416), .A(n15415), .ZN(n15417) );
  AOI211_X1 U18518 ( .C1(n15419), .C2(n16360), .A(n15418), .B(n15417), .ZN(
        n15420) );
  OAI21_X1 U18519 ( .B1(n16271), .B2(n16383), .A(n15420), .ZN(P2_U3038) );
  OAI22_X1 U18520 ( .A1(n11795), .A2(n19746), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15421), .ZN(n15423) );
  OAI22_X1 U18521 ( .A1(n19106), .A2(n16319), .B1(n16309), .B2(n19113), .ZN(
        n15422) );
  AOI211_X1 U18522 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n16355), .A(
        n15423), .B(n15422), .ZN(n15426) );
  NAND2_X1 U18523 ( .A1(n15424), .A2(n16358), .ZN(n15425) );
  OAI211_X1 U18524 ( .C1(n15427), .C2(n16373), .A(n15426), .B(n15425), .ZN(
        P2_U3042) );
  INV_X1 U18525 ( .A(n16374), .ZN(n15432) );
  OAI22_X1 U18526 ( .A1(n16309), .A2(n15429), .B1(n15428), .B2(n16319), .ZN(
        n15430) );
  AOI211_X1 U18527 ( .C1(n15432), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15431), .B(n15430), .ZN(n15438) );
  AOI22_X1 U18528 ( .A1(n16360), .A2(n15434), .B1(n16358), .B2(n15433), .ZN(
        n15437) );
  OAI211_X1 U18529 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16376), .B(n15435), .ZN(n15436) );
  NAND3_X1 U18530 ( .A1(n15438), .A2(n15437), .A3(n15436), .ZN(P2_U3045) );
  OAI221_X1 U18531 ( .B1(n19094), .B2(n15439), .C1(n9591), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(P2_STATE2_REG_1__SCAN_IN), .ZN(
        n15470) );
  INV_X1 U18532 ( .A(n11766), .ZN(n15441) );
  NAND2_X1 U18533 ( .A1(n15441), .A2(n15440), .ZN(n15452) );
  MUX2_X1 U18534 ( .A(n15452), .B(n12307), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15442) );
  AOI21_X1 U18535 ( .B1(n16368), .B2(n15467), .A(n15442), .ZN(n16384) );
  OAI21_X1 U18536 ( .B1(n16384), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13505), 
        .ZN(n15444) );
  AOI22_X1 U18537 ( .A1(n15470), .A2(n15444), .B1(n15443), .B2(n16428), .ZN(
        n15446) );
  NAND2_X1 U18538 ( .A1(n15474), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15445) );
  OAI21_X1 U18539 ( .B1(n15446), .B2(n15474), .A(n15445), .ZN(P2_U3601) );
  AOI21_X1 U18540 ( .B1(n19094), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15447), .ZN(n15469) );
  INV_X1 U18541 ( .A(n15469), .ZN(n15456) );
  NAND2_X1 U18542 ( .A1(n15448), .A2(n15467), .ZN(n15454) );
  XNOR2_X1 U18543 ( .A(n15449), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15451) );
  AOI22_X1 U18544 ( .A1(n15452), .A2(n15451), .B1(n15450), .B2(n12307), .ZN(
        n15453) );
  NAND2_X1 U18545 ( .A1(n15454), .A2(n15453), .ZN(n16387) );
  AOI22_X1 U18546 ( .A1(n19823), .A2(n16428), .B1(n18952), .B2(n16387), .ZN(
        n15455) );
  OAI21_X1 U18547 ( .B1(n15470), .B2(n15456), .A(n15455), .ZN(n15457) );
  MUX2_X1 U18548 ( .A(n15457), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15474), .Z(P2_U3600) );
  AOI21_X1 U18549 ( .B1(n15460), .B2(n15459), .A(n15458), .ZN(n15466) );
  OAI22_X1 U18550 ( .A1(n15464), .A2(n15463), .B1(n15461), .B2(n15462), .ZN(
        n15465) );
  AOI211_X1 U18551 ( .C1(n9592), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        n16391) );
  INV_X1 U18552 ( .A(n16391), .ZN(n16412) );
  AOI22_X1 U18553 ( .A1(n19812), .A2(n16428), .B1(n18952), .B2(n16412), .ZN(
        n15468) );
  OAI21_X1 U18554 ( .B1(n15470), .B2(n15469), .A(n15468), .ZN(n15471) );
  MUX2_X1 U18555 ( .A(n15471), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15474), .Z(P2_U3599) );
  NOR4_X1 U18556 ( .A1(n15473), .A2(n15472), .A3(n19801), .A4(n15526), .ZN(
        n15475) );
  MUX2_X1 U18557 ( .A(n15475), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n15474), .Z(P2_U3595) );
  NOR3_X1 U18558 ( .A1(n19707), .A2(n19252), .A3(n19552), .ZN(n15478) );
  NOR2_X1 U18559 ( .A1(n19552), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19428) );
  NOR2_X1 U18560 ( .A1(n15478), .A2(n19428), .ZN(n15482) );
  NOR2_X1 U18561 ( .A1(n15479), .A2(n19809), .ZN(n19702) );
  NAND2_X1 U18562 ( .A1(n19809), .A2(n19817), .ZN(n19253) );
  OR2_X1 U18563 ( .A1(n19253), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19256) );
  NOR2_X1 U18564 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19256), .ZN(
        n19246) );
  NOR2_X1 U18565 ( .A1(n19702), .A2(n19246), .ZN(n15485) );
  INV_X1 U18566 ( .A(n15480), .ZN(n15483) );
  OAI21_X1 U18567 ( .B1(n15483), .B2(n19246), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15481) );
  INV_X1 U18568 ( .A(n15482), .ZN(n15486) );
  AOI211_X1 U18569 ( .C1(n15483), .C2(n12070), .A(n19246), .B(n19799), .ZN(
        n15484) );
  AOI22_X1 U18570 ( .A1(n19662), .A2(n19252), .B1(n19652), .B2(n19246), .ZN(
        n15488) );
  NAND2_X1 U18571 ( .A1(n19605), .A2(n19707), .ZN(n15487) );
  OAI211_X1 U18572 ( .C1(n19251), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        n15490) );
  AOI21_X1 U18573 ( .B1(n19653), .B2(n19247), .A(n15490), .ZN(n15491) );
  INV_X1 U18574 ( .A(n15491), .ZN(P2_U3048) );
  NOR2_X2 U18575 ( .A1(n15492), .A2(n19463), .ZN(n19697) );
  INV_X1 U18576 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16533) );
  INV_X1 U18577 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18305) );
  OAI22_X2 U18578 ( .A1(n16533), .A2(n15564), .B1(n18305), .B2(n15563), .ZN(
        n19698) );
  AND2_X1 U18579 ( .A1(n15494), .A2(n15558), .ZN(n19696) );
  AOI22_X1 U18580 ( .A1(n19698), .A2(n19252), .B1(n19246), .B2(n19696), .ZN(
        n15496) );
  INV_X1 U18581 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18307) );
  INV_X1 U18582 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16519) );
  NAND2_X1 U18583 ( .A1(n19635), .A2(n19707), .ZN(n15495) );
  OAI211_X1 U18584 ( .C1(n19251), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15498) );
  AOI21_X1 U18585 ( .B1(n19697), .B2(n19247), .A(n15498), .ZN(n15499) );
  INV_X1 U18586 ( .A(n15499), .ZN(P2_U3054) );
  NOR2_X1 U18587 ( .A1(n19494), .A2(n19253), .ZN(n19296) );
  AOI21_X1 U18588 ( .B1(n15503), .B2(n12070), .A(n19296), .ZN(n15501) );
  NOR2_X1 U18589 ( .A1(n19497), .A2(n19253), .ZN(n15504) );
  AOI221_X1 U18590 ( .B1(n19299), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19298), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n15504), .ZN(n15500) );
  MUX2_X1 U18591 ( .A(n15501), .B(n15500), .S(n19799), .Z(n15502) );
  INV_X1 U18592 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18593 ( .A1(n19299), .A2(n19662), .B1(n19298), .B2(n19605), .ZN(
        n15508) );
  OAI21_X1 U18594 ( .B1(n15503), .B2(n19296), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15506) );
  INV_X1 U18595 ( .A(n15504), .ZN(n15505) );
  NAND2_X1 U18596 ( .A1(n15506), .A2(n15505), .ZN(n19297) );
  AOI22_X1 U18597 ( .A1(n19297), .A2(n19653), .B1(n19652), .B2(n19296), .ZN(
        n15507) );
  OAI211_X1 U18598 ( .C1(n19303), .C2(n15509), .A(n15508), .B(n15507), .ZN(
        P2_U3064) );
  INV_X1 U18599 ( .A(n19253), .ZN(n15510) );
  NAND2_X1 U18600 ( .A1(n15511), .A2(n15510), .ZN(n15560) );
  INV_X1 U18601 ( .A(n15516), .ZN(n15512) );
  OAI21_X1 U18602 ( .B1(n15512), .B2(n16425), .A(n12070), .ZN(n15515) );
  OAI21_X1 U18603 ( .B1(n19399), .B2(n19800), .A(n19799), .ZN(n15517) );
  NOR2_X1 U18604 ( .A1(n19827), .A2(n19253), .ZN(n15513) );
  NOR2_X1 U18605 ( .A1(n15517), .A2(n15513), .ZN(n15514) );
  AOI21_X1 U18606 ( .B1(n15516), .B2(n15560), .A(n16425), .ZN(n15519) );
  NOR3_X1 U18607 ( .A1(n19827), .A2(n19253), .A3(n15517), .ZN(n15518) );
  INV_X1 U18608 ( .A(n19653), .ZN(n19614) );
  INV_X1 U18609 ( .A(n19652), .ZN(n15520) );
  OAI22_X1 U18610 ( .A1(n15561), .A2(n19614), .B1(n15520), .B2(n15560), .ZN(
        n15521) );
  AOI21_X1 U18611 ( .B1(n19605), .B2(n19299), .A(n15521), .ZN(n15523) );
  NAND2_X1 U18612 ( .A1(n19662), .A2(n19330), .ZN(n15522) );
  OAI211_X1 U18613 ( .C1(n15568), .C2(n15524), .A(n15523), .B(n15522), .ZN(
        P2_U3072) );
  INV_X1 U18614 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18273) );
  INV_X1 U18615 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16527) );
  NOR2_X2 U18616 ( .A1(n15525), .A2(n19463), .ZN(n19667) );
  INV_X1 U18617 ( .A(n19667), .ZN(n19618) );
  NAND2_X1 U18618 ( .A1(n15526), .A2(n15558), .ZN(n19230) );
  OAI22_X1 U18619 ( .A1(n15561), .A2(n19618), .B1(n15560), .B2(n19230), .ZN(
        n15527) );
  AOI21_X1 U18620 ( .B1(n19615), .B2(n19299), .A(n15527), .ZN(n15529) );
  INV_X1 U18621 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16542) );
  INV_X1 U18622 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18271) );
  OAI22_X2 U18623 ( .A1(n16542), .A2(n15564), .B1(n18271), .B2(n15563), .ZN(
        n19668) );
  NAND2_X1 U18624 ( .A1(n19668), .A2(n19330), .ZN(n15528) );
  OAI211_X1 U18625 ( .C1(n15568), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        P2_U3073) );
  INV_X1 U18626 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18280) );
  NOR2_X2 U18627 ( .A1(n15531), .A2(n19463), .ZN(n19673) );
  INV_X1 U18628 ( .A(n19673), .ZN(n19622) );
  NAND2_X1 U18629 ( .A1(n11297), .A2(n15558), .ZN(n19233) );
  OAI22_X1 U18630 ( .A1(n15561), .A2(n19622), .B1(n15560), .B2(n19233), .ZN(
        n15532) );
  AOI21_X1 U18631 ( .B1(n19619), .B2(n19299), .A(n15532), .ZN(n15534) );
  INV_X1 U18632 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16540) );
  INV_X1 U18633 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18278) );
  OAI22_X2 U18634 ( .A1(n16540), .A2(n15564), .B1(n18278), .B2(n15563), .ZN(
        n19674) );
  NAND2_X1 U18635 ( .A1(n19674), .A2(n19330), .ZN(n15533) );
  OAI211_X1 U18636 ( .C1(n15568), .C2(n15535), .A(n15534), .B(n15533), .ZN(
        P2_U3074) );
  INV_X1 U18637 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16524) );
  INV_X1 U18638 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18285) );
  NOR2_X2 U18639 ( .A1(n15536), .A2(n19463), .ZN(n19679) );
  INV_X1 U18640 ( .A(n19679), .ZN(n19626) );
  NAND2_X1 U18641 ( .A1(n15537), .A2(n15558), .ZN(n19236) );
  OAI22_X1 U18642 ( .A1(n15561), .A2(n19626), .B1(n15560), .B2(n19236), .ZN(
        n15538) );
  AOI21_X1 U18643 ( .B1(n19623), .B2(n19299), .A(n15538), .ZN(n15540) );
  INV_X1 U18644 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16538) );
  INV_X1 U18645 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18288) );
  OAI22_X2 U18646 ( .A1(n16538), .A2(n15564), .B1(n18288), .B2(n15563), .ZN(
        n19680) );
  NAND2_X1 U18647 ( .A1(n19680), .A2(n19330), .ZN(n15539) );
  OAI211_X1 U18648 ( .C1(n15568), .C2(n15541), .A(n15540), .B(n15539), .ZN(
        P2_U3075) );
  INV_X1 U18649 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18292) );
  NOR2_X2 U18650 ( .A1(n15542), .A2(n19463), .ZN(n19685) );
  INV_X1 U18651 ( .A(n19685), .ZN(n19630) );
  NAND2_X1 U18652 ( .A1(n15543), .A2(n15558), .ZN(n19239) );
  OAI22_X1 U18653 ( .A1(n15561), .A2(n19630), .B1(n15560), .B2(n19239), .ZN(
        n15544) );
  AOI21_X1 U18654 ( .B1(n19627), .B2(n19299), .A(n15544), .ZN(n15546) );
  INV_X1 U18655 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18294) );
  OAI22_X2 U18656 ( .A1(n16536), .A2(n15564), .B1(n18294), .B2(n15563), .ZN(
        n19686) );
  NAND2_X1 U18657 ( .A1(n19686), .A2(n19330), .ZN(n15545) );
  OAI211_X1 U18658 ( .C1(n15568), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        P2_U3076) );
  INV_X1 U18659 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16521) );
  INV_X1 U18660 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18298) );
  NOR2_X2 U18661 ( .A1(n15548), .A2(n19463), .ZN(n19691) );
  INV_X1 U18662 ( .A(n19691), .ZN(n19634) );
  NAND2_X1 U18663 ( .A1(n11720), .A2(n15558), .ZN(n19242) );
  OAI22_X1 U18664 ( .A1(n15561), .A2(n19634), .B1(n15560), .B2(n19242), .ZN(
        n15549) );
  AOI21_X1 U18665 ( .B1(n19631), .B2(n19299), .A(n15549), .ZN(n15551) );
  INV_X1 U18666 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20774) );
  INV_X1 U18667 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18301) );
  OAI22_X2 U18668 ( .A1(n20774), .A2(n15564), .B1(n18301), .B2(n15563), .ZN(
        n19692) );
  NAND2_X1 U18669 ( .A1(n19692), .A2(n19330), .ZN(n15550) );
  OAI211_X1 U18670 ( .C1(n15568), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        P2_U3077) );
  INV_X1 U18671 ( .A(n19697), .ZN(n19638) );
  INV_X1 U18672 ( .A(n19696), .ZN(n15553) );
  OAI22_X1 U18673 ( .A1(n15561), .A2(n19638), .B1(n15553), .B2(n15560), .ZN(
        n15554) );
  AOI21_X1 U18674 ( .B1(n19635), .B2(n19299), .A(n15554), .ZN(n15556) );
  NAND2_X1 U18675 ( .A1(n19698), .A2(n19330), .ZN(n15555) );
  OAI211_X1 U18676 ( .C1(n15568), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        P2_U3078) );
  INV_X1 U18677 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15567) );
  INV_X1 U18678 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18312) );
  NAND2_X1 U18679 ( .A1(n16229), .A2(n19655), .ZN(n19646) );
  NAND2_X1 U18680 ( .A1(n9603), .A2(n15558), .ZN(n19245) );
  OAI22_X1 U18681 ( .A1(n15561), .A2(n19646), .B1(n15560), .B2(n19245), .ZN(
        n15562) );
  AOI21_X1 U18682 ( .B1(n19641), .B2(n19299), .A(n15562), .ZN(n15566) );
  INV_X1 U18683 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16531) );
  INV_X1 U18684 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18317) );
  OAI22_X2 U18685 ( .A1(n16531), .A2(n15564), .B1(n18317), .B2(n15563), .ZN(
        n19706) );
  NAND2_X1 U18686 ( .A1(n19706), .A2(n19330), .ZN(n15565) );
  OAI211_X1 U18687 ( .C1(n15568), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        P2_U3079) );
  INV_X1 U18688 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16692) );
  INV_X1 U18689 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17042) );
  INV_X1 U18690 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17004) );
  INV_X1 U18691 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17162) );
  NAND2_X1 U18692 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n17217) );
  NAND4_X1 U18693 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n15571)
         );
  INV_X1 U18694 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16940) );
  NOR3_X1 U18695 ( .A1(n16940), .A2(n17294), .A3(n17293), .ZN(n15659) );
  NAND3_X1 U18696 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n17278) );
  INV_X1 U18697 ( .A(n17278), .ZN(n15569) );
  NAND4_X1 U18698 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n15659), .A4(n15569), .ZN(n15570) );
  NOR4_X1 U18699 ( .A1(n17162), .A2(n17217), .A3(n15571), .A4(n15570), .ZN(
        n17147) );
  NAND4_X1 U18700 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n17305), .A4(n17147), .ZN(n17111) );
  NOR2_X1 U18701 ( .A1(n16766), .A2(n17111), .ZN(n17123) );
  NAND2_X1 U18702 ( .A1(n18316), .A2(n17123), .ZN(n17107) );
  NOR2_X1 U18703 ( .A1(n15572), .A2(n17107), .ZN(n17095) );
  NAND4_X1 U18704 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17095), .ZN(n17057) );
  NOR2_X1 U18705 ( .A1(n17004), .A2(n17057), .ZN(n17062) );
  NAND2_X1 U18706 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17062), .ZN(n17047) );
  NOR3_X1 U18707 ( .A1(n16692), .A2(n17042), .A3(n17047), .ZN(n17046) );
  NAND2_X1 U18708 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17046), .ZN(n17041) );
  AOI21_X1 U18709 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17300), .A(n17046), .ZN(
        n15573) );
  INV_X1 U18710 ( .A(n15573), .ZN(n15646) );
  AOI22_X1 U18711 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U18712 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U18713 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15575) );
  AOI22_X1 U18714 ( .A1(n17239), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15574) );
  NAND4_X1 U18715 ( .A1(n15577), .A2(n15576), .A3(n15575), .A4(n15574), .ZN(
        n15583) );
  AOI22_X1 U18716 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15581) );
  AOI22_X1 U18717 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U18718 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U18719 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15578) );
  NAND4_X1 U18720 ( .A1(n15581), .A2(n15580), .A3(n15579), .A4(n15578), .ZN(
        n15582) );
  NOR2_X1 U18721 ( .A1(n15583), .A2(n15582), .ZN(n15645) );
  AOI22_X1 U18722 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U18723 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U18724 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15585) );
  AOI22_X1 U18725 ( .A1(n17239), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15584) );
  NAND4_X1 U18726 ( .A1(n15587), .A2(n15586), .A3(n15585), .A4(n15584), .ZN(
        n15593) );
  AOI22_X1 U18727 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15591) );
  AOI22_X1 U18728 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15590) );
  AOI22_X1 U18729 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18730 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15588) );
  NAND4_X1 U18731 ( .A1(n15591), .A2(n15590), .A3(n15589), .A4(n15588), .ZN(
        n15592) );
  NOR2_X1 U18732 ( .A1(n15593), .A2(n15592), .ZN(n17049) );
  AOI22_X1 U18733 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U18734 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15596) );
  AOI22_X1 U18735 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U18736 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15594) );
  NAND4_X1 U18737 ( .A1(n15597), .A2(n15596), .A3(n15595), .A4(n15594), .ZN(
        n15603) );
  AOI22_X1 U18738 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U18739 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17260), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U18740 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U18741 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15598) );
  NAND4_X1 U18742 ( .A1(n15601), .A2(n15600), .A3(n15599), .A4(n15598), .ZN(
        n15602) );
  NOR2_X1 U18743 ( .A1(n15603), .A2(n15602), .ZN(n17059) );
  AOI22_X1 U18744 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18745 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15613) );
  INV_X1 U18746 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U18747 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15604) );
  OAI21_X1 U18748 ( .B1(n17241), .B2(n18270), .A(n15604), .ZN(n15611) );
  AOI22_X1 U18749 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15609) );
  AOI22_X1 U18750 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U18751 ( .A1(n17239), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U18752 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15606) );
  NAND4_X1 U18753 ( .A1(n15609), .A2(n15608), .A3(n15607), .A4(n15606), .ZN(
        n15610) );
  AOI211_X1 U18754 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n15611), .B(n15610), .ZN(n15612) );
  NAND3_X1 U18755 ( .A1(n15614), .A2(n15613), .A3(n15612), .ZN(n17066) );
  AOI22_X1 U18756 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n15780), .ZN(n15624) );
  AOI22_X1 U18757 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17020), .ZN(n15623) );
  INV_X1 U18758 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U18759 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17238), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15615) );
  OAI21_X1 U18760 ( .B1(n9642), .B2(n18320), .A(n15615), .ZN(n15621) );
  AOI22_X1 U18761 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17269), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17237), .ZN(n15619) );
  AOI22_X1 U18762 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17244), .B1(
        n17260), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18763 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17271), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17242), .ZN(n15617) );
  AOI22_X1 U18764 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17239), .ZN(n15616) );
  NAND4_X1 U18765 ( .A1(n15619), .A2(n15618), .A3(n15617), .A4(n15616), .ZN(
        n15620) );
  AOI211_X1 U18766 ( .C1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .C2(n9596), .A(
        n15621), .B(n15620), .ZN(n15622) );
  NAND3_X1 U18767 ( .A1(n15624), .A2(n15623), .A3(n15622), .ZN(n17067) );
  NAND2_X1 U18768 ( .A1(n17066), .A2(n17067), .ZN(n17065) );
  NOR2_X1 U18769 ( .A1(n17059), .A2(n17065), .ZN(n17058) );
  AOI22_X1 U18770 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U18771 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15633) );
  AOI22_X1 U18772 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U18773 ( .B1(n17241), .B2(n18284), .A(n15625), .ZN(n15631) );
  AOI22_X1 U18774 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18775 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18776 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18777 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15626) );
  NAND4_X1 U18778 ( .A1(n15629), .A2(n15628), .A3(n15627), .A4(n15626), .ZN(
        n15630) );
  AOI211_X1 U18779 ( .C1(n17238), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15631), .B(n15630), .ZN(n15632) );
  NAND3_X1 U18780 ( .A1(n15634), .A2(n15633), .A3(n15632), .ZN(n17054) );
  NAND2_X1 U18781 ( .A1(n17058), .A2(n17054), .ZN(n17053) );
  NOR2_X1 U18782 ( .A1(n17049), .A2(n17053), .ZN(n17048) );
  AOI22_X1 U18783 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15644) );
  AOI22_X1 U18784 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15643) );
  INV_X1 U18785 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U18786 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15635) );
  OAI21_X1 U18787 ( .B1(n17241), .B2(n18297), .A(n15635), .ZN(n15641) );
  AOI22_X1 U18788 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15639) );
  AOI22_X1 U18789 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15638) );
  AOI22_X1 U18790 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18791 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15636) );
  NAND4_X1 U18792 ( .A1(n15639), .A2(n15638), .A3(n15637), .A4(n15636), .ZN(
        n15640) );
  AOI211_X1 U18793 ( .C1(n17262), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15641), .B(n15640), .ZN(n15642) );
  NAND3_X1 U18794 ( .A1(n15644), .A2(n15643), .A3(n15642), .ZN(n17044) );
  NAND2_X1 U18795 ( .A1(n17048), .A2(n17044), .ZN(n17043) );
  NOR2_X1 U18796 ( .A1(n15645), .A2(n17043), .ZN(n17039) );
  AOI21_X1 U18797 ( .B1(n15645), .B2(n17043), .A(n17039), .ZN(n17324) );
  AOI22_X1 U18798 ( .A1(n17041), .A2(n15646), .B1(n17324), .B2(n17303), .ZN(
        n15647) );
  INV_X1 U18799 ( .A(n15647), .ZN(P3_U2675) );
  AOI22_X1 U18800 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17260), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18801 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15651) );
  AOI22_X1 U18802 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15650) );
  AOI22_X1 U18803 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15649) );
  NAND4_X1 U18804 ( .A1(n15652), .A2(n15651), .A3(n15650), .A4(n15649), .ZN(
        n15658) );
  AOI22_X1 U18805 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18806 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18807 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U18808 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15653) );
  NAND4_X1 U18809 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15657) );
  NOR2_X1 U18810 ( .A1(n15658), .A2(n15657), .ZN(n17402) );
  INV_X1 U18811 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U18812 ( .A1(n17305), .A2(n15659), .ZN(n17289) );
  NOR2_X1 U18813 ( .A1(n17278), .A2(n17289), .ZN(n17285) );
  NAND2_X1 U18814 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17285), .ZN(n17254) );
  NOR3_X1 U18815 ( .A1(n16863), .A2(n17217), .A3(n17254), .ZN(n17220) );
  NAND2_X1 U18816 ( .A1(n18316), .A2(n17220), .ZN(n17205) );
  NOR2_X1 U18817 ( .A1(n16851), .A2(n17205), .ZN(n15660) );
  NAND3_X1 U18818 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17220), .ZN(n17189) );
  OAI211_X1 U18819 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n15660), .A(n17189), .B(
        n17300), .ZN(n15661) );
  OAI21_X1 U18820 ( .B1(n17402), .B2(n17300), .A(n15661), .ZN(P3_U2690) );
  NAND2_X1 U18821 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18748), .ZN(n18323) );
  NOR2_X1 U18822 ( .A1(n17270), .A2(n15662), .ZN(n18253) );
  AOI221_X1 U18823 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18885), .C1(n18938), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18900), .ZN(n15663) );
  INV_X1 U18824 ( .A(n15663), .ZN(n18266) );
  INV_X1 U18825 ( .A(n15664), .ZN(n15665) );
  OAI211_X1 U18826 ( .C1(n18871), .C2(n18253), .A(n18394), .B(n15665), .ZN(
        n18260) );
  NAND2_X1 U18827 ( .A1(n18323), .A2(n18260), .ZN(n15668) );
  INV_X1 U18828 ( .A(n15668), .ZN(n15667) );
  NAND3_X1 U18829 ( .A1(n18938), .A2(n18872), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18620) );
  INV_X1 U18830 ( .A(n18260), .ZN(n18256) );
  NAND2_X1 U18831 ( .A1(n18938), .A2(n18872), .ZN(n16610) );
  NAND2_X1 U18832 ( .A1(n18884), .A2(n16610), .ZN(n18254) );
  NOR2_X1 U18833 ( .A1(n18885), .A2(n16612), .ZN(n17834) );
  INV_X1 U18834 ( .A(n17834), .ZN(n17891) );
  NOR2_X1 U18835 ( .A1(n18748), .A2(n18872), .ZN(n18261) );
  AOI21_X1 U18836 ( .B1(n18254), .B2(n17891), .A(n18261), .ZN(n15670) );
  OR3_X1 U18837 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18256), .A3(
        n15670), .ZN(n15666) );
  OAI221_X1 U18838 ( .B1(n18750), .B2(n15667), .C1(n18750), .C2(n18620), .A(
        n15666), .ZN(P3_U2864) );
  NAND2_X1 U18839 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18439) );
  INV_X1 U18840 ( .A(n18254), .ZN(n18922) );
  NOR2_X1 U18841 ( .A1(n18922), .A2(n17834), .ZN(n15669) );
  AOI221_X1 U18842 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18439), .C1(n15669), 
        .C2(n18439), .A(n15668), .ZN(n18259) );
  AOI221_X1 U18843 ( .B1(n18620), .B2(n18750), .C1(n18620), .C2(n15670), .A(
        n18256), .ZN(n15671) );
  INV_X1 U18844 ( .A(n15671), .ZN(n18257) );
  AOI22_X1 U18845 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18259), .B1(
        n18257), .B2(n18755), .ZN(P3_U2865) );
  NAND2_X1 U18846 ( .A1(n15673), .A2(n15672), .ZN(n18940) );
  NAND2_X1 U18847 ( .A1(n18729), .A2(n15675), .ZN(n18726) );
  INV_X1 U18848 ( .A(n15676), .ZN(n15679) );
  INV_X1 U18849 ( .A(n15677), .ZN(n15678) );
  NAND3_X1 U18850 ( .A1(n15679), .A2(n16445), .A3(n15678), .ZN(n15680) );
  NAND2_X1 U18851 ( .A1(n15681), .A2(n15680), .ZN(n18720) );
  NOR2_X1 U18852 ( .A1(n18274), .A2(n15682), .ZN(n15688) );
  NAND2_X1 U18853 ( .A1(n15688), .A2(n15683), .ZN(n15815) );
  INV_X1 U18854 ( .A(n15684), .ZN(n15686) );
  OAI21_X1 U18855 ( .B1(n15686), .B2(n15685), .A(n18710), .ZN(n18705) );
  OAI21_X1 U18856 ( .B1(n18281), .B2(n16445), .A(n18792), .ZN(n15687) );
  OAI21_X1 U18857 ( .B1(n15688), .B2(n15687), .A(n18919), .ZN(n16613) );
  NOR3_X1 U18858 ( .A1(n15691), .A2(n16614), .A3(n16613), .ZN(n15690) );
  AOI211_X1 U18859 ( .C1(n15691), .C2(n18707), .A(n15690), .B(n15689), .ZN(
        n15692) );
  OAI21_X1 U18860 ( .B1(n15815), .B2(n18705), .A(n15692), .ZN(n15693) );
  INV_X1 U18861 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20878) );
  INV_X1 U18862 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18070) );
  NOR2_X1 U18863 ( .A1(n20878), .A2(n18070), .ZN(n17715) );
  INV_X1 U18864 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17709) );
  INV_X1 U18865 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17995) );
  INV_X1 U18866 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18034) );
  INV_X1 U18867 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17994) );
  NOR2_X1 U18868 ( .A1(n18034), .A2(n17994), .ZN(n18021) );
  INV_X1 U18869 ( .A(n18021), .ZN(n17996) );
  NOR3_X1 U18870 ( .A1(n17709), .A2(n17995), .A3(n17996), .ZN(n17661) );
  AND2_X1 U18871 ( .A1(n17661), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15840) );
  NAND2_X1 U18872 ( .A1(n17715), .A2(n15840), .ZN(n17640) );
  NOR2_X1 U18873 ( .A1(n18144), .A2(n18137), .ZN(n18123) );
  NAND2_X1 U18874 ( .A1(n18123), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18125) );
  INV_X1 U18875 ( .A(n18125), .ZN(n18106) );
  NAND2_X1 U18876 ( .A1(n18106), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18088) );
  INV_X1 U18877 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17774) );
  INV_X1 U18878 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18093) );
  OR2_X1 U18879 ( .A1(n18092), .A2(n18093), .ZN(n18075) );
  INV_X1 U18880 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18082) );
  NOR2_X1 U18881 ( .A1(n18075), .A2(n18082), .ZN(n18041) );
  INV_X1 U18882 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18173) );
  INV_X1 U18883 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18206) );
  INV_X1 U18884 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18187) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18198) );
  NOR3_X1 U18886 ( .A1(n18206), .A2(n18187), .A3(n18198), .ZN(n18156) );
  NAND2_X1 U18887 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18156), .ZN(
        n18170) );
  NOR2_X1 U18888 ( .A1(n18173), .A2(n18170), .ZN(n18153) );
  NAND2_X1 U18889 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18153), .ZN(
        n18074) );
  NAND2_X1 U18890 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18155) );
  NOR2_X1 U18891 ( .A1(n18074), .A2(n18155), .ZN(n18062) );
  NAND2_X1 U18892 ( .A1(n18041), .A2(n18062), .ZN(n18043) );
  NOR2_X1 U18893 ( .A1(n17640), .A2(n18043), .ZN(n15695) );
  NAND2_X1 U18894 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15695), .ZN(
        n17997) );
  INV_X1 U18895 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17991) );
  INV_X1 U18896 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17938) );
  NAND2_X1 U18897 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17941) );
  NOR3_X1 U18898 ( .A1(n17991), .A2(n17938), .A3(n17941), .ZN(n15694) );
  NAND2_X1 U18899 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15694), .ZN(
        n16499) );
  OAI21_X1 U18900 ( .B1(n17997), .B2(n16499), .A(n18743), .ZN(n15697) );
  INV_X1 U18901 ( .A(n17715), .ZN(n18048) );
  AOI21_X1 U18902 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18154) );
  NOR2_X1 U18903 ( .A1(n18154), .A2(n18074), .ZN(n18061) );
  NAND2_X1 U18904 ( .A1(n18041), .A2(n18061), .ZN(n18004) );
  NOR2_X1 U18905 ( .A1(n18048), .A2(n18004), .ZN(n18044) );
  NAND2_X1 U18906 ( .A1(n15840), .A2(n18044), .ZN(n17979) );
  INV_X1 U18907 ( .A(n15694), .ZN(n16457) );
  OAI21_X1 U18908 ( .B1(n17979), .B2(n16457), .A(n18717), .ZN(n17942) );
  INV_X1 U18909 ( .A(n15695), .ZN(n17939) );
  OAI21_X1 U18910 ( .B1(n16457), .B2(n17939), .A(n18726), .ZN(n15696) );
  NAND4_X1 U18911 ( .A1(n18231), .A2(n15697), .A3(n17942), .A4(n15696), .ZN(
        n15900) );
  AOI21_X1 U18912 ( .B1(n18126), .B2(n10178), .A(n15900), .ZN(n16507) );
  OAI21_X1 U18913 ( .B1(n18158), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16507), .ZN(n15833) );
  NAND2_X1 U18914 ( .A1(n18706), .A2(n18231), .ZN(n18251) );
  NAND2_X1 U18915 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16472) );
  INV_X1 U18916 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15848) );
  NOR2_X1 U18917 ( .A1(n16472), .A2(n15848), .ZN(n16446) );
  INV_X1 U18918 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U18919 ( .A1(n17640), .A2(n17991), .ZN(n17633) );
  NAND2_X1 U18920 ( .A1(n17633), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17961) );
  INV_X1 U18921 ( .A(n17961), .ZN(n17963) );
  AOI22_X1 U18922 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15701) );
  AOI22_X1 U18923 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15700) );
  AOI22_X1 U18924 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U18925 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15698) );
  NAND4_X1 U18926 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        n15707) );
  AOI22_X1 U18927 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15705) );
  AOI22_X1 U18928 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U18929 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18930 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15702) );
  NAND4_X1 U18931 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15706) );
  AOI22_X1 U18932 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15717) );
  AOI22_X1 U18933 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U18934 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15708) );
  OAI21_X1 U18935 ( .B1(n17178), .B2(n18297), .A(n15708), .ZN(n15714) );
  AOI22_X1 U18936 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15712) );
  AOI22_X1 U18937 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15711) );
  AOI22_X1 U18938 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18939 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15709) );
  NAND4_X1 U18940 ( .A1(n15712), .A2(n15711), .A3(n15710), .A4(n15709), .ZN(
        n15713) );
  AOI211_X1 U18941 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15714), .B(n15713), .ZN(n15715) );
  NAND3_X1 U18942 ( .A1(n15717), .A2(n15716), .A3(n15715), .ZN(n17441) );
  AOI22_X1 U18943 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17260), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U18944 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18945 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U18946 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15718) );
  NAND4_X1 U18947 ( .A1(n15721), .A2(n15720), .A3(n15719), .A4(n15718), .ZN(
        n15727) );
  AOI22_X1 U18948 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U18949 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U18950 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15723) );
  AOI22_X1 U18951 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15722) );
  NAND4_X1 U18952 ( .A1(n15725), .A2(n15724), .A3(n15723), .A4(n15722), .ZN(
        n15726) );
  INV_X1 U18953 ( .A(n17445), .ZN(n15788) );
  AOI22_X1 U18954 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15735) );
  AOI22_X1 U18955 ( .A1(n15753), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U18956 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U18957 ( .A1(n15741), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15740), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U18958 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15729), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U18959 ( .A1(n15737), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U18960 ( .A1(n15736), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15738), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15730) );
  INV_X1 U18961 ( .A(n15817), .ZN(n17450) );
  AOI22_X1 U18962 ( .A1(n15736), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18963 ( .A1(n15729), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18964 ( .A1(n15753), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15738), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U18965 ( .A1(n15740), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15739), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15745) );
  AOI22_X1 U18966 ( .A1(n15751), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15741), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U18967 ( .A1(n15742), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15752), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15743) );
  NAND4_X1 U18968 ( .A1(n15746), .A2(n15745), .A3(n15744), .A4(n15743), .ZN(
        n15747) );
  AOI22_X1 U18969 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U18970 ( .A1(n15780), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15761) );
  AOI22_X1 U18971 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15729), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15750) );
  OAI21_X1 U18972 ( .B1(n17178), .B2(n18270), .A(n15750), .ZN(n15759) );
  AOI22_X1 U18973 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18974 ( .A1(n15751), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15736), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15756) );
  AOI22_X1 U18975 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15752), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U18976 ( .A1(n15753), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15754) );
  NAND4_X1 U18977 ( .A1(n15757), .A2(n15756), .A3(n15755), .A4(n15754), .ZN(
        n15758) );
  AOI211_X1 U18978 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15759), .B(n15758), .ZN(n15760) );
  NAND3_X1 U18979 ( .A1(n15762), .A2(n15761), .A3(n15760), .ZN(n17930) );
  NAND2_X1 U18980 ( .A1(n17455), .A2(n17930), .ZN(n15789) );
  NAND2_X1 U18981 ( .A1(n17450), .A2(n15789), .ZN(n15787) );
  AOI22_X1 U18982 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U18983 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15765) );
  AOI22_X1 U18984 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U18985 ( .A1(n15780), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15763) );
  NAND4_X1 U18986 ( .A1(n15766), .A2(n15765), .A3(n15764), .A4(n15763), .ZN(
        n15772) );
  AOI22_X1 U18987 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15770) );
  AOI22_X1 U18988 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15769) );
  AOI22_X1 U18989 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U18990 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15767) );
  NAND4_X1 U18991 ( .A1(n15770), .A2(n15769), .A3(n15768), .A4(n15767), .ZN(
        n15771) );
  INV_X1 U18992 ( .A(n17437), .ZN(n15785) );
  NAND2_X1 U18993 ( .A1(n15784), .A2(n15785), .ZN(n15802) );
  NOR2_X1 U18994 ( .A1(n17433), .A2(n15802), .ZN(n15806) );
  AOI22_X1 U18995 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15783) );
  AOI22_X1 U18996 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18997 ( .A1(n17239), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15773) );
  OAI21_X1 U18998 ( .B1(n17178), .B2(n18320), .A(n15773), .ZN(n15779) );
  AOI22_X1 U18999 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15777) );
  AOI22_X1 U19000 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U19001 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15775) );
  AOI22_X1 U19002 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15774) );
  NAND4_X1 U19003 ( .A1(n15777), .A2(n15776), .A3(n15775), .A4(n15774), .ZN(
        n15778) );
  AOI211_X1 U19004 ( .C1(n15780), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15779), .B(n15778), .ZN(n15781) );
  NAND2_X1 U19005 ( .A1(n15806), .A2(n16505), .ZN(n15807) );
  XOR2_X1 U19006 ( .A(n15785), .B(n15784), .Z(n15786) );
  XOR2_X1 U19007 ( .A(n18198), .B(n15786), .Z(n17869) );
  XNOR2_X1 U19008 ( .A(n15788), .B(n15787), .ZN(n15797) );
  NOR2_X1 U19009 ( .A1(n18187), .A2(n15797), .ZN(n15798) );
  XNOR2_X1 U19010 ( .A(n15817), .B(n15789), .ZN(n15790) );
  INV_X1 U19011 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18234) );
  NOR2_X1 U19012 ( .A1(n15790), .A2(n18234), .ZN(n15796) );
  XOR2_X1 U19013 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15790), .Z(
        n17913) );
  INV_X1 U19014 ( .A(n17455), .ZN(n15792) );
  INV_X1 U19015 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18902) );
  NOR2_X1 U19016 ( .A1(n15792), .A2(n18902), .ZN(n15794) );
  INV_X1 U19017 ( .A(n17930), .ZN(n15793) );
  NAND3_X1 U19018 ( .A1(n15793), .A2(n15792), .A3(n18902), .ZN(n15791) );
  OAI221_X1 U19019 ( .B1(n15794), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15793), .C2(n15792), .A(n15791), .ZN(n17912) );
  NOR2_X1 U19020 ( .A1(n17913), .A2(n17912), .ZN(n15795) );
  NOR2_X1 U19021 ( .A1(n15796), .A2(n15795), .ZN(n17901) );
  XOR2_X1 U19022 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15797), .Z(
        n17900) );
  NOR2_X1 U19023 ( .A1(n17901), .A2(n17900), .ZN(n17899) );
  NOR2_X1 U19024 ( .A1(n15798), .A2(n17899), .ZN(n17883) );
  XNOR2_X1 U19025 ( .A(n17441), .B(n15799), .ZN(n17884) );
  NOR2_X1 U19026 ( .A1(n17883), .A2(n17884), .ZN(n15800) );
  NAND2_X1 U19027 ( .A1(n17883), .A2(n17884), .ZN(n17882) );
  OAI21_X1 U19028 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15800), .A(
        n17882), .ZN(n17868) );
  XNOR2_X1 U19029 ( .A(n17433), .B(n15802), .ZN(n15804) );
  NOR2_X1 U19030 ( .A1(n15803), .A2(n15804), .ZN(n15805) );
  INV_X1 U19031 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18188) );
  XNOR2_X1 U19032 ( .A(n15804), .B(n15803), .ZN(n17862) );
  NOR2_X1 U19033 ( .A1(n15805), .A2(n17861), .ZN(n15808) );
  XOR2_X1 U19034 ( .A(n17430), .B(n15806), .Z(n15809) );
  NAND2_X1 U19035 ( .A1(n15808), .A2(n15809), .ZN(n17850) );
  NOR2_X1 U19036 ( .A1(n15807), .A2(n15811), .ZN(n15813) );
  INV_X1 U19037 ( .A(n15807), .ZN(n15812) );
  OR2_X1 U19038 ( .A1(n15809), .A2(n15808), .ZN(n17851) );
  OAI21_X1 U19039 ( .B1(n15812), .B2(n15811), .A(n17851), .ZN(n15810) );
  INV_X1 U19040 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18161) );
  NAND2_X1 U19041 ( .A1(n17963), .A2(n18080), .ZN(n17621) );
  NOR2_X1 U19042 ( .A1(n17964), .A2(n17621), .ZN(n17620) );
  NAND2_X1 U19043 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17620), .ZN(
        n17580) );
  INV_X1 U19044 ( .A(n17580), .ZN(n17944) );
  NAND2_X1 U19045 ( .A1(n16446), .A2(n17944), .ZN(n16459) );
  NAND2_X1 U19046 ( .A1(n17430), .A2(n18247), .ZN(n18040) );
  INV_X1 U19047 ( .A(n18040), .ZN(n18164) );
  NAND2_X1 U19048 ( .A1(n17455), .A2(n15817), .ZN(n15819) );
  NAND2_X1 U19049 ( .A1(n15821), .A2(n17441), .ZN(n15823) );
  XNOR2_X1 U19050 ( .A(n15826), .B(n17433), .ZN(n15824) );
  NOR2_X1 U19051 ( .A1(n15824), .A2(n18188), .ZN(n15825) );
  INV_X1 U19052 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18886) );
  NOR2_X1 U19053 ( .A1(n17455), .A2(n18886), .ZN(n15816) );
  NAND2_X1 U19054 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17930), .ZN(
        n17929) );
  XOR2_X1 U19055 ( .A(n17455), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17921) );
  XNOR2_X1 U19056 ( .A(n15819), .B(n17445), .ZN(n17898) );
  XNOR2_X1 U19057 ( .A(n15821), .B(n17441), .ZN(n17887) );
  XNOR2_X1 U19058 ( .A(n15823), .B(n17437), .ZN(n17872) );
  XOR2_X1 U19059 ( .A(n15824), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(
        n17859) );
  OAI21_X1 U19060 ( .B1(n15827), .B2(n16505), .A(n17829), .ZN(n15829) );
  NOR2_X1 U19061 ( .A1(n15828), .A2(n15829), .ZN(n15830) );
  XNOR2_X1 U19062 ( .A(n15829), .B(n15828), .ZN(n17849) );
  NOR2_X1 U19063 ( .A1(n18173), .A2(n17849), .ZN(n17848) );
  INV_X1 U19064 ( .A(n18041), .ZN(n18016) );
  NAND2_X1 U19065 ( .A1(n18073), .A2(n17963), .ZN(n17609) );
  NAND2_X1 U19066 ( .A1(n16471), .A2(n16446), .ZN(n16458) );
  AOI22_X1 U19067 ( .A1(n18236), .A2(n16459), .B1(n18164), .B2(n16458), .ZN(
        n15902) );
  INV_X1 U19068 ( .A(n15902), .ZN(n15832) );
  AOI21_X1 U19069 ( .B1(n18181), .B2(n15833), .A(n15832), .ZN(n15849) );
  NAND3_X1 U19070 ( .A1(n16505), .A2(n18225), .A3(n18231), .ZN(n18169) );
  NOR2_X1 U19071 ( .A1(n17818), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17716) );
  NAND2_X1 U19072 ( .A1(n17716), .A2(n18034), .ZN(n15834) );
  NOR2_X1 U19073 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15834), .ZN(
        n17672) );
  NAND2_X1 U19074 ( .A1(n17672), .A2(n17995), .ZN(n17662) );
  NOR4_X1 U19075 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15835) );
  INV_X1 U19076 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18113) );
  NAND2_X1 U19077 ( .A1(n15837), .A2(n15838), .ZN(n17730) );
  NAND2_X1 U19078 ( .A1(n17715), .A2(n17730), .ZN(n17670) );
  NOR2_X1 U19079 ( .A1(n15842), .A2(n17829), .ZN(n17622) );
  NAND2_X1 U19080 ( .A1(n17829), .A2(n17623), .ZN(n15841) );
  NAND2_X1 U19081 ( .A1(n17818), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16500) );
  OAI21_X1 U19082 ( .B1(n17586), .B2(n16500), .A(n15897), .ZN(n15843) );
  XOR2_X1 U19083 ( .A(n15843), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16478) );
  NOR3_X1 U19084 ( .A1(n17961), .A2(n17941), .A3(n18248), .ZN(n16487) );
  NAND2_X1 U19085 ( .A1(n17430), .A2(n18225), .ZN(n18072) );
  NOR2_X1 U19086 ( .A1(n18228), .A2(n18002), .ZN(n15844) );
  AOI21_X1 U19087 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18743), .A(
        n18726), .ZN(n18215) );
  OAI22_X1 U19088 ( .A1(n18738), .A2(n18004), .B1(n18215), .B2(n18043), .ZN(
        n17962) );
  INV_X1 U19089 ( .A(n17986), .ZN(n15845) );
  NAND2_X1 U19090 ( .A1(n16487), .A2(n15845), .ZN(n17947) );
  NOR3_X1 U19091 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16472), .A3(
        n17947), .ZN(n15846) );
  AOI21_X1 U19092 ( .B1(n18150), .B2(n16478), .A(n15846), .ZN(n15847) );
  NAND2_X1 U19093 ( .A1(n9593), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16485) );
  OAI211_X1 U19094 ( .C1(n15849), .C2(n15848), .A(n15847), .B(n16485), .ZN(
        P3_U2833) );
  OAI21_X1 U19095 ( .B1(n9717), .B2(n15850), .A(n19098), .ZN(n15851) );
  OAI22_X1 U19096 ( .A1(n15852), .A2(n15851), .B1(n19109), .B2(n13512), .ZN(
        n15853) );
  AOI21_X1 U19097 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19103), .A(
        n15853), .ZN(n15858) );
  AOI222_X1 U19098 ( .A1(n15856), .A2(n19104), .B1(n19115), .B2(n15855), .C1(
        n19070), .C2(n15854), .ZN(n15857) );
  OAI211_X1 U19099 ( .C1(n19772), .C2(n19091), .A(n15858), .B(n15857), .ZN(
        P2_U2833) );
  INV_X1 U19100 ( .A(n15859), .ZN(n15861) );
  NOR3_X1 U19101 ( .A1(n15861), .A2(n15860), .A3(n20509), .ZN(n15867) );
  INV_X1 U19102 ( .A(n15867), .ZN(n15865) );
  INV_X1 U19103 ( .A(n15862), .ZN(n15863) );
  OAI211_X1 U19104 ( .C1(n10622), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15866) );
  OAI21_X1 U19105 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15867), .A(
        n15866), .ZN(n15868) );
  AOI222_X1 U19106 ( .A1(n15869), .A2(n15868), .B1(n15869), .B2(n10625), .C1(
        n15868), .C2(n10625), .ZN(n15873) );
  INV_X1 U19107 ( .A(n15873), .ZN(n15871) );
  OAI21_X1 U19108 ( .B1(n15871), .B2(n20474), .A(n15870), .ZN(n15872) );
  OAI21_X1 U19109 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15873), .A(
        n15872), .ZN(n15883) );
  INV_X1 U19110 ( .A(n15874), .ZN(n15882) );
  INV_X1 U19111 ( .A(n15875), .ZN(n15879) );
  OAI21_X1 U19112 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15876), .ZN(n15878) );
  NAND4_X1 U19113 ( .A1(n15880), .A2(n15879), .A3(n15878), .A4(n15877), .ZN(
        n15881) );
  AOI211_X1 U19114 ( .C1(n15883), .C2(n20094), .A(n15882), .B(n15881), .ZN(
        n15896) );
  NOR3_X1 U19115 ( .A1(n15885), .A2(n15907), .A3(n15884), .ZN(n15886) );
  AOI221_X1 U19116 ( .B1(n15888), .B2(n15887), .C1(n20741), .C2(n15887), .A(
        n15886), .ZN(n16179) );
  OAI221_X1 U19117 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15896), 
        .A(n16179), .ZN(n16186) );
  NOR2_X1 U19118 ( .A1(n16176), .A2(n20722), .ZN(n15889) );
  NOR2_X1 U19119 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15889), .ZN(n15893) );
  AOI21_X1 U19120 ( .B1(n15905), .B2(n10675), .A(n15890), .ZN(n15891) );
  NAND2_X1 U19121 ( .A1(n16186), .A2(n15891), .ZN(n15892) );
  AOI22_X1 U19122 ( .A1(n16186), .A2(n15893), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15892), .ZN(n15894) );
  OAI211_X1 U19123 ( .C1(n15896), .C2(n19849), .A(n15895), .B(n15894), .ZN(
        P1_U3161) );
  INV_X1 U19124 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U19125 ( .A1(n16446), .A2(n16460), .ZN(n16469) );
  INV_X1 U19126 ( .A(n16449), .ZN(n15898) );
  NOR2_X1 U19127 ( .A1(n16448), .A2(n15898), .ZN(n15899) );
  AOI21_X1 U19128 ( .B1(n15899), .B2(n16460), .A(n16451), .ZN(n16466) );
  NOR2_X1 U19129 ( .A1(n18158), .A2(n18248), .ZN(n18240) );
  INV_X1 U19130 ( .A(n16446), .ZN(n15901) );
  AOI22_X1 U19131 ( .A1(n18240), .A2(n15901), .B1(n18181), .B2(n15900), .ZN(
        n16490) );
  AOI21_X1 U19132 ( .B1(n16490), .B2(n15902), .A(n16460), .ZN(n15903) );
  AOI21_X1 U19133 ( .B1(n18150), .B2(n16466), .A(n15903), .ZN(n15904) );
  NAND2_X1 U19134 ( .A1(n9593), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16461) );
  OAI211_X1 U19135 ( .C1(n17947), .C2(n16469), .A(n15904), .B(n16461), .ZN(
        P3_U2832) );
  NAND2_X1 U19136 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15905), .ZN(n20662) );
  INV_X1 U19137 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20661) );
  NOR2_X1 U19138 ( .A1(n20668), .A2(n20661), .ZN(n20665) );
  INV_X1 U19139 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20825) );
  INV_X1 U19140 ( .A(HOLD), .ZN(n19731) );
  NOR2_X1 U19141 ( .A1(n20825), .A2(n19731), .ZN(n20657) );
  OAI22_X1 U19142 ( .A1(n20665), .A2(n20657), .B1(n20670), .B2(n19731), .ZN(
        n15906) );
  NAND3_X1 U19143 ( .A1(n15907), .A2(n20662), .A3(n15906), .ZN(P1_U3195) );
  AND2_X1 U19144 ( .A1(n19986), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19145 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15909) );
  NOR2_X1 U19146 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15908) );
  NOR2_X1 U19147 ( .A1(n16435), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19715) );
  AND2_X1 U19148 ( .A1(n19733), .A2(n19715), .ZN(n16418) );
  NOR4_X1 U19149 ( .A1(n15909), .A2(n15908), .A3(n16418), .A4(n16434), .ZN(
        P2_U3178) );
  INV_X1 U19150 ( .A(n19843), .ZN(n15910) );
  AOI221_X1 U19151 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16434), .C1(n15910), .C2(
        n16434), .A(n19655), .ZN(n19834) );
  INV_X1 U19152 ( .A(n19834), .ZN(n19835) );
  NOR2_X1 U19153 ( .A1(n15911), .A2(n19835), .ZN(P2_U3047) );
  OAI221_X1 U19154 ( .B1(n15914), .B2(n15913), .C1(n15914), .C2(n15912), .A(
        n18923), .ZN(n17309) );
  INV_X1 U19155 ( .A(n17309), .ZN(n15915) );
  INV_X1 U19156 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17533) );
  NAND2_X1 U19157 ( .A1(n18316), .A2(n15915), .ZN(n17358) );
  NAND2_X1 U19158 ( .A1(n17449), .A2(n17460), .ZN(n17459) );
  AOI22_X1 U19159 ( .A1(n17457), .A2(BUF2_REG_0__SCAN_IN), .B1(n17456), .B2(
        n17930), .ZN(n15916) );
  OAI221_X1 U19160 ( .B1(n17459), .B2(n17533), .C1(n17459), .C2(n17358), .A(
        n15916), .ZN(P3_U2735) );
  AOI22_X1 U19161 ( .A1(n15917), .A2(n19879), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n19934), .ZN(n15925) );
  AOI21_X1 U19162 ( .B1(n15918), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15920) );
  OAI22_X1 U19163 ( .A1(n15921), .A2(n15943), .B1(n15920), .B2(n15919), .ZN(
        n15922) );
  AOI21_X1 U19164 ( .B1(n19914), .B2(n15923), .A(n15922), .ZN(n15924) );
  OAI211_X1 U19165 ( .C1(n15926), .C2(n19926), .A(n15925), .B(n15924), .ZN(
        P1_U2817) );
  NOR2_X1 U19166 ( .A1(n19926), .A2(n15927), .ZN(n15930) );
  NOR3_X1 U19167 ( .A1(n19890), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n15928), 
        .ZN(n15929) );
  AOI211_X1 U19168 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n19934), .A(n15930), .B(
        n15929), .ZN(n15932) );
  NAND2_X1 U19169 ( .A1(n15942), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15931) );
  OAI211_X1 U19170 ( .C1(n15933), .C2(n15943), .A(n15932), .B(n15931), .ZN(
        n15934) );
  AOI21_X1 U19171 ( .B1(n15935), .B2(n19879), .A(n15934), .ZN(n15936) );
  OAI21_X1 U19172 ( .B1(n19939), .B2(n15937), .A(n15936), .ZN(P1_U2819) );
  AND2_X1 U19173 ( .A1(n19923), .A2(n15938), .ZN(n15941) );
  OAI22_X1 U19174 ( .A1(n15939), .A2(n19926), .B1(n20792), .B2(n16011), .ZN(
        n15940) );
  AOI221_X1 U19175 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n15942), .C1(n15941), 
        .C2(n15942), .A(n15940), .ZN(n15946) );
  OAI22_X1 U19176 ( .A1(n16021), .A2(n15943), .B1(n19939), .B2(n16019), .ZN(
        n15944) );
  INV_X1 U19177 ( .A(n15944), .ZN(n15945) );
  OAI211_X1 U19178 ( .C1(n15947), .C2(n19948), .A(n15946), .B(n15945), .ZN(
        P1_U2820) );
  NOR3_X1 U19179 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15948), .A3(n19873), 
        .ZN(n15953) );
  AOI22_X1 U19180 ( .A1(n15949), .A2(n19879), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n19934), .ZN(n15950) );
  OAI211_X1 U19181 ( .C1(n15951), .C2(n19926), .A(n15950), .B(n20068), .ZN(
        n15952) );
  AOI211_X1 U19182 ( .C1(n15954), .C2(n19904), .A(n15953), .B(n15952), .ZN(
        n15959) );
  AOI21_X1 U19183 ( .B1(n15955), .B2(n15956), .A(n15982), .ZN(n15977) );
  INV_X1 U19184 ( .A(n15956), .ZN(n15957) );
  NOR3_X1 U19185 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15957), .A3(n15974), 
        .ZN(n15961) );
  OAI21_X1 U19186 ( .B1(n15977), .B2(n15961), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15958) );
  OAI211_X1 U19187 ( .C1(n15960), .C2(n19939), .A(n15959), .B(n15958), .ZN(
        P1_U2821) );
  AOI21_X1 U19188 ( .B1(n19879), .B2(n15962), .A(n15961), .ZN(n15969) );
  AOI22_X1 U19189 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19901), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n19934), .ZN(n15968) );
  AOI21_X1 U19190 ( .B1(n15977), .B2(P1_REIP_REG_18__SCAN_IN), .A(n20021), 
        .ZN(n15967) );
  NOR2_X1 U19191 ( .A1(n15963), .A2(n19939), .ZN(n15964) );
  AOI21_X1 U19192 ( .B1(n15965), .B2(n19904), .A(n15964), .ZN(n15966) );
  NAND4_X1 U19193 ( .A1(n15969), .A2(n15968), .A3(n15967), .A4(n15966), .ZN(
        P1_U2822) );
  OAI22_X1 U19194 ( .A1(n15971), .A2(n19926), .B1(n15970), .B2(n16011), .ZN(
        n15972) );
  AOI211_X1 U19195 ( .C1(n19879), .C2(n15973), .A(n20021), .B(n15972), .ZN(
        n15980) );
  OAI21_X1 U19196 ( .B1(n15975), .B2(n15974), .A(n20691), .ZN(n15976) );
  AOI22_X1 U19197 ( .A1(n15978), .A2(n19904), .B1(n15977), .B2(n15976), .ZN(
        n15979) );
  OAI211_X1 U19198 ( .C1(n19939), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        P1_U2823) );
  AND2_X1 U19199 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15990) );
  OAI211_X1 U19200 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15991), .B(n16016), .ZN(n15989) );
  NOR2_X1 U19201 ( .A1(n20685), .A2(n20686), .ZN(n15984) );
  AOI21_X1 U19202 ( .B1(n15984), .B2(n15983), .A(n15982), .ZN(n15998) );
  AOI22_X1 U19203 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n19934), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n15998), .ZN(n15985) );
  OAI21_X1 U19204 ( .B1(n16038), .B2(n19948), .A(n15985), .ZN(n15986) );
  AOI211_X1 U19205 ( .C1(n19901), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20021), .B(n15986), .ZN(n15988) );
  AOI22_X1 U19206 ( .A1(n16035), .A2(n19904), .B1(n19914), .B2(n16096), .ZN(
        n15987) );
  OAI211_X1 U19207 ( .C1(n15990), .C2(n15989), .A(n15988), .B(n15987), .ZN(
        P1_U2824) );
  NAND2_X1 U19208 ( .A1(n15991), .A2(n16016), .ZN(n15997) );
  AOI22_X1 U19209 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n19934), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n15998), .ZN(n15994) );
  OAI21_X1 U19210 ( .B1(n19948), .B2(n16045), .A(n20068), .ZN(n15992) );
  AOI21_X1 U19211 ( .B1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19901), .A(
        n15992), .ZN(n15993) );
  OAI211_X1 U19212 ( .C1(n19939), .C2(n16101), .A(n15994), .B(n15993), .ZN(
        n15995) );
  AOI21_X1 U19213 ( .B1(n16047), .B2(n19904), .A(n15995), .ZN(n15996) );
  OAI21_X1 U19214 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15997), .A(n15996), 
        .ZN(P1_U2825) );
  AOI22_X1 U19215 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19901), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n19934), .ZN(n16003) );
  AOI21_X1 U19216 ( .B1(n16109), .B2(n19914), .A(n20021), .ZN(n16002) );
  AOI22_X1 U19217 ( .A1(n16059), .A2(n19904), .B1(n19879), .B2(n16058), .ZN(
        n16001) );
  OAI221_X1 U19218 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(P1_REIP_REG_13__SCAN_IN), .C1(P1_REIP_REG_14__SCAN_IN), .C2(n15999), .A(n15998), .ZN(n16000) );
  NAND4_X1 U19219 ( .A1(n16003), .A2(n16002), .A3(n16001), .A4(n16000), .ZN(
        P1_U2826) );
  AOI21_X1 U19220 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16016), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16009) );
  OAI22_X1 U19221 ( .A1(n20808), .A2(n19926), .B1(n16026), .B2(n16011), .ZN(
        n16004) );
  AOI211_X1 U19222 ( .C1(n16024), .C2(n19914), .A(n20021), .B(n16004), .ZN(
        n16007) );
  INV_X1 U19223 ( .A(n16005), .ZN(n16062) );
  AOI22_X1 U19224 ( .A1(n16063), .A2(n19879), .B1(n19904), .B2(n16062), .ZN(
        n16006) );
  OAI211_X1 U19225 ( .C1(n16009), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        P1_U2828) );
  AOI21_X1 U19226 ( .B1(n19901), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20021), .ZN(n16010) );
  INV_X1 U19227 ( .A(n16010), .ZN(n16014) );
  OAI22_X1 U19228 ( .A1(n16012), .A2(n16011), .B1(n19939), .B2(n16123), .ZN(
        n16013) );
  AOI211_X1 U19229 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16015), .A(n16014), 
        .B(n16013), .ZN(n16018) );
  AOI22_X1 U19230 ( .A1(n16075), .A2(n19904), .B1(n16016), .B2(n16122), .ZN(
        n16017) );
  OAI211_X1 U19231 ( .C1(n16078), .C2(n19948), .A(n16018), .B(n16017), .ZN(
        P1_U2829) );
  OAI22_X1 U19232 ( .A1(n16021), .A2(n16020), .B1(n19954), .B2(n16019), .ZN(
        n16022) );
  INV_X1 U19233 ( .A(n16022), .ZN(n16023) );
  OAI21_X1 U19234 ( .B1(n13839), .B2(n20792), .A(n16023), .ZN(P1_U2852) );
  AOI22_X1 U19235 ( .A1(n16062), .A2(n19956), .B1(n19950), .B2(n16024), .ZN(
        n16025) );
  OAI21_X1 U19236 ( .B1(n13839), .B2(n16026), .A(n16025), .ZN(P1_U2860) );
  AOI22_X1 U19237 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16037) );
  INV_X1 U19238 ( .A(n14027), .ZN(n16030) );
  INV_X1 U19239 ( .A(n16027), .ZN(n16029) );
  AOI21_X1 U19240 ( .B1(n16030), .B2(n16029), .A(n16028), .ZN(n16039) );
  INV_X1 U19241 ( .A(n16031), .ZN(n16032) );
  NAND3_X1 U19242 ( .A1(n16039), .A2(n16032), .A3(n16040), .ZN(n16041) );
  NAND2_X1 U19243 ( .A1(n16041), .A2(n16040), .ZN(n16034) );
  XNOR2_X1 U19244 ( .A(n16034), .B(n16033), .ZN(n16097) );
  AOI22_X1 U19245 ( .A1(n16097), .A2(n20029), .B1(n20028), .B2(n16035), .ZN(
        n16036) );
  OAI211_X1 U19246 ( .C1(n20033), .C2(n16038), .A(n16037), .B(n16036), .ZN(
        P1_U2983) );
  INV_X1 U19247 ( .A(n16039), .ZN(n16044) );
  OAI21_X1 U19248 ( .B1(n13547), .B2(n16055), .A(n16040), .ZN(n16043) );
  INV_X1 U19249 ( .A(n16041), .ZN(n16042) );
  AOI21_X1 U19250 ( .B1(n16044), .B2(n16043), .A(n16042), .ZN(n16102) );
  AOI22_X1 U19251 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16049) );
  INV_X1 U19252 ( .A(n16045), .ZN(n16046) );
  AOI22_X1 U19253 ( .A1(n16047), .A2(n20028), .B1(n16064), .B2(n16046), .ZN(
        n16048) );
  OAI211_X1 U19254 ( .C1(n16102), .C2(n16067), .A(n16049), .B(n16048), .ZN(
        P1_U2984) );
  NAND3_X1 U19255 ( .A1(n16052), .A2(n16051), .A3(n16050), .ZN(n16054) );
  NAND2_X1 U19256 ( .A1(n16054), .A2(n16053), .ZN(n16057) );
  XNOR2_X1 U19257 ( .A(n16055), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16056) );
  XNOR2_X1 U19258 ( .A(n16057), .B(n16056), .ZN(n16108) );
  AOI22_X1 U19259 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U19260 ( .A1(n16059), .A2(n20028), .B1(n16064), .B2(n16058), .ZN(
        n16060) );
  OAI211_X1 U19261 ( .C1(n16108), .C2(n16067), .A(n16061), .B(n16060), .ZN(
        P1_U2985) );
  AOI22_X1 U19262 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U19263 ( .A1(n16064), .A2(n16063), .B1(n20028), .B2(n16062), .ZN(
        n16065) );
  OAI211_X1 U19264 ( .C1(n16068), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        P1_U2987) );
  AOI22_X1 U19265 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U19266 ( .A1(n16069), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16072) );
  NOR2_X1 U19267 ( .A1(n14027), .A2(n16136), .ZN(n16071) );
  MUX2_X1 U19268 ( .A(n16072), .B(n16071), .S(n16070), .Z(n16074) );
  XNOR2_X1 U19269 ( .A(n16074), .B(n16073), .ZN(n16125) );
  AOI22_X1 U19270 ( .A1(n20029), .A2(n16125), .B1(n20028), .B2(n16075), .ZN(
        n16076) );
  OAI211_X1 U19271 ( .C1(n20033), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        P1_U2988) );
  AOI22_X1 U19272 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16081) );
  AOI22_X1 U19273 ( .A1(n16079), .A2(n20029), .B1(n20028), .B2(n19888), .ZN(
        n16080) );
  OAI211_X1 U19274 ( .C1(n20033), .C2(n19896), .A(n16081), .B(n16080), .ZN(
        P1_U2992) );
  AOI22_X1 U19275 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16086) );
  XNOR2_X1 U19276 ( .A(n16083), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16084) );
  XNOR2_X1 U19277 ( .A(n16082), .B(n16084), .ZN(n16155) );
  AOI22_X1 U19278 ( .A1(n16155), .A2(n20029), .B1(n20028), .B2(n19951), .ZN(
        n16085) );
  OAI211_X1 U19279 ( .C1(n20033), .C2(n19907), .A(n16086), .B(n16085), .ZN(
        P1_U2993) );
  AOI22_X1 U19280 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16092) );
  OAI21_X1 U19281 ( .B1(n16089), .B2(n16088), .A(n16087), .ZN(n16090) );
  INV_X1 U19282 ( .A(n16090), .ZN(n16165) );
  AOI22_X1 U19283 ( .A1(n16165), .A2(n20029), .B1(n20028), .B2(n19918), .ZN(
        n16091) );
  OAI211_X1 U19284 ( .C1(n20033), .C2(n19921), .A(n16092), .B(n16091), .ZN(
        P1_U2994) );
  AOI21_X1 U19285 ( .B1(n13547), .B2(n16100), .A(n16093), .ZN(n16095) );
  AOI22_X1 U19286 ( .A1(n20021), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n16095), 
        .B2(n16094), .ZN(n16099) );
  AOI22_X1 U19287 ( .A1(n16097), .A2(n20075), .B1(n20071), .B2(n16096), .ZN(
        n16098) );
  OAI211_X1 U19288 ( .C1(n16107), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P1_U3015) );
  OAI22_X1 U19289 ( .A1(n16102), .A2(n20085), .B1(n20083), .B2(n16101), .ZN(
        n16103) );
  AOI21_X1 U19290 ( .B1(n16104), .B2(n13547), .A(n16103), .ZN(n16106) );
  NAND2_X1 U19291 ( .A1(n20021), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16105) );
  OAI211_X1 U19292 ( .C1(n16107), .C2(n13547), .A(n16106), .B(n16105), .ZN(
        P1_U3016) );
  OR2_X1 U19293 ( .A1(n16108), .A2(n20085), .ZN(n16111) );
  NAND2_X1 U19294 ( .A1(n20071), .A2(n16109), .ZN(n16110) );
  AND2_X1 U19295 ( .A1(n16111), .A2(n16110), .ZN(n16119) );
  NAND2_X1 U19296 ( .A1(n20021), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16118) );
  OAI21_X1 U19297 ( .B1(n16113), .B2(n16112), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16117) );
  NAND3_X1 U19298 ( .A1(n16115), .A2(n16114), .A3(n16120), .ZN(n16116) );
  NAND4_X1 U19299 ( .A1(n16119), .A2(n16118), .A3(n16117), .A4(n16116), .ZN(
        P1_U3017) );
  NAND2_X1 U19300 ( .A1(n16121), .A2(n16120), .ZN(n16128) );
  OAI22_X1 U19301 ( .A1(n20083), .A2(n16123), .B1(n16122), .B2(n20068), .ZN(
        n16124) );
  AOI21_X1 U19302 ( .B1(n16125), .B2(n20075), .A(n16124), .ZN(n16126) );
  OAI221_X1 U19303 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16128), 
        .C1(n16073), .C2(n16127), .A(n16126), .ZN(P1_U3020) );
  AOI21_X1 U19304 ( .B1(n20071), .B2(n16130), .A(n16129), .ZN(n16135) );
  AOI22_X1 U19305 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n10604), .B2(n16136), .ZN(
        n16132) );
  AOI22_X1 U19306 ( .A1(n16133), .A2(n20075), .B1(n16132), .B2(n16131), .ZN(
        n16134) );
  OAI211_X1 U19307 ( .C1(n16137), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        P1_U3021) );
  AOI21_X1 U19308 ( .B1(n20071), .B2(n16139), .A(n16138), .ZN(n16147) );
  AOI22_X1 U19309 ( .A1(n16141), .A2(n20075), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16140), .ZN(n16146) );
  INV_X1 U19310 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16144) );
  INV_X1 U19311 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16143) );
  OAI221_X1 U19312 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16144), .C2(n16143), .A(
        n16142), .ZN(n16145) );
  NAND3_X1 U19313 ( .A1(n16147), .A2(n16146), .A3(n16145), .ZN(P1_U3023) );
  AOI21_X1 U19314 ( .B1(n10016), .B2(n16149), .A(n16148), .ZN(n16151) );
  OR2_X1 U19315 ( .A1(n16151), .A2(n16150), .ZN(n19902) );
  INV_X1 U19316 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n16152) );
  OAI22_X1 U19317 ( .A1(n20083), .A2(n19902), .B1(n20068), .B2(n16152), .ZN(
        n16153) );
  INV_X1 U19318 ( .A(n16153), .ZN(n16157) );
  AOI22_X1 U19319 ( .A1(n16155), .A2(n20075), .B1(n16154), .B2(n16158), .ZN(
        n16156) );
  OAI211_X1 U19320 ( .C1(n16159), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        P1_U3025) );
  INV_X1 U19321 ( .A(n16160), .ZN(n16169) );
  INV_X1 U19322 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n16161) );
  OAI22_X1 U19323 ( .A1(n20083), .A2(n16162), .B1(n20068), .B2(n16161), .ZN(
        n16163) );
  INV_X1 U19324 ( .A(n16163), .ZN(n16167) );
  INV_X1 U19325 ( .A(n20049), .ZN(n20039) );
  AOI22_X1 U19326 ( .A1(n16165), .A2(n20075), .B1(n16164), .B2(n20039), .ZN(
        n16166) );
  OAI211_X1 U19327 ( .C1(n16169), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        P1_U3026) );
  NAND3_X1 U19328 ( .A1(n19935), .A2(n16171), .A3(n16170), .ZN(n16174) );
  OAI22_X1 U19329 ( .A1(n16175), .A2(n16174), .B1(n16173), .B2(n16172), .ZN(
        P1_U3468) );
  AOI21_X1 U19330 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16186), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16183) );
  AOI21_X1 U19331 ( .B1(n20355), .B2(n20741), .A(n16176), .ZN(n16182) );
  NAND4_X1 U19332 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n10675), .A4(n20741), .ZN(n16177) );
  AND2_X1 U19333 ( .A1(n16178), .A2(n16177), .ZN(n20651) );
  AOI21_X1 U19334 ( .B1(n20651), .B2(n16180), .A(n16179), .ZN(n16181) );
  NOR3_X1 U19335 ( .A1(n16183), .A2(n16182), .A3(n16181), .ZN(P1_U3162) );
  INV_X1 U19336 ( .A(n16184), .ZN(n16185) );
  OAI221_X1 U19337 ( .B1(n20355), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20355), 
        .C2(n16186), .A(n16185), .ZN(P1_U3466) );
  NOR2_X1 U19338 ( .A1(n16187), .A2(n19107), .ZN(n16188) );
  AOI21_X1 U19339 ( .B1(n16189), .B2(n19115), .A(n16188), .ZN(n16202) );
  INV_X1 U19340 ( .A(n16192), .ZN(n16199) );
  AOI22_X1 U19341 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19112), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19103), .ZN(n16193) );
  OAI21_X1 U19342 ( .B1(n16194), .B2(n19075), .A(n16193), .ZN(n16195) );
  INV_X1 U19343 ( .A(n16195), .ZN(n16197) );
  NAND2_X1 U19344 ( .A1(n16197), .A2(n16196), .ZN(n16198) );
  NAND2_X1 U19345 ( .A1(n16202), .A2(n16201), .ZN(P2_U2825) );
  AOI211_X1 U19346 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n19717), .ZN(
        n16214) );
  INV_X1 U19347 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16208) );
  AOI22_X1 U19348 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19112), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19087), .ZN(n16206) );
  OAI21_X1 U19349 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n16209) );
  AOI21_X1 U19350 ( .B1(n16210), .B2(n19104), .A(n16209), .ZN(n16211) );
  OAI21_X1 U19351 ( .B1(n16212), .B2(n19021), .A(n16211), .ZN(n16213) );
  AOI211_X1 U19352 ( .C1(n19070), .C2(n16215), .A(n16214), .B(n16213), .ZN(
        n16216) );
  INV_X1 U19353 ( .A(n16216), .ZN(P2_U2826) );
  AOI22_X1 U19354 ( .A1(n16217), .A2(n19104), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n19112), .ZN(n16228) );
  AOI22_X1 U19355 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19103), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19087), .ZN(n16227) );
  INV_X1 U19356 ( .A(n16218), .ZN(n16220) );
  AOI22_X1 U19357 ( .A1(n16220), .A2(n19115), .B1(n16219), .B2(n19070), .ZN(
        n16226) );
  AOI21_X1 U19358 ( .B1(n16223), .B2(n16222), .A(n16221), .ZN(n16224) );
  NAND2_X1 U19359 ( .A1(n19098), .A2(n16224), .ZN(n16225) );
  NAND4_X1 U19360 ( .A1(n16228), .A2(n16227), .A3(n16226), .A4(n16225), .ZN(
        P2_U2827) );
  AOI22_X1 U19361 ( .A1(n16230), .A2(n16229), .B1(n19131), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16237) );
  AOI22_X1 U19362 ( .A1(n19130), .A2(BUF2_REG_23__SCAN_IN), .B1(n19132), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16236) );
  INV_X1 U19363 ( .A(n16231), .ZN(n16232) );
  AOI22_X1 U19364 ( .A1(n16234), .A2(n16233), .B1(n19129), .B2(n16232), .ZN(
        n16235) );
  NAND3_X1 U19365 ( .A1(n16237), .A2(n16236), .A3(n16235), .ZN(P2_U2896) );
  AOI22_X1 U19366 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19215), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19111), .ZN(n16240) );
  AOI22_X1 U19367 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19111), .B1(n16295), 
        .B2(n16241), .ZN(n16251) );
  AOI21_X1 U19368 ( .B1(n16244), .B2(n16243), .A(n16242), .ZN(n16312) );
  NAND2_X1 U19369 ( .A1(n16246), .A2(n16245), .ZN(n16248) );
  XOR2_X1 U19370 ( .A(n16248), .B(n16247), .Z(n16307) );
  AOI222_X1 U19371 ( .A1(n16312), .A2(n19216), .B1(n16302), .B2(n16307), .C1(
        n19227), .C2(n16249), .ZN(n16250) );
  OAI211_X1 U19372 ( .C1(n16252), .C2(n16305), .A(n16251), .B(n16250), .ZN(
        P2_U3001) );
  AOI22_X1 U19373 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19111), .B1(n16295), 
        .B2(n19064), .ZN(n16261) );
  NAND2_X1 U19374 ( .A1(n9712), .A2(n16254), .ZN(n16255) );
  XNOR2_X1 U19375 ( .A(n16253), .B(n16255), .ZN(n16339) );
  NAND2_X1 U19376 ( .A1(n16258), .A2(n16257), .ZN(n16342) );
  INV_X1 U19377 ( .A(n16342), .ZN(n16259) );
  AOI222_X1 U19378 ( .A1(n16339), .A2(n16302), .B1(n19227), .B2(n19071), .C1(
        n19216), .C2(n16259), .ZN(n16260) );
  OAI211_X1 U19379 ( .C1(n16262), .C2(n16305), .A(n16261), .B(n16260), .ZN(
        P2_U3003) );
  AOI22_X1 U19380 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19111), .B1(n16295), 
        .B2(n16263), .ZN(n16268) );
  AOI222_X1 U19381 ( .A1(n16266), .A2(n19216), .B1(n16302), .B2(n16265), .C1(
        n19227), .C2(n16264), .ZN(n16267) );
  OAI211_X1 U19382 ( .C1(n16269), .C2(n16305), .A(n16268), .B(n16267), .ZN(
        P2_U3005) );
  AOI22_X1 U19383 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19111), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19215), .ZN(n16274) );
  OAI22_X1 U19384 ( .A1(n16271), .A2(n16287), .B1(n16270), .B2(n19218), .ZN(
        n16272) );
  AOI21_X1 U19385 ( .B1(n19227), .B2(n19097), .A(n16272), .ZN(n16273) );
  OAI211_X1 U19386 ( .C1(n19224), .C2(n19095), .A(n16274), .B(n16273), .ZN(
        P2_U3006) );
  AOI22_X1 U19387 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19111), .B1(n16295), 
        .B2(n16275), .ZN(n16284) );
  NAND2_X1 U19388 ( .A1(n16277), .A2(n16276), .ZN(n16278) );
  XNOR2_X1 U19389 ( .A(n15405), .B(n16278), .ZN(n16350) );
  XNOR2_X1 U19390 ( .A(n16279), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16280) );
  XNOR2_X1 U19391 ( .A(n16281), .B(n16280), .ZN(n16353) );
  INV_X1 U19392 ( .A(n16353), .ZN(n16282) );
  AOI222_X1 U19393 ( .A1(n16350), .A2(n16302), .B1(n19227), .B2(n16349), .C1(
        n19216), .C2(n16282), .ZN(n16283) );
  OAI211_X1 U19394 ( .C1(n16285), .C2(n16305), .A(n16284), .B(n16283), .ZN(
        P2_U3007) );
  AOI22_X1 U19395 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19111), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19215), .ZN(n16292) );
  OAI22_X1 U19396 ( .A1(n16288), .A2(n16287), .B1(n19218), .B2(n16286), .ZN(
        n16289) );
  AOI21_X1 U19397 ( .B1(n19227), .B2(n16290), .A(n16289), .ZN(n16291) );
  OAI211_X1 U19398 ( .C1(n19224), .C2(n16293), .A(n16292), .B(n16291), .ZN(
        P2_U3008) );
  AOI22_X1 U19399 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19111), .B1(n16295), 
        .B2(n16294), .ZN(n16304) );
  XOR2_X1 U19400 ( .A(n16297), .B(n16296), .Z(n16361) );
  NAND2_X1 U19401 ( .A1(n16299), .A2(n16298), .ZN(n16300) );
  XNOR2_X1 U19402 ( .A(n16301), .B(n16300), .ZN(n16359) );
  AOI222_X1 U19403 ( .A1(n16361), .A2(n16302), .B1(n16359), .B2(n19216), .C1(
        n19227), .C2(n16357), .ZN(n16303) );
  OAI211_X1 U19404 ( .C1(n16306), .C2(n16305), .A(n16304), .B(n16303), .ZN(
        P2_U3009) );
  AOI22_X1 U19405 ( .A1(n16321), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16371), .B2(n19137), .ZN(n16318) );
  INV_X1 U19406 ( .A(n16307), .ZN(n16310) );
  OAI22_X1 U19407 ( .A1(n16310), .A2(n16373), .B1(n16309), .B2(n16308), .ZN(
        n16311) );
  AOI21_X1 U19408 ( .B1(n16358), .B2(n16312), .A(n16311), .ZN(n16317) );
  NAND2_X1 U19409 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19111), .ZN(n16316) );
  INV_X1 U19410 ( .A(n16313), .ZN(n16323) );
  OAI211_X1 U19411 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16323), .B(n16314), .ZN(
        n16315) );
  NAND4_X1 U19412 ( .A1(n16318), .A2(n16317), .A3(n16316), .A4(n16315), .ZN(
        P2_U3033) );
  OAI22_X1 U19413 ( .A1(n16319), .A2(n19061), .B1(n19755), .B2(n19089), .ZN(
        n16320) );
  AOI221_X1 U19414 ( .B1(n16323), .B2(n16322), .C1(n16321), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16320), .ZN(n16326) );
  AOI22_X1 U19415 ( .A1(n16324), .A2(n16360), .B1(n16369), .B2(n19057), .ZN(
        n16325) );
  OAI211_X1 U19416 ( .C1(n16383), .C2(n16327), .A(n16326), .B(n16325), .ZN(
        P2_U3034) );
  AOI21_X1 U19417 ( .B1(n16330), .B2(n16329), .A(n16328), .ZN(n19141) );
  NAND2_X1 U19418 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19111), .ZN(n16335) );
  INV_X1 U19419 ( .A(n16331), .ZN(n16332) );
  OAI211_X1 U19420 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16333), .B(n16332), .ZN(
        n16334) );
  OAI211_X1 U19421 ( .C1(n16337), .C2(n16336), .A(n16335), .B(n16334), .ZN(
        n16338) );
  AOI21_X1 U19422 ( .B1(n16371), .B2(n19141), .A(n16338), .ZN(n16341) );
  AOI22_X1 U19423 ( .A1(n16339), .A2(n16360), .B1(n16369), .B2(n19071), .ZN(
        n16340) );
  OAI211_X1 U19424 ( .C1(n16383), .C2(n16342), .A(n16341), .B(n16340), .ZN(
        P2_U3035) );
  NAND2_X1 U19425 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19111), .ZN(n16343) );
  OAI221_X1 U19426 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16346), .C1(
        n16345), .C2(n16344), .A(n16343), .ZN(n16347) );
  AOI21_X1 U19427 ( .B1(n16348), .B2(n16371), .A(n16347), .ZN(n16352) );
  AOI22_X1 U19428 ( .A1(n16350), .A2(n16360), .B1(n16369), .B2(n16349), .ZN(
        n16351) );
  OAI211_X1 U19429 ( .C1(n16383), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        P2_U3039) );
  INV_X1 U19430 ( .A(n16354), .ZN(n16356) );
  AOI22_X1 U19431 ( .A1(n16356), .A2(n16371), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16355), .ZN(n16367) );
  AOI222_X1 U19432 ( .A1(n16361), .A2(n16360), .B1(n16359), .B2(n16358), .C1(
        n16369), .C2(n16357), .ZN(n16366) );
  NAND2_X1 U19433 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19111), .ZN(n16365) );
  OAI211_X1 U19434 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16363), .B(n16362), .ZN(n16364) );
  NAND4_X1 U19435 ( .A1(n16367), .A2(n16366), .A3(n16365), .A4(n16364), .ZN(
        P2_U3041) );
  AOI22_X1 U19436 ( .A1(n16371), .A2(n16370), .B1(n16369), .B2(n16368), .ZN(
        n16379) );
  OAI22_X1 U19437 ( .A1(n16374), .A2(n12087), .B1(n16373), .B2(n16372), .ZN(
        n16375) );
  INV_X1 U19438 ( .A(n16375), .ZN(n16378) );
  NAND2_X1 U19439 ( .A1(n16376), .A2(n12087), .ZN(n16377) );
  AND3_X1 U19440 ( .A1(n16379), .A2(n16378), .A3(n16377), .ZN(n16381) );
  OAI211_X1 U19441 ( .C1(n16383), .C2(n16382), .A(n16381), .B(n16380), .ZN(
        P2_U3046) );
  INV_X1 U19442 ( .A(n16387), .ZN(n16385) );
  OAI211_X1 U19443 ( .C1(n16385), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16384), .ZN(n16386) );
  OAI21_X1 U19444 ( .B1(n16387), .B2(n19827), .A(n16386), .ZN(n16388) );
  AOI211_X1 U19445 ( .C1(n16391), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16413), .B(n16388), .ZN(n16393) );
  INV_X1 U19446 ( .A(n16413), .ZN(n16389) );
  MUX2_X1 U19447 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16390), .S(
        n16389), .Z(n16411) );
  NOR2_X1 U19448 ( .A1(n16391), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16392) );
  OR3_X1 U19449 ( .A1(n16393), .A2(n16411), .A3(n16392), .ZN(n16394) );
  AOI22_X1 U19450 ( .A1(n16394), .A2(n19809), .B1(n16393), .B2(n16411), .ZN(
        n16416) );
  INV_X1 U19451 ( .A(n16395), .ZN(n16396) );
  AOI22_X1 U19452 ( .A1(n16401), .A2(n16398), .B1(n16397), .B2(n16396), .ZN(
        n16399) );
  OAI21_X1 U19453 ( .B1(n16401), .B2(n16400), .A(n16399), .ZN(n19838) );
  OAI21_X1 U19454 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16402), .ZN(n16406) );
  NAND3_X1 U19455 ( .A1(n16404), .A2(n16421), .A3(n16403), .ZN(n16405) );
  OAI211_X1 U19456 ( .C1(n16408), .C2(n16407), .A(n16406), .B(n16405), .ZN(
        n16409) );
  AOI211_X1 U19457 ( .C1(n16413), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19838), .B(n16409), .ZN(n16415) );
  NAND2_X1 U19458 ( .A1(n16413), .A2(n11550), .ZN(n16410) );
  OAI211_X1 U19459 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        n16414) );
  OAI211_X1 U19460 ( .C1(n16416), .C2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16415), .B(n16414), .ZN(n16419) );
  INV_X1 U19461 ( .A(n16419), .ZN(n16433) );
  AOI211_X1 U19462 ( .C1(n16434), .C2(n19843), .A(n16418), .B(n16417), .ZN(
        n16432) );
  OAI21_X1 U19463 ( .B1(n16419), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16423) );
  NAND3_X1 U19464 ( .A1(n11767), .A2(n16421), .A3(n16420), .ZN(n16422) );
  NAND2_X1 U19465 ( .A1(n16423), .A2(n16422), .ZN(n16424) );
  OAI21_X1 U19466 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16428), .A(n16427), 
        .ZN(n16430) );
  NAND2_X1 U19467 ( .A1(n19719), .A2(n19733), .ZN(n16429) );
  AOI22_X1 U19468 ( .A1(n19719), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16430), 
        .B2(n16429), .ZN(n16431) );
  OAI211_X1 U19469 ( .C1(n16433), .C2(n19146), .A(n16432), .B(n16431), .ZN(
        P2_U3176) );
  INV_X1 U19470 ( .A(n19719), .ZN(n16437) );
  AOI21_X1 U19471 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16435), .A(n16434), 
        .ZN(n16436) );
  OAI21_X1 U19472 ( .B1(n12070), .B2(n16437), .A(n16436), .ZN(P2_U3593) );
  INV_X1 U19473 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18887) );
  NAND3_X1 U19474 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16446), .A3(
        n16471), .ZN(n16438) );
  XNOR2_X1 U19475 ( .A(n18887), .B(n16438), .ZN(n16498) );
  NAND2_X1 U19476 ( .A1(n18765), .A2(n16440), .ZN(n17935) );
  INV_X1 U19477 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18858) );
  NOR2_X1 U19478 ( .A1(n18858), .A2(n18181), .ZN(n16492) );
  NAND2_X1 U19479 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16482), .ZN(
        n16441) );
  NAND2_X1 U19480 ( .A1(n18928), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17932) );
  OR2_X1 U19481 ( .A1(n16441), .A2(n17777), .ZN(n16463) );
  XNOR2_X1 U19482 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16443) );
  NOR2_X1 U19483 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17613), .ZN(
        n16480) );
  INV_X1 U19484 ( .A(n16479), .ZN(n16637) );
  NAND2_X1 U19485 ( .A1(n18653), .A2(n16441), .ZN(n16442) );
  OAI211_X1 U19486 ( .C1(n16637), .C2(n17932), .A(n16442), .B(n17931), .ZN(
        n16481) );
  NOR2_X1 U19487 ( .A1(n16480), .A2(n16481), .ZN(n16462) );
  OAI22_X1 U19488 ( .A1(n16463), .A2(n16443), .B1(n16462), .B2(n16654), .ZN(
        n16444) );
  AOI211_X1 U19489 ( .C1(n17772), .C2(n16986), .A(n16492), .B(n16444), .ZN(
        n16456) );
  NAND3_X1 U19490 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16446), .A3(
        n18887), .ZN(n16489) );
  OAI21_X1 U19491 ( .B1(n16460), .B2(n16459), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16447) );
  OAI21_X1 U19492 ( .B1(n16489), .B2(n17580), .A(n16447), .ZN(n16494) );
  AOI21_X1 U19493 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18887), .A(
        n16452), .ZN(n16450) );
  NOR2_X1 U19494 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18887), .ZN(
        n16493) );
  AOI21_X1 U19495 ( .B1(n16450), .B2(n16449), .A(n16493), .ZN(n16454) );
  AOI22_X1 U19496 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17818), .B1(
        n17829), .B2(n18887), .ZN(n16453) );
  OAI211_X1 U19497 ( .C1(n16498), .C2(n17751), .A(n16456), .B(n16455), .ZN(
        P3_U2799) );
  NOR3_X1 U19498 ( .A1(n17640), .A2(n16457), .A3(n17741), .ZN(n17595) );
  INV_X1 U19499 ( .A(n17595), .ZN(n16470) );
  XNOR2_X1 U19500 ( .A(n10061), .B(n9705), .ZN(n16657) );
  NAND2_X1 U19501 ( .A1(n17841), .A2(n16458), .ZN(n16475) );
  NAND2_X1 U19502 ( .A1(n9589), .A2(n16459), .ZN(n16473) );
  AOI21_X1 U19503 ( .B1(n16475), .B2(n16473), .A(n16460), .ZN(n16465) );
  OAI221_X1 U19504 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16463), .C1(
        n10061), .C2(n16462), .A(n16461), .ZN(n16464) );
  AOI211_X1 U19505 ( .C1(n17772), .C2(n16657), .A(n16465), .B(n16464), .ZN(
        n16468) );
  NAND2_X1 U19506 ( .A1(n17824), .A2(n16466), .ZN(n16467) );
  OAI211_X1 U19507 ( .C1(n16470), .C2(n16469), .A(n16468), .B(n16467), .ZN(
        P3_U2800) );
  INV_X1 U19508 ( .A(n16471), .ZN(n17946) );
  NOR2_X1 U19509 ( .A1(n17946), .A2(n16472), .ZN(n16506) );
  NOR2_X1 U19510 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16506), .ZN(
        n16476) );
  NOR2_X1 U19511 ( .A1(n16472), .A2(n17580), .ZN(n16508) );
  NOR2_X1 U19512 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16508), .ZN(
        n16474) );
  OAI22_X1 U19513 ( .A1(n16476), .A2(n16475), .B1(n16474), .B2(n16473), .ZN(
        n16477) );
  AOI21_X1 U19514 ( .B1(n17824), .B2(n16478), .A(n16477), .ZN(n16486) );
  AOI21_X1 U19515 ( .B1(n16667), .B2(n16479), .A(n9705), .ZN(n16666) );
  OAI21_X1 U19516 ( .B1(n16480), .B2(n17772), .A(n16666), .ZN(n16484) );
  OAI221_X1 U19517 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18653), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16482), .A(n16481), .ZN(
        n16483) );
  NAND4_X1 U19518 ( .A1(n16486), .A2(n16485), .A3(n16484), .A4(n16483), .ZN(
        P3_U2801) );
  NAND2_X1 U19519 ( .A1(n16487), .A2(n17962), .ZN(n16488) );
  OAI22_X1 U19520 ( .A1(n16490), .A2(n18887), .B1(n16489), .B2(n16488), .ZN(
        n16491) );
  AOI211_X1 U19521 ( .C1(n16493), .C2(n18240), .A(n16492), .B(n16491), .ZN(
        n16497) );
  AOI22_X1 U19522 ( .A1(n18150), .A2(n16495), .B1(n18236), .B2(n16494), .ZN(
        n16496) );
  OAI211_X1 U19523 ( .C1(n16498), .C2(n18040), .A(n16497), .B(n16496), .ZN(
        P3_U2831) );
  NOR2_X1 U19524 ( .A1(n17986), .A2(n18248), .ZN(n18014) );
  NOR3_X1 U19525 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17640), .A3(
        n16499), .ZN(n17578) );
  AOI22_X1 U19526 ( .A1(n9593), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18014), 
        .B2(n17578), .ZN(n16513) );
  AOI21_X1 U19527 ( .B1(n17818), .B2(n17586), .A(n17585), .ZN(n17577) );
  NAND2_X1 U19528 ( .A1(n9637), .A2(n16500), .ZN(n17576) );
  NOR2_X1 U19529 ( .A1(n17577), .A2(n17576), .ZN(n17575) );
  NOR3_X1 U19530 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17575), .A3(
        n16503), .ZN(n16501) );
  OAI221_X1 U19531 ( .B1(n16501), .B2(n17585), .C1(n16501), .C2(n17576), .A(
        n18150), .ZN(n16512) );
  INV_X1 U19532 ( .A(n17575), .ZN(n16502) );
  OAI21_X1 U19533 ( .B1(n17586), .B2(n16503), .A(n16502), .ZN(n16504) );
  AOI221_X1 U19534 ( .B1(n17430), .B2(n16506), .C1(n16505), .C2(n16504), .A(
        n18712), .ZN(n16510) );
  OAI21_X1 U19535 ( .B1(n16508), .B2(n18228), .A(n16507), .ZN(n16509) );
  OAI211_X1 U19536 ( .C1(n16510), .C2(n16509), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18181), .ZN(n16511) );
  NAND3_X1 U19537 ( .A1(n16513), .A2(n16512), .A3(n16511), .ZN(P3_U2834) );
  NOR3_X1 U19538 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16515) );
  NOR4_X1 U19539 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16514) );
  NAND4_X1 U19540 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16515), .A3(n16514), .A4(
        U215), .ZN(U213) );
  INV_X1 U19541 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16601) );
  NOR2_X2 U19542 ( .A1(n16565), .A2(n16516), .ZN(n16567) );
  INV_X1 U19543 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16602) );
  OAI222_X1 U19544 ( .A1(U212), .A2(n16601), .B1(n16558), .B2(n16517), .C1(
        U214), .C2(n16602), .ZN(U216) );
  AOI22_X1 U19545 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16556), .ZN(n16518) );
  OAI21_X1 U19546 ( .B1(n16519), .B2(n16558), .A(n16518), .ZN(U217) );
  AOI22_X1 U19547 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16556), .ZN(n16520) );
  OAI21_X1 U19548 ( .B1(n16521), .B2(n16558), .A(n16520), .ZN(U218) );
  AOI22_X1 U19549 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16556), .ZN(n16522) );
  OAI21_X1 U19550 ( .B1(n13859), .B2(n16558), .A(n16522), .ZN(U219) );
  AOI22_X1 U19551 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16556), .ZN(n16523) );
  OAI21_X1 U19552 ( .B1(n16524), .B2(n16558), .A(n16523), .ZN(U220) );
  AOI22_X1 U19553 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16556), .ZN(n16525) );
  OAI21_X1 U19554 ( .B1(n13868), .B2(n16558), .A(n16525), .ZN(U221) );
  AOI22_X1 U19555 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16556), .ZN(n16526) );
  OAI21_X1 U19556 ( .B1(n16527), .B2(n16558), .A(n16526), .ZN(U222) );
  AOI22_X1 U19557 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16556), .ZN(n16528) );
  OAI21_X1 U19558 ( .B1(n16529), .B2(n16558), .A(n16528), .ZN(U223) );
  AOI22_X1 U19559 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16556), .ZN(n16530) );
  OAI21_X1 U19560 ( .B1(n16531), .B2(n16558), .A(n16530), .ZN(U224) );
  AOI22_X1 U19561 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16556), .ZN(n16532) );
  OAI21_X1 U19562 ( .B1(n16533), .B2(n16558), .A(n16532), .ZN(U225) );
  AOI22_X1 U19563 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16556), .ZN(n16534) );
  OAI21_X1 U19564 ( .B1(n20774), .B2(n16558), .A(n16534), .ZN(U226) );
  AOI22_X1 U19565 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16556), .ZN(n16535) );
  OAI21_X1 U19566 ( .B1(n16536), .B2(n16558), .A(n16535), .ZN(U227) );
  AOI22_X1 U19567 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16556), .ZN(n16537) );
  OAI21_X1 U19568 ( .B1(n16538), .B2(n16558), .A(n16537), .ZN(U228) );
  AOI22_X1 U19569 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16556), .ZN(n16539) );
  OAI21_X1 U19570 ( .B1(n16540), .B2(n16558), .A(n16539), .ZN(U229) );
  AOI22_X1 U19571 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16556), .ZN(n16541) );
  OAI21_X1 U19572 ( .B1(n16542), .B2(n16558), .A(n16541), .ZN(U230) );
  AOI22_X1 U19573 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16556), .ZN(n16543) );
  OAI21_X1 U19574 ( .B1(n16544), .B2(n16558), .A(n16543), .ZN(U231) );
  INV_X1 U19575 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U19576 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16565), .ZN(n16545) );
  OAI21_X1 U19577 ( .B1(n20889), .B2(U212), .A(n16545), .ZN(U232) );
  INV_X1 U19578 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U19579 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16565), .ZN(n16546) );
  OAI21_X1 U19580 ( .B1(n20798), .B2(U212), .A(n16546), .ZN(U233) );
  AOI22_X1 U19581 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16556), .ZN(n16547) );
  OAI21_X1 U19582 ( .B1(n16548), .B2(n16558), .A(n16547), .ZN(U234) );
  INV_X1 U19583 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19584 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16565), .ZN(n16549) );
  OAI21_X1 U19585 ( .B1(n16581), .B2(U212), .A(n16549), .ZN(U235) );
  AOI22_X1 U19586 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16556), .ZN(n16550) );
  OAI21_X1 U19587 ( .B1(n16551), .B2(n16558), .A(n16550), .ZN(U236) );
  INV_X1 U19588 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16579) );
  AOI22_X1 U19589 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16565), .ZN(n16552) );
  OAI21_X1 U19590 ( .B1(n16579), .B2(U212), .A(n16552), .ZN(U237) );
  INV_X1 U19591 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U19592 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16565), .ZN(n16553) );
  OAI21_X1 U19593 ( .B1(n16554), .B2(U212), .A(n16553), .ZN(U238) );
  INV_X1 U19594 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U19595 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16567), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16556), .ZN(n16555) );
  OAI21_X1 U19596 ( .B1(n20822), .B2(U214), .A(n16555), .ZN(U239) );
  INV_X1 U19597 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U19598 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16565), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16556), .ZN(n16557) );
  OAI21_X1 U19599 ( .B1(n16559), .B2(n16558), .A(n16557), .ZN(U240) );
  INV_X1 U19600 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16575) );
  AOI22_X1 U19601 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16565), .ZN(n16560) );
  OAI21_X1 U19602 ( .B1(n16575), .B2(U212), .A(n16560), .ZN(U241) );
  INV_X1 U19603 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16574) );
  AOI22_X1 U19604 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16565), .ZN(n16561) );
  OAI21_X1 U19605 ( .B1(n16574), .B2(U212), .A(n16561), .ZN(U242) );
  INV_X1 U19606 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16573) );
  AOI22_X1 U19607 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16565), .ZN(n16562) );
  OAI21_X1 U19608 ( .B1(n16573), .B2(U212), .A(n16562), .ZN(U243) );
  INV_X1 U19609 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16572) );
  AOI22_X1 U19610 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16565), .ZN(n16563) );
  OAI21_X1 U19611 ( .B1(n16572), .B2(U212), .A(n16563), .ZN(U244) );
  INV_X1 U19612 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16571) );
  AOI22_X1 U19613 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16565), .ZN(n16564) );
  OAI21_X1 U19614 ( .B1(n16571), .B2(U212), .A(n16564), .ZN(U245) );
  INV_X1 U19615 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16570) );
  AOI22_X1 U19616 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16565), .ZN(n16566) );
  OAI21_X1 U19617 ( .B1(n16570), .B2(U212), .A(n16566), .ZN(U246) );
  INV_X1 U19618 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U19619 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16567), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16565), .ZN(n16568) );
  OAI21_X1 U19620 ( .B1(n16569), .B2(U212), .A(n16568), .ZN(U247) );
  INV_X1 U19621 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U19622 ( .A1(n20772), .A2(n16569), .B1(n18264), .B2(U215), .ZN(U251) );
  INV_X1 U19623 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18272) );
  AOI22_X1 U19624 ( .A1(n20772), .A2(n16570), .B1(n18272), .B2(U215), .ZN(U252) );
  INV_X1 U19625 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U19626 ( .A1(n20772), .A2(n16571), .B1(n18279), .B2(U215), .ZN(U253) );
  INV_X1 U19627 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U19628 ( .A1(n20772), .A2(n16572), .B1(n18286), .B2(U215), .ZN(U254) );
  INV_X1 U19629 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U19630 ( .A1(n16593), .A2(n16573), .B1(n20858), .B2(U215), .ZN(U255) );
  INV_X1 U19631 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18299) );
  AOI22_X1 U19632 ( .A1(n16593), .A2(n16574), .B1(n18299), .B2(U215), .ZN(U256) );
  INV_X1 U19633 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U19634 ( .A1(n16593), .A2(n16575), .B1(n18306), .B2(U215), .ZN(U257) );
  OAI22_X1 U19635 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n20772), .ZN(n16576) );
  INV_X1 U19636 ( .A(n16576), .ZN(U258) );
  OAI22_X1 U19637 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16593), .ZN(n16577) );
  INV_X1 U19638 ( .A(n16577), .ZN(U259) );
  OAI22_X1 U19639 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n20772), .ZN(n16578) );
  INV_X1 U19640 ( .A(n16578), .ZN(U260) );
  INV_X1 U19641 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U19642 ( .A1(n20772), .A2(n16579), .B1(n17418), .B2(U215), .ZN(U261) );
  INV_X1 U19643 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n20812) );
  INV_X1 U19644 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n16580) );
  AOI22_X1 U19645 ( .A1(n20772), .A2(n20812), .B1(n16580), .B2(U215), .ZN(U262) );
  INV_X1 U19646 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U19647 ( .A1(n20772), .A2(n16581), .B1(n17410), .B2(U215), .ZN(U263) );
  OAI22_X1 U19648 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n20772), .ZN(n16582) );
  INV_X1 U19649 ( .A(n16582), .ZN(U264) );
  OAI22_X1 U19650 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n20772), .ZN(n16583) );
  INV_X1 U19651 ( .A(n16583), .ZN(U265) );
  OAI22_X1 U19652 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n20772), .ZN(n16584) );
  INV_X1 U19653 ( .A(n16584), .ZN(U266) );
  OAI22_X1 U19654 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20772), .ZN(n16585) );
  INV_X1 U19655 ( .A(n16585), .ZN(U267) );
  OAI22_X1 U19656 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20772), .ZN(n16586) );
  INV_X1 U19657 ( .A(n16586), .ZN(U268) );
  OAI22_X1 U19658 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20772), .ZN(n16587) );
  INV_X1 U19659 ( .A(n16587), .ZN(U269) );
  OAI22_X1 U19660 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16593), .ZN(n16588) );
  INV_X1 U19661 ( .A(n16588), .ZN(U270) );
  OAI22_X1 U19662 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16593), .ZN(n16589) );
  INV_X1 U19663 ( .A(n16589), .ZN(U271) );
  OAI22_X1 U19664 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16593), .ZN(n16590) );
  INV_X1 U19665 ( .A(n16590), .ZN(U272) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16593), .ZN(n16591) );
  INV_X1 U19667 ( .A(n16591), .ZN(U273) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16593), .ZN(n16592) );
  INV_X1 U19669 ( .A(n16592), .ZN(U275) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16593), .ZN(n16594) );
  INV_X1 U19671 ( .A(n16594), .ZN(U276) );
  OAI22_X1 U19672 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20772), .ZN(n16595) );
  INV_X1 U19673 ( .A(n16595), .ZN(U277) );
  OAI22_X1 U19674 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20772), .ZN(n16596) );
  INV_X1 U19675 ( .A(n16596), .ZN(U278) );
  OAI22_X1 U19676 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20772), .ZN(n16597) );
  INV_X1 U19677 ( .A(n16597), .ZN(U279) );
  OAI22_X1 U19678 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20772), .ZN(n16598) );
  INV_X1 U19679 ( .A(n16598), .ZN(U280) );
  OAI22_X1 U19680 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20772), .ZN(n16599) );
  INV_X1 U19681 ( .A(n16599), .ZN(U281) );
  AOI22_X1 U19682 ( .A1(n20772), .A2(n16601), .B1(n18312), .B2(U215), .ZN(U282) );
  INV_X1 U19683 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16600) );
  AOI222_X1 U19684 ( .A1(n16602), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16601), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16600), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16603) );
  INV_X2 U19685 ( .A(n16605), .ZN(n16604) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18820) );
  INV_X1 U19687 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19688 ( .A1(n16604), .A2(n18820), .B1(n19753), .B2(n16605), .ZN(
        U347) );
  INV_X1 U19689 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18818) );
  INV_X1 U19690 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19691 ( .A1(n16604), .A2(n18818), .B1(n19752), .B2(n16605), .ZN(
        U348) );
  INV_X1 U19692 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18815) );
  INV_X1 U19693 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19694 ( .A1(n16604), .A2(n18815), .B1(n19751), .B2(n16605), .ZN(
        U349) );
  INV_X1 U19695 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18814) );
  INV_X1 U19696 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19697 ( .A1(n16604), .A2(n18814), .B1(n19750), .B2(n16605), .ZN(
        U350) );
  INV_X1 U19698 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18812) );
  INV_X1 U19699 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19700 ( .A1(n16604), .A2(n18812), .B1(n19749), .B2(n16605), .ZN(
        U351) );
  INV_X1 U19701 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18810) );
  INV_X1 U19702 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19703 ( .A1(n16604), .A2(n18810), .B1(n19748), .B2(n16605), .ZN(
        U352) );
  INV_X1 U19704 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18808) );
  INV_X1 U19705 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19706 ( .A1(n16604), .A2(n18808), .B1(n19747), .B2(n16605), .ZN(
        U353) );
  INV_X1 U19707 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18806) );
  AOI22_X1 U19708 ( .A1(n16604), .A2(n18806), .B1(n19744), .B2(n16605), .ZN(
        U354) );
  INV_X1 U19709 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18859) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19711 ( .A1(n16604), .A2(n18859), .B1(n19788), .B2(n16605), .ZN(
        U355) );
  INV_X1 U19712 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18856) );
  INV_X1 U19713 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19714 ( .A1(n16604), .A2(n18856), .B1(n19785), .B2(n16605), .ZN(
        U356) );
  INV_X1 U19715 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18853) );
  INV_X1 U19716 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19717 ( .A1(n16604), .A2(n18853), .B1(n19784), .B2(n16605), .ZN(
        U357) );
  INV_X1 U19718 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18852) );
  INV_X1 U19719 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19720 ( .A1(n16604), .A2(n18852), .B1(n19781), .B2(n16605), .ZN(
        U358) );
  INV_X1 U19721 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18850) );
  INV_X1 U19722 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19723 ( .A1(n16604), .A2(n18850), .B1(n19780), .B2(n16605), .ZN(
        U359) );
  INV_X1 U19724 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18848) );
  INV_X1 U19725 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19726 ( .A1(n16604), .A2(n18848), .B1(n19778), .B2(n16605), .ZN(
        U360) );
  INV_X1 U19727 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18846) );
  INV_X1 U19728 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19776) );
  AOI22_X1 U19729 ( .A1(n16604), .A2(n18846), .B1(n19776), .B2(n16605), .ZN(
        U361) );
  INV_X1 U19730 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18843) );
  INV_X1 U19731 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19732 ( .A1(n16604), .A2(n18843), .B1(n19774), .B2(n16605), .ZN(
        U362) );
  INV_X1 U19733 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18842) );
  INV_X1 U19734 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U19735 ( .A1(n16604), .A2(n18842), .B1(n20846), .B2(n16605), .ZN(
        U363) );
  INV_X1 U19736 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18840) );
  INV_X1 U19737 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19738 ( .A1(n16604), .A2(n18840), .B1(n19771), .B2(n16605), .ZN(
        U364) );
  INV_X1 U19739 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18804) );
  INV_X1 U19740 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19741 ( .A1(n16604), .A2(n18804), .B1(n19742), .B2(n16605), .ZN(
        U365) );
  INV_X1 U19742 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18839) );
  INV_X1 U19743 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19744 ( .A1(n16604), .A2(n18839), .B1(n19769), .B2(n16605), .ZN(
        U366) );
  INV_X1 U19745 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18837) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19747 ( .A1(n16604), .A2(n18837), .B1(n19767), .B2(n16605), .ZN(
        U367) );
  INV_X1 U19748 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18835) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19750 ( .A1(n16604), .A2(n18835), .B1(n19765), .B2(n16605), .ZN(
        U368) );
  INV_X1 U19751 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18832) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U19753 ( .A1(n16604), .A2(n18832), .B1(n19763), .B2(n16605), .ZN(
        U369) );
  INV_X1 U19754 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18831) );
  INV_X1 U19755 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19756 ( .A1(n16604), .A2(n18831), .B1(n19762), .B2(n16605), .ZN(
        U370) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18829) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U19759 ( .A1(n16604), .A2(n18829), .B1(n19760), .B2(n16605), .ZN(
        U371) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18826) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U19762 ( .A1(n16604), .A2(n18826), .B1(n19758), .B2(n16605), .ZN(
        U372) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18825) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U19765 ( .A1(n16604), .A2(n18825), .B1(n19757), .B2(n16605), .ZN(
        U373) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18824) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19756) );
  AOI22_X1 U19768 ( .A1(n16604), .A2(n18824), .B1(n19756), .B2(n16605), .ZN(
        U374) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18822) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19771 ( .A1(n16604), .A2(n18822), .B1(n19754), .B2(n16605), .ZN(
        U375) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18802) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19774 ( .A1(n16604), .A2(n18802), .B1(n19741), .B2(n16605), .ZN(
        U376) );
  INV_X1 U19775 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18801) );
  NAND2_X1 U19776 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18801), .ZN(n18790) );
  AOI21_X1 U19777 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n18790), .A(n18935), 
        .ZN(n18869) );
  AOI21_X1 U19778 ( .B1(P3_ADS_N_REG_SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), 
        .A(n18869), .ZN(n16606) );
  INV_X1 U19779 ( .A(n16606), .ZN(P3_U2633) );
  INV_X1 U19780 ( .A(n18778), .ZN(n16609) );
  OAI21_X1 U19781 ( .B1(n16616), .B2(n16607), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16608) );
  OAI21_X1 U19782 ( .B1(n16610), .B2(n16609), .A(n16608), .ZN(P3_U2634) );
  AOI21_X1 U19783 ( .B1(n18799), .B2(n18801), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16611) );
  AOI22_X1 U19784 ( .A1(n18935), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16611), 
        .B2(n18936), .ZN(P3_U2635) );
  NOR2_X1 U19785 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18786) );
  OAI21_X1 U19786 ( .B1(n18786), .B2(BS16), .A(n18869), .ZN(n18867) );
  OAI21_X1 U19787 ( .B1(n18869), .B2(n16612), .A(n18867), .ZN(P3_U2636) );
  INV_X1 U19788 ( .A(n16613), .ZN(n16615) );
  NOR3_X1 U19789 ( .A1(n16616), .A2(n16615), .A3(n16614), .ZN(n18713) );
  NOR2_X1 U19790 ( .A1(n18713), .A2(n18773), .ZN(n18917) );
  OAI21_X1 U19791 ( .B1(n18917), .B2(n16618), .A(n16617), .ZN(P3_U2637) );
  NOR4_X1 U19792 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16622) );
  NOR4_X1 U19793 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16621) );
  NOR4_X1 U19794 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16620) );
  NOR4_X1 U19795 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_23__SCAN_IN), .A3(P3_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n16619) );
  NAND4_X1 U19796 ( .A1(n16622), .A2(n16621), .A3(n16620), .A4(n16619), .ZN(
        n16628) );
  NOR4_X1 U19797 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16626) );
  INV_X1 U19798 ( .A(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20809) );
  INV_X1 U19799 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20859) );
  NAND2_X1 U19800 ( .A1(n20809), .A2(n20859), .ZN(n20759) );
  AOI21_X1 U19801 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(n20759), .ZN(n16625) );
  NOR4_X1 U19802 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16624) );
  NOR4_X1 U19803 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16623) );
  NAND4_X1 U19804 ( .A1(n16626), .A2(n16625), .A3(n16624), .A4(n16623), .ZN(
        n16627) );
  NOR2_X1 U19805 ( .A1(n16628), .A2(n16627), .ZN(n18911) );
  INV_X1 U19806 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16630) );
  NOR3_X1 U19807 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16631) );
  OAI21_X1 U19808 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16631), .A(n18911), .ZN(
        n16629) );
  OAI21_X1 U19809 ( .B1(n18911), .B2(n16630), .A(n16629), .ZN(P3_U2638) );
  INV_X1 U19810 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18907) );
  INV_X1 U19811 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18868) );
  AOI21_X1 U19812 ( .B1(n18907), .B2(n18868), .A(n16631), .ZN(n16633) );
  INV_X1 U19813 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16632) );
  INV_X1 U19814 ( .A(n18911), .ZN(n18914) );
  AOI22_X1 U19815 ( .A1(n18911), .A2(n16633), .B1(n16632), .B2(n18914), .ZN(
        P3_U2639) );
  INV_X1 U19816 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18860) );
  INV_X1 U19817 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18845) );
  INV_X1 U19818 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18844) );
  NAND3_X1 U19819 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16634), .A3(
        P3_REIP_REG_22__SCAN_IN), .ZN(n16736) );
  NOR2_X1 U19820 ( .A1(n18844), .A2(n16736), .ZN(n16710) );
  NAND2_X1 U19821 ( .A1(n16635), .A2(n16710), .ZN(n16725) );
  NOR2_X1 U19822 ( .A1(n18845), .A2(n16725), .ZN(n16648) );
  NAND2_X1 U19823 ( .A1(n16971), .A2(n16648), .ZN(n16711) );
  NAND2_X1 U19824 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16646) );
  NOR2_X1 U19825 ( .A1(n16711), .A2(n16646), .ZN(n16686) );
  NAND4_X1 U19826 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16686), .ZN(n16650) );
  NOR3_X1 U19827 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18860), .A3(n16650), 
        .ZN(n16636) );
  AOI21_X1 U19828 ( .B1(n16976), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16636), .ZN(
        n16653) );
  INV_X1 U19829 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17094) );
  NAND2_X1 U19830 ( .A1(n16751), .A2(n17094), .ZN(n16750) );
  INV_X1 U19831 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20806) );
  NAND2_X1 U19832 ( .A1(n16738), .A2(n20806), .ZN(n16733) );
  NOR2_X1 U19833 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16733), .ZN(n16706) );
  INV_X1 U19834 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17005) );
  NAND2_X1 U19835 ( .A1(n16706), .A2(n17005), .ZN(n16699) );
  NOR2_X1 U19836 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16699), .ZN(n16698) );
  NAND2_X1 U19837 ( .A1(n16698), .A2(n16692), .ZN(n16691) );
  NOR2_X1 U19838 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16691), .ZN(n16677) );
  INV_X1 U19839 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16673) );
  NAND2_X1 U19840 ( .A1(n16677), .A2(n16673), .ZN(n16655) );
  NOR2_X1 U19841 ( .A1(n16995), .A2(n16655), .ZN(n16661) );
  INV_X1 U19842 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17034) );
  INV_X1 U19843 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20814) );
  NAND3_X1 U19844 ( .A1(n17610), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16642) );
  NOR2_X1 U19845 ( .A1(n17615), .A2(n16642), .ZN(n17569) );
  INV_X1 U19846 ( .A(n17569), .ZN(n16640) );
  NOR2_X1 U19847 ( .A1(n20814), .A2(n16640), .ZN(n16639) );
  NAND2_X1 U19848 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16639), .ZN(
        n16638) );
  AOI21_X1 U19849 ( .B1(n17572), .B2(n16638), .A(n16637), .ZN(n17574) );
  OAI21_X1 U19850 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16639), .A(
        n16638), .ZN(n17589) );
  INV_X1 U19851 ( .A(n17589), .ZN(n16688) );
  AOI21_X1 U19852 ( .B1(n20814), .B2(n16640), .A(n16639), .ZN(n17600) );
  INV_X1 U19853 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17630) );
  NOR2_X1 U19854 ( .A1(n17630), .A2(n16642), .ZN(n16641) );
  OAI21_X1 U19855 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16641), .A(
        n16640), .ZN(n17618) );
  INV_X1 U19856 ( .A(n17618), .ZN(n16709) );
  AOI21_X1 U19857 ( .B1(n17630), .B2(n16642), .A(n16641), .ZN(n17627) );
  INV_X1 U19858 ( .A(n17610), .ZN(n17598) );
  NOR2_X1 U19859 ( .A1(n17598), .A2(n17927), .ZN(n17611) );
  OAI21_X1 U19860 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17611), .A(
        n16642), .ZN(n17648) );
  INV_X1 U19861 ( .A(n17648), .ZN(n16728) );
  INV_X1 U19862 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17658) );
  NAND2_X1 U19863 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16644), .ZN(
        n16643) );
  AOI21_X1 U19864 ( .B1(n17658), .B2(n16643), .A(n17611), .ZN(n17660) );
  INV_X1 U19865 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17676) );
  XNOR2_X1 U19866 ( .A(n17676), .B(n16644), .ZN(n17679) );
  NOR2_X1 U19867 ( .A1(n16645), .A2(n9694), .ZN(n16749) );
  NOR2_X1 U19868 ( .A1(n17679), .A2(n16749), .ZN(n16748) );
  NOR2_X1 U19869 ( .A1(n16748), .A2(n9694), .ZN(n16742) );
  NOR2_X1 U19870 ( .A1(n17660), .A2(n16742), .ZN(n16741) );
  NOR2_X1 U19871 ( .A1(n16741), .A2(n9694), .ZN(n16727) );
  NOR2_X1 U19872 ( .A1(n16728), .A2(n16727), .ZN(n16726) );
  NOR2_X1 U19873 ( .A1(n16726), .A2(n9694), .ZN(n16719) );
  NOR2_X1 U19874 ( .A1(n17627), .A2(n16719), .ZN(n16718) );
  NOR2_X1 U19875 ( .A1(n16718), .A2(n9694), .ZN(n16708) );
  NOR2_X1 U19876 ( .A1(n16709), .A2(n16708), .ZN(n16707) );
  NOR2_X1 U19877 ( .A1(n16687), .A2(n9694), .ZN(n16679) );
  NOR2_X1 U19878 ( .A1(n17574), .A2(n16679), .ZN(n16678) );
  NOR2_X1 U19879 ( .A1(n16678), .A2(n9694), .ZN(n16665) );
  NOR2_X1 U19880 ( .A1(n16666), .A2(n16665), .ZN(n16664) );
  NOR2_X1 U19881 ( .A1(n9694), .A2(n18781), .ZN(n16977) );
  INV_X1 U19882 ( .A(n16977), .ZN(n16818) );
  NAND3_X1 U19883 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16649) );
  INV_X1 U19884 ( .A(n16646), .ZN(n16647) );
  OAI221_X1 U19885 ( .B1(n16989), .B2(n16648), .C1(n16989), .C2(n16647), .A(
        n16999), .ZN(n16703) );
  AOI21_X1 U19886 ( .B1(n16971), .B2(n16649), .A(n16703), .ZN(n16676) );
  NOR2_X1 U19887 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16650), .ZN(n16659) );
  INV_X1 U19888 ( .A(n16659), .ZN(n16651) );
  AOI21_X1 U19889 ( .B1(n16676), .B2(n16651), .A(n18858), .ZN(n16652) );
  NAND2_X1 U19890 ( .A1(n16965), .A2(n16655), .ZN(n16671) );
  XOR2_X1 U19891 ( .A(n16657), .B(n16656), .Z(n16660) );
  OAI22_X1 U19892 ( .A1(n16676), .A2(n18860), .B1(n10061), .B2(n16987), .ZN(
        n16658) );
  AOI211_X1 U19893 ( .C1(n16660), .C2(n16951), .A(n16659), .B(n16658), .ZN(
        n16663) );
  OAI21_X1 U19894 ( .B1(n16976), .B2(n16661), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16662) );
  OAI211_X1 U19895 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16671), .A(n16663), .B(
        n16662), .ZN(P3_U2641) );
  INV_X1 U19896 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18855) );
  AOI211_X1 U19897 ( .C1(n16666), .C2(n16665), .A(n16664), .B(n18781), .ZN(
        n16670) );
  NAND3_X1 U19898 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16686), .ZN(n16668) );
  OAI22_X1 U19899 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16668), .B1(n16667), 
        .B2(n16987), .ZN(n16669) );
  AOI211_X1 U19900 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16976), .A(n16670), .B(
        n16669), .ZN(n16675) );
  INV_X1 U19901 ( .A(n16671), .ZN(n16672) );
  OAI21_X1 U19902 ( .B1(n16677), .B2(n16673), .A(n16672), .ZN(n16674) );
  OAI211_X1 U19903 ( .C1(n16676), .C2(n18855), .A(n16675), .B(n16674), .ZN(
        P3_U2642) );
  AOI22_X1 U19904 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16963), .B1(
        n16976), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16685) );
  AOI211_X1 U19905 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16691), .A(n16677), .B(
        n16995), .ZN(n16681) );
  AOI211_X1 U19906 ( .C1(n17574), .C2(n16679), .A(n16678), .B(n18781), .ZN(
        n16680) );
  AOI211_X1 U19907 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16703), .A(n16681), 
        .B(n16680), .ZN(n16684) );
  NAND2_X1 U19908 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16682) );
  OAI211_X1 U19909 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16686), .B(n16682), .ZN(n16683) );
  NAND3_X1 U19910 ( .A1(n16685), .A2(n16684), .A3(n16683), .ZN(P3_U2643) );
  INV_X1 U19911 ( .A(n16686), .ZN(n16695) );
  AOI211_X1 U19912 ( .C1(n16688), .C2(n9699), .A(n16687), .B(n18781), .ZN(
        n16690) );
  OAI22_X1 U19913 ( .A1(n17592), .A2(n16987), .B1(n16996), .B2(n16692), .ZN(
        n16689) );
  AOI211_X1 U19914 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16703), .A(n16690), 
        .B(n16689), .ZN(n16694) );
  OAI211_X1 U19915 ( .C1(n16698), .C2(n16692), .A(n16965), .B(n16691), .ZN(
        n16693) );
  OAI211_X1 U19916 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16695), .A(n16694), 
        .B(n16693), .ZN(P3_U2644) );
  AOI22_X1 U19917 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16963), .B1(
        n16976), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16705) );
  INV_X1 U19918 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18847) );
  INV_X1 U19919 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18849) );
  OAI21_X1 U19920 ( .B1(n18847), .B2(n16711), .A(n18849), .ZN(n16702) );
  AOI211_X1 U19921 ( .C1(n17600), .C2(n16697), .A(n16696), .B(n18781), .ZN(
        n16701) );
  AOI211_X1 U19922 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16699), .A(n16698), .B(
        n16995), .ZN(n16700) );
  AOI211_X1 U19923 ( .C1(n16703), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        n16704) );
  NAND2_X1 U19924 ( .A1(n16705), .A2(n16704), .ZN(P3_U2645) );
  OR2_X1 U19925 ( .A1(n16995), .A2(n16706), .ZN(n16717) );
  AOI21_X1 U19926 ( .B1(n16965), .B2(n16706), .A(n16976), .ZN(n16716) );
  AOI211_X1 U19927 ( .C1(n16709), .C2(n16708), .A(n16707), .B(n18781), .ZN(
        n16714) );
  AOI21_X1 U19928 ( .B1(n16710), .B2(n16759), .A(n16758), .ZN(n16732) );
  AOI21_X1 U19929 ( .B1(n16971), .B2(n18845), .A(n16732), .ZN(n16712) );
  AOI22_X1 U19930 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16712), .B1(n16711), 
        .B2(n18847), .ZN(n16713) );
  AOI211_X1 U19931 ( .C1(n16963), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16714), .B(n16713), .ZN(n16715) );
  OAI221_X1 U19932 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16717), .C1(n17005), 
        .C2(n16716), .A(n16715), .ZN(P3_U2646) );
  NAND2_X1 U19933 ( .A1(n16971), .A2(n18845), .ZN(n16724) );
  AOI22_X1 U19934 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16963), .B1(
        n16976), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16723) );
  AOI21_X1 U19935 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16733), .A(n16717), .ZN(
        n16721) );
  AOI211_X1 U19936 ( .C1(n17627), .C2(n16719), .A(n16718), .B(n18781), .ZN(
        n16720) );
  AOI211_X1 U19937 ( .C1(n16732), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16721), 
        .B(n16720), .ZN(n16722) );
  OAI211_X1 U19938 ( .C1(n16725), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        P3_U2647) );
  NAND2_X1 U19939 ( .A1(n16786), .A2(n18844), .ZN(n16737) );
  AOI211_X1 U19940 ( .C1(n16728), .C2(n16727), .A(n16726), .B(n18781), .ZN(
        n16731) );
  OAI22_X1 U19941 ( .A1(n16729), .A2(n16987), .B1(n16996), .B2(n20806), .ZN(
        n16730) );
  AOI211_X1 U19942 ( .C1(n16732), .C2(P3_REIP_REG_23__SCAN_IN), .A(n16731), 
        .B(n16730), .ZN(n16735) );
  OAI211_X1 U19943 ( .C1(n16738), .C2(n20806), .A(n16965), .B(n16733), .ZN(
        n16734) );
  OAI211_X1 U19944 ( .C1(n16737), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P3_U2648) );
  AOI211_X1 U19945 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16750), .A(n16738), .B(
        n16995), .ZN(n16739) );
  AOI21_X1 U19946 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16976), .A(n16739), .ZN(
        n16746) );
  INV_X1 U19947 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20827) );
  INV_X1 U19948 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18841) );
  NAND2_X1 U19949 ( .A1(n16740), .A2(n16778), .ZN(n16757) );
  AOI221_X1 U19950 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n20827), .C2(n18841), .A(n16757), .ZN(n16744) );
  AOI211_X1 U19951 ( .C1(n17660), .C2(n16742), .A(n16741), .B(n18781), .ZN(
        n16743) );
  AOI211_X1 U19952 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16747), .A(n16744), 
        .B(n16743), .ZN(n16745) );
  OAI211_X1 U19953 ( .C1(n17658), .C2(n16987), .A(n16746), .B(n16745), .ZN(
        P3_U2649) );
  INV_X1 U19954 ( .A(n16747), .ZN(n16756) );
  AOI211_X1 U19955 ( .C1(n17679), .C2(n16749), .A(n16748), .B(n18781), .ZN(
        n16754) );
  OAI211_X1 U19956 ( .C1(n16751), .C2(n17094), .A(n16965), .B(n16750), .ZN(
        n16752) );
  OAI21_X1 U19957 ( .B1(n17094), .B2(n16996), .A(n16752), .ZN(n16753) );
  AOI211_X1 U19958 ( .C1(n16963), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16754), .B(n16753), .ZN(n16755) );
  OAI221_X1 U19959 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16757), .C1(n20827), 
        .C2(n16756), .A(n16755), .ZN(P3_U2650) );
  AOI21_X1 U19960 ( .B1(n16760), .B2(n16759), .A(n16758), .ZN(n16789) );
  AOI21_X1 U19961 ( .B1(n16778), .B2(n18834), .A(n16789), .ZN(n16770) );
  INV_X1 U19962 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17713) );
  INV_X1 U19963 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16796) );
  NOR2_X1 U19964 ( .A1(n16796), .A2(n16805), .ZN(n16782) );
  NAND2_X1 U19965 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16782), .ZN(
        n16781) );
  NOR2_X1 U19966 ( .A1(n17713), .A2(n16781), .ZN(n16761) );
  OAI21_X1 U19967 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16761), .A(
        n17653), .ZN(n17703) );
  INV_X1 U19968 ( .A(n16781), .ZN(n17699) );
  NAND2_X1 U19969 ( .A1(n16800), .A2(n17699), .ZN(n16774) );
  OAI21_X1 U19970 ( .B1(n17713), .B2(n16774), .A(n16986), .ZN(n16763) );
  OAI21_X1 U19971 ( .B1(n17703), .B2(n16763), .A(n16951), .ZN(n16762) );
  AOI21_X1 U19972 ( .B1(n17703), .B2(n16763), .A(n16762), .ZN(n16768) );
  OAI211_X1 U19973 ( .C1(n16772), .C2(n16766), .A(n16965), .B(n16764), .ZN(
        n16765) );
  OAI211_X1 U19974 ( .C1(n16996), .C2(n16766), .A(n18181), .B(n16765), .ZN(
        n16767) );
  AOI211_X1 U19975 ( .C1(n16963), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16768), .B(n16767), .ZN(n16769) );
  OAI221_X1 U19976 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n16771), .C1(n18836), 
        .C2(n16770), .A(n16769), .ZN(P3_U2652) );
  AOI211_X1 U19977 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16790), .A(n16772), .B(
        n16995), .ZN(n16773) );
  AOI211_X1 U19978 ( .C1(n16976), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9593), .B(
        n16773), .ZN(n16780) );
  AOI22_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16781), .B1(
        n17699), .B2(n17713), .ZN(n17710) );
  NAND2_X1 U19980 ( .A1(n16986), .A2(n16774), .ZN(n16776) );
  OAI21_X1 U19981 ( .B1(n17710), .B2(n16776), .A(n16951), .ZN(n16775) );
  AOI21_X1 U19982 ( .B1(n17710), .B2(n16776), .A(n16775), .ZN(n16777) );
  AOI221_X1 U19983 ( .B1(n16789), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16778), 
        .C2(n18834), .A(n16777), .ZN(n16779) );
  OAI211_X1 U19984 ( .C1(n17713), .C2(n16987), .A(n16780), .B(n16779), .ZN(
        P3_U2653) );
  AOI22_X1 U19985 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16963), .B1(
        n16976), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16794) );
  OAI21_X1 U19986 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16782), .A(
        n16781), .ZN(n17721) );
  AOI21_X1 U19987 ( .B1(n16796), .B2(n16805), .A(n16782), .ZN(n16783) );
  INV_X1 U19988 ( .A(n16783), .ZN(n17737) );
  OAI21_X1 U19989 ( .B1(n16800), .B2(n9694), .A(n17737), .ZN(n16801) );
  NAND2_X1 U19990 ( .A1(n16986), .A2(n16801), .ZN(n16785) );
  OAI21_X1 U19991 ( .B1(n17721), .B2(n16785), .A(n16951), .ZN(n16784) );
  AOI21_X1 U19992 ( .B1(n17721), .B2(n16785), .A(n16784), .ZN(n16788) );
  INV_X1 U19993 ( .A(n16786), .ZN(n16807) );
  NOR4_X1 U19994 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18830), .A3(n18828), 
        .A4(n16807), .ZN(n16787) );
  AOI211_X1 U19995 ( .C1(n16789), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16788), 
        .B(n16787), .ZN(n16793) );
  OAI211_X1 U19996 ( .C1(n16795), .C2(n16791), .A(n16965), .B(n16790), .ZN(
        n16792) );
  NAND4_X1 U19997 ( .A1(n16794), .A2(n16793), .A3(n18181), .A4(n16792), .ZN(
        P3_U2654) );
  OAI21_X1 U19998 ( .B1(n18828), .B2(n16822), .A(n16997), .ZN(n16806) );
  NOR3_X1 U19999 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18828), .A3(n16807), 
        .ZN(n16799) );
  AOI211_X1 U20000 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16810), .A(n16795), .B(
        n16995), .ZN(n16798) );
  OAI22_X1 U20001 ( .A1(n16796), .A2(n16987), .B1(n16996), .B2(n17162), .ZN(
        n16797) );
  NOR4_X1 U20002 ( .A1(n9593), .A2(n16799), .A3(n16798), .A4(n16797), .ZN(
        n16803) );
  OR2_X1 U20003 ( .A1(n9694), .A2(n16800), .ZN(n16804) );
  OAI211_X1 U20004 ( .C1(n17737), .C2(n16804), .A(n16951), .B(n16801), .ZN(
        n16802) );
  OAI211_X1 U20005 ( .C1(n18830), .C2(n16806), .A(n16803), .B(n16802), .ZN(
        P3_U2655) );
  AOI22_X1 U20006 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16963), .B1(
        n16976), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16816) );
  NOR2_X1 U20007 ( .A1(n18781), .A2(n16804), .ZN(n16809) );
  OAI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17732), .A(
        n16805), .ZN(n17742) );
  AOI21_X1 U20009 ( .B1(n18828), .B2(n16807), .A(n16806), .ZN(n16808) );
  AOI211_X1 U20010 ( .C1(n16809), .C2(n17742), .A(n9593), .B(n16808), .ZN(
        n16815) );
  OAI211_X1 U20011 ( .C1(n16817), .C2(n16811), .A(n16965), .B(n16810), .ZN(
        n16814) );
  INV_X1 U20012 ( .A(n17742), .ZN(n16812) );
  AOI21_X1 U20013 ( .B1(n16986), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18781), .ZN(n16992) );
  OAI211_X1 U20014 ( .C1(n17732), .C2(n9694), .A(n16812), .B(n16992), .ZN(
        n16813) );
  NAND4_X1 U20015 ( .A1(n16816), .A2(n16815), .A3(n16814), .A4(n16813), .ZN(
        P3_U2656) );
  INV_X1 U20016 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17190) );
  AOI211_X1 U20017 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16840), .A(n16817), .B(
        n16995), .ZN(n16827) );
  AOI21_X1 U20018 ( .B1(n10043), .B2(n16820), .A(n17732), .ZN(n17762) );
  NOR2_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17927), .ZN(
        n16979) );
  AOI21_X1 U20020 ( .B1(n17758), .B2(n16979), .A(n16818), .ZN(n16819) );
  INV_X1 U20021 ( .A(n16819), .ZN(n16832) );
  INV_X1 U20022 ( .A(n16820), .ZN(n16831) );
  OAI211_X1 U20023 ( .C1(n16831), .C2(n9694), .A(n17762), .B(n16992), .ZN(
        n16825) );
  NOR2_X1 U20024 ( .A1(n16989), .A2(n16821), .ZN(n16823) );
  OAI211_X1 U20025 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n16823), .A(n16822), 
        .B(n16997), .ZN(n16824) );
  OAI211_X1 U20026 ( .C1(n17762), .C2(n16832), .A(n16825), .B(n16824), .ZN(
        n16826) );
  AOI211_X1 U20027 ( .C1(n16963), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16827), .B(n16826), .ZN(n16828) );
  OAI211_X1 U20028 ( .C1(n16996), .C2(n17190), .A(n16828), .B(n18181), .ZN(
        P3_U2657) );
  NAND3_X1 U20029 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n16830) );
  NAND2_X1 U20030 ( .A1(n16829), .A2(n16999), .ZN(n16870) );
  OAI21_X1 U20031 ( .B1(n16830), .B2(n16870), .A(n16997), .ZN(n16859) );
  OAI21_X1 U20032 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16989), .A(n16859), 
        .ZN(n16839) );
  NAND2_X1 U20033 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17770), .ZN(
        n16847) );
  AOI21_X1 U20034 ( .B1(n16844), .B2(n16847), .A(n16831), .ZN(n17771) );
  OAI22_X1 U20035 ( .A1(n17771), .A2(n16832), .B1(n16996), .B2(n16841), .ZN(
        n16838) );
  NAND2_X1 U20036 ( .A1(n16971), .A2(n16833), .ZN(n16836) );
  INV_X1 U20037 ( .A(n16847), .ZN(n16834) );
  OAI211_X1 U20038 ( .C1(n16834), .C2(n9694), .A(n17771), .B(n16992), .ZN(
        n16835) );
  OAI211_X1 U20039 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16836), .A(n18181), 
        .B(n16835), .ZN(n16837) );
  AOI211_X1 U20040 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16839), .A(n16838), 
        .B(n16837), .ZN(n16843) );
  OAI211_X1 U20041 ( .C1(n16845), .C2(n16841), .A(n16965), .B(n16840), .ZN(
        n16842) );
  OAI211_X1 U20042 ( .C1(n16987), .C2(n16844), .A(n16843), .B(n16842), .ZN(
        P3_U2658) );
  AOI211_X1 U20043 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16862), .A(n16845), .B(
        n16995), .ZN(n16846) );
  AOI21_X1 U20044 ( .B1(n16963), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16846), .ZN(n16855) );
  OAI21_X1 U20045 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17770), .A(
        n16847), .ZN(n17796) );
  INV_X1 U20046 ( .A(n16979), .ZN(n16978) );
  OAI21_X1 U20047 ( .B1(n17776), .B2(n16978), .A(n16986), .ZN(n16848) );
  XOR2_X1 U20048 ( .A(n17796), .B(n16848), .Z(n16853) );
  NAND2_X1 U20049 ( .A1(n16971), .A2(n18823), .ZN(n16849) );
  OAI22_X1 U20050 ( .A1(n16996), .A2(n16851), .B1(n16850), .B2(n16849), .ZN(
        n16852) );
  AOI211_X1 U20051 ( .C1(n16951), .C2(n16853), .A(n9593), .B(n16852), .ZN(
        n16854) );
  OAI211_X1 U20052 ( .C1(n18823), .C2(n16859), .A(n16855), .B(n16854), .ZN(
        P3_U2659) );
  INV_X1 U20053 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16866) );
  INV_X1 U20054 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18819) );
  INV_X1 U20055 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18817) );
  NOR2_X1 U20056 ( .A1(n18819), .A2(n18817), .ZN(n16856) );
  NOR3_X1 U20057 ( .A1(n16989), .A2(n18816), .A3(n16894), .ZN(n16877) );
  AOI21_X1 U20058 ( .B1(n16856), .B2(n16877), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16860) );
  INV_X1 U20059 ( .A(n16867), .ZN(n17798) );
  NOR2_X1 U20060 ( .A1(n17833), .A2(n17927), .ZN(n16917) );
  NAND2_X1 U20061 ( .A1(n17798), .A2(n16917), .ZN(n16881) );
  INV_X1 U20062 ( .A(n16881), .ZN(n16869) );
  NAND2_X1 U20063 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16869), .ZN(
        n16868) );
  AOI21_X1 U20064 ( .B1(n16866), .B2(n16868), .A(n17770), .ZN(n17801) );
  AOI21_X1 U20065 ( .B1(n9724), .B2(n16979), .A(n9694), .ZN(n16857) );
  XNOR2_X1 U20066 ( .A(n17801), .B(n16857), .ZN(n16858) );
  OAI22_X1 U20067 ( .A1(n16860), .A2(n16859), .B1(n18781), .B2(n16858), .ZN(
        n16861) );
  AOI211_X1 U20068 ( .C1(n16976), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9593), .B(
        n16861), .ZN(n16865) );
  OAI211_X1 U20069 ( .C1(n16871), .C2(n16863), .A(n16965), .B(n16862), .ZN(
        n16864) );
  OAI211_X1 U20070 ( .C1(n16987), .C2(n16866), .A(n16865), .B(n16864), .ZN(
        P3_U2660) );
  OAI21_X1 U20071 ( .B1(n17833), .B2(n16978), .A(n16986), .ZN(n16918) );
  INV_X1 U20072 ( .A(n16918), .ZN(n16905) );
  AOI21_X1 U20073 ( .B1(n16986), .B2(n16867), .A(n16905), .ZN(n16885) );
  OAI21_X1 U20074 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16869), .A(
        n16868), .ZN(n17816) );
  XNOR2_X1 U20075 ( .A(n16885), .B(n17816), .ZN(n16880) );
  NAND2_X1 U20076 ( .A1(n16997), .A2(n16870), .ZN(n16898) );
  NAND2_X1 U20077 ( .A1(n16877), .A2(n18817), .ZN(n16883) );
  AOI21_X1 U20078 ( .B1(n16898), .B2(n16883), .A(n18819), .ZN(n16876) );
  AOI211_X1 U20079 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16872), .A(n16871), .B(
        n16995), .ZN(n16875) );
  INV_X1 U20080 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17234) );
  OAI22_X1 U20081 ( .A1(n16873), .A2(n16987), .B1(n16996), .B2(n17234), .ZN(
        n16874) );
  NOR4_X1 U20082 ( .A1(n9593), .A2(n16876), .A3(n16875), .A4(n16874), .ZN(
        n16879) );
  NAND3_X1 U20083 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16877), .A3(n18819), 
        .ZN(n16878) );
  OAI211_X1 U20084 ( .C1(n18781), .C2(n16880), .A(n16879), .B(n16878), .ZN(
        P3_U2661) );
  AND2_X1 U20085 ( .A1(n17831), .A2(n16917), .ZN(n16896) );
  OAI21_X1 U20086 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16896), .A(
        n16881), .ZN(n17820) );
  NOR2_X1 U20087 ( .A1(n18781), .A2(n16986), .ZN(n16943) );
  INV_X1 U20088 ( .A(n16943), .ZN(n16982) );
  NOR2_X1 U20089 ( .A1(n16886), .A2(n16995), .ZN(n16893) );
  AOI21_X1 U20090 ( .B1(n16893), .B2(n17233), .A(n9593), .ZN(n16891) );
  NOR2_X1 U20091 ( .A1(n17833), .A2(n16978), .ZN(n16882) );
  OAI221_X1 U20092 ( .B1(n17820), .B2(n17831), .C1(n17820), .C2(n16882), .A(
        n16951), .ZN(n16884) );
  OAI21_X1 U20093 ( .B1(n16885), .B2(n16884), .A(n16883), .ZN(n16889) );
  AOI21_X1 U20094 ( .B1(n16965), .B2(n16886), .A(n16976), .ZN(n16887) );
  OAI22_X1 U20095 ( .A1(n17233), .A2(n16887), .B1(n18817), .B2(n16898), .ZN(
        n16888) );
  AOI211_X1 U20096 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16963), .A(
        n16889), .B(n16888), .ZN(n16890) );
  OAI211_X1 U20097 ( .C1(n17820), .C2(n16982), .A(n16891), .B(n16890), .ZN(
        P3_U2662) );
  NAND2_X1 U20098 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16907), .ZN(n16892) );
  AOI22_X1 U20099 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16963), .B1(
        n16893), .B2(n16892), .ZN(n16903) );
  NOR2_X1 U20100 ( .A1(n16989), .A2(n16894), .ZN(n16895) );
  AOI22_X1 U20101 ( .A1(n16976), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n16895), .B2(
        n18816), .ZN(n16902) );
  INV_X1 U20102 ( .A(n17833), .ZN(n17830) );
  NAND3_X1 U20103 ( .A1(n17830), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16904) );
  AOI21_X1 U20104 ( .B1(n17835), .B2(n16904), .A(n16896), .ZN(n17838) );
  OAI21_X1 U20105 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16904), .A(
        n16986), .ZN(n16897) );
  XNOR2_X1 U20106 ( .A(n17838), .B(n16897), .ZN(n16900) );
  INV_X1 U20107 ( .A(n16898), .ZN(n16899) );
  AOI22_X1 U20108 ( .A1(n16951), .A2(n16900), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16899), .ZN(n16901) );
  NAND4_X1 U20109 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n18181), .ZN(
        P3_U2663) );
  AOI21_X1 U20110 ( .B1(n16971), .B2(n16916), .A(n16969), .ZN(n16933) );
  OAI21_X1 U20111 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16989), .A(n16933), .ZN(
        n16911) );
  OAI21_X1 U20112 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16917), .A(
        n16904), .ZN(n17855) );
  INV_X1 U20113 ( .A(n17855), .ZN(n16906) );
  AOI221_X1 U20114 ( .B1(n16906), .B2(n16905), .C1(n17855), .C2(n16918), .A(
        n18781), .ZN(n16910) );
  OAI211_X1 U20115 ( .C1(n16915), .C2(n20874), .A(n16965), .B(n16907), .ZN(
        n16908) );
  OAI211_X1 U20116 ( .C1(n16996), .C2(n20874), .A(n18181), .B(n16908), .ZN(
        n16909) );
  AOI211_X1 U20117 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16911), .A(n16910), .B(
        n16909), .ZN(n16914) );
  INV_X1 U20118 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18813) );
  NAND3_X1 U20119 ( .A1(n16971), .A2(n16912), .A3(n18813), .ZN(n16913) );
  OAI211_X1 U20120 ( .C1(n16987), .C2(n17847), .A(n16914), .B(n16913), .ZN(
        P3_U2664) );
  AOI211_X1 U20121 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16936), .A(n16915), .B(
        n16995), .ZN(n16926) );
  INV_X1 U20122 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16924) );
  INV_X1 U20123 ( .A(n16916), .ZN(n16929) );
  NOR2_X1 U20124 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16989), .ZN(n16920) );
  NAND2_X1 U20125 ( .A1(n17876), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16928) );
  AOI21_X1 U20126 ( .B1(n16924), .B2(n16928), .A(n16917), .ZN(n17857) );
  NOR3_X1 U20127 ( .A1(n17857), .A2(n18781), .A3(n16918), .ZN(n16919) );
  AOI211_X1 U20128 ( .C1(n16929), .C2(n16920), .A(n9593), .B(n16919), .ZN(
        n16923) );
  OAI211_X1 U20129 ( .C1(n16924), .C2(n9694), .A(n17857), .B(n16992), .ZN(
        n16922) );
  OAI211_X1 U20130 ( .C1(n16987), .C2(n16924), .A(n16923), .B(n16922), .ZN(
        n16925) );
  AOI211_X1 U20131 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16976), .A(n16926), .B(
        n16925), .ZN(n16927) );
  OAI21_X1 U20132 ( .B1(n16933), .B2(n18811), .A(n16927), .ZN(P3_U2665) );
  NOR2_X1 U20133 ( .A1(n17874), .A2(n17927), .ZN(n16939) );
  OAI21_X1 U20134 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16939), .A(
        n16928), .ZN(n17881) );
  OAI21_X1 U20135 ( .B1(n17874), .B2(n16978), .A(n16986), .ZN(n16945) );
  XOR2_X1 U20136 ( .A(n17881), .B(n16945), .Z(n16935) );
  INV_X1 U20137 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18809) );
  NOR2_X1 U20138 ( .A1(n16929), .A2(n16989), .ZN(n16930) );
  AOI22_X1 U20139 ( .A1(n16976), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n16931), .B2(
        n16930), .ZN(n16932) );
  OAI211_X1 U20140 ( .C1(n16933), .C2(n18809), .A(n16932), .B(n18181), .ZN(
        n16934) );
  AOI21_X1 U20141 ( .B1(n16951), .B2(n16935), .A(n16934), .ZN(n16938) );
  OAI211_X1 U20142 ( .C1(n16946), .C2(n17281), .A(n16965), .B(n16936), .ZN(
        n16937) );
  OAI211_X1 U20143 ( .C1(n16987), .C2(n17875), .A(n16938), .B(n16937), .ZN(
        P3_U2666) );
  AOI21_X1 U20144 ( .B1(n16971), .B2(n16954), .A(n16969), .ZN(n16960) );
  INV_X1 U20145 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16944) );
  NAND2_X1 U20146 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16956) );
  AOI21_X1 U20147 ( .B1(n16944), .B2(n16956), .A(n16939), .ZN(n17893) );
  NOR3_X1 U20148 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16989), .A3(n16954), .ZN(
        n16942) );
  OAI22_X1 U20149 ( .A1(n16944), .A2(n16987), .B1(n16996), .B2(n16940), .ZN(
        n16941) );
  AOI211_X1 U20150 ( .C1(n16943), .C2(n17893), .A(n16942), .B(n16941), .ZN(
        n16953) );
  NAND2_X1 U20151 ( .A1(n17892), .A2(n16944), .ZN(n17889) );
  OAI22_X1 U20152 ( .A1(n17893), .A2(n16945), .B1(n16978), .B2(n17889), .ZN(
        n16950) );
  AOI211_X1 U20153 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16964), .A(n16946), .B(
        n16995), .ZN(n16949) );
  NOR2_X1 U20154 ( .A1(n17462), .A2(n16947), .ZN(n18943) );
  INV_X1 U20155 ( .A(n18943), .ZN(n17002) );
  OAI221_X1 U20156 ( .B1(n17002), .B2(n17178), .C1(n17002), .C2(n18716), .A(
        n18181), .ZN(n16948) );
  AOI211_X1 U20157 ( .C1(n16951), .C2(n16950), .A(n16949), .B(n16948), .ZN(
        n16952) );
  OAI211_X1 U20158 ( .C1(n16960), .C2(n18807), .A(n16953), .B(n16952), .ZN(
        P3_U2667) );
  NAND2_X1 U20159 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16970) );
  NAND2_X1 U20160 ( .A1(n16971), .A2(n16954), .ZN(n16955) );
  NOR2_X1 U20161 ( .A1(n18905), .A2(n18734), .ZN(n18724) );
  OAI21_X1 U20162 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18724), .A(
        n17178), .ZN(n18874) );
  OAI22_X1 U20163 ( .A1(n16970), .A2(n16955), .B1(n17002), .B2(n18874), .ZN(
        n16962) );
  INV_X1 U20164 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18805) );
  NOR2_X1 U20165 ( .A1(n17918), .A2(n17927), .ZN(n16957) );
  OAI21_X1 U20166 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16957), .A(
        n16956), .ZN(n17908) );
  OAI21_X1 U20167 ( .B1(n17918), .B2(n16978), .A(n16986), .ZN(n16958) );
  XNOR2_X1 U20168 ( .A(n17908), .B(n16958), .ZN(n16959) );
  OAI22_X1 U20169 ( .A1(n16960), .A2(n18805), .B1(n18781), .B2(n16959), .ZN(
        n16961) );
  AOI211_X1 U20170 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n16963), .A(
        n16962), .B(n16961), .ZN(n16967) );
  OAI211_X1 U20171 ( .C1(n16968), .C2(n17294), .A(n16965), .B(n16964), .ZN(
        n16966) );
  OAI211_X1 U20172 ( .C1(n17294), .C2(n16996), .A(n16967), .B(n16966), .ZN(
        P3_U2668) );
  AOI22_X1 U20173 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17927), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17918), .ZN(n17914) );
  NAND2_X1 U20174 ( .A1(n17306), .A2(n17301), .ZN(n16984) );
  AOI211_X1 U20175 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16984), .A(n16968), .B(
        n16995), .ZN(n16975) );
  AOI21_X1 U20176 ( .B1(n18892), .B2(n18740), .A(n18724), .ZN(n18888) );
  AOI22_X1 U20177 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16969), .B1(n18888), 
        .B2(n18943), .ZN(n16973) );
  OAI211_X1 U20178 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16971), .B(n16970), .ZN(n16972) );
  OAI211_X1 U20179 ( .C1(n16987), .C2(n17918), .A(n16973), .B(n16972), .ZN(
        n16974) );
  AOI211_X1 U20180 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16976), .A(n16975), .B(
        n16974), .ZN(n16981) );
  OAI221_X1 U20181 ( .B1(n16979), .B2(n17914), .C1(n16978), .C2(n17918), .A(
        n16977), .ZN(n16980) );
  OAI211_X1 U20182 ( .C1(n16982), .C2(n17914), .A(n16981), .B(n16980), .ZN(
        P3_U2669) );
  NAND2_X1 U20183 ( .A1(n16983), .A2(n18740), .ZN(n18893) );
  OAI21_X1 U20184 ( .B1(n17301), .B2(n17306), .A(n16984), .ZN(n17302) );
  OAI22_X1 U20185 ( .A1(n16995), .A2(n17302), .B1(n18907), .B2(n16999), .ZN(
        n16985) );
  INV_X1 U20186 ( .A(n16985), .ZN(n16994) );
  NAND2_X1 U20187 ( .A1(n16986), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16988) );
  OAI21_X1 U20188 ( .B1(n18781), .B2(n16988), .A(n16987), .ZN(n16991) );
  OAI22_X1 U20189 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16989), .B1(n16996), 
        .B2(n17301), .ZN(n16990) );
  AOI221_X1 U20190 ( .B1(n16992), .B2(n17927), .C1(n16991), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16990), .ZN(n16993) );
  OAI211_X1 U20191 ( .C1(n18893), .C2(n17002), .A(n16994), .B(n16993), .ZN(
        P3_U2670) );
  NAND2_X1 U20192 ( .A1(n16996), .A2(n16995), .ZN(n16998) );
  AOI22_X1 U20193 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16998), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16997), .ZN(n17001) );
  NAND3_X1 U20194 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18884), .A3(
        n16999), .ZN(n17000) );
  OAI211_X1 U20195 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17002), .A(
        n17001), .B(n17000), .ZN(P3_U2671) );
  INV_X1 U20196 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17063) );
  NOR3_X1 U20197 ( .A1(n20806), .A2(n17063), .A3(n17094), .ZN(n17007) );
  NAND2_X1 U20198 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .ZN(n17003) );
  NAND2_X1 U20199 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17123), .ZN(n17093) );
  NOR4_X1 U20200 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17093), .ZN(
        n17006) );
  NAND4_X1 U20201 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(n17007), .A4(n17006), .ZN(n17033) );
  NOR2_X1 U20202 ( .A1(n17034), .A2(n17033), .ZN(n17032) );
  NAND2_X1 U20203 ( .A1(n17300), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17009) );
  NAND2_X1 U20204 ( .A1(n17032), .A2(n18316), .ZN(n17008) );
  OAI22_X1 U20205 ( .A1(n17032), .A2(n17009), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17008), .ZN(P3_U2672) );
  AOI22_X1 U20206 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20207 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20208 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17010) );
  OAI21_X1 U20209 ( .B1(n9642), .B2(n20811), .A(n17010), .ZN(n17016) );
  AOI22_X1 U20210 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20211 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20212 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20213 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20214 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  AOI211_X1 U20215 ( .C1(n17262), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17017) );
  NAND3_X1 U20216 ( .A1(n17019), .A2(n17018), .A3(n17017), .ZN(n17038) );
  NAND2_X1 U20217 ( .A1(n17039), .A2(n17038), .ZN(n17037) );
  AOI22_X1 U20218 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n15780), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17259), .ZN(n17024) );
  AOI22_X1 U20219 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17270), .ZN(n17023) );
  AOI22_X1 U20220 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17020), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20221 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17269), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17239), .ZN(n17021) );
  NAND4_X1 U20222 ( .A1(n17024), .A2(n17023), .A3(n17022), .A4(n17021), .ZN(
        n17030) );
  AOI22_X1 U20223 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9596), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20224 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17237), .ZN(n17027) );
  AOI22_X1 U20225 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20226 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20227 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17029) );
  NOR2_X1 U20228 ( .A1(n17030), .A2(n17029), .ZN(n17031) );
  XOR2_X1 U20229 ( .A(n17037), .B(n17031), .Z(n17314) );
  AOI211_X1 U20230 ( .C1(n17034), .C2(n17033), .A(n17032), .B(n17303), .ZN(
        n17035) );
  AOI21_X1 U20231 ( .B1(n17303), .B2(n17314), .A(n17035), .ZN(n17036) );
  INV_X1 U20232 ( .A(n17036), .ZN(P3_U2673) );
  OAI21_X1 U20233 ( .B1(n17039), .B2(n17038), .A(n17037), .ZN(n17323) );
  NAND3_X1 U20234 ( .A1(n17041), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17300), 
        .ZN(n17040) );
  OAI221_X1 U20235 ( .B1(n17041), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17300), 
        .C2(n17323), .A(n17040), .ZN(P3_U2674) );
  NOR2_X1 U20236 ( .A1(n17042), .A2(n17047), .ZN(n17052) );
  AOI21_X1 U20237 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17300), .A(n17052), .ZN(
        n17045) );
  OAI21_X1 U20238 ( .B1(n17048), .B2(n17044), .A(n17043), .ZN(n17333) );
  OAI22_X1 U20239 ( .A1(n17046), .A2(n17045), .B1(n17333), .B2(n17300), .ZN(
        P3_U2676) );
  INV_X1 U20240 ( .A(n17047), .ZN(n17056) );
  AOI21_X1 U20241 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17300), .A(n17056), .ZN(
        n17051) );
  AOI21_X1 U20242 ( .B1(n17049), .B2(n17053), .A(n17048), .ZN(n17334) );
  INV_X1 U20243 ( .A(n17334), .ZN(n17050) );
  OAI22_X1 U20244 ( .A1(n17052), .A2(n17051), .B1(n17050), .B2(n17300), .ZN(
        P3_U2677) );
  AOI21_X1 U20245 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17300), .A(n17062), .ZN(
        n17055) );
  OAI21_X1 U20246 ( .B1(n17058), .B2(n17054), .A(n17053), .ZN(n17344) );
  OAI22_X1 U20247 ( .A1(n17056), .A2(n17055), .B1(n17344), .B2(n17300), .ZN(
        P3_U2678) );
  INV_X1 U20248 ( .A(n17057), .ZN(n17069) );
  AOI21_X1 U20249 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17300), .A(n17069), .ZN(
        n17061) );
  AOI21_X1 U20250 ( .B1(n17059), .B2(n17065), .A(n17058), .ZN(n17345) );
  INV_X1 U20251 ( .A(n17345), .ZN(n17060) );
  OAI22_X1 U20252 ( .A1(n17062), .A2(n17061), .B1(n17060), .B2(n17300), .ZN(
        P3_U2679) );
  NAND2_X1 U20253 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17095), .ZN(n17082) );
  NOR2_X1 U20254 ( .A1(n17063), .A2(n17082), .ZN(n17064) );
  AOI21_X1 U20255 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17300), .A(n17064), .ZN(
        n17068) );
  OAI21_X1 U20256 ( .B1(n17067), .B2(n17066), .A(n17065), .ZN(n17354) );
  OAI22_X1 U20257 ( .A1(n17069), .A2(n17068), .B1(n17300), .B2(n17354), .ZN(
        P3_U2680) );
  AOI22_X1 U20258 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20259 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20260 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17070) );
  OAI21_X1 U20261 ( .B1(n17207), .B2(n20811), .A(n17070), .ZN(n17076) );
  AOI22_X1 U20262 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20263 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20264 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20265 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17071) );
  NAND4_X1 U20266 ( .A1(n17074), .A2(n17073), .A3(n17072), .A4(n17071), .ZN(
        n17075) );
  AOI211_X1 U20267 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17076), .B(n17075), .ZN(n17077) );
  NAND3_X1 U20268 ( .A1(n17079), .A2(n17078), .A3(n17077), .ZN(n17356) );
  INV_X1 U20269 ( .A(n17356), .ZN(n17081) );
  NAND3_X1 U20270 ( .A1(n17082), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17300), 
        .ZN(n17080) );
  OAI221_X1 U20271 ( .B1(n17082), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17300), 
        .C2(n17081), .A(n17080), .ZN(P3_U2681) );
  AOI22_X1 U20272 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20273 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20274 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20275 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20276 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17092) );
  AOI22_X1 U20277 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U20278 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20279 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20280 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17087) );
  NAND4_X1 U20281 ( .A1(n17090), .A2(n17089), .A3(n17088), .A4(n17087), .ZN(
        n17091) );
  NOR2_X1 U20282 ( .A1(n17092), .A2(n17091), .ZN(n17363) );
  AND2_X1 U20283 ( .A1(n17300), .A2(n17093), .ZN(n17108) );
  AOI22_X1 U20284 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17108), .B1(n17095), 
        .B2(n17094), .ZN(n17096) );
  OAI21_X1 U20285 ( .B1(n17363), .B2(n17300), .A(n17096), .ZN(P3_U2682) );
  AOI22_X1 U20286 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20287 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20288 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20289 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17097) );
  NAND4_X1 U20290 ( .A1(n17100), .A2(n17099), .A3(n17098), .A4(n17097), .ZN(
        n17106) );
  AOI22_X1 U20291 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20292 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20293 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20294 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17101) );
  NAND4_X1 U20295 ( .A1(n17104), .A2(n17103), .A3(n17102), .A4(n17101), .ZN(
        n17105) );
  NOR2_X1 U20296 ( .A1(n17106), .A2(n17105), .ZN(n17368) );
  INV_X1 U20297 ( .A(n17107), .ZN(n17109) );
  OAI21_X1 U20298 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17109), .A(n17108), .ZN(
        n17110) );
  OAI21_X1 U20299 ( .B1(n17368), .B2(n17300), .A(n17110), .ZN(P3_U2683) );
  INV_X1 U20300 ( .A(n17111), .ZN(n17136) );
  OAI21_X1 U20301 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17136), .A(n17300), .ZN(
        n17122) );
  AOI22_X1 U20302 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20303 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20304 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20305 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17112) );
  NAND4_X1 U20306 ( .A1(n17115), .A2(n17114), .A3(n17113), .A4(n17112), .ZN(
        n17121) );
  AOI22_X1 U20307 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20308 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20309 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20310 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17116) );
  NAND4_X1 U20311 ( .A1(n17119), .A2(n17118), .A3(n17117), .A4(n17116), .ZN(
        n17120) );
  NOR2_X1 U20312 ( .A1(n17121), .A2(n17120), .ZN(n17376) );
  OAI22_X1 U20313 ( .A1(n17123), .A2(n17122), .B1(n17376), .B2(n17300), .ZN(
        P3_U2684) );
  INV_X1 U20314 ( .A(n17147), .ZN(n17124) );
  NOR2_X1 U20315 ( .A1(n17124), .A2(n17307), .ZN(n17149) );
  AOI22_X1 U20316 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17300), .B1(
        P3_EBX_REG_17__SCAN_IN), .B2(n17149), .ZN(n17135) );
  AOI22_X1 U20317 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20318 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20319 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20320 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20321 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17134) );
  AOI22_X1 U20322 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20323 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20324 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20325 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20326 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  NOR2_X1 U20327 ( .A1(n17134), .A2(n17133), .ZN(n17381) );
  OAI22_X1 U20328 ( .A1(n17136), .A2(n17135), .B1(n17381), .B2(n17300), .ZN(
        P3_U2685) );
  AOI22_X1 U20329 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20330 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20331 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20332 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17137) );
  NAND4_X1 U20333 ( .A1(n17140), .A2(n17139), .A3(n17138), .A4(n17137), .ZN(
        n17146) );
  AOI22_X1 U20334 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20335 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20336 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20337 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17141) );
  NAND4_X1 U20338 ( .A1(n17144), .A2(n17143), .A3(n17142), .A4(n17141), .ZN(
        n17145) );
  NOR2_X1 U20339 ( .A1(n17146), .A2(n17145), .ZN(n17386) );
  NOR2_X1 U20340 ( .A1(n17424), .A2(n17147), .ZN(n17151) );
  NAND2_X1 U20341 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17305), .ZN(n17148) );
  OAI22_X1 U20342 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17149), .B1(n17151), 
        .B2(n17148), .ZN(n17150) );
  OAI21_X1 U20343 ( .B1(n17386), .B2(n17300), .A(n17150), .ZN(P3_U2686) );
  INV_X1 U20344 ( .A(n17151), .ZN(n17164) );
  INV_X1 U20345 ( .A(n17189), .ZN(n17191) );
  NAND3_X1 U20346 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17191), .ZN(n17163) );
  AOI22_X1 U20347 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20348 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20349 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20350 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17152) );
  NAND4_X1 U20351 ( .A1(n17155), .A2(n17154), .A3(n17153), .A4(n17152), .ZN(
        n17161) );
  AOI22_X1 U20352 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20353 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20354 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17157) );
  AOI22_X1 U20355 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17156) );
  NAND4_X1 U20356 ( .A1(n17159), .A2(n17158), .A3(n17157), .A4(n17156), .ZN(
        n17160) );
  NOR2_X1 U20357 ( .A1(n17161), .A2(n17160), .ZN(n17392) );
  NAND2_X1 U20358 ( .A1(n17300), .A2(n17163), .ZN(n17175) );
  OAI222_X1 U20359 ( .A1(n17164), .A2(n17163), .B1(n17300), .B2(n17392), .C1(
        n17162), .C2(n17175), .ZN(P3_U2687) );
  AOI21_X1 U20360 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17191), .A(
        P3_EBX_REG_15__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20361 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20362 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17271), .ZN(n17167) );
  AOI22_X1 U20363 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20364 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17165) );
  NAND4_X1 U20365 ( .A1(n17168), .A2(n17167), .A3(n17166), .A4(n17165), .ZN(
        n17174) );
  AOI22_X1 U20366 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17269), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17270), .ZN(n17172) );
  AOI22_X1 U20367 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17242), .ZN(n17171) );
  AOI22_X1 U20368 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17244), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17237), .ZN(n17170) );
  AOI22_X1 U20369 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17268), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n15780), .ZN(n17169) );
  NAND4_X1 U20370 ( .A1(n17172), .A2(n17171), .A3(n17170), .A4(n17169), .ZN(
        n17173) );
  NOR2_X1 U20371 ( .A1(n17174), .A2(n17173), .ZN(n17395) );
  OAI22_X1 U20372 ( .A1(n17176), .A2(n17175), .B1(n17395), .B2(n17300), .ZN(
        P3_U2688) );
  AOI22_X1 U20373 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20374 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20375 ( .A1(n17242), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17177) );
  OAI21_X1 U20376 ( .B1(n17178), .B2(n20811), .A(n17177), .ZN(n17184) );
  AOI22_X1 U20377 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20378 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17262), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20379 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20380 ( .A1(n15780), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17179) );
  NAND4_X1 U20381 ( .A1(n17182), .A2(n17181), .A3(n17180), .A4(n17179), .ZN(
        n17183) );
  AOI211_X1 U20382 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17184), .B(n17183), .ZN(n17186) );
  NAND3_X1 U20383 ( .A1(n17188), .A2(n17187), .A3(n17186), .ZN(n17397) );
  INV_X1 U20384 ( .A(n17397), .ZN(n17193) );
  OAI221_X1 U20385 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17191), .C1(n17190), 
        .C2(n17189), .A(n17300), .ZN(n17192) );
  OAI21_X1 U20386 ( .B1(n17193), .B2(n17300), .A(n17192), .ZN(P3_U2689) );
  AOI22_X1 U20387 ( .A1(n15648), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20388 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20389 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20390 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17194) );
  NAND4_X1 U20391 ( .A1(n17197), .A2(n17196), .A3(n17195), .A4(n17194), .ZN(
        n17203) );
  AOI22_X1 U20392 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20393 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20394 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20395 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17198) );
  NAND4_X1 U20396 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        n17202) );
  NOR2_X1 U20397 ( .A1(n17203), .A2(n17202), .ZN(n17407) );
  NAND3_X1 U20398 ( .A1(n17205), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17300), 
        .ZN(n17204) );
  OAI221_X1 U20399 ( .B1(n17205), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17300), 
        .C2(n17407), .A(n17204), .ZN(P3_U2691) );
  AOI22_X1 U20400 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20401 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17215) );
  INV_X1 U20402 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U20403 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17206) );
  OAI21_X1 U20404 ( .B1(n17207), .B2(n18291), .A(n17206), .ZN(n17213) );
  AOI22_X1 U20405 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20406 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20407 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20408 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17208) );
  NAND4_X1 U20409 ( .A1(n17211), .A2(n17210), .A3(n17209), .A4(n17208), .ZN(
        n17212) );
  AOI211_X1 U20410 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17213), .B(n17212), .ZN(n17214) );
  NAND3_X1 U20411 ( .A1(n17216), .A2(n17215), .A3(n17214), .ZN(n17411) );
  INV_X1 U20412 ( .A(n17411), .ZN(n17221) );
  NOR2_X1 U20413 ( .A1(n17217), .A2(n17254), .ZN(n17218) );
  OAI21_X1 U20414 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17218), .A(n17300), .ZN(
        n17219) );
  OAI22_X1 U20415 ( .A1(n17221), .A2(n17300), .B1(n17220), .B2(n17219), .ZN(
        P3_U2692) );
  AOI22_X1 U20416 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20417 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20418 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20419 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17222) );
  NAND4_X1 U20420 ( .A1(n17225), .A2(n17224), .A3(n17223), .A4(n17222), .ZN(
        n17231) );
  AOI22_X1 U20421 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20422 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20423 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20424 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17226) );
  NAND4_X1 U20425 ( .A1(n17229), .A2(n17228), .A3(n17227), .A4(n17226), .ZN(
        n17230) );
  NOR2_X1 U20426 ( .A1(n17231), .A2(n17230), .ZN(n17415) );
  NOR2_X1 U20427 ( .A1(n17233), .A2(n17254), .ZN(n17232) );
  NOR2_X1 U20428 ( .A1(n17303), .A2(n17232), .ZN(n17255) );
  NOR3_X1 U20429 ( .A1(n17424), .A2(n17233), .A3(n17254), .ZN(n17235) );
  AOI22_X1 U20430 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17255), .B1(n17235), 
        .B2(n17234), .ZN(n17236) );
  OAI21_X1 U20431 ( .B1(n17415), .B2(n17300), .A(n17236), .ZN(P3_U2693) );
  AOI22_X1 U20432 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17271), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U20433 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20434 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U20435 ( .B1(n17241), .B2(n20791), .A(n17240), .ZN(n17250) );
  AOI22_X1 U20436 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17242), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20437 ( .A1(n17243), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20438 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20439 ( .A1(n17244), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17245) );
  NAND4_X1 U20440 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        n17249) );
  AOI211_X1 U20441 ( .C1(n15648), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n17250), .B(n17249), .ZN(n17251) );
  NAND3_X1 U20442 ( .A1(n17253), .A2(n17252), .A3(n17251), .ZN(n17419) );
  INV_X1 U20443 ( .A(n17419), .ZN(n17258) );
  INV_X1 U20444 ( .A(n17254), .ZN(n17256) );
  OAI21_X1 U20445 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17256), .A(n17255), .ZN(
        n17257) );
  OAI21_X1 U20446 ( .B1(n17258), .B2(n17300), .A(n17257), .ZN(P3_U2694) );
  AOI22_X1 U20447 ( .A1(n17260), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17259), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20448 ( .A1(n17261), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U20449 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U20450 ( .A1(n17263), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17264) );
  NAND4_X1 U20451 ( .A1(n17267), .A2(n17266), .A3(n17265), .A4(n17264), .ZN(
        n17277) );
  AOI22_X1 U20452 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15780), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20453 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20454 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20455 ( .A1(n17271), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17270), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17272) );
  NAND4_X1 U20456 ( .A1(n17275), .A2(n17274), .A3(n17273), .A4(n17272), .ZN(
        n17276) );
  NOR2_X1 U20457 ( .A1(n17277), .A2(n17276), .ZN(n17428) );
  NOR2_X1 U20458 ( .A1(n17303), .A2(n17285), .ZN(n17282) );
  NOR2_X1 U20459 ( .A1(n17424), .A2(n17289), .ZN(n17296) );
  NOR2_X1 U20460 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17278), .ZN(n17279) );
  AOI22_X1 U20461 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17282), .B1(n17296), .B2(
        n17279), .ZN(n17280) );
  OAI21_X1 U20462 ( .B1(n17428), .B2(n17300), .A(n17280), .ZN(P3_U2695) );
  NOR3_X1 U20463 ( .A1(n17424), .A2(n17281), .A3(n17289), .ZN(n17287) );
  NAND2_X1 U20464 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17287), .ZN(n17284) );
  AOI22_X1 U20465 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17303), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17282), .ZN(n17283) );
  OAI21_X1 U20466 ( .B1(n17285), .B2(n17284), .A(n17283), .ZN(P3_U2696) );
  INV_X1 U20467 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18311) );
  NOR2_X1 U20468 ( .A1(n17303), .A2(n17287), .ZN(n17290) );
  INV_X1 U20469 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20470 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17290), .B1(n17287), .B2(
        n17286), .ZN(n17288) );
  OAI21_X1 U20471 ( .B1(n18311), .B2(n17300), .A(n17288), .ZN(P3_U2697) );
  INV_X1 U20472 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18304) );
  INV_X1 U20473 ( .A(n17289), .ZN(n17291) );
  OAI21_X1 U20474 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17291), .A(n17290), .ZN(
        n17292) );
  OAI21_X1 U20475 ( .B1(n17300), .B2(n18304), .A(n17292), .ZN(P3_U2698) );
  NOR3_X1 U20476 ( .A1(n17294), .A2(n17293), .A3(n17307), .ZN(n17299) );
  AOI21_X1 U20477 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17300), .A(n17299), .ZN(
        n17295) );
  OAI22_X1 U20478 ( .A1(n17296), .A2(n17295), .B1(n18297), .B2(n17300), .ZN(
        P3_U2699) );
  AOI21_X1 U20479 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17300), .A(n17297), .ZN(
        n17298) );
  OAI22_X1 U20480 ( .A1(n17299), .A2(n17298), .B1(n18291), .B2(n17300), .ZN(
        P3_U2700) );
  INV_X1 U20481 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18277) );
  OAI222_X1 U20482 ( .A1(n17307), .A2(n17302), .B1(n17301), .B2(n17305), .C1(
        n18277), .C2(n17300), .ZN(P3_U2702) );
  NAND2_X1 U20483 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17303), .ZN(
        n17304) );
  OAI221_X1 U20484 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17307), .C1(n17306), 
        .C2(n17305), .A(n17304), .ZN(P3_U2703) );
  INV_X1 U20485 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17527) );
  INV_X1 U20486 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17523) );
  INV_X1 U20487 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17568) );
  NAND4_X1 U20488 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20489 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n17308) );
  INV_X1 U20490 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17558) );
  INV_X1 U20491 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17555) );
  INV_X1 U20492 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17549) );
  NAND2_X1 U20493 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17396) );
  NOR4_X1 U20494 ( .A1(n17558), .A2(n17555), .A3(n17549), .A4(n17396), .ZN(
        n17310) );
  NAND2_X1 U20495 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n17355) );
  NAND2_X1 U20496 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17351), .ZN(n17350) );
  NAND2_X1 U20497 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17335), .ZN(n17330) );
  INV_X1 U20498 ( .A(n17320), .ZN(n17316) );
  NAND2_X1 U20499 ( .A1(n17316), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17387), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17311), .ZN(n17312) );
  OAI21_X1 U20501 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17313), .A(n17312), .ZN(
        P3_U2704) );
  INV_X1 U20502 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20503 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17387), .B1(n17456), .B2(
        n17314), .ZN(n17318) );
  NOR2_X2 U20504 ( .A1(n17315), .A2(n17449), .ZN(n17388) );
  AOI22_X1 U20505 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17388), .B1(n17316), .B2(
        n17531), .ZN(n17317) );
  OAI211_X1 U20506 ( .C1(n17319), .C2(n17531), .A(n17318), .B(n17317), .ZN(
        P3_U2705) );
  AOI22_X1 U20507 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17387), .ZN(n17322) );
  OAI211_X1 U20508 ( .C1(n17325), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17449), .B(
        n17320), .ZN(n17321) );
  OAI211_X1 U20509 ( .C1(n17323), .C2(n17451), .A(n17322), .B(n17321), .ZN(
        P3_U2706) );
  INV_X1 U20510 ( .A(n17387), .ZN(n17367) );
  AOI22_X1 U20511 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17388), .B1(n17456), .B2(
        n17324), .ZN(n17329) );
  INV_X1 U20512 ( .A(n17330), .ZN(n17327) );
  INV_X1 U20513 ( .A(n17325), .ZN(n17326) );
  OAI211_X1 U20514 ( .C1(n17327), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17449), .B(
        n17326), .ZN(n17328) );
  OAI211_X1 U20515 ( .C1(n17367), .C2(n18292), .A(n17329), .B(n17328), .ZN(
        P3_U2707) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17387), .ZN(n17332) );
  OAI211_X1 U20517 ( .C1(n17335), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17449), .B(
        n17330), .ZN(n17331) );
  OAI211_X1 U20518 ( .C1(n17333), .C2(n17451), .A(n17332), .B(n17331), .ZN(
        P3_U2708) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17388), .B1(n17456), .B2(
        n17334), .ZN(n17339) );
  INV_X1 U20520 ( .A(n17340), .ZN(n17337) );
  INV_X1 U20521 ( .A(n17335), .ZN(n17336) );
  OAI211_X1 U20522 ( .C1(n17337), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17449), .B(
        n17336), .ZN(n17338) );
  OAI211_X1 U20523 ( .C1(n17367), .C2(n18280), .A(n17339), .B(n17338), .ZN(
        P3_U2709) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17387), .ZN(n17343) );
  OAI211_X1 U20525 ( .C1(n17341), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17449), .B(
        n17340), .ZN(n17342) );
  OAI211_X1 U20526 ( .C1(n17344), .C2(n17451), .A(n17343), .B(n17342), .ZN(
        P3_U2710) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17388), .B1(n17456), .B2(
        n17345), .ZN(n17349) );
  OAI211_X1 U20528 ( .C1(n17347), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17449), .B(
        n17346), .ZN(n17348) );
  OAI211_X1 U20529 ( .C1(n17367), .C2(n18265), .A(n17349), .B(n17348), .ZN(
        P3_U2711) );
  AOI22_X1 U20530 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17387), .ZN(n17353) );
  OAI211_X1 U20531 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17351), .A(n17449), .B(
        n17350), .ZN(n17352) );
  OAI211_X1 U20532 ( .C1(n17354), .C2(n17451), .A(n17353), .B(n17352), .ZN(
        P3_U2712) );
  INV_X1 U20533 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17508) );
  INV_X1 U20534 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17506) );
  INV_X1 U20535 ( .A(n17378), .ZN(n17382) );
  INV_X1 U20536 ( .A(n17373), .ZN(n17377) );
  NOR2_X1 U20537 ( .A1(n17355), .A2(n17377), .ZN(n17357) );
  NAND2_X1 U20538 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17357), .ZN(n17362) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17387), .B1(n17456), .B2(
        n17356), .ZN(n17361) );
  INV_X1 U20540 ( .A(n17357), .ZN(n17366) );
  NAND2_X1 U20541 ( .A1(n17449), .A2(n17366), .ZN(n17371) );
  OAI21_X1 U20542 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17358), .A(n17371), .ZN(
        n17359) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17388), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17359), .ZN(n17360) );
  OAI211_X1 U20544 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17362), .A(n17361), .B(
        n17360), .ZN(P3_U2713) );
  INV_X1 U20545 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17513) );
  OAI22_X1 U20546 ( .A1(n17363), .A2(n17451), .B1(n18301), .B2(n17367), .ZN(
        n17364) );
  AOI21_X1 U20547 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17388), .A(n17364), .ZN(
        n17365) );
  OAI221_X1 U20548 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17366), .C1(n17513), 
        .C2(n17371), .A(n17365), .ZN(P3_U2714) );
  NAND2_X1 U20549 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17373), .ZN(n17372) );
  INV_X1 U20550 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17511) );
  OAI22_X1 U20551 ( .A1(n17368), .A2(n17451), .B1(n18294), .B2(n17367), .ZN(
        n17369) );
  AOI21_X1 U20552 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17388), .A(n17369), .ZN(
        n17370) );
  OAI221_X1 U20553 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17372), .C1(n17511), 
        .C2(n17371), .A(n17370), .ZN(P3_U2715) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17387), .ZN(n17375) );
  OAI211_X1 U20555 ( .C1(n17373), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17449), .B(
        n17372), .ZN(n17374) );
  OAI211_X1 U20556 ( .C1(n17376), .C2(n17451), .A(n17375), .B(n17374), .ZN(
        P3_U2716) );
  AOI22_X1 U20557 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17387), .ZN(n17380) );
  OAI211_X1 U20558 ( .C1(n17378), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17449), .B(
        n17377), .ZN(n17379) );
  OAI211_X1 U20559 ( .C1(n17381), .C2(n17451), .A(n17380), .B(n17379), .ZN(
        P3_U2717) );
  AOI22_X1 U20560 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17387), .ZN(n17385) );
  INV_X1 U20561 ( .A(n17389), .ZN(n17383) );
  OAI211_X1 U20562 ( .C1(n17383), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17449), .B(
        n17382), .ZN(n17384) );
  OAI211_X1 U20563 ( .C1(n17386), .C2(n17451), .A(n17385), .B(n17384), .ZN(
        P3_U2718) );
  AOI22_X1 U20564 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17388), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17387), .ZN(n17391) );
  OAI211_X1 U20565 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n9652), .A(n17449), .B(
        n17389), .ZN(n17390) );
  OAI211_X1 U20566 ( .C1(n17392), .C2(n17451), .A(n17391), .B(n17390), .ZN(
        P3_U2719) );
  AOI21_X1 U20567 ( .B1(n17568), .B2(n17398), .A(n9652), .ZN(n17393) );
  AOI22_X1 U20568 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17457), .B1(n17393), .B2(
        n17449), .ZN(n17394) );
  OAI21_X1 U20569 ( .B1(n17395), .B2(n17451), .A(n17394), .ZN(P3_U2720) );
  NAND3_X1 U20570 ( .A1(n18316), .A2(n17423), .A3(P3_EAX_REG_8__SCAN_IN), .ZN(
        n17422) );
  OR2_X1 U20571 ( .A1(n17396), .A2(n17422), .ZN(n17413) );
  NOR2_X1 U20572 ( .A1(n17555), .A2(n17413), .ZN(n17406) );
  NAND2_X1 U20573 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17409), .ZN(n17401) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17457), .B1(n17456), .B2(
        n17397), .ZN(n17400) );
  NAND3_X1 U20575 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17449), .A3(n17398), 
        .ZN(n17399) );
  OAI211_X1 U20576 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17401), .A(n17400), .B(
        n17399), .ZN(P3_U2721) );
  INV_X1 U20577 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17405) );
  INV_X1 U20578 ( .A(n17401), .ZN(n17404) );
  AOI21_X1 U20579 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17449), .A(n17409), .ZN(
        n17403) );
  OAI222_X1 U20580 ( .A1(n17454), .A2(n17405), .B1(n17404), .B2(n17403), .C1(
        n17451), .C2(n17402), .ZN(P3_U2722) );
  AOI21_X1 U20581 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17449), .A(n17406), .ZN(
        n17408) );
  OAI222_X1 U20582 ( .A1(n17454), .A2(n17410), .B1(n17409), .B2(n17408), .C1(
        n17451), .C2(n17407), .ZN(P3_U2723) );
  NAND2_X1 U20583 ( .A1(n17449), .A2(n17413), .ZN(n17417) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17457), .B1(n17456), .B2(
        n17411), .ZN(n17412) );
  OAI221_X1 U20585 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17413), .C1(n17555), 
        .C2(n17417), .A(n17412), .ZN(P3_U2724) );
  INV_X1 U20586 ( .A(n17422), .ZN(n17414) );
  AOI21_X1 U20587 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17414), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17416) );
  OAI222_X1 U20588 ( .A1(n17454), .A2(n17418), .B1(n17417), .B2(n17416), .C1(
        n17451), .C2(n17415), .ZN(P3_U2725) );
  NAND3_X1 U20589 ( .A1(n17449), .A2(P3_EAX_REG_9__SCAN_IN), .A3(n17422), .ZN(
        n17421) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17457), .B1(n17456), .B2(
        n17419), .ZN(n17420) );
  OAI211_X1 U20591 ( .C1(P3_EAX_REG_9__SCAN_IN), .C2(n17422), .A(n17421), .B(
        n17420), .ZN(P3_U2726) );
  INV_X1 U20592 ( .A(n17423), .ZN(n17425) );
  NOR2_X1 U20593 ( .A1(n17424), .A2(n17425), .ZN(n17432) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17457), .B1(n17432), .B2(
        n17549), .ZN(n17427) );
  NAND3_X1 U20595 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17449), .A3(n17425), .ZN(
        n17426) );
  OAI211_X1 U20596 ( .C1(n17428), .C2(n17451), .A(n17427), .B(n17426), .ZN(
        P3_U2727) );
  INV_X1 U20597 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18313) );
  INV_X1 U20598 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17535) );
  NOR2_X1 U20599 ( .A1(n17535), .A2(n17460), .ZN(n17448) );
  INV_X1 U20600 ( .A(n17448), .ZN(n17440) );
  NOR2_X1 U20601 ( .A1(n17429), .A2(n17440), .ZN(n17438) );
  AOI22_X1 U20602 ( .A1(n17438), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17449), .ZN(n17431) );
  OAI222_X1 U20603 ( .A1(n17454), .A2(n18313), .B1(n17432), .B2(n17431), .C1(
        n17451), .C2(n17430), .ZN(P3_U2728) );
  AOI21_X1 U20604 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17449), .A(n17438), .ZN(
        n17435) );
  AND2_X1 U20605 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17438), .ZN(n17434) );
  OAI222_X1 U20606 ( .A1(n17454), .A2(n18306), .B1(n17435), .B2(n17434), .C1(
        n17451), .C2(n17433), .ZN(P3_U2729) );
  NAND3_X1 U20607 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n17436) );
  NOR2_X1 U20608 ( .A1(n17436), .A2(n17440), .ZN(n17443) );
  AOI21_X1 U20609 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17449), .A(n17443), .ZN(
        n17439) );
  OAI222_X1 U20610 ( .A1(n17454), .A2(n18299), .B1(n17439), .B2(n17438), .C1(
        n17451), .C2(n17437), .ZN(P3_U2730) );
  INV_X1 U20611 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17537) );
  NOR2_X1 U20612 ( .A1(n17537), .A2(n17440), .ZN(n17453) );
  AOI22_X1 U20613 ( .A1(n17453), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17449), .ZN(n17444) );
  INV_X1 U20614 ( .A(n17441), .ZN(n17442) );
  OAI222_X1 U20615 ( .A1(n17454), .A2(n20858), .B1(n17444), .B2(n17443), .C1(
        n17451), .C2(n17442), .ZN(P3_U2731) );
  AND2_X1 U20616 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17453), .ZN(n17447) );
  AOI21_X1 U20617 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17449), .A(n17453), .ZN(
        n17446) );
  OAI222_X1 U20618 ( .A1(n18286), .A2(n17454), .B1(n17447), .B2(n17446), .C1(
        n17451), .C2(n17445), .ZN(P3_U2732) );
  AOI21_X1 U20619 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17449), .A(n17448), .ZN(
        n17452) );
  OAI222_X1 U20620 ( .A1(n18279), .A2(n17454), .B1(n17453), .B2(n17452), .C1(
        n17451), .C2(n17450), .ZN(P3_U2733) );
  AOI22_X1 U20621 ( .A1(n17457), .A2(BUF2_REG_1__SCAN_IN), .B1(n17456), .B2(
        n17455), .ZN(n17458) );
  OAI221_X1 U20622 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17460), .C1(n17535), 
        .C2(n17459), .A(n17458), .ZN(P3_U2734) );
  AND2_X1 U20623 ( .A1(n17489), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20624 ( .A1(n17463), .A2(n17462), .ZN(n17479) );
  AOI22_X1 U20625 ( .A1(n18920), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20626 ( .B1(n17531), .B2(n17479), .A(n17464), .ZN(P3_U2737) );
  INV_X1 U20627 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U20628 ( .A1(n18920), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20629 ( .B1(n17529), .B2(n17479), .A(n17465), .ZN(P3_U2738) );
  AOI22_X1 U20630 ( .A1(n18920), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20631 ( .B1(n17527), .B2(n17479), .A(n17466), .ZN(P3_U2739) );
  INV_X1 U20632 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20633 ( .A1(n18920), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20634 ( .B1(n17525), .B2(n17479), .A(n17467), .ZN(P3_U2740) );
  AOI22_X1 U20635 ( .A1(n18920), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20636 ( .B1(n17523), .B2(n17479), .A(n17468), .ZN(P3_U2741) );
  INV_X1 U20637 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17521) );
  AOI22_X1 U20638 ( .A1(n18920), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20639 ( .B1(n17521), .B2(n17479), .A(n17469), .ZN(P3_U2742) );
  INV_X1 U20640 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20641 ( .A1(n18920), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U20642 ( .B1(n17519), .B2(n17479), .A(n17470), .ZN(P3_U2743) );
  INV_X1 U20643 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17517) );
  CLKBUF_X1 U20644 ( .A(n18920), .Z(n17497) );
  AOI22_X1 U20645 ( .A1(n17497), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20646 ( .B1(n17517), .B2(n17479), .A(n17471), .ZN(P3_U2744) );
  INV_X1 U20647 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17515) );
  AOI22_X1 U20648 ( .A1(n17497), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U20649 ( .B1(n17515), .B2(n17479), .A(n17472), .ZN(P3_U2745) );
  AOI22_X1 U20650 ( .A1(n17497), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20651 ( .B1(n17513), .B2(n17479), .A(n17473), .ZN(P3_U2746) );
  AOI22_X1 U20652 ( .A1(n17497), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20653 ( .B1(n17511), .B2(n17479), .A(n17474), .ZN(P3_U2747) );
  INV_X1 U20654 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U20655 ( .A1(n17497), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20656 ( .B1(n20892), .B2(n17479), .A(n17475), .ZN(P3_U2748) );
  AOI22_X1 U20657 ( .A1(n17497), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17476) );
  OAI21_X1 U20658 ( .B1(n17508), .B2(n17479), .A(n17476), .ZN(P3_U2749) );
  AOI22_X1 U20659 ( .A1(n17497), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20660 ( .B1(n17506), .B2(n17479), .A(n17477), .ZN(P3_U2750) );
  INV_X1 U20661 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U20662 ( .A1(n17497), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20663 ( .B1(n17504), .B2(n17479), .A(n17478), .ZN(P3_U2751) );
  AOI22_X1 U20664 ( .A1(n17497), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17480) );
  OAI21_X1 U20665 ( .B1(n17568), .B2(n17499), .A(n17480), .ZN(P3_U2752) );
  INV_X1 U20666 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20667 ( .A1(n17497), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20668 ( .B1(n17563), .B2(n17499), .A(n17481), .ZN(P3_U2753) );
  INV_X1 U20669 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17560) );
  AOI22_X1 U20670 ( .A1(n17497), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17482) );
  OAI21_X1 U20671 ( .B1(n17560), .B2(n17499), .A(n17482), .ZN(P3_U2754) );
  AOI22_X1 U20672 ( .A1(n17497), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20673 ( .B1(n17558), .B2(n17499), .A(n17483), .ZN(P3_U2755) );
  AOI22_X1 U20674 ( .A1(n17497), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17484) );
  OAI21_X1 U20675 ( .B1(n17555), .B2(n17499), .A(n17484), .ZN(P3_U2756) );
  INV_X1 U20676 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17553) );
  AOI22_X1 U20677 ( .A1(n17497), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17485) );
  OAI21_X1 U20678 ( .B1(n17553), .B2(n17499), .A(n17485), .ZN(P3_U2757) );
  INV_X1 U20679 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20680 ( .A1(n17497), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17486) );
  OAI21_X1 U20681 ( .B1(n17551), .B2(n17499), .A(n17486), .ZN(P3_U2758) );
  AOI22_X1 U20682 ( .A1(n17497), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20683 ( .B1(n17549), .B2(n17499), .A(n17487), .ZN(P3_U2759) );
  INV_X1 U20684 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17547) );
  AOI22_X1 U20685 ( .A1(n17497), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17488) );
  OAI21_X1 U20686 ( .B1(n17547), .B2(n17499), .A(n17488), .ZN(P3_U2760) );
  INV_X1 U20687 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17545) );
  AOI22_X1 U20688 ( .A1(n17497), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17489), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17490) );
  OAI21_X1 U20689 ( .B1(n17545), .B2(n17499), .A(n17490), .ZN(P3_U2761) );
  INV_X1 U20690 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20691 ( .A1(n17497), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20692 ( .B1(n17543), .B2(n17499), .A(n17491), .ZN(P3_U2762) );
  INV_X1 U20693 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20694 ( .A1(n17497), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17492) );
  OAI21_X1 U20695 ( .B1(n17541), .B2(n17499), .A(n17492), .ZN(P3_U2763) );
  INV_X1 U20696 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20697 ( .A1(n17497), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20698 ( .B1(n17539), .B2(n17499), .A(n17493), .ZN(P3_U2764) );
  AOI22_X1 U20699 ( .A1(n17497), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20700 ( .B1(n17537), .B2(n17499), .A(n17494), .ZN(P3_U2765) );
  AOI22_X1 U20701 ( .A1(n17497), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17495) );
  OAI21_X1 U20702 ( .B1(n17535), .B2(n17499), .A(n17495), .ZN(P3_U2766) );
  AOI22_X1 U20703 ( .A1(n17497), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17496), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20704 ( .B1(n17533), .B2(n17499), .A(n17498), .ZN(P3_U2767) );
  OAI211_X1 U20705 ( .C1(n18274), .C2(n18919), .A(n17502), .B(n17501), .ZN(
        n17556) );
  AOI22_X1 U20706 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17564), .ZN(n17503) );
  OAI21_X1 U20707 ( .B1(n17504), .B2(n17567), .A(n17503), .ZN(P3_U2768) );
  AOI22_X1 U20708 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17564), .ZN(n17505) );
  OAI21_X1 U20709 ( .B1(n17506), .B2(n17567), .A(n17505), .ZN(P3_U2769) );
  AOI22_X1 U20710 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17564), .ZN(n17507) );
  OAI21_X1 U20711 ( .B1(n17508), .B2(n17567), .A(n17507), .ZN(P3_U2770) );
  AOI22_X1 U20712 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17564), .ZN(n17509) );
  OAI21_X1 U20713 ( .B1(n20892), .B2(n17567), .A(n17509), .ZN(P3_U2771) );
  AOI22_X1 U20714 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17564), .ZN(n17510) );
  OAI21_X1 U20715 ( .B1(n17511), .B2(n17567), .A(n17510), .ZN(P3_U2772) );
  AOI22_X1 U20716 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17564), .ZN(n17512) );
  OAI21_X1 U20717 ( .B1(n17513), .B2(n17567), .A(n17512), .ZN(P3_U2773) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17564), .ZN(n17514) );
  OAI21_X1 U20719 ( .B1(n17515), .B2(n17567), .A(n17514), .ZN(P3_U2774) );
  AOI22_X1 U20720 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17564), .ZN(n17516) );
  OAI21_X1 U20721 ( .B1(n17517), .B2(n17567), .A(n17516), .ZN(P3_U2775) );
  AOI22_X1 U20722 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17564), .ZN(n17518) );
  OAI21_X1 U20723 ( .B1(n17519), .B2(n17567), .A(n17518), .ZN(P3_U2776) );
  AOI22_X1 U20724 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17564), .ZN(n17520) );
  OAI21_X1 U20725 ( .B1(n17521), .B2(n17567), .A(n17520), .ZN(P3_U2777) );
  AOI22_X1 U20726 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17564), .ZN(n17522) );
  OAI21_X1 U20727 ( .B1(n17523), .B2(n17567), .A(n17522), .ZN(P3_U2778) );
  AOI22_X1 U20728 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17565), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17564), .ZN(n17524) );
  OAI21_X1 U20729 ( .B1(n17525), .B2(n17567), .A(n17524), .ZN(P3_U2779) );
  AOI22_X1 U20730 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17564), .ZN(n17526) );
  OAI21_X1 U20731 ( .B1(n17527), .B2(n17567), .A(n17526), .ZN(P3_U2780) );
  AOI22_X1 U20732 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17564), .ZN(n17528) );
  OAI21_X1 U20733 ( .B1(n17529), .B2(n17567), .A(n17528), .ZN(P3_U2781) );
  AOI22_X1 U20734 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17561), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17564), .ZN(n17530) );
  OAI21_X1 U20735 ( .B1(n17531), .B2(n17567), .A(n17530), .ZN(P3_U2782) );
  AOI22_X1 U20736 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17564), .ZN(n17532) );
  OAI21_X1 U20737 ( .B1(n17533), .B2(n17567), .A(n17532), .ZN(P3_U2783) );
  AOI22_X1 U20738 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17564), .ZN(n17534) );
  OAI21_X1 U20739 ( .B1(n17535), .B2(n17567), .A(n17534), .ZN(P3_U2784) );
  AOI22_X1 U20740 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17564), .ZN(n17536) );
  OAI21_X1 U20741 ( .B1(n17537), .B2(n17567), .A(n17536), .ZN(P3_U2785) );
  AOI22_X1 U20742 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17556), .ZN(n17538) );
  OAI21_X1 U20743 ( .B1(n17539), .B2(n17567), .A(n17538), .ZN(P3_U2786) );
  AOI22_X1 U20744 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17556), .ZN(n17540) );
  OAI21_X1 U20745 ( .B1(n17541), .B2(n17567), .A(n17540), .ZN(P3_U2787) );
  AOI22_X1 U20746 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17556), .ZN(n17542) );
  OAI21_X1 U20747 ( .B1(n17543), .B2(n17567), .A(n17542), .ZN(P3_U2788) );
  AOI22_X1 U20748 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17556), .ZN(n17544) );
  OAI21_X1 U20749 ( .B1(n17545), .B2(n17567), .A(n17544), .ZN(P3_U2789) );
  AOI22_X1 U20750 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17556), .ZN(n17546) );
  OAI21_X1 U20751 ( .B1(n17547), .B2(n17567), .A(n17546), .ZN(P3_U2790) );
  AOI22_X1 U20752 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17556), .ZN(n17548) );
  OAI21_X1 U20753 ( .B1(n17549), .B2(n17567), .A(n17548), .ZN(P3_U2791) );
  AOI22_X1 U20754 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17556), .ZN(n17550) );
  OAI21_X1 U20755 ( .B1(n17551), .B2(n17567), .A(n17550), .ZN(P3_U2792) );
  AOI22_X1 U20756 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17565), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17556), .ZN(n17552) );
  OAI21_X1 U20757 ( .B1(n17553), .B2(n17567), .A(n17552), .ZN(P3_U2793) );
  AOI22_X1 U20758 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17556), .ZN(n17554) );
  OAI21_X1 U20759 ( .B1(n17555), .B2(n17567), .A(n17554), .ZN(P3_U2794) );
  AOI22_X1 U20760 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17556), .ZN(n17557) );
  OAI21_X1 U20761 ( .B1(n17558), .B2(n17567), .A(n17557), .ZN(P3_U2795) );
  AOI22_X1 U20762 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17565), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17564), .ZN(n17559) );
  OAI21_X1 U20763 ( .B1(n17560), .B2(n17567), .A(n17559), .ZN(P3_U2796) );
  AOI22_X1 U20764 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17561), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17564), .ZN(n17562) );
  OAI21_X1 U20765 ( .B1(n17563), .B2(n17567), .A(n17562), .ZN(P3_U2797) );
  AOI22_X1 U20766 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17565), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17564), .ZN(n17566) );
  OAI21_X1 U20767 ( .B1(n17568), .B2(n17567), .A(n17566), .ZN(P3_U2798) );
  OAI21_X1 U20768 ( .B1(n17569), .B2(n17932), .A(n17931), .ZN(n17570) );
  AOI21_X1 U20769 ( .B1(n17834), .B2(n17571), .A(n17570), .ZN(n17608) );
  OAI21_X1 U20770 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17613), .A(
        n17608), .ZN(n17591) );
  NOR2_X1 U20771 ( .A1(n17777), .A2(n17571), .ZN(n17593) );
  XOR2_X1 U20772 ( .A(n17572), .B(n17592), .Z(n17573) );
  AOI22_X1 U20773 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17591), .B1(
        n17593), .B2(n17573), .ZN(n17584) );
  AOI22_X1 U20774 ( .A1(n9593), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17772), 
        .B2(n17574), .ZN(n17583) );
  AOI21_X1 U20775 ( .B1(n17577), .B2(n17576), .A(n17575), .ZN(n17579) );
  AOI22_X1 U20776 ( .A1(n17824), .A2(n17579), .B1(n17578), .B2(n17666), .ZN(
        n17582) );
  AOI22_X1 U20777 ( .A1(n17841), .A2(n17946), .B1(n9589), .B2(n17580), .ZN(
        n17603) );
  NAND2_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17603), .ZN(
        n17594) );
  OAI211_X1 U20779 ( .C1(n17841), .C2(n9589), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17594), .ZN(n17581) );
  NAND4_X1 U20780 ( .A1(n17584), .A2(n17583), .A3(n17582), .A4(n17581), .ZN(
        P3_U2802) );
  INV_X1 U20781 ( .A(n17585), .ZN(n17587) );
  NAND2_X1 U20782 ( .A1(n17587), .A2(n17586), .ZN(n17588) );
  XOR2_X1 U20783 ( .A(n17829), .B(n17588), .Z(n17952) );
  INV_X1 U20784 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18851) );
  OAI22_X1 U20785 ( .A1(n18181), .A2(n18851), .B1(n17797), .B2(n17589), .ZN(
        n17590) );
  AOI221_X1 U20786 ( .B1(n17593), .B2(n17592), .C1(n17591), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17590), .ZN(n17597) );
  OAI21_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17595), .A(
        n17594), .ZN(n17596) );
  OAI211_X1 U20788 ( .C1(n17952), .C2(n17844), .A(n17597), .B(n17596), .ZN(
        P3_U2803) );
  NOR2_X1 U20789 ( .A1(n18395), .A2(n17598), .ZN(n17645) );
  AOI21_X1 U20790 ( .B1(n17599), .B2(n17645), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U20791 ( .A1(n17797), .A2(n17613), .ZN(n17923) );
  AOI22_X1 U20792 ( .A1(n9593), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17600), 
        .B2(n17923), .ZN(n17606) );
  NOR3_X1 U20793 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17964), .A3(
        n17961), .ZN(n17956) );
  INV_X1 U20794 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17953) );
  AOI21_X1 U20795 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17602), .A(
        n17601), .ZN(n17959) );
  OAI22_X1 U20796 ( .A1(n17603), .A2(n17953), .B1(n17959), .B2(n17844), .ZN(
        n17604) );
  AOI21_X1 U20797 ( .B1(n17666), .B2(n17956), .A(n17604), .ZN(n17605) );
  OAI211_X1 U20798 ( .C1(n17608), .C2(n17607), .A(n17606), .B(n17605), .ZN(
        P3_U2804) );
  XOR2_X1 U20799 ( .A(n17609), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17973) );
  NAND2_X1 U20800 ( .A1(n17610), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17614) );
  OAI21_X1 U20801 ( .B1(n17611), .B2(n17932), .A(n17931), .ZN(n17612) );
  AOI21_X1 U20802 ( .B1(n18653), .B2(n17614), .A(n17612), .ZN(n17647) );
  OAI21_X1 U20803 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17613), .A(
        n17647), .ZN(n17629) );
  NOR2_X1 U20804 ( .A1(n17777), .A2(n17614), .ZN(n17631) );
  OAI211_X1 U20805 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17631), .B(n17615), .ZN(n17617) );
  NOR2_X1 U20806 ( .A1(n18181), .A2(n18847), .ZN(n17968) );
  INV_X1 U20807 ( .A(n17968), .ZN(n17616) );
  OAI211_X1 U20808 ( .C1(n17797), .C2(n17618), .A(n17617), .B(n17616), .ZN(
        n17619) );
  AOI21_X1 U20809 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17629), .A(
        n17619), .ZN(n17626) );
  AOI21_X1 U20810 ( .B1(n17964), .B2(n17621), .A(n17620), .ZN(n17970) );
  AOI21_X1 U20811 ( .B1(n17623), .B2(n17829), .A(n17622), .ZN(n17624) );
  XOR2_X1 U20812 ( .A(n17624), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17969) );
  AOI22_X1 U20813 ( .A1(n9589), .A2(n17970), .B1(n17824), .B2(n17969), .ZN(
        n17625) );
  OAI211_X1 U20814 ( .C1(n17751), .C2(n17973), .A(n17626), .B(n17625), .ZN(
        P3_U2805) );
  INV_X1 U20815 ( .A(n17627), .ZN(n17639) );
  NOR2_X1 U20816 ( .A1(n18181), .A2(n18845), .ZN(n17628) );
  AOI221_X1 U20817 ( .B1(n17631), .B2(n17630), .C1(n17629), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17628), .ZN(n17638) );
  INV_X1 U20818 ( .A(n17633), .ZN(n17632) );
  NOR2_X1 U20819 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17632), .ZN(
        n17974) );
  NAND2_X1 U20820 ( .A1(n18073), .A2(n17633), .ZN(n17975) );
  NAND2_X1 U20821 ( .A1(n17633), .A2(n18080), .ZN(n17976) );
  AOI22_X1 U20822 ( .A1(n17841), .A2(n17975), .B1(n9589), .B2(n17976), .ZN(
        n17651) );
  AOI21_X1 U20823 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17635), .A(
        n17634), .ZN(n17984) );
  OAI22_X1 U20824 ( .A1(n17651), .A2(n17938), .B1(n17984), .B2(n17844), .ZN(
        n17636) );
  AOI21_X1 U20825 ( .B1(n17666), .B2(n17974), .A(n17636), .ZN(n17637) );
  OAI211_X1 U20826 ( .C1(n17797), .C2(n17639), .A(n17638), .B(n17637), .ZN(
        P3_U2806) );
  INV_X1 U20827 ( .A(n17640), .ZN(n17641) );
  NAND2_X1 U20828 ( .A1(n17641), .A2(n17666), .ZN(n17652) );
  AOI22_X1 U20829 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17829), .B1(
        n17642), .B2(n17662), .ZN(n17643) );
  NAND2_X1 U20830 ( .A1(n17683), .A2(n17643), .ZN(n17644) );
  XOR2_X1 U20831 ( .A(n17644), .B(n17991), .Z(n17988) );
  NOR2_X1 U20832 ( .A1(n18181), .A2(n18844), .ZN(n17987) );
  NOR2_X1 U20833 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17645), .ZN(
        n17646) );
  OAI22_X1 U20834 ( .A1(n17915), .A2(n17648), .B1(n17647), .B2(n17646), .ZN(
        n17649) );
  AOI211_X1 U20835 ( .C1(n17988), .C2(n17824), .A(n17987), .B(n17649), .ZN(
        n17650) );
  OAI221_X1 U20836 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17652), 
        .C1(n17991), .C2(n17651), .A(n17650), .ZN(P3_U2807) );
  INV_X1 U20837 ( .A(n17932), .ZN(n17768) );
  AOI22_X1 U20838 ( .A1(n17768), .A2(n17653), .B1(n17834), .B2(n17655), .ZN(
        n17654) );
  NAND2_X1 U20839 ( .A1(n17654), .A2(n17931), .ZN(n17693) );
  AOI21_X1 U20840 ( .B1(n17687), .B2(n17685), .A(n17693), .ZN(n17675) );
  OR2_X1 U20841 ( .A1(n17655), .A2(n17777), .ZN(n17677) );
  OAI21_X1 U20842 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17656), .ZN(n17657) );
  OAI22_X1 U20843 ( .A1(n17675), .A2(n17658), .B1(n17677), .B2(n17657), .ZN(
        n17659) );
  AOI21_X1 U20844 ( .B1(n17772), .B2(n17660), .A(n17659), .ZN(n17669) );
  NOR2_X1 U20845 ( .A1(n17841), .A2(n9589), .ZN(n17694) );
  NAND2_X1 U20846 ( .A1(n17715), .A2(n17661), .ZN(n17993) );
  INV_X1 U20847 ( .A(n17993), .ZN(n17665) );
  INV_X1 U20848 ( .A(n18073), .ZN(n18001) );
  AOI22_X1 U20849 ( .A1(n17841), .A2(n18001), .B1(n9589), .B2(n18002), .ZN(
        n17740) );
  OAI21_X1 U20850 ( .B1(n17694), .B2(n17665), .A(n17740), .ZN(n17680) );
  INV_X1 U20851 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17998) );
  INV_X1 U20852 ( .A(n17662), .ZN(n17663) );
  OAI221_X1 U20853 ( .B1(n17663), .B2(n17665), .C1(n17663), .C2(n17730), .A(
        n17683), .ZN(n17664) );
  XOR2_X1 U20854 ( .A(n17998), .B(n17664), .Z(n18010) );
  AOI22_X1 U20855 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17680), .B1(
        n17824), .B2(n18010), .ZN(n17668) );
  NAND2_X1 U20856 ( .A1(n9593), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18011) );
  NAND3_X1 U20857 ( .A1(n17666), .A2(n17665), .A3(n17998), .ZN(n17667) );
  NAND4_X1 U20858 ( .A1(n17669), .A2(n17668), .A3(n18011), .A4(n17667), .ZN(
        P3_U2808) );
  NOR3_X1 U20859 ( .A1(n17829), .A2(n17709), .A3(n17670), .ZN(n17697) );
  INV_X1 U20860 ( .A(n17671), .ZN(n17717) );
  AOI22_X1 U20861 ( .A1(n18021), .A2(n17697), .B1(n17717), .B2(n17672), .ZN(
        n17673) );
  XOR2_X1 U20862 ( .A(n17673), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n18025) );
  NAND2_X1 U20863 ( .A1(n9593), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17674) );
  OAI221_X1 U20864 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17677), .C1(
        n17676), .C2(n17675), .A(n17674), .ZN(n17678) );
  AOI21_X1 U20865 ( .B1(n17772), .B2(n17679), .A(n17678), .ZN(n17682) );
  NOR2_X1 U20866 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17996), .ZN(
        n18015) );
  NOR2_X1 U20867 ( .A1(n18048), .A2(n17709), .ZN(n18017) );
  INV_X1 U20868 ( .A(n18017), .ZN(n18003) );
  NOR2_X1 U20869 ( .A1(n17741), .A2(n18003), .ZN(n17705) );
  AOI22_X1 U20870 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17680), .B1(
        n18015), .B2(n17705), .ZN(n17681) );
  OAI211_X1 U20871 ( .C1(n18025), .C2(n17844), .A(n17682), .B(n17681), .ZN(
        P3_U2809) );
  OAI221_X1 U20872 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17716), 
        .C1(n18034), .C2(n17697), .A(n17683), .ZN(n17684) );
  XOR2_X1 U20873 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17684), .Z(
        n18033) );
  OAI21_X1 U20874 ( .B1(n17686), .B2(n18395), .A(n17685), .ZN(n17692) );
  NOR2_X1 U20875 ( .A1(n18181), .A2(n18838), .ZN(n17691) );
  INV_X1 U20876 ( .A(n17688), .ZN(n17689) );
  AOI21_X1 U20877 ( .B1(n17797), .B2(n17613), .A(n17689), .ZN(n17690) );
  AOI211_X1 U20878 ( .C1(n17693), .C2(n17692), .A(n17691), .B(n17690), .ZN(
        n17696) );
  NOR2_X1 U20879 ( .A1(n18034), .A2(n18003), .ZN(n18005) );
  OAI21_X1 U20880 ( .B1(n17694), .B2(n18005), .A(n17740), .ZN(n17706) );
  NOR2_X1 U20881 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18034), .ZN(
        n18026) );
  AOI22_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17706), .B1(
        n18026), .B2(n17705), .ZN(n17695) );
  OAI211_X1 U20883 ( .C1(n17844), .C2(n18033), .A(n17696), .B(n17695), .ZN(
        P3_U2810) );
  AOI21_X1 U20884 ( .B1(n17717), .B2(n17716), .A(n17697), .ZN(n17698) );
  XOR2_X1 U20885 ( .A(n17698), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18039) );
  AOI21_X1 U20886 ( .B1(n17834), .B2(n17700), .A(n17903), .ZN(n17722) );
  OAI21_X1 U20887 ( .B1(n17699), .B2(n17932), .A(n17722), .ZN(n17712) );
  NOR2_X1 U20888 ( .A1(n17777), .A2(n17700), .ZN(n17714) );
  OAI211_X1 U20889 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17714), .B(n17701), .ZN(n17702) );
  NAND2_X1 U20890 ( .A1(n9593), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18037) );
  OAI211_X1 U20891 ( .C1(n17797), .C2(n17703), .A(n17702), .B(n18037), .ZN(
        n17704) );
  AOI21_X1 U20892 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17712), .A(
        n17704), .ZN(n17708) );
  AOI22_X1 U20893 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17706), .B1(
        n17705), .B2(n18034), .ZN(n17707) );
  OAI211_X1 U20894 ( .C1(n18039), .C2(n17844), .A(n17708), .B(n17707), .ZN(
        P3_U2811) );
  NAND2_X1 U20895 ( .A1(n17715), .A2(n17709), .ZN(n18054) );
  NAND2_X1 U20896 ( .A1(n9593), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18052) );
  OAI21_X1 U20897 ( .B1(n17797), .B2(n17710), .A(n18052), .ZN(n17711) );
  AOI221_X1 U20898 ( .B1(n17714), .B2(n17713), .C1(n17712), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17711), .ZN(n17720) );
  OAI21_X1 U20899 ( .B1(n17715), .B2(n17741), .A(n17740), .ZN(n17727) );
  AOI21_X1 U20900 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17818), .A(
        n17716), .ZN(n17718) );
  XOR2_X1 U20901 ( .A(n17718), .B(n17717), .Z(n18050) );
  AOI22_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17727), .B1(
        n17824), .B2(n18050), .ZN(n17719) );
  OAI211_X1 U20903 ( .C1(n17741), .C2(n18054), .A(n17720), .B(n17719), .ZN(
        P3_U2812) );
  NAND2_X1 U20904 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n20878), .ZN(
        n18060) );
  AOI21_X1 U20905 ( .B1(n18653), .B2(n9721), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17723) );
  OAI22_X1 U20906 ( .A1(n17723), .A2(n17722), .B1(n17915), .B2(n17721), .ZN(
        n17724) );
  AOI21_X1 U20907 ( .B1(n9593), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17724), .ZN(
        n17729) );
  OAI21_X1 U20908 ( .B1(n17726), .B2(n20878), .A(n17725), .ZN(n18057) );
  AOI22_X1 U20909 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17727), .B1(
        n17824), .B2(n18057), .ZN(n17728) );
  OAI211_X1 U20910 ( .C1(n17741), .C2(n18060), .A(n17729), .B(n17728), .ZN(
        P3_U2813) );
  NAND2_X1 U20911 ( .A1(n17818), .A2(n17747), .ZN(n17817) );
  OAI22_X1 U20912 ( .A1(n17818), .A2(n17730), .B1(n17817), .B2(n18016), .ZN(
        n17731) );
  XOR2_X1 U20913 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17731), .Z(
        n18067) );
  AOI21_X1 U20914 ( .B1(n17834), .B2(n17733), .A(n17903), .ZN(n17760) );
  OAI21_X1 U20915 ( .B1(n17732), .B2(n17932), .A(n17760), .ZN(n17744) );
  AOI22_X1 U20916 ( .A1(n9593), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17744), .ZN(n17736) );
  NOR2_X1 U20917 ( .A1(n17777), .A2(n17733), .ZN(n17746) );
  OAI211_X1 U20918 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17746), .B(n17734), .ZN(n17735) );
  OAI211_X1 U20919 ( .C1(n17737), .C2(n17797), .A(n17736), .B(n17735), .ZN(
        n17738) );
  AOI21_X1 U20920 ( .B1(n17824), .B2(n18067), .A(n17738), .ZN(n17739) );
  OAI221_X1 U20921 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17741), 
        .C1(n18070), .C2(n17740), .A(n17739), .ZN(P3_U2814) );
  AND2_X1 U20922 ( .A1(n18082), .A2(n18081), .ZN(n17756) );
  NAND2_X1 U20923 ( .A1(n9589), .A2(n18002), .ZN(n17755) );
  INV_X1 U20924 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17745) );
  OAI22_X1 U20925 ( .A1(n18181), .A2(n18828), .B1(n17797), .B2(n17742), .ZN(
        n17743) );
  AOI221_X1 U20926 ( .B1(n17746), .B2(n17745), .C1(n17744), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17743), .ZN(n17754) );
  NAND3_X1 U20927 ( .A1(n17747), .A2(n18106), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17748) );
  NAND3_X1 U20928 ( .A1(n9673), .A2(n17829), .A3(n18144), .ZN(n17808) );
  NOR2_X1 U20929 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17808), .ZN(
        n17802) );
  INV_X1 U20930 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18127) );
  NAND2_X1 U20931 ( .A1(n17802), .A2(n18127), .ZN(n17788) );
  AOI22_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17748), .B1(
        n17788), .B2(n17774), .ZN(n17749) );
  OAI221_X1 U20933 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18093), 
        .C1(n18113), .C2(n17818), .A(n17749), .ZN(n17750) );
  XOR2_X1 U20934 ( .A(n18082), .B(n17750), .Z(n18084) );
  NOR2_X1 U20935 ( .A1(n18073), .A2(n17751), .ZN(n17752) );
  OAI21_X1 U20936 ( .B1(n18075), .B2(n18119), .A(n18082), .ZN(n18078) );
  AOI22_X1 U20937 ( .A1(n17824), .A2(n18084), .B1(n17752), .B2(n18078), .ZN(
        n17753) );
  OAI211_X1 U20938 ( .C1(n17756), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        P3_U2815) );
  OAI21_X1 U20939 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17757), .A(
        n18081), .ZN(n18100) );
  AOI21_X1 U20940 ( .B1(n18653), .B2(n17758), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17759) );
  OAI22_X1 U20941 ( .A1(n17760), .A2(n17759), .B1(n18181), .B2(n18827), .ZN(
        n17761) );
  AOI21_X1 U20942 ( .B1(n17762), .B2(n17923), .A(n17761), .ZN(n17767) );
  NOR2_X1 U20943 ( .A1(n18119), .A2(n18075), .ZN(n17763) );
  AOI221_X1 U20944 ( .B1(n18092), .B2(n18093), .C1(n18119), .C2(n18093), .A(
        n17763), .ZN(n18097) );
  NAND2_X1 U20945 ( .A1(n18113), .A2(n17774), .ZN(n17764) );
  OAI22_X1 U20946 ( .A1(n18092), .A2(n17817), .B1(n17764), .B2(n17788), .ZN(
        n17765) );
  XOR2_X1 U20947 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17765), .Z(
        n18096) );
  AOI22_X1 U20948 ( .A1(n17841), .A2(n18097), .B1(n17824), .B2(n18096), .ZN(
        n17766) );
  OAI211_X1 U20949 ( .C1(n17937), .C2(n18100), .A(n17767), .B(n17766), .ZN(
        P3_U2816) );
  AOI21_X1 U20950 ( .B1(n17834), .B2(n17776), .A(n17768), .ZN(n17769) );
  OAI21_X1 U20951 ( .B1(n17770), .B2(n17769), .A(n17931), .ZN(n17784) );
  AOI22_X1 U20952 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17784), .B1(
        n17772), .B2(n17771), .ZN(n17782) );
  NOR2_X1 U20953 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18088), .ZN(
        n18101) );
  OR2_X1 U20954 ( .A1(n18125), .A2(n17817), .ZN(n17789) );
  AOI22_X1 U20955 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17789), .B1(
        n17788), .B2(n18113), .ZN(n17773) );
  XOR2_X1 U20956 ( .A(n17774), .B(n17773), .Z(n18110) );
  OR2_X1 U20957 ( .A1(n18119), .A2(n18088), .ZN(n18102) );
  OR2_X1 U20958 ( .A1(n18088), .A2(n18121), .ZN(n18103) );
  AOI22_X1 U20959 ( .A1(n17841), .A2(n18102), .B1(n9589), .B2(n18103), .ZN(
        n17791) );
  OAI22_X1 U20960 ( .A1(n18110), .A2(n17844), .B1(n17791), .B2(n17774), .ZN(
        n17775) );
  AOI21_X1 U20961 ( .B1(n18101), .B2(n17787), .A(n17775), .ZN(n17781) );
  NAND2_X1 U20962 ( .A1(n9593), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17780) );
  NOR2_X1 U20963 ( .A1(n17777), .A2(n17776), .ZN(n17786) );
  OAI211_X1 U20964 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17786), .B(n17778), .ZN(n17779) );
  NAND4_X1 U20965 ( .A1(n17782), .A2(n17781), .A3(n17780), .A4(n17779), .ZN(
        P3_U2817) );
  NOR2_X1 U20966 ( .A1(n18181), .A2(n18823), .ZN(n17783) );
  AOI221_X1 U20967 ( .B1(n17786), .B2(n17785), .C1(n17784), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17783), .ZN(n17795) );
  INV_X1 U20968 ( .A(n17787), .ZN(n17827) );
  NOR2_X1 U20969 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17827), .ZN(
        n17793) );
  NAND2_X1 U20970 ( .A1(n17789), .A2(n17788), .ZN(n17790) );
  XOR2_X1 U20971 ( .A(n17790), .B(n18113), .Z(n18117) );
  OAI22_X1 U20972 ( .A1(n17791), .A2(n18113), .B1(n18117), .B2(n17844), .ZN(
        n17792) );
  AOI21_X1 U20973 ( .B1(n17793), .B2(n18106), .A(n17792), .ZN(n17794) );
  OAI211_X1 U20974 ( .C1(n17797), .C2(n17796), .A(n17795), .B(n17794), .ZN(
        P3_U2818) );
  NAND2_X1 U20975 ( .A1(n18123), .A2(n18127), .ZN(n18133) );
  NOR2_X1 U20976 ( .A1(n18395), .A2(n17833), .ZN(n17866) );
  AND2_X1 U20977 ( .A1(n17798), .A2(n17866), .ZN(n17822) );
  NAND2_X1 U20978 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17822), .ZN(
        n17807) );
  INV_X1 U20979 ( .A(n17928), .ZN(n17856) );
  NAND3_X1 U20980 ( .A1(n17856), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17807), .ZN(n17799) );
  NAND2_X1 U20981 ( .A1(n9593), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18131) );
  OAI211_X1 U20982 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17807), .A(
        n17799), .B(n18131), .ZN(n17800) );
  AOI21_X1 U20983 ( .B1(n17801), .B2(n17923), .A(n17800), .ZN(n17806) );
  AOI22_X1 U20984 ( .A1(n17841), .A2(n18119), .B1(n9589), .B2(n18121), .ZN(
        n17826) );
  OAI21_X1 U20985 ( .B1(n18123), .B2(n17827), .A(n17826), .ZN(n17814) );
  NOR2_X1 U20986 ( .A1(n18144), .A2(n17817), .ZN(n17803) );
  AOI21_X1 U20987 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17803), .A(
        n17802), .ZN(n17804) );
  XOR2_X1 U20988 ( .A(n18127), .B(n17804), .Z(n18130) );
  AOI22_X1 U20989 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17814), .B1(
        n17824), .B2(n18130), .ZN(n17805) );
  OAI211_X1 U20990 ( .C1(n17827), .C2(n18133), .A(n17806), .B(n17805), .ZN(
        P3_U2819) );
  OAI21_X1 U20991 ( .B1(n17827), .B2(n18144), .A(n18137), .ZN(n17813) );
  INV_X1 U20992 ( .A(n17807), .ZN(n17811) );
  AOI21_X1 U20993 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17856), .A(
        n17822), .ZN(n17810) );
  OAI21_X1 U20994 ( .B1(n18144), .B2(n17817), .A(n17808), .ZN(n17809) );
  XOR2_X1 U20995 ( .A(n17809), .B(n18137), .Z(n18141) );
  OAI22_X1 U20996 ( .A1(n17811), .A2(n17810), .B1(n18141), .B2(n17844), .ZN(
        n17812) );
  AOI21_X1 U20997 ( .B1(n17814), .B2(n17813), .A(n17812), .ZN(n17815) );
  NAND2_X1 U20998 ( .A1(n9593), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18139) );
  OAI211_X1 U20999 ( .C1(n17915), .C2(n17816), .A(n17815), .B(n18139), .ZN(
        P3_U2820) );
  XOR2_X1 U21000 ( .A(n17819), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18149) );
  NOR2_X1 U21001 ( .A1(n18181), .A2(n18817), .ZN(n18148) );
  AOI22_X1 U21002 ( .A1(n17831), .A2(n17866), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17856), .ZN(n17821) );
  OAI22_X1 U21003 ( .A1(n17822), .A2(n17821), .B1(n17915), .B2(n17820), .ZN(
        n17823) );
  AOI211_X1 U21004 ( .C1(n17824), .C2(n18149), .A(n18148), .B(n17823), .ZN(
        n17825) );
  OAI221_X1 U21005 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17827), .C1(
        n18144), .C2(n17826), .A(n17825), .ZN(P3_U2821) );
  OAI21_X1 U21006 ( .B1(n18165), .B2(n17829), .A(n17828), .ZN(n18168) );
  NAND2_X1 U21007 ( .A1(n17830), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17832) );
  AOI211_X1 U21008 ( .C1(n17835), .C2(n17832), .A(n17831), .B(n18395), .ZN(
        n17837) );
  AOI21_X1 U21009 ( .B1(n17834), .B2(n17833), .A(n17903), .ZN(n17845) );
  OAI22_X1 U21010 ( .A1(n17845), .A2(n17835), .B1(n18181), .B2(n18816), .ZN(
        n17836) );
  AOI211_X1 U21011 ( .C1(n17838), .C2(n17923), .A(n17837), .B(n17836), .ZN(
        n17843) );
  AOI21_X1 U21012 ( .B1(n17840), .B2(n18161), .A(n17839), .ZN(n18163) );
  AOI22_X1 U21013 ( .A1(n17841), .A2(n18165), .B1(n9589), .B2(n18163), .ZN(
        n17842) );
  OAI211_X1 U21014 ( .C1(n17844), .C2(n18168), .A(n17843), .B(n17842), .ZN(
        P3_U2822) );
  INV_X1 U21015 ( .A(n17845), .ZN(n17846) );
  NOR2_X1 U21016 ( .A1(n18181), .A2(n18813), .ZN(n18177) );
  AOI221_X1 U21017 ( .B1(n17866), .B2(n17847), .C1(n17846), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18177), .ZN(n17854) );
  AOI21_X1 U21018 ( .B1(n18173), .B2(n17849), .A(n17848), .ZN(n18178) );
  NAND2_X1 U21019 ( .A1(n17851), .A2(n17850), .ZN(n17852) );
  XOR2_X1 U21020 ( .A(n17852), .B(n18173), .Z(n18176) );
  AOI22_X1 U21021 ( .A1(n17920), .A2(n18178), .B1(n9589), .B2(n18176), .ZN(
        n17853) );
  OAI211_X1 U21022 ( .C1(n17915), .C2(n17855), .A(n17854), .B(n17853), .ZN(
        P3_U2823) );
  AOI22_X1 U21023 ( .A1(n18653), .A2(n17876), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17856), .ZN(n17865) );
  AOI22_X1 U21024 ( .A1(n9593), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17857), .B2(
        n17923), .ZN(n17864) );
  AOI21_X1 U21025 ( .B1(n17860), .B2(n17859), .A(n17858), .ZN(n18185) );
  AOI21_X1 U21026 ( .B1(n18188), .B2(n17862), .A(n17861), .ZN(n18184) );
  AOI22_X1 U21027 ( .A1(n17920), .A2(n18185), .B1(n9589), .B2(n18184), .ZN(
        n17863) );
  OAI211_X1 U21028 ( .C1(n17866), .C2(n17865), .A(n17864), .B(n17863), .ZN(
        P3_U2824) );
  AOI21_X1 U21029 ( .B1(n17869), .B2(n17868), .A(n17867), .ZN(n18192) );
  AOI22_X1 U21030 ( .A1(n9589), .A2(n18192), .B1(n9593), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17880) );
  OAI21_X1 U21031 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n17873) );
  XOR2_X1 U21032 ( .A(n17873), .B(n18198), .Z(n18194) );
  AOI221_X1 U21033 ( .B1(n17903), .B2(n17875), .C1(n17874), .C2(n17875), .A(
        n17928), .ZN(n17878) );
  NAND2_X1 U21034 ( .A1(n18653), .A2(n17876), .ZN(n17877) );
  AOI22_X1 U21035 ( .A1(n17920), .A2(n18194), .B1(n17878), .B2(n17877), .ZN(
        n17879) );
  OAI211_X1 U21036 ( .C1(n17915), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        P3_U2825) );
  OAI21_X1 U21037 ( .B1(n17884), .B2(n17883), .A(n17882), .ZN(n17885) );
  XOR2_X1 U21038 ( .A(n17885), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18201) );
  AOI21_X1 U21039 ( .B1(n17888), .B2(n17887), .A(n17886), .ZN(n18203) );
  OAI22_X1 U21040 ( .A1(n18181), .A2(n18807), .B1(n18395), .B2(n17889), .ZN(
        n17890) );
  AOI21_X1 U21041 ( .B1(n17920), .B2(n18203), .A(n17890), .ZN(n17895) );
  OAI21_X1 U21042 ( .B1(n17892), .B2(n17891), .A(n17931), .ZN(n17905) );
  AOI22_X1 U21043 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17905), .B1(
        n17893), .B2(n17923), .ZN(n17894) );
  OAI211_X1 U21044 ( .C1(n17937), .C2(n18201), .A(n17895), .B(n17894), .ZN(
        P3_U2826) );
  AOI21_X1 U21045 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n18208) );
  AOI22_X1 U21046 ( .A1(n17920), .A2(n18208), .B1(n9593), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17907) );
  AOI21_X1 U21047 ( .B1(n17901), .B2(n17900), .A(n17899), .ZN(n18209) );
  OAI21_X1 U21048 ( .B1(n17903), .B2(n17918), .A(n17902), .ZN(n17904) );
  AOI22_X1 U21049 ( .A1(n9589), .A2(n18209), .B1(n17905), .B2(n17904), .ZN(
        n17906) );
  OAI211_X1 U21050 ( .C1(n17915), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2827) );
  AOI21_X1 U21051 ( .B1(n17911), .B2(n17910), .A(n17909), .ZN(n18224) );
  INV_X1 U21052 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18803) );
  NOR2_X1 U21053 ( .A1(n18181), .A2(n18803), .ZN(n18229) );
  XNOR2_X1 U21054 ( .A(n17913), .B(n17912), .ZN(n18227) );
  OAI22_X1 U21055 ( .A1(n17915), .A2(n17914), .B1(n17937), .B2(n18227), .ZN(
        n17916) );
  AOI211_X1 U21056 ( .C1(n17920), .C2(n18224), .A(n18229), .B(n17916), .ZN(
        n17917) );
  OAI221_X1 U21057 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18395), .C1(
        n17918), .C2(n17931), .A(n17917), .ZN(P3_U2828) );
  AOI21_X1 U21058 ( .B1(n17929), .B2(n17921), .A(n17919), .ZN(n18237) );
  AOI22_X1 U21059 ( .A1(n17920), .A2(n18237), .B1(n9593), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17926) );
  NOR2_X1 U21060 ( .A1(n17930), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17922) );
  XNOR2_X1 U21061 ( .A(n17922), .B(n17921), .ZN(n18235) );
  AOI22_X1 U21062 ( .A1(n9589), .A2(n18235), .B1(n17927), .B2(n17923), .ZN(
        n17925) );
  OAI211_X1 U21063 ( .C1(n17928), .C2(n17927), .A(n17926), .B(n17925), .ZN(
        P3_U2829) );
  OAI21_X1 U21064 ( .B1(n17930), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17929), .ZN(n17936) );
  INV_X1 U21065 ( .A(n17936), .ZN(n18252) );
  NAND3_X1 U21066 ( .A1(n18885), .A2(n17932), .A3(n17931), .ZN(n17933) );
  AOI22_X1 U21067 ( .A1(n9593), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17933), .ZN(n17934) );
  OAI221_X1 U21068 ( .B1(n18252), .B2(n17937), .C1(n17936), .C2(n17935), .A(
        n17934), .ZN(P3_U2830) );
  NAND2_X1 U21069 ( .A1(n18181), .A2(n18248), .ZN(n18233) );
  NOR2_X1 U21070 ( .A1(n17991), .A2(n17938), .ZN(n17940) );
  NOR2_X1 U21071 ( .A1(n9588), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18217) );
  NOR2_X1 U21072 ( .A1(n18217), .A2(n17939), .ZN(n17978) );
  NAND2_X1 U21073 ( .A1(n18745), .A2(n9588), .ZN(n18218) );
  INV_X1 U21074 ( .A(n18218), .ZN(n18049) );
  AOI21_X1 U21075 ( .B1(n17940), .B2(n17978), .A(n18049), .ZN(n17960) );
  AOI22_X1 U21076 ( .A1(n18726), .A2(n17964), .B1(n18743), .B2(n17941), .ZN(
        n17943) );
  OAI211_X1 U21077 ( .C1(n17944), .C2(n18228), .A(n17943), .B(n17942), .ZN(
        n17945) );
  OAI211_X1 U21078 ( .C1(n18745), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17954), .ZN(n17949) );
  OAI21_X1 U21079 ( .B1(n18248), .B2(n10178), .A(n17947), .ZN(n17948) );
  AOI22_X1 U21080 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18239), .B1(
        n17949), .B2(n17948), .ZN(n17951) );
  NAND2_X1 U21081 ( .A1(n9593), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17950) );
  OAI211_X1 U21082 ( .C1(n17952), .C2(n18169), .A(n17951), .B(n17950), .ZN(
        P3_U2835) );
  AOI211_X1 U21083 ( .C1(n18231), .C2(n17954), .A(n9593), .B(n17953), .ZN(
        n17955) );
  AOI21_X1 U21084 ( .B1(n17956), .B2(n18014), .A(n17955), .ZN(n17958) );
  NAND2_X1 U21085 ( .A1(n9593), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17957) );
  OAI211_X1 U21086 ( .C1(n17959), .C2(n18169), .A(n17958), .B(n17957), .ZN(
        P3_U2836) );
  AOI221_X1 U21087 ( .B1(n17961), .B2(n18717), .C1(n18004), .C2(n18717), .A(
        n17960), .ZN(n17966) );
  NAND2_X1 U21088 ( .A1(n17963), .A2(n17962), .ZN(n17965) );
  AOI221_X1 U21089 ( .B1(n17966), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17965), .C2(n17964), .A(n18248), .ZN(n17967) );
  AOI211_X1 U21090 ( .C1(n18239), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17968), .B(n17967), .ZN(n17972) );
  AOI22_X1 U21091 ( .A1(n18236), .A2(n17970), .B1(n18150), .B2(n17969), .ZN(
        n17971) );
  OAI211_X1 U21092 ( .C1(n18040), .C2(n17973), .A(n17972), .B(n17971), .ZN(
        P3_U2837) );
  AOI22_X1 U21093 ( .A1(n9593), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18014), 
        .B2(n17974), .ZN(n17983) );
  INV_X1 U21094 ( .A(n18158), .ZN(n18065) );
  AOI22_X1 U21095 ( .A1(n18706), .A2(n17976), .B1(n18120), .B2(n17975), .ZN(
        n17977) );
  OAI211_X1 U21096 ( .C1(n18049), .C2(n17978), .A(n17977), .B(n18233), .ZN(
        n17981) );
  AOI211_X1 U21097 ( .C1(n18717), .C2(n17979), .A(n17991), .B(n17981), .ZN(
        n17980) );
  NOR2_X1 U21098 ( .A1(n9593), .A2(n17980), .ZN(n17985) );
  OAI211_X1 U21099 ( .C1(n18065), .C2(n17981), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17985), .ZN(n17982) );
  OAI211_X1 U21100 ( .C1(n17984), .C2(n18169), .A(n17983), .B(n17982), .ZN(
        P3_U2838) );
  INV_X1 U21101 ( .A(n17985), .ZN(n17992) );
  NOR2_X1 U21102 ( .A1(n17986), .A2(n17993), .ZN(n18009) );
  NAND3_X1 U21103 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18009), .A3(
        n18233), .ZN(n17990) );
  AOI21_X1 U21104 ( .B1(n17988), .B2(n18150), .A(n17987), .ZN(n17989) );
  OAI221_X1 U21105 ( .B1(n17992), .B2(n17991), .C1(n17992), .C2(n17990), .A(
        n17989), .ZN(P3_U2839) );
  NOR2_X1 U21106 ( .A1(n18706), .A2(n18120), .ZN(n18122) );
  INV_X1 U21107 ( .A(n18122), .ZN(n18047) );
  AOI22_X1 U21108 ( .A1(n18726), .A2(n17994), .B1(n17993), .B2(n18047), .ZN(
        n18020) );
  AOI22_X1 U21109 ( .A1(n18717), .A2(n17996), .B1(n18126), .B2(n17995), .ZN(
        n18000) );
  OAI21_X1 U21110 ( .B1(n17998), .B2(n18743), .A(n17997), .ZN(n17999) );
  NAND3_X1 U21111 ( .A1(n18020), .A2(n18000), .A3(n17999), .ZN(n18008) );
  AOI22_X1 U21112 ( .A1(n18706), .A2(n18002), .B1(n18120), .B2(n18001), .ZN(
        n18042) );
  OAI21_X1 U21113 ( .B1(n18004), .B2(n18003), .A(n18717), .ZN(n18007) );
  INV_X1 U21114 ( .A(n18005), .ZN(n18027) );
  OAI21_X1 U21115 ( .B1(n18043), .B2(n18027), .A(n18726), .ZN(n18006) );
  NAND3_X1 U21116 ( .A1(n18042), .A2(n18007), .A3(n18006), .ZN(n18018) );
  OAI22_X1 U21117 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18009), .B1(
        n18008), .B2(n18018), .ZN(n18013) );
  AOI22_X1 U21118 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18239), .B1(
        n18150), .B2(n18010), .ZN(n18012) );
  OAI211_X1 U21119 ( .C1(n18248), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        P3_U2840) );
  AND2_X1 U21120 ( .A1(n18014), .A2(n18017), .ZN(n18035) );
  AOI22_X1 U21121 ( .A1(n9593), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18035), 
        .B2(n18015), .ZN(n18024) );
  NOR2_X1 U21122 ( .A1(n18717), .A2(n18743), .ZN(n18238) );
  NAND2_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18062), .ZN(
        n18143) );
  NOR2_X1 U21124 ( .A1(n18016), .A2(n18143), .ZN(n18064) );
  AOI21_X1 U21125 ( .B1(n18017), .B2(n18064), .A(n9588), .ZN(n18019) );
  NOR3_X1 U21126 ( .A1(n18019), .A2(n18018), .A3(n18248), .ZN(n18029) );
  OAI211_X1 U21127 ( .C1(n18021), .C2(n18238), .A(n18029), .B(n18020), .ZN(
        n18022) );
  NAND3_X1 U21128 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18181), .A3(
        n18022), .ZN(n18023) );
  OAI211_X1 U21129 ( .C1(n18025), .C2(n18169), .A(n18024), .B(n18023), .ZN(
        P3_U2841) );
  AOI22_X1 U21130 ( .A1(n9593), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18035), 
        .B2(n18026), .ZN(n18032) );
  NAND2_X1 U21131 ( .A1(n18047), .A2(n18027), .ZN(n18028) );
  AOI21_X1 U21132 ( .B1(n18029), .B2(n18028), .A(n9593), .ZN(n18036) );
  NOR3_X1 U21133 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18238), .A3(
        n18938), .ZN(n18030) );
  OAI21_X1 U21134 ( .B1(n18036), .B2(n18030), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18031) );
  OAI211_X1 U21135 ( .C1(n18033), .C2(n18169), .A(n18032), .B(n18031), .ZN(
        P3_U2842) );
  AOI22_X1 U21136 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18036), .B1(
        n18035), .B2(n18034), .ZN(n18038) );
  OAI211_X1 U21137 ( .C1(n18039), .C2(n18169), .A(n18038), .B(n18037), .ZN(
        P3_U2843) );
  OAI22_X1 U21138 ( .A1(n18154), .A2(n18738), .B1(n18215), .B2(n18155), .ZN(
        n18211) );
  INV_X1 U21139 ( .A(n18211), .ZN(n18171) );
  NOR2_X1 U21140 ( .A1(n18248), .A2(n18171), .ZN(n18199) );
  INV_X1 U21141 ( .A(n18199), .ZN(n18186) );
  OAI222_X1 U21142 ( .A1(n18186), .A2(n18074), .B1(n18251), .B2(n18121), .C1(
        n18119), .C2(n18040), .ZN(n18111) );
  NAND2_X1 U21143 ( .A1(n18041), .A2(n18111), .ZN(n18071) );
  NAND2_X1 U21144 ( .A1(n18231), .A2(n18042), .ZN(n18066) );
  NOR3_X1 U21145 ( .A1(n18217), .A2(n18043), .A3(n18070), .ZN(n18045) );
  OAI22_X1 U21146 ( .A1(n18049), .A2(n18045), .B1(n18044), .B2(n18738), .ZN(
        n18046) );
  AOI211_X1 U21147 ( .C1(n18048), .C2(n18047), .A(n18066), .B(n18046), .ZN(
        n18055) );
  AOI221_X1 U21148 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18055), 
        .C1(n18049), .C2(n18055), .A(n9593), .ZN(n18051) );
  AOI22_X1 U21149 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18051), .B1(
        n18150), .B2(n18050), .ZN(n18053) );
  OAI211_X1 U21150 ( .C1(n18071), .C2(n18054), .A(n18053), .B(n18052), .ZN(
        P3_U2844) );
  NOR3_X1 U21151 ( .A1(n9593), .A2(n18055), .A3(n20878), .ZN(n18056) );
  AOI21_X1 U21152 ( .B1(n18150), .B2(n18057), .A(n18056), .ZN(n18059) );
  NAND2_X1 U21153 ( .A1(n9593), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18058) );
  OAI211_X1 U21154 ( .C1(n18060), .C2(n18071), .A(n18059), .B(n18058), .ZN(
        P3_U2845) );
  OAI22_X1 U21155 ( .A1(n18745), .A2(n18062), .B1(n18061), .B2(n18738), .ZN(
        n18118) );
  AOI21_X1 U21156 ( .B1(n18126), .B2(n18075), .A(n18118), .ZN(n18063) );
  OAI211_X1 U21157 ( .C1(n18064), .C2(n9588), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18063), .ZN(n18077) );
  OAI221_X1 U21158 ( .B1(n18066), .B2(n18065), .C1(n18066), .C2(n18077), .A(
        n18181), .ZN(n18069) );
  AOI22_X1 U21159 ( .A1(n9593), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18150), 
        .B2(n18067), .ZN(n18068) );
  OAI221_X1 U21160 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18071), 
        .C1(n18070), .C2(n18069), .A(n18068), .ZN(P3_U2846) );
  NOR2_X1 U21161 ( .A1(n18073), .A2(n18072), .ZN(n18079) );
  OR2_X1 U21162 ( .A1(n18074), .A2(n18171), .ZN(n18091) );
  OAI21_X1 U21163 ( .B1(n18075), .B2(n18091), .A(n18082), .ZN(n18076) );
  AOI22_X1 U21164 ( .A1(n18079), .A2(n18078), .B1(n18077), .B2(n18076), .ZN(
        n18087) );
  AOI22_X1 U21165 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18239), .B1(
        n9593), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18086) );
  AOI211_X1 U21166 ( .C1(n18082), .C2(n18081), .A(n18080), .B(n18251), .ZN(
        n18083) );
  AOI21_X1 U21167 ( .B1(n18084), .B2(n18150), .A(n18083), .ZN(n18085) );
  OAI211_X1 U21168 ( .C1(n18087), .C2(n18248), .A(n18086), .B(n18085), .ZN(
        P3_U2847) );
  AOI221_X1 U21169 ( .B1(n18088), .B2(n18743), .C1(n18143), .C2(n18743), .A(
        n18118), .ZN(n18105) );
  OAI21_X1 U21170 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18238), .A(
        n18105), .ZN(n18089) );
  AOI211_X1 U21171 ( .C1(n18126), .C2(n18092), .A(n18093), .B(n18089), .ZN(
        n18090) );
  AOI221_X1 U21172 ( .B1(n18092), .B2(n18093), .C1(n18091), .C2(n18093), .A(
        n18090), .ZN(n18095) );
  OAI22_X1 U21173 ( .A1(n18093), .A2(n18233), .B1(n18181), .B2(n18827), .ZN(
        n18094) );
  AOI21_X1 U21174 ( .B1(n18231), .B2(n18095), .A(n18094), .ZN(n18099) );
  AOI22_X1 U21175 ( .A1(n18164), .A2(n18097), .B1(n18150), .B2(n18096), .ZN(
        n18098) );
  OAI211_X1 U21176 ( .C1(n18251), .C2(n18100), .A(n18099), .B(n18098), .ZN(
        P3_U2848) );
  AOI22_X1 U21177 ( .A1(n9593), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18101), 
        .B2(n18111), .ZN(n18109) );
  INV_X1 U21178 ( .A(n18126), .ZN(n18135) );
  AOI22_X1 U21179 ( .A1(n18706), .A2(n18103), .B1(n18120), .B2(n18102), .ZN(
        n18104) );
  OAI211_X1 U21180 ( .C1(n18135), .C2(n18106), .A(n18105), .B(n18104), .ZN(
        n18114) );
  OAI21_X1 U21181 ( .B1(n18135), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18231), .ZN(n18107) );
  OAI211_X1 U21182 ( .C1(n18114), .C2(n18107), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18181), .ZN(n18108) );
  OAI211_X1 U21183 ( .C1(n18110), .C2(n18169), .A(n18109), .B(n18108), .ZN(
        P3_U2849) );
  AOI22_X1 U21184 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18239), .B1(
        n9593), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n18116) );
  INV_X1 U21185 ( .A(n18111), .ZN(n18152) );
  OAI22_X1 U21186 ( .A1(n18152), .A2(n18125), .B1(n18113), .B2(n18248), .ZN(
        n18112) );
  OAI21_X1 U21187 ( .B1(n18114), .B2(n18113), .A(n18112), .ZN(n18115) );
  OAI211_X1 U21188 ( .C1(n18117), .C2(n18169), .A(n18116), .B(n18115), .ZN(
        P3_U2850) );
  OR2_X1 U21189 ( .A1(n18743), .A2(n18118), .ZN(n18142) );
  AOI22_X1 U21190 ( .A1(n18706), .A2(n18121), .B1(n18120), .B2(n18119), .ZN(
        n18146) );
  OAI211_X1 U21191 ( .C1(n18123), .C2(n18122), .A(n18146), .B(n18233), .ZN(
        n18124) );
  AOI221_X1 U21192 ( .B1(n18144), .B2(n18142), .C1(n18143), .C2(n18142), .A(
        n18124), .ZN(n18134) );
  AOI22_X1 U21193 ( .A1(n18126), .A2(n18125), .B1(n18743), .B2(n18137), .ZN(
        n18128) );
  AOI211_X1 U21194 ( .C1(n18134), .C2(n18128), .A(n9593), .B(n18127), .ZN(
        n18129) );
  AOI21_X1 U21195 ( .B1(n18150), .B2(n18130), .A(n18129), .ZN(n18132) );
  OAI211_X1 U21196 ( .C1(n18152), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        P3_U2851) );
  AOI221_X1 U21197 ( .B1(n18135), .B2(n18134), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18134), .A(n9593), .ZN(n18138) );
  OAI21_X1 U21198 ( .B1(n18144), .B2(n18152), .A(n18137), .ZN(n18136) );
  OAI21_X1 U21199 ( .B1(n18138), .B2(n18137), .A(n18136), .ZN(n18140) );
  OAI211_X1 U21200 ( .C1(n18141), .C2(n18169), .A(n18140), .B(n18139), .ZN(
        P3_U2852) );
  AOI21_X1 U21201 ( .B1(n18143), .B2(n18142), .A(n18248), .ZN(n18145) );
  AOI211_X1 U21202 ( .C1(n18146), .C2(n18145), .A(n9593), .B(n18144), .ZN(
        n18147) );
  AOI211_X1 U21203 ( .C1(n18150), .C2(n18149), .A(n18148), .B(n18147), .ZN(
        n18151) );
  OAI21_X1 U21204 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18152), .A(
        n18151), .ZN(P3_U2853) );
  AND2_X1 U21205 ( .A1(n18153), .A2(n18199), .ZN(n18162) );
  AND2_X1 U21206 ( .A1(n18717), .A2(n18154), .ZN(n18223) );
  AOI211_X1 U21207 ( .C1(n18218), .C2(n18155), .A(n18223), .B(n18217), .ZN(
        n18200) );
  OAI21_X1 U21208 ( .B1(n18158), .B2(n18156), .A(n18200), .ZN(n18182) );
  OAI21_X1 U21209 ( .B1(n18158), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18157) );
  OAI21_X1 U21210 ( .B1(n18182), .B2(n18157), .A(n18231), .ZN(n18172) );
  OAI21_X1 U21211 ( .B1(n18158), .B2(n18172), .A(n18233), .ZN(n18160) );
  NOR2_X1 U21212 ( .A1(n18181), .A2(n18816), .ZN(n18159) );
  AOI221_X1 U21213 ( .B1(n18162), .B2(n18161), .C1(n18160), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18159), .ZN(n18167) );
  AOI22_X1 U21214 ( .A1(n18165), .A2(n18164), .B1(n18236), .B2(n18163), .ZN(
        n18166) );
  OAI211_X1 U21215 ( .C1(n18169), .C2(n18168), .A(n18167), .B(n18166), .ZN(
        P3_U2854) );
  OAI21_X1 U21216 ( .B1(n18171), .B2(n18170), .A(n18173), .ZN(n18175) );
  OAI21_X1 U21217 ( .B1(n18233), .B2(n18173), .A(n18172), .ZN(n18174) );
  AOI22_X1 U21218 ( .A1(n18236), .A2(n18176), .B1(n18175), .B2(n18174), .ZN(
        n18180) );
  AOI21_X1 U21219 ( .B1(n18178), .B2(n18247), .A(n18177), .ZN(n18179) );
  NAND2_X1 U21220 ( .A1(n18180), .A2(n18179), .ZN(P3_U2855) );
  OAI21_X1 U21221 ( .B1(n18248), .B2(n18182), .A(n18181), .ZN(n18197) );
  OAI22_X1 U21222 ( .A1(n18188), .A2(n18197), .B1(n18181), .B2(n18811), .ZN(
        n18183) );
  INV_X1 U21223 ( .A(n18183), .ZN(n18191) );
  AOI22_X1 U21224 ( .A1(n18247), .A2(n18185), .B1(n18236), .B2(n18184), .ZN(
        n18190) );
  NOR3_X1 U21225 ( .A1(n18206), .A2(n18187), .A3(n18186), .ZN(n18193) );
  NAND3_X1 U21226 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18193), .A3(
        n18188), .ZN(n18189) );
  NAND3_X1 U21227 ( .A1(n18191), .A2(n18190), .A3(n18189), .ZN(P3_U2856) );
  AOI22_X1 U21228 ( .A1(n9593), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18236), .B2(
        n18192), .ZN(n18196) );
  AOI22_X1 U21229 ( .A1(n18194), .A2(n18247), .B1(n18193), .B2(n18198), .ZN(
        n18195) );
  OAI211_X1 U21230 ( .C1(n18198), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        P3_U2857) );
  NAND2_X1 U21231 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18199), .ZN(
        n18207) );
  NAND2_X1 U21232 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18200), .ZN(
        n18210) );
  AOI21_X1 U21233 ( .B1(n18240), .B2(n18210), .A(n18239), .ZN(n18205) );
  OAI22_X1 U21234 ( .A1(n18181), .A2(n18807), .B1(n18251), .B2(n18201), .ZN(
        n18202) );
  AOI21_X1 U21235 ( .B1(n18247), .B2(n18203), .A(n18202), .ZN(n18204) );
  OAI221_X1 U21236 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18207), .C1(
        n18206), .C2(n18205), .A(n18204), .ZN(P3_U2858) );
  AOI22_X1 U21237 ( .A1(n9593), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18247), .B2(
        n18208), .ZN(n18214) );
  AOI22_X1 U21238 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18239), .B1(
        n18236), .B2(n18209), .ZN(n18213) );
  OAI211_X1 U21239 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18211), .A(
        n18231), .B(n18210), .ZN(n18212) );
  NAND3_X1 U21240 ( .A1(n18214), .A2(n18213), .A3(n18212), .ZN(P3_U2859) );
  NOR2_X1 U21241 ( .A1(n18886), .A2(n18215), .ZN(n18221) );
  NOR3_X1 U21242 ( .A1(n18738), .A2(n18886), .A3(n18902), .ZN(n18216) );
  AOI211_X1 U21243 ( .C1(n18218), .C2(n18886), .A(n18217), .B(n18216), .ZN(
        n18219) );
  INV_X1 U21244 ( .A(n18219), .ZN(n18220) );
  MUX2_X1 U21245 ( .A(n18221), .B(n18220), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18222) );
  AOI211_X1 U21246 ( .C1(n18225), .C2(n18224), .A(n18223), .B(n18222), .ZN(
        n18226) );
  OAI21_X1 U21247 ( .B1(n18228), .B2(n18227), .A(n18226), .ZN(n18230) );
  AOI21_X1 U21248 ( .B1(n18231), .B2(n18230), .A(n18229), .ZN(n18232) );
  OAI21_X1 U21249 ( .B1(n18234), .B2(n18233), .A(n18232), .ZN(P3_U2860) );
  AOI22_X1 U21250 ( .A1(n18247), .A2(n18237), .B1(n18236), .B2(n18235), .ZN(
        n18244) );
  NAND2_X1 U21251 ( .A1(n9593), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18243) );
  NOR3_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18238), .A3(
        n18248), .ZN(n18245) );
  OAI21_X1 U21253 ( .B1(n18239), .B2(n18245), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18242) );
  OAI211_X1 U21254 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18726), .A(
        n18240), .B(n18886), .ZN(n18241) );
  NAND4_X1 U21255 ( .A1(n18244), .A2(n18243), .A3(n18242), .A4(n18241), .ZN(
        P3_U2861) );
  INV_X1 U21256 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18913) );
  NOR2_X1 U21257 ( .A1(n18181), .A2(n18913), .ZN(n18246) );
  AOI211_X1 U21258 ( .C1(n18247), .C2(n18252), .A(n18246), .B(n18245), .ZN(
        n18250) );
  OAI211_X1 U21259 ( .C1(n18726), .C2(n18248), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18181), .ZN(n18249) );
  OAI211_X1 U21260 ( .C1(n18252), .C2(n18251), .A(n18250), .B(n18249), .ZN(
        P3_U2862) );
  OAI211_X1 U21261 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18253), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18766)
         );
  OAI21_X1 U21262 ( .B1(n18256), .B2(n18254), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18255) );
  OAI221_X1 U21263 ( .B1(n18256), .B2(n18766), .C1(n18256), .C2(n18323), .A(
        n18255), .ZN(P3_U2863) );
  INV_X1 U21264 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18758) );
  NAND2_X1 U21265 ( .A1(n18758), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18418) );
  INV_X1 U21266 ( .A(n18418), .ZN(n18463) );
  NAND2_X1 U21267 ( .A1(n18755), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18529) );
  INV_X1 U21268 ( .A(n18529), .ZN(n18553) );
  NOR2_X1 U21269 ( .A1(n18463), .A2(n18553), .ZN(n18258) );
  OAI22_X1 U21270 ( .A1(n18259), .A2(n18758), .B1(n18258), .B2(n18257), .ZN(
        P3_U2866) );
  NOR2_X1 U21271 ( .A1(n18759), .A2(n18260), .ZN(P3_U2867) );
  NOR3_X1 U21272 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18755), .A3(
        n18758), .ZN(n18652) );
  NAND2_X1 U21273 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18652), .ZN(
        n18618) );
  INV_X1 U21274 ( .A(n18618), .ZN(n18697) );
  NOR2_X1 U21275 ( .A1(n18758), .A2(n18439), .ZN(n18651) );
  INV_X1 U21276 ( .A(n18651), .ZN(n18646) );
  NOR2_X2 U21277 ( .A1(n18646), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18624) );
  NOR2_X1 U21278 ( .A1(n18697), .A2(n18624), .ZN(n18619) );
  NOR2_X2 U21279 ( .A1(n18748), .A2(n18646), .ZN(n18645) );
  NAND2_X1 U21280 ( .A1(n18750), .A2(n18748), .ZN(n18751) );
  NAND2_X1 U21281 ( .A1(n18755), .A2(n18758), .ZN(n18349) );
  NOR2_X1 U21282 ( .A1(n18751), .A2(n18349), .ZN(n18373) );
  CLKBUF_X1 U21283 ( .A(n18373), .Z(n18390) );
  NOR2_X1 U21284 ( .A1(n18645), .A2(n18390), .ZN(n18351) );
  OAI22_X1 U21285 ( .A1(n18620), .A2(n18619), .B1(n18351), .B2(n18261), .ZN(
        n18262) );
  INV_X1 U21286 ( .A(n18394), .ZN(n18623) );
  AND2_X1 U21287 ( .A1(n18262), .A2(n18623), .ZN(n18321) );
  NOR2_X2 U21288 ( .A1(n18395), .A2(n18263), .ZN(n18654) );
  NOR2_X2 U21289 ( .A1(n18394), .A2(n18264), .ZN(n18648) );
  NOR2_X1 U21290 ( .A1(n18647), .A2(n18351), .ZN(n18314) );
  AOI22_X1 U21291 ( .A1(n18624), .A2(n18654), .B1(n18648), .B2(n18314), .ZN(
        n18269) );
  NOR2_X2 U21292 ( .A1(n18265), .A2(n18395), .ZN(n18649) );
  NAND2_X1 U21293 ( .A1(n18267), .A2(n18266), .ZN(n18315) );
  NOR2_X1 U21294 ( .A1(n18925), .A2(n18315), .ZN(n18322) );
  AOI22_X1 U21295 ( .A1(n18697), .A2(n18649), .B1(n18390), .B2(n18322), .ZN(
        n18268) );
  OAI211_X1 U21296 ( .C1(n18321), .C2(n18270), .A(n18269), .B(n18268), .ZN(
        P3_U2868) );
  NOR2_X2 U21297 ( .A1(n18395), .A2(n18271), .ZN(n18660) );
  NOR2_X2 U21298 ( .A1(n18394), .A2(n18272), .ZN(n18658) );
  AOI22_X1 U21299 ( .A1(n18624), .A2(n18660), .B1(n18314), .B2(n18658), .ZN(
        n18276) );
  NOR2_X2 U21300 ( .A1(n18273), .A2(n18395), .ZN(n18659) );
  NOR2_X1 U21301 ( .A1(n18274), .A2(n18315), .ZN(n18326) );
  AOI22_X1 U21302 ( .A1(n18697), .A2(n18659), .B1(n18373), .B2(n18326), .ZN(
        n18275) );
  OAI211_X1 U21303 ( .C1(n18321), .C2(n18277), .A(n18276), .B(n18275), .ZN(
        P3_U2869) );
  NOR2_X2 U21304 ( .A1(n18395), .A2(n18278), .ZN(n18665) );
  NOR2_X2 U21305 ( .A1(n18394), .A2(n18279), .ZN(n18664) );
  AOI22_X1 U21306 ( .A1(n18624), .A2(n18665), .B1(n18314), .B2(n18664), .ZN(
        n18283) );
  NOR2_X2 U21307 ( .A1(n18280), .A2(n18395), .ZN(n18666) );
  NOR2_X1 U21308 ( .A1(n18281), .A2(n18315), .ZN(n18329) );
  AOI22_X1 U21309 ( .A1(n18697), .A2(n18666), .B1(n18373), .B2(n18329), .ZN(
        n18282) );
  OAI211_X1 U21310 ( .C1(n18321), .C2(n18284), .A(n18283), .B(n18282), .ZN(
        P3_U2870) );
  NOR2_X2 U21311 ( .A1(n18285), .A2(n18395), .ZN(n18671) );
  NOR2_X2 U21312 ( .A1(n18394), .A2(n18286), .ZN(n18670) );
  AOI22_X1 U21313 ( .A1(n18697), .A2(n18671), .B1(n18314), .B2(n18670), .ZN(
        n18290) );
  NOR2_X1 U21314 ( .A1(n18287), .A2(n18315), .ZN(n18332) );
  NOR2_X2 U21315 ( .A1(n18395), .A2(n18288), .ZN(n18672) );
  AOI22_X1 U21316 ( .A1(n18373), .A2(n18332), .B1(n18624), .B2(n18672), .ZN(
        n18289) );
  OAI211_X1 U21317 ( .C1(n18321), .C2(n18291), .A(n18290), .B(n18289), .ZN(
        P3_U2871) );
  NOR2_X2 U21318 ( .A1(n18292), .A2(n18395), .ZN(n18678) );
  NOR2_X2 U21319 ( .A1(n20858), .A2(n18394), .ZN(n18676) );
  AOI22_X1 U21320 ( .A1(n18697), .A2(n18678), .B1(n18314), .B2(n18676), .ZN(
        n18296) );
  NOR2_X1 U21321 ( .A1(n18293), .A2(n18315), .ZN(n18335) );
  NOR2_X2 U21322 ( .A1(n18294), .A2(n18395), .ZN(n18677) );
  AOI22_X1 U21323 ( .A1(n18373), .A2(n18335), .B1(n18624), .B2(n18677), .ZN(
        n18295) );
  OAI211_X1 U21324 ( .C1(n18321), .C2(n18297), .A(n18296), .B(n18295), .ZN(
        P3_U2872) );
  NOR2_X2 U21325 ( .A1(n18298), .A2(n18395), .ZN(n18684) );
  NOR2_X2 U21326 ( .A1(n18299), .A2(n18394), .ZN(n18682) );
  AOI22_X1 U21327 ( .A1(n18697), .A2(n18684), .B1(n18314), .B2(n18682), .ZN(
        n18303) );
  NOR2_X1 U21328 ( .A1(n18300), .A2(n18315), .ZN(n18338) );
  NOR2_X2 U21329 ( .A1(n18301), .A2(n18395), .ZN(n18683) );
  AOI22_X1 U21330 ( .A1(n18390), .A2(n18338), .B1(n18624), .B2(n18683), .ZN(
        n18302) );
  OAI211_X1 U21331 ( .C1(n18321), .C2(n18304), .A(n18303), .B(n18302), .ZN(
        P3_U2873) );
  NOR2_X2 U21332 ( .A1(n18305), .A2(n18395), .ZN(n18690) );
  NOR2_X2 U21333 ( .A1(n18306), .A2(n18394), .ZN(n18688) );
  AOI22_X1 U21334 ( .A1(n18624), .A2(n18690), .B1(n18314), .B2(n18688), .ZN(
        n18310) );
  NOR2_X2 U21335 ( .A1(n18307), .A2(n18395), .ZN(n18689) );
  NOR2_X1 U21336 ( .A1(n18308), .A2(n18315), .ZN(n18341) );
  AOI22_X1 U21337 ( .A1(n18697), .A2(n18689), .B1(n18373), .B2(n18341), .ZN(
        n18309) );
  OAI211_X1 U21338 ( .C1(n18321), .C2(n18311), .A(n18310), .B(n18309), .ZN(
        P3_U2874) );
  NOR2_X2 U21339 ( .A1(n18395), .A2(n18312), .ZN(n18699) );
  NOR2_X2 U21340 ( .A1(n18313), .A2(n18394), .ZN(n18695) );
  AOI22_X1 U21341 ( .A1(n18697), .A2(n18699), .B1(n18314), .B2(n18695), .ZN(
        n18319) );
  NOR2_X1 U21342 ( .A1(n18316), .A2(n18315), .ZN(n18344) );
  NOR2_X2 U21343 ( .A1(n18317), .A2(n18395), .ZN(n18696) );
  AOI22_X1 U21344 ( .A1(n18390), .A2(n18344), .B1(n18624), .B2(n18696), .ZN(
        n18318) );
  OAI211_X1 U21345 ( .C1(n18321), .C2(n18320), .A(n18319), .B(n18318), .ZN(
        P3_U2875) );
  INV_X1 U21346 ( .A(n18349), .ZN(n18372) );
  NOR2_X1 U21347 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18748), .ZN(
        n18507) );
  NAND2_X1 U21348 ( .A1(n18372), .A2(n18507), .ZN(n18350) );
  NAND2_X1 U21349 ( .A1(n18750), .A2(n18776), .ZN(n18508) );
  NOR2_X1 U21350 ( .A1(n18349), .A2(n18508), .ZN(n18345) );
  AOI22_X1 U21351 ( .A1(n18645), .A2(n18654), .B1(n18648), .B2(n18345), .ZN(
        n18325) );
  AND2_X1 U21352 ( .A1(n18623), .A2(n18323), .ZN(n18650) );
  AND2_X1 U21353 ( .A1(n18750), .A2(n18650), .ZN(n18596) );
  AOI22_X1 U21354 ( .A1(n18653), .A2(n18651), .B1(n18372), .B2(n18596), .ZN(
        n18346) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18346), .B1(
        n18649), .B2(n18624), .ZN(n18324) );
  OAI211_X1 U21356 ( .C1(n18657), .C2(n18350), .A(n18325), .B(n18324), .ZN(
        P3_U2876) );
  INV_X1 U21357 ( .A(n18326), .ZN(n18663) );
  AOI22_X1 U21358 ( .A1(n18624), .A2(n18659), .B1(n18658), .B2(n18345), .ZN(
        n18328) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18346), .B1(
        n18645), .B2(n18660), .ZN(n18327) );
  OAI211_X1 U21360 ( .C1(n18663), .C2(n18350), .A(n18328), .B(n18327), .ZN(
        P3_U2877) );
  INV_X1 U21361 ( .A(n18329), .ZN(n18669) );
  AOI22_X1 U21362 ( .A1(n18624), .A2(n18666), .B1(n18664), .B2(n18345), .ZN(
        n18331) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18346), .B1(
        n18645), .B2(n18665), .ZN(n18330) );
  OAI211_X1 U21364 ( .C1(n18669), .C2(n18350), .A(n18331), .B(n18330), .ZN(
        P3_U2878) );
  INV_X1 U21365 ( .A(n18332), .ZN(n18675) );
  AOI22_X1 U21366 ( .A1(n18645), .A2(n18672), .B1(n18670), .B2(n18345), .ZN(
        n18334) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18346), .B1(
        n18624), .B2(n18671), .ZN(n18333) );
  OAI211_X1 U21368 ( .C1(n18675), .C2(n18350), .A(n18334), .B(n18333), .ZN(
        P3_U2879) );
  AOI22_X1 U21369 ( .A1(n18645), .A2(n18677), .B1(n18676), .B2(n18345), .ZN(
        n18337) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18346), .B1(
        n18624), .B2(n18678), .ZN(n18336) );
  OAI211_X1 U21371 ( .C1(n18681), .C2(n18350), .A(n18337), .B(n18336), .ZN(
        P3_U2880) );
  INV_X1 U21372 ( .A(n18338), .ZN(n18687) );
  AOI22_X1 U21373 ( .A1(n18645), .A2(n18683), .B1(n18682), .B2(n18345), .ZN(
        n18340) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18346), .B1(
        n18624), .B2(n18684), .ZN(n18339) );
  OAI211_X1 U21375 ( .C1(n18687), .C2(n18350), .A(n18340), .B(n18339), .ZN(
        P3_U2881) );
  INV_X1 U21376 ( .A(n18341), .ZN(n18693) );
  AOI22_X1 U21377 ( .A1(n18624), .A2(n18689), .B1(n18688), .B2(n18345), .ZN(
        n18343) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18346), .B1(
        n18645), .B2(n18690), .ZN(n18342) );
  OAI211_X1 U21379 ( .C1(n18693), .C2(n18350), .A(n18343), .B(n18342), .ZN(
        P3_U2882) );
  INV_X1 U21380 ( .A(n18344), .ZN(n18703) );
  AOI22_X1 U21381 ( .A1(n18624), .A2(n18699), .B1(n18695), .B2(n18345), .ZN(
        n18348) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18346), .B1(
        n18645), .B2(n18696), .ZN(n18347) );
  OAI211_X1 U21383 ( .C1(n18703), .C2(n18350), .A(n18348), .B(n18347), .ZN(
        P3_U2883) );
  NOR2_X1 U21384 ( .A1(n18750), .A2(n18349), .ZN(n18419) );
  NAND2_X1 U21385 ( .A1(n18419), .A2(n18748), .ZN(n18371) );
  INV_X1 U21386 ( .A(n18350), .ZN(n18413) );
  NOR2_X1 U21387 ( .A1(n18413), .A2(n18435), .ZN(n18396) );
  NOR2_X1 U21388 ( .A1(n18647), .A2(n18396), .ZN(n18367) );
  AOI22_X1 U21389 ( .A1(n18649), .A2(n18645), .B1(n18648), .B2(n18367), .ZN(
        n18354) );
  OAI21_X1 U21390 ( .B1(n18351), .B2(n18620), .A(n18396), .ZN(n18352) );
  OAI211_X1 U21391 ( .C1(n18435), .C2(n18872), .A(n18623), .B(n18352), .ZN(
        n18368) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18368), .B1(
        n18373), .B2(n18654), .ZN(n18353) );
  OAI211_X1 U21393 ( .C1(n18657), .C2(n18371), .A(n18354), .B(n18353), .ZN(
        P3_U2884) );
  AOI22_X1 U21394 ( .A1(n18645), .A2(n18659), .B1(n18658), .B2(n18367), .ZN(
        n18356) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18368), .B1(
        n18390), .B2(n18660), .ZN(n18355) );
  OAI211_X1 U21396 ( .C1(n18663), .C2(n18371), .A(n18356), .B(n18355), .ZN(
        P3_U2885) );
  AOI22_X1 U21397 ( .A1(n18390), .A2(n18665), .B1(n18664), .B2(n18367), .ZN(
        n18358) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18368), .B1(
        n18645), .B2(n18666), .ZN(n18357) );
  OAI211_X1 U21399 ( .C1(n18669), .C2(n18371), .A(n18358), .B(n18357), .ZN(
        P3_U2886) );
  AOI22_X1 U21400 ( .A1(n18390), .A2(n18672), .B1(n18670), .B2(n18367), .ZN(
        n18360) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18368), .B1(
        n18645), .B2(n18671), .ZN(n18359) );
  OAI211_X1 U21402 ( .C1(n18675), .C2(n18371), .A(n18360), .B(n18359), .ZN(
        P3_U2887) );
  AOI22_X1 U21403 ( .A1(n18645), .A2(n18678), .B1(n18676), .B2(n18367), .ZN(
        n18362) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18368), .B1(
        n18373), .B2(n18677), .ZN(n18361) );
  OAI211_X1 U21405 ( .C1(n18681), .C2(n18371), .A(n18362), .B(n18361), .ZN(
        P3_U2888) );
  AOI22_X1 U21406 ( .A1(n18390), .A2(n18683), .B1(n18682), .B2(n18367), .ZN(
        n18364) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18368), .B1(
        n18645), .B2(n18684), .ZN(n18363) );
  OAI211_X1 U21408 ( .C1(n18687), .C2(n18371), .A(n18364), .B(n18363), .ZN(
        P3_U2889) );
  AOI22_X1 U21409 ( .A1(n18645), .A2(n18689), .B1(n18688), .B2(n18367), .ZN(
        n18366) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18368), .B1(
        n18373), .B2(n18690), .ZN(n18365) );
  OAI211_X1 U21411 ( .C1(n18693), .C2(n18371), .A(n18366), .B(n18365), .ZN(
        P3_U2890) );
  AOI22_X1 U21412 ( .A1(n18390), .A2(n18696), .B1(n18695), .B2(n18367), .ZN(
        n18370) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18368), .B1(
        n18645), .B2(n18699), .ZN(n18369) );
  OAI211_X1 U21414 ( .C1(n18703), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2891) );
  NAND2_X1 U21415 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18419), .ZN(
        n18393) );
  AOI21_X1 U21416 ( .B1(n18750), .B2(n18620), .A(n18394), .ZN(n18464) );
  OAI211_X1 U21417 ( .C1(n18458), .C2(n18872), .A(n18372), .B(n18464), .ZN(
        n18389) );
  AND2_X1 U21418 ( .A1(n18776), .A2(n18419), .ZN(n18388) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18389), .B1(
        n18648), .B2(n18388), .ZN(n18375) );
  AOI22_X1 U21420 ( .A1(n18649), .A2(n18373), .B1(n18654), .B2(n18413), .ZN(
        n18374) );
  OAI211_X1 U21421 ( .C1(n18657), .C2(n18393), .A(n18375), .B(n18374), .ZN(
        P3_U2892) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18389), .B1(
        n18658), .B2(n18388), .ZN(n18377) );
  AOI22_X1 U21423 ( .A1(n18390), .A2(n18659), .B1(n18660), .B2(n18413), .ZN(
        n18376) );
  OAI211_X1 U21424 ( .C1(n18663), .C2(n18393), .A(n18377), .B(n18376), .ZN(
        P3_U2893) );
  AOI22_X1 U21425 ( .A1(n18665), .A2(n18413), .B1(n18664), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18389), .B1(
        n18390), .B2(n18666), .ZN(n18378) );
  OAI211_X1 U21427 ( .C1(n18669), .C2(n18393), .A(n18379), .B(n18378), .ZN(
        P3_U2894) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18389), .B1(
        n18670), .B2(n18388), .ZN(n18381) );
  AOI22_X1 U21429 ( .A1(n18390), .A2(n18671), .B1(n18672), .B2(n18413), .ZN(
        n18380) );
  OAI211_X1 U21430 ( .C1(n18675), .C2(n18393), .A(n18381), .B(n18380), .ZN(
        P3_U2895) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18389), .B1(
        n18676), .B2(n18388), .ZN(n18383) );
  AOI22_X1 U21432 ( .A1(n18390), .A2(n18678), .B1(n18677), .B2(n18413), .ZN(
        n18382) );
  OAI211_X1 U21433 ( .C1(n18681), .C2(n18393), .A(n18383), .B(n18382), .ZN(
        P3_U2896) );
  AOI22_X1 U21434 ( .A1(n18683), .A2(n18413), .B1(n18682), .B2(n18388), .ZN(
        n18385) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18389), .B1(
        n18390), .B2(n18684), .ZN(n18384) );
  OAI211_X1 U21436 ( .C1(n18687), .C2(n18393), .A(n18385), .B(n18384), .ZN(
        P3_U2897) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18389), .B1(
        n18688), .B2(n18388), .ZN(n18387) );
  AOI22_X1 U21438 ( .A1(n18390), .A2(n18689), .B1(n18690), .B2(n18413), .ZN(
        n18386) );
  OAI211_X1 U21439 ( .C1(n18693), .C2(n18393), .A(n18387), .B(n18386), .ZN(
        P3_U2898) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18389), .B1(
        n18695), .B2(n18388), .ZN(n18392) );
  AOI22_X1 U21441 ( .A1(n18390), .A2(n18699), .B1(n18696), .B2(n18413), .ZN(
        n18391) );
  OAI211_X1 U21442 ( .C1(n18703), .C2(n18393), .A(n18392), .B(n18391), .ZN(
        P3_U2899) );
  NOR2_X2 U21443 ( .A1(n18751), .A2(n18418), .ZN(n18480) );
  INV_X1 U21444 ( .A(n18480), .ZN(n18417) );
  NOR2_X1 U21445 ( .A1(n18458), .A2(n18480), .ZN(n18441) );
  NOR2_X1 U21446 ( .A1(n18647), .A2(n18441), .ZN(n18412) );
  AOI22_X1 U21447 ( .A1(n18649), .A2(n18413), .B1(n18648), .B2(n18412), .ZN(
        n18399) );
  OAI22_X1 U21448 ( .A1(n18396), .A2(n18395), .B1(n18441), .B2(n18394), .ZN(
        n18397) );
  OAI21_X1 U21449 ( .B1(n18480), .B2(n18872), .A(n18397), .ZN(n18414) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18414), .B1(
        n18654), .B2(n18435), .ZN(n18398) );
  OAI211_X1 U21451 ( .C1(n18657), .C2(n18417), .A(n18399), .B(n18398), .ZN(
        P3_U2900) );
  AOI22_X1 U21452 ( .A1(n18660), .A2(n18435), .B1(n18658), .B2(n18412), .ZN(
        n18401) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18414), .B1(
        n18659), .B2(n18413), .ZN(n18400) );
  OAI211_X1 U21454 ( .C1(n18663), .C2(n18417), .A(n18401), .B(n18400), .ZN(
        P3_U2901) );
  AOI22_X1 U21455 ( .A1(n18666), .A2(n18413), .B1(n18664), .B2(n18412), .ZN(
        n18403) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18414), .B1(
        n18665), .B2(n18435), .ZN(n18402) );
  OAI211_X1 U21457 ( .C1(n18669), .C2(n18417), .A(n18403), .B(n18402), .ZN(
        P3_U2902) );
  AOI22_X1 U21458 ( .A1(n18671), .A2(n18413), .B1(n18670), .B2(n18412), .ZN(
        n18405) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18414), .B1(
        n18672), .B2(n18435), .ZN(n18404) );
  OAI211_X1 U21460 ( .C1(n18675), .C2(n18417), .A(n18405), .B(n18404), .ZN(
        P3_U2903) );
  AOI22_X1 U21461 ( .A1(n18676), .A2(n18412), .B1(n18678), .B2(n18413), .ZN(
        n18407) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18414), .B1(
        n18677), .B2(n18435), .ZN(n18406) );
  OAI211_X1 U21463 ( .C1(n18681), .C2(n18417), .A(n18407), .B(n18406), .ZN(
        P3_U2904) );
  AOI22_X1 U21464 ( .A1(n18683), .A2(n18435), .B1(n18682), .B2(n18412), .ZN(
        n18409) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18414), .B1(
        n18684), .B2(n18413), .ZN(n18408) );
  OAI211_X1 U21466 ( .C1(n18687), .C2(n18417), .A(n18409), .B(n18408), .ZN(
        P3_U2905) );
  AOI22_X1 U21467 ( .A1(n18690), .A2(n18435), .B1(n18688), .B2(n18412), .ZN(
        n18411) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18414), .B1(
        n18689), .B2(n18413), .ZN(n18410) );
  OAI211_X1 U21469 ( .C1(n18693), .C2(n18417), .A(n18411), .B(n18410), .ZN(
        P3_U2906) );
  AOI22_X1 U21470 ( .A1(n18699), .A2(n18413), .B1(n18695), .B2(n18412), .ZN(
        n18416) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18414), .B1(
        n18696), .B2(n18435), .ZN(n18415) );
  OAI211_X1 U21472 ( .C1(n18703), .C2(n18417), .A(n18416), .B(n18415), .ZN(
        P3_U2907) );
  NAND2_X1 U21473 ( .A1(n18507), .A2(n18463), .ZN(n18440) );
  NOR2_X1 U21474 ( .A1(n18508), .A2(n18418), .ZN(n18434) );
  AOI22_X1 U21475 ( .A1(n18654), .A2(n18458), .B1(n18648), .B2(n18434), .ZN(
        n18421) );
  AOI22_X1 U21476 ( .A1(n18653), .A2(n18419), .B1(n18596), .B2(n18463), .ZN(
        n18436) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18436), .B1(
        n18649), .B2(n18435), .ZN(n18420) );
  OAI211_X1 U21478 ( .C1(n18657), .C2(n18440), .A(n18421), .B(n18420), .ZN(
        P3_U2908) );
  AOI22_X1 U21479 ( .A1(n18660), .A2(n18458), .B1(n18658), .B2(n18434), .ZN(
        n18423) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18436), .B1(
        n18659), .B2(n18435), .ZN(n18422) );
  OAI211_X1 U21481 ( .C1(n18663), .C2(n18440), .A(n18423), .B(n18422), .ZN(
        P3_U2909) );
  AOI22_X1 U21482 ( .A1(n18665), .A2(n18458), .B1(n18664), .B2(n18434), .ZN(
        n18425) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18436), .B1(
        n18666), .B2(n18435), .ZN(n18424) );
  OAI211_X1 U21484 ( .C1(n18669), .C2(n18440), .A(n18425), .B(n18424), .ZN(
        P3_U2910) );
  AOI22_X1 U21485 ( .A1(n18671), .A2(n18435), .B1(n18670), .B2(n18434), .ZN(
        n18427) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18436), .B1(
        n18672), .B2(n18458), .ZN(n18426) );
  OAI211_X1 U21487 ( .C1(n18675), .C2(n18440), .A(n18427), .B(n18426), .ZN(
        P3_U2911) );
  AOI22_X1 U21488 ( .A1(n18676), .A2(n18434), .B1(n18678), .B2(n18435), .ZN(
        n18429) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18436), .B1(
        n18677), .B2(n18458), .ZN(n18428) );
  OAI211_X1 U21490 ( .C1(n18681), .C2(n18440), .A(n18429), .B(n18428), .ZN(
        P3_U2912) );
  AOI22_X1 U21491 ( .A1(n18682), .A2(n18434), .B1(n18684), .B2(n18435), .ZN(
        n18431) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18436), .B1(
        n18683), .B2(n18458), .ZN(n18430) );
  OAI211_X1 U21493 ( .C1(n18687), .C2(n18440), .A(n18431), .B(n18430), .ZN(
        P3_U2913) );
  AOI22_X1 U21494 ( .A1(n18690), .A2(n18458), .B1(n18688), .B2(n18434), .ZN(
        n18433) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18436), .B1(
        n18689), .B2(n18435), .ZN(n18432) );
  OAI211_X1 U21496 ( .C1(n18693), .C2(n18440), .A(n18433), .B(n18432), .ZN(
        P3_U2914) );
  AOI22_X1 U21497 ( .A1(n18699), .A2(n18435), .B1(n18695), .B2(n18434), .ZN(
        n18438) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18436), .B1(
        n18696), .B2(n18458), .ZN(n18437) );
  OAI211_X1 U21499 ( .C1(n18703), .C2(n18440), .A(n18438), .B(n18437), .ZN(
        P3_U2915) );
  NOR2_X1 U21500 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18439), .ZN(
        n18509) );
  NAND2_X1 U21501 ( .A1(n18509), .A2(n18748), .ZN(n18462) );
  INV_X1 U21502 ( .A(n18440), .ZN(n18502) );
  INV_X1 U21503 ( .A(n18462), .ZN(n18525) );
  NOR2_X1 U21504 ( .A1(n18502), .A2(n18525), .ZN(n18485) );
  NOR2_X1 U21505 ( .A1(n18647), .A2(n18485), .ZN(n18457) );
  AOI22_X1 U21506 ( .A1(n18654), .A2(n18480), .B1(n18648), .B2(n18457), .ZN(
        n18444) );
  OAI21_X1 U21507 ( .B1(n18441), .B2(n18620), .A(n18485), .ZN(n18442) );
  OAI211_X1 U21508 ( .C1(n18525), .C2(n18872), .A(n18623), .B(n18442), .ZN(
        n18459) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18459), .B1(
        n18649), .B2(n18458), .ZN(n18443) );
  OAI211_X1 U21510 ( .C1(n18657), .C2(n18462), .A(n18444), .B(n18443), .ZN(
        P3_U2916) );
  AOI22_X1 U21511 ( .A1(n18660), .A2(n18480), .B1(n18658), .B2(n18457), .ZN(
        n18446) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18459), .B1(
        n18659), .B2(n18458), .ZN(n18445) );
  OAI211_X1 U21513 ( .C1(n18663), .C2(n18462), .A(n18446), .B(n18445), .ZN(
        P3_U2917) );
  AOI22_X1 U21514 ( .A1(n18665), .A2(n18480), .B1(n18664), .B2(n18457), .ZN(
        n18448) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18459), .B1(
        n18666), .B2(n18458), .ZN(n18447) );
  OAI211_X1 U21516 ( .C1(n18669), .C2(n18462), .A(n18448), .B(n18447), .ZN(
        P3_U2918) );
  AOI22_X1 U21517 ( .A1(n18671), .A2(n18458), .B1(n18670), .B2(n18457), .ZN(
        n18450) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18459), .B1(
        n18672), .B2(n18480), .ZN(n18449) );
  OAI211_X1 U21519 ( .C1(n18675), .C2(n18462), .A(n18450), .B(n18449), .ZN(
        P3_U2919) );
  AOI22_X1 U21520 ( .A1(n18676), .A2(n18457), .B1(n18678), .B2(n18458), .ZN(
        n18452) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18459), .B1(
        n18677), .B2(n18480), .ZN(n18451) );
  OAI211_X1 U21522 ( .C1(n18681), .C2(n18462), .A(n18452), .B(n18451), .ZN(
        P3_U2920) );
  AOI22_X1 U21523 ( .A1(n18682), .A2(n18457), .B1(n18684), .B2(n18458), .ZN(
        n18454) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18459), .B1(
        n18683), .B2(n18480), .ZN(n18453) );
  OAI211_X1 U21525 ( .C1(n18687), .C2(n18462), .A(n18454), .B(n18453), .ZN(
        P3_U2921) );
  AOI22_X1 U21526 ( .A1(n18690), .A2(n18480), .B1(n18688), .B2(n18457), .ZN(
        n18456) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18459), .B1(
        n18689), .B2(n18458), .ZN(n18455) );
  OAI211_X1 U21528 ( .C1(n18693), .C2(n18462), .A(n18456), .B(n18455), .ZN(
        P3_U2922) );
  AOI22_X1 U21529 ( .A1(n18699), .A2(n18458), .B1(n18695), .B2(n18457), .ZN(
        n18461) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18459), .B1(
        n18696), .B2(n18480), .ZN(n18460) );
  OAI211_X1 U21531 ( .C1(n18703), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        P3_U2923) );
  NAND2_X1 U21532 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18509), .ZN(
        n18484) );
  AND2_X1 U21533 ( .A1(n18776), .A2(n18509), .ZN(n18479) );
  AOI22_X1 U21534 ( .A1(n18654), .A2(n18502), .B1(n18648), .B2(n18479), .ZN(
        n18466) );
  INV_X1 U21535 ( .A(n18484), .ZN(n18548) );
  OAI211_X1 U21536 ( .C1(n18548), .C2(n18872), .A(n18464), .B(n18463), .ZN(
        n18481) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18481), .B1(
        n18649), .B2(n18480), .ZN(n18465) );
  OAI211_X1 U21538 ( .C1(n18657), .C2(n18484), .A(n18466), .B(n18465), .ZN(
        P3_U2924) );
  AOI22_X1 U21539 ( .A1(n18660), .A2(n18502), .B1(n18658), .B2(n18479), .ZN(
        n18468) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18481), .B1(
        n18659), .B2(n18480), .ZN(n18467) );
  OAI211_X1 U21541 ( .C1(n18663), .C2(n18484), .A(n18468), .B(n18467), .ZN(
        P3_U2925) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18481), .B1(
        n18664), .B2(n18479), .ZN(n18470) );
  AOI22_X1 U21543 ( .A1(n18666), .A2(n18480), .B1(n18665), .B2(n18502), .ZN(
        n18469) );
  OAI211_X1 U21544 ( .C1(n18669), .C2(n18484), .A(n18470), .B(n18469), .ZN(
        P3_U2926) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18481), .B1(
        n18670), .B2(n18479), .ZN(n18472) );
  AOI22_X1 U21546 ( .A1(n18672), .A2(n18502), .B1(n18671), .B2(n18480), .ZN(
        n18471) );
  OAI211_X1 U21547 ( .C1(n18675), .C2(n18484), .A(n18472), .B(n18471), .ZN(
        P3_U2927) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18481), .B1(
        n18676), .B2(n18479), .ZN(n18474) );
  AOI22_X1 U21549 ( .A1(n18677), .A2(n18502), .B1(n18678), .B2(n18480), .ZN(
        n18473) );
  OAI211_X1 U21550 ( .C1(n18681), .C2(n18484), .A(n18474), .B(n18473), .ZN(
        P3_U2928) );
  AOI22_X1 U21551 ( .A1(n18683), .A2(n18502), .B1(n18682), .B2(n18479), .ZN(
        n18476) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18481), .B1(
        n18684), .B2(n18480), .ZN(n18475) );
  OAI211_X1 U21553 ( .C1(n18687), .C2(n18484), .A(n18476), .B(n18475), .ZN(
        P3_U2929) );
  AOI22_X1 U21554 ( .A1(n18690), .A2(n18502), .B1(n18688), .B2(n18479), .ZN(
        n18478) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18481), .B1(
        n18689), .B2(n18480), .ZN(n18477) );
  OAI211_X1 U21556 ( .C1(n18693), .C2(n18484), .A(n18478), .B(n18477), .ZN(
        P3_U2930) );
  AOI22_X1 U21557 ( .A1(n18696), .A2(n18502), .B1(n18695), .B2(n18479), .ZN(
        n18483) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18481), .B1(
        n18699), .B2(n18480), .ZN(n18482) );
  OAI211_X1 U21559 ( .C1(n18703), .C2(n18484), .A(n18483), .B(n18482), .ZN(
        P3_U2931) );
  NOR2_X2 U21560 ( .A1(n18751), .A2(n18529), .ZN(n18569) );
  INV_X1 U21561 ( .A(n18569), .ZN(n18506) );
  NOR2_X1 U21562 ( .A1(n18548), .A2(n18569), .ZN(n18531) );
  NOR2_X1 U21563 ( .A1(n18647), .A2(n18531), .ZN(n18501) );
  AOI22_X1 U21564 ( .A1(n18654), .A2(n18525), .B1(n18648), .B2(n18501), .ZN(
        n18488) );
  OAI21_X1 U21565 ( .B1(n18485), .B2(n18620), .A(n18531), .ZN(n18486) );
  OAI211_X1 U21566 ( .C1(n18569), .C2(n18872), .A(n18623), .B(n18486), .ZN(
        n18503) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18503), .B1(
        n18649), .B2(n18502), .ZN(n18487) );
  OAI211_X1 U21568 ( .C1(n18657), .C2(n18506), .A(n18488), .B(n18487), .ZN(
        P3_U2932) );
  AOI22_X1 U21569 ( .A1(n18660), .A2(n18525), .B1(n18658), .B2(n18501), .ZN(
        n18490) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18503), .B1(
        n18659), .B2(n18502), .ZN(n18489) );
  OAI211_X1 U21571 ( .C1(n18663), .C2(n18506), .A(n18490), .B(n18489), .ZN(
        P3_U2933) );
  AOI22_X1 U21572 ( .A1(n18665), .A2(n18525), .B1(n18664), .B2(n18501), .ZN(
        n18492) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18503), .B1(
        n18666), .B2(n18502), .ZN(n18491) );
  OAI211_X1 U21574 ( .C1(n18669), .C2(n18506), .A(n18492), .B(n18491), .ZN(
        P3_U2934) );
  AOI22_X1 U21575 ( .A1(n18671), .A2(n18502), .B1(n18670), .B2(n18501), .ZN(
        n18494) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18503), .B1(
        n18672), .B2(n18525), .ZN(n18493) );
  OAI211_X1 U21577 ( .C1(n18675), .C2(n18506), .A(n18494), .B(n18493), .ZN(
        P3_U2935) );
  AOI22_X1 U21578 ( .A1(n18676), .A2(n18501), .B1(n18678), .B2(n18502), .ZN(
        n18496) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18503), .B1(
        n18677), .B2(n18525), .ZN(n18495) );
  OAI211_X1 U21580 ( .C1(n18681), .C2(n18506), .A(n18496), .B(n18495), .ZN(
        P3_U2936) );
  AOI22_X1 U21581 ( .A1(n18682), .A2(n18501), .B1(n18684), .B2(n18502), .ZN(
        n18498) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18503), .B1(
        n18683), .B2(n18525), .ZN(n18497) );
  OAI211_X1 U21583 ( .C1(n18687), .C2(n18506), .A(n18498), .B(n18497), .ZN(
        P3_U2937) );
  AOI22_X1 U21584 ( .A1(n18690), .A2(n18525), .B1(n18688), .B2(n18501), .ZN(
        n18500) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18503), .B1(
        n18689), .B2(n18502), .ZN(n18499) );
  OAI211_X1 U21586 ( .C1(n18693), .C2(n18506), .A(n18500), .B(n18499), .ZN(
        P3_U2938) );
  AOI22_X1 U21587 ( .A1(n18699), .A2(n18502), .B1(n18695), .B2(n18501), .ZN(
        n18505) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18503), .B1(
        n18696), .B2(n18525), .ZN(n18504) );
  OAI211_X1 U21589 ( .C1(n18703), .C2(n18506), .A(n18505), .B(n18504), .ZN(
        P3_U2939) );
  NAND2_X1 U21590 ( .A1(n18507), .A2(n18553), .ZN(n18530) );
  NOR2_X1 U21591 ( .A1(n18508), .A2(n18529), .ZN(n18524) );
  AOI22_X1 U21592 ( .A1(n18654), .A2(n18548), .B1(n18648), .B2(n18524), .ZN(
        n18511) );
  AOI22_X1 U21593 ( .A1(n18653), .A2(n18509), .B1(n18596), .B2(n18553), .ZN(
        n18526) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18526), .B1(
        n18649), .B2(n18525), .ZN(n18510) );
  OAI211_X1 U21595 ( .C1(n18657), .C2(n18530), .A(n18511), .B(n18510), .ZN(
        P3_U2940) );
  AOI22_X1 U21596 ( .A1(n18660), .A2(n18548), .B1(n18658), .B2(n18524), .ZN(
        n18513) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18526), .B1(
        n18659), .B2(n18525), .ZN(n18512) );
  OAI211_X1 U21598 ( .C1(n18663), .C2(n18530), .A(n18513), .B(n18512), .ZN(
        P3_U2941) );
  AOI22_X1 U21599 ( .A1(n18666), .A2(n18525), .B1(n18664), .B2(n18524), .ZN(
        n18515) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18526), .B1(
        n18665), .B2(n18548), .ZN(n18514) );
  OAI211_X1 U21601 ( .C1(n18669), .C2(n18530), .A(n18515), .B(n18514), .ZN(
        P3_U2942) );
  AOI22_X1 U21602 ( .A1(n18671), .A2(n18525), .B1(n18670), .B2(n18524), .ZN(
        n18517) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18526), .B1(
        n18672), .B2(n18548), .ZN(n18516) );
  OAI211_X1 U21604 ( .C1(n18675), .C2(n18530), .A(n18517), .B(n18516), .ZN(
        P3_U2943) );
  AOI22_X1 U21605 ( .A1(n18676), .A2(n18524), .B1(n18678), .B2(n18525), .ZN(
        n18519) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18526), .B1(
        n18677), .B2(n18548), .ZN(n18518) );
  OAI211_X1 U21607 ( .C1(n18681), .C2(n18530), .A(n18519), .B(n18518), .ZN(
        P3_U2944) );
  AOI22_X1 U21608 ( .A1(n18683), .A2(n18548), .B1(n18682), .B2(n18524), .ZN(
        n18521) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18526), .B1(
        n18684), .B2(n18525), .ZN(n18520) );
  OAI211_X1 U21610 ( .C1(n18687), .C2(n18530), .A(n18521), .B(n18520), .ZN(
        P3_U2945) );
  AOI22_X1 U21611 ( .A1(n18690), .A2(n18548), .B1(n18688), .B2(n18524), .ZN(
        n18523) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18526), .B1(
        n18689), .B2(n18525), .ZN(n18522) );
  OAI211_X1 U21613 ( .C1(n18693), .C2(n18530), .A(n18523), .B(n18522), .ZN(
        P3_U2946) );
  AOI22_X1 U21614 ( .A1(n18699), .A2(n18525), .B1(n18695), .B2(n18524), .ZN(
        n18528) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18526), .B1(
        n18696), .B2(n18548), .ZN(n18527) );
  OAI211_X1 U21616 ( .C1(n18703), .C2(n18530), .A(n18528), .B(n18527), .ZN(
        P3_U2947) );
  NOR2_X1 U21617 ( .A1(n18750), .A2(n18529), .ZN(n18598) );
  NAND2_X1 U21618 ( .A1(n18598), .A2(n18748), .ZN(n18552) );
  INV_X1 U21619 ( .A(n18530), .ZN(n18591) );
  NOR2_X1 U21620 ( .A1(n18591), .A2(n18614), .ZN(n18574) );
  NOR2_X1 U21621 ( .A1(n18647), .A2(n18574), .ZN(n18547) );
  AOI22_X1 U21622 ( .A1(n18654), .A2(n18569), .B1(n18648), .B2(n18547), .ZN(
        n18534) );
  OAI21_X1 U21623 ( .B1(n18531), .B2(n18620), .A(n18574), .ZN(n18532) );
  OAI211_X1 U21624 ( .C1(n18614), .C2(n18872), .A(n18623), .B(n18532), .ZN(
        n18549) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18549), .B1(
        n18649), .B2(n18548), .ZN(n18533) );
  OAI211_X1 U21626 ( .C1(n18657), .C2(n18552), .A(n18534), .B(n18533), .ZN(
        P3_U2948) );
  AOI22_X1 U21627 ( .A1(n18660), .A2(n18569), .B1(n18658), .B2(n18547), .ZN(
        n18536) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18549), .B1(
        n18659), .B2(n18548), .ZN(n18535) );
  OAI211_X1 U21629 ( .C1(n18663), .C2(n18552), .A(n18536), .B(n18535), .ZN(
        P3_U2949) );
  AOI22_X1 U21630 ( .A1(n18666), .A2(n18548), .B1(n18664), .B2(n18547), .ZN(
        n18538) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18549), .B1(
        n18665), .B2(n18569), .ZN(n18537) );
  OAI211_X1 U21632 ( .C1(n18669), .C2(n18552), .A(n18538), .B(n18537), .ZN(
        P3_U2950) );
  AOI22_X1 U21633 ( .A1(n18672), .A2(n18569), .B1(n18670), .B2(n18547), .ZN(
        n18540) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18549), .B1(
        n18671), .B2(n18548), .ZN(n18539) );
  OAI211_X1 U21635 ( .C1(n18675), .C2(n18552), .A(n18540), .B(n18539), .ZN(
        P3_U2951) );
  AOI22_X1 U21636 ( .A1(n18676), .A2(n18547), .B1(n18678), .B2(n18548), .ZN(
        n18542) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18549), .B1(
        n18677), .B2(n18569), .ZN(n18541) );
  OAI211_X1 U21638 ( .C1(n18681), .C2(n18552), .A(n18542), .B(n18541), .ZN(
        P3_U2952) );
  AOI22_X1 U21639 ( .A1(n18683), .A2(n18569), .B1(n18682), .B2(n18547), .ZN(
        n18544) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18549), .B1(
        n18684), .B2(n18548), .ZN(n18543) );
  OAI211_X1 U21641 ( .C1(n18687), .C2(n18552), .A(n18544), .B(n18543), .ZN(
        P3_U2953) );
  AOI22_X1 U21642 ( .A1(n18689), .A2(n18548), .B1(n18688), .B2(n18547), .ZN(
        n18546) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18549), .B1(
        n18690), .B2(n18569), .ZN(n18545) );
  OAI211_X1 U21644 ( .C1(n18693), .C2(n18552), .A(n18546), .B(n18545), .ZN(
        P3_U2954) );
  AOI22_X1 U21645 ( .A1(n18699), .A2(n18548), .B1(n18695), .B2(n18547), .ZN(
        n18551) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18549), .B1(
        n18696), .B2(n18569), .ZN(n18550) );
  OAI211_X1 U21647 ( .C1(n18703), .C2(n18552), .A(n18551), .B(n18550), .ZN(
        P3_U2955) );
  NAND2_X1 U21648 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18598), .ZN(
        n18573) );
  AND2_X1 U21649 ( .A1(n18776), .A2(n18598), .ZN(n18568) );
  AOI22_X1 U21650 ( .A1(n18649), .A2(n18569), .B1(n18648), .B2(n18568), .ZN(
        n18555) );
  AOI22_X1 U21651 ( .A1(n18653), .A2(n18553), .B1(n18650), .B2(n18598), .ZN(
        n18570) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18570), .B1(
        n18654), .B2(n18591), .ZN(n18554) );
  OAI211_X1 U21653 ( .C1(n18657), .C2(n18573), .A(n18555), .B(n18554), .ZN(
        P3_U2956) );
  AOI22_X1 U21654 ( .A1(n18660), .A2(n18591), .B1(n18658), .B2(n18568), .ZN(
        n18557) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18570), .B1(
        n18659), .B2(n18569), .ZN(n18556) );
  OAI211_X1 U21656 ( .C1(n18663), .C2(n18573), .A(n18557), .B(n18556), .ZN(
        P3_U2957) );
  AOI22_X1 U21657 ( .A1(n18665), .A2(n18591), .B1(n18664), .B2(n18568), .ZN(
        n18559) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18570), .B1(
        n18666), .B2(n18569), .ZN(n18558) );
  OAI211_X1 U21659 ( .C1(n18669), .C2(n18573), .A(n18559), .B(n18558), .ZN(
        P3_U2958) );
  AOI22_X1 U21660 ( .A1(n18672), .A2(n18591), .B1(n18670), .B2(n18568), .ZN(
        n18561) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18570), .B1(
        n18671), .B2(n18569), .ZN(n18560) );
  OAI211_X1 U21662 ( .C1(n18675), .C2(n18573), .A(n18561), .B(n18560), .ZN(
        P3_U2959) );
  AOI22_X1 U21663 ( .A1(n18676), .A2(n18568), .B1(n18678), .B2(n18569), .ZN(
        n18563) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18570), .B1(
        n18677), .B2(n18591), .ZN(n18562) );
  OAI211_X1 U21665 ( .C1(n18681), .C2(n18573), .A(n18563), .B(n18562), .ZN(
        P3_U2960) );
  AOI22_X1 U21666 ( .A1(n18682), .A2(n18568), .B1(n18684), .B2(n18569), .ZN(
        n18565) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18570), .B1(
        n18683), .B2(n18591), .ZN(n18564) );
  OAI211_X1 U21668 ( .C1(n18687), .C2(n18573), .A(n18565), .B(n18564), .ZN(
        P3_U2961) );
  AOI22_X1 U21669 ( .A1(n18690), .A2(n18591), .B1(n18688), .B2(n18568), .ZN(
        n18567) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18570), .B1(
        n18689), .B2(n18569), .ZN(n18566) );
  OAI211_X1 U21671 ( .C1(n18693), .C2(n18573), .A(n18567), .B(n18566), .ZN(
        P3_U2962) );
  AOI22_X1 U21672 ( .A1(n18699), .A2(n18569), .B1(n18695), .B2(n18568), .ZN(
        n18572) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18570), .B1(
        n18696), .B2(n18591), .ZN(n18571) );
  OAI211_X1 U21674 ( .C1(n18703), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2963) );
  NAND2_X1 U21675 ( .A1(n18652), .A2(n18748), .ZN(n18595) );
  INV_X1 U21676 ( .A(n18573), .ZN(n18640) );
  INV_X1 U21677 ( .A(n18595), .ZN(n18698) );
  NOR2_X1 U21678 ( .A1(n18640), .A2(n18698), .ZN(n18621) );
  NOR2_X1 U21679 ( .A1(n18647), .A2(n18621), .ZN(n18590) );
  AOI22_X1 U21680 ( .A1(n18654), .A2(n18614), .B1(n18648), .B2(n18590), .ZN(
        n18577) );
  OAI21_X1 U21681 ( .B1(n18574), .B2(n18620), .A(n18621), .ZN(n18575) );
  OAI211_X1 U21682 ( .C1(n18698), .C2(n18872), .A(n18623), .B(n18575), .ZN(
        n18592) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18592), .B1(
        n18649), .B2(n18591), .ZN(n18576) );
  OAI211_X1 U21684 ( .C1(n18657), .C2(n18595), .A(n18577), .B(n18576), .ZN(
        P3_U2964) );
  AOI22_X1 U21685 ( .A1(n18659), .A2(n18591), .B1(n18658), .B2(n18590), .ZN(
        n18579) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18592), .B1(
        n18660), .B2(n18614), .ZN(n18578) );
  OAI211_X1 U21687 ( .C1(n18663), .C2(n18595), .A(n18579), .B(n18578), .ZN(
        P3_U2965) );
  AOI22_X1 U21688 ( .A1(n18666), .A2(n18591), .B1(n18664), .B2(n18590), .ZN(
        n18581) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18592), .B1(
        n18665), .B2(n18614), .ZN(n18580) );
  OAI211_X1 U21690 ( .C1(n18669), .C2(n18595), .A(n18581), .B(n18580), .ZN(
        P3_U2966) );
  AOI22_X1 U21691 ( .A1(n18671), .A2(n18591), .B1(n18670), .B2(n18590), .ZN(
        n18583) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18592), .B1(
        n18672), .B2(n18614), .ZN(n18582) );
  OAI211_X1 U21693 ( .C1(n18675), .C2(n18595), .A(n18583), .B(n18582), .ZN(
        P3_U2967) );
  AOI22_X1 U21694 ( .A1(n18677), .A2(n18614), .B1(n18676), .B2(n18590), .ZN(
        n18585) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18592), .B1(
        n18678), .B2(n18591), .ZN(n18584) );
  OAI211_X1 U21696 ( .C1(n18681), .C2(n18595), .A(n18585), .B(n18584), .ZN(
        P3_U2968) );
  AOI22_X1 U21697 ( .A1(n18682), .A2(n18590), .B1(n18684), .B2(n18591), .ZN(
        n18587) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18592), .B1(
        n18683), .B2(n18614), .ZN(n18586) );
  OAI211_X1 U21699 ( .C1(n18687), .C2(n18595), .A(n18587), .B(n18586), .ZN(
        P3_U2969) );
  AOI22_X1 U21700 ( .A1(n18689), .A2(n18591), .B1(n18688), .B2(n18590), .ZN(
        n18589) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18592), .B1(
        n18690), .B2(n18614), .ZN(n18588) );
  OAI211_X1 U21702 ( .C1(n18693), .C2(n18595), .A(n18589), .B(n18588), .ZN(
        P3_U2970) );
  AOI22_X1 U21703 ( .A1(n18696), .A2(n18614), .B1(n18695), .B2(n18590), .ZN(
        n18594) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18592), .B1(
        n18699), .B2(n18591), .ZN(n18593) );
  OAI211_X1 U21705 ( .C1(n18703), .C2(n18595), .A(n18594), .B(n18593), .ZN(
        P3_U2971) );
  AND2_X1 U21706 ( .A1(n18776), .A2(n18652), .ZN(n18613) );
  AOI22_X1 U21707 ( .A1(n18654), .A2(n18640), .B1(n18648), .B2(n18613), .ZN(
        n18600) );
  NOR2_X1 U21708 ( .A1(n18755), .A2(n18758), .ZN(n18597) );
  AOI22_X1 U21709 ( .A1(n18653), .A2(n18598), .B1(n18597), .B2(n18596), .ZN(
        n18615) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18615), .B1(
        n18649), .B2(n18614), .ZN(n18599) );
  OAI211_X1 U21711 ( .C1(n18618), .C2(n18657), .A(n18600), .B(n18599), .ZN(
        P3_U2972) );
  AOI22_X1 U21712 ( .A1(n18659), .A2(n18614), .B1(n18658), .B2(n18613), .ZN(
        n18602) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18615), .B1(
        n18660), .B2(n18640), .ZN(n18601) );
  OAI211_X1 U21714 ( .C1(n18618), .C2(n18663), .A(n18602), .B(n18601), .ZN(
        P3_U2973) );
  AOI22_X1 U21715 ( .A1(n18665), .A2(n18640), .B1(n18664), .B2(n18613), .ZN(
        n18604) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18615), .B1(
        n18666), .B2(n18614), .ZN(n18603) );
  OAI211_X1 U21717 ( .C1(n18618), .C2(n18669), .A(n18604), .B(n18603), .ZN(
        P3_U2974) );
  AOI22_X1 U21718 ( .A1(n18672), .A2(n18640), .B1(n18670), .B2(n18613), .ZN(
        n18606) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18615), .B1(
        n18671), .B2(n18614), .ZN(n18605) );
  OAI211_X1 U21720 ( .C1(n18618), .C2(n18675), .A(n18606), .B(n18605), .ZN(
        P3_U2975) );
  AOI22_X1 U21721 ( .A1(n18677), .A2(n18640), .B1(n18676), .B2(n18613), .ZN(
        n18608) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18615), .B1(
        n18678), .B2(n18614), .ZN(n18607) );
  OAI211_X1 U21723 ( .C1(n18618), .C2(n18681), .A(n18608), .B(n18607), .ZN(
        P3_U2976) );
  AOI22_X1 U21724 ( .A1(n18683), .A2(n18640), .B1(n18682), .B2(n18613), .ZN(
        n18610) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18615), .B1(
        n18684), .B2(n18614), .ZN(n18609) );
  OAI211_X1 U21726 ( .C1(n18618), .C2(n18687), .A(n18610), .B(n18609), .ZN(
        P3_U2977) );
  AOI22_X1 U21727 ( .A1(n18690), .A2(n18640), .B1(n18688), .B2(n18613), .ZN(
        n18612) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18615), .B1(
        n18689), .B2(n18614), .ZN(n18611) );
  OAI211_X1 U21729 ( .C1(n18618), .C2(n18693), .A(n18612), .B(n18611), .ZN(
        P3_U2978) );
  AOI22_X1 U21730 ( .A1(n18699), .A2(n18614), .B1(n18695), .B2(n18613), .ZN(
        n18617) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18615), .B1(
        n18696), .B2(n18640), .ZN(n18616) );
  OAI211_X1 U21732 ( .C1(n18618), .C2(n18703), .A(n18617), .B(n18616), .ZN(
        P3_U2979) );
  INV_X1 U21733 ( .A(n18624), .ZN(n18644) );
  NOR2_X1 U21734 ( .A1(n18647), .A2(n18619), .ZN(n18639) );
  AOI22_X1 U21735 ( .A1(n18649), .A2(n18640), .B1(n18648), .B2(n18639), .ZN(
        n18626) );
  OAI21_X1 U21736 ( .B1(n18621), .B2(n18620), .A(n18619), .ZN(n18622) );
  OAI211_X1 U21737 ( .C1(n18624), .C2(n18872), .A(n18623), .B(n18622), .ZN(
        n18641) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18641), .B1(
        n18654), .B2(n18698), .ZN(n18625) );
  OAI211_X1 U21739 ( .C1(n18644), .C2(n18657), .A(n18626), .B(n18625), .ZN(
        P3_U2980) );
  AOI22_X1 U21740 ( .A1(n18660), .A2(n18698), .B1(n18658), .B2(n18639), .ZN(
        n18628) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18641), .B1(
        n18659), .B2(n18640), .ZN(n18627) );
  OAI211_X1 U21742 ( .C1(n18644), .C2(n18663), .A(n18628), .B(n18627), .ZN(
        P3_U2981) );
  AOI22_X1 U21743 ( .A1(n18665), .A2(n18698), .B1(n18664), .B2(n18639), .ZN(
        n18630) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18641), .B1(
        n18666), .B2(n18640), .ZN(n18629) );
  OAI211_X1 U21745 ( .C1(n18644), .C2(n18669), .A(n18630), .B(n18629), .ZN(
        P3_U2982) );
  AOI22_X1 U21746 ( .A1(n18671), .A2(n18640), .B1(n18670), .B2(n18639), .ZN(
        n18632) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18641), .B1(
        n18672), .B2(n18698), .ZN(n18631) );
  OAI211_X1 U21748 ( .C1(n18644), .C2(n18675), .A(n18632), .B(n18631), .ZN(
        P3_U2983) );
  AOI22_X1 U21749 ( .A1(n18677), .A2(n18698), .B1(n18676), .B2(n18639), .ZN(
        n18634) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18641), .B1(
        n18678), .B2(n18640), .ZN(n18633) );
  OAI211_X1 U21751 ( .C1(n18644), .C2(n18681), .A(n18634), .B(n18633), .ZN(
        P3_U2984) );
  AOI22_X1 U21752 ( .A1(n18683), .A2(n18698), .B1(n18682), .B2(n18639), .ZN(
        n18636) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18641), .B1(
        n18684), .B2(n18640), .ZN(n18635) );
  OAI211_X1 U21754 ( .C1(n18644), .C2(n18687), .A(n18636), .B(n18635), .ZN(
        P3_U2985) );
  AOI22_X1 U21755 ( .A1(n18690), .A2(n18698), .B1(n18688), .B2(n18639), .ZN(
        n18638) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18641), .B1(
        n18689), .B2(n18640), .ZN(n18637) );
  OAI211_X1 U21757 ( .C1(n18644), .C2(n18693), .A(n18638), .B(n18637), .ZN(
        P3_U2986) );
  AOI22_X1 U21758 ( .A1(n18696), .A2(n18698), .B1(n18695), .B2(n18639), .ZN(
        n18643) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18641), .B1(
        n18699), .B2(n18640), .ZN(n18642) );
  OAI211_X1 U21760 ( .C1(n18644), .C2(n18703), .A(n18643), .B(n18642), .ZN(
        P3_U2987) );
  INV_X1 U21761 ( .A(n18645), .ZN(n18704) );
  NOR2_X1 U21762 ( .A1(n18647), .A2(n18646), .ZN(n18694) );
  AOI22_X1 U21763 ( .A1(n18649), .A2(n18698), .B1(n18648), .B2(n18694), .ZN(
        n18656) );
  AOI22_X1 U21764 ( .A1(n18653), .A2(n18652), .B1(n18651), .B2(n18650), .ZN(
        n18700) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18700), .B1(
        n18697), .B2(n18654), .ZN(n18655) );
  OAI211_X1 U21766 ( .C1(n18704), .C2(n18657), .A(n18656), .B(n18655), .ZN(
        P3_U2988) );
  AOI22_X1 U21767 ( .A1(n18659), .A2(n18698), .B1(n18658), .B2(n18694), .ZN(
        n18662) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18700), .B1(
        n18697), .B2(n18660), .ZN(n18661) );
  OAI211_X1 U21769 ( .C1(n18704), .C2(n18663), .A(n18662), .B(n18661), .ZN(
        P3_U2989) );
  AOI22_X1 U21770 ( .A1(n18697), .A2(n18665), .B1(n18664), .B2(n18694), .ZN(
        n18668) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18700), .B1(
        n18666), .B2(n18698), .ZN(n18667) );
  OAI211_X1 U21772 ( .C1(n18704), .C2(n18669), .A(n18668), .B(n18667), .ZN(
        P3_U2990) );
  AOI22_X1 U21773 ( .A1(n18671), .A2(n18698), .B1(n18670), .B2(n18694), .ZN(
        n18674) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18700), .B1(
        n18697), .B2(n18672), .ZN(n18673) );
  OAI211_X1 U21775 ( .C1(n18704), .C2(n18675), .A(n18674), .B(n18673), .ZN(
        P3_U2991) );
  AOI22_X1 U21776 ( .A1(n18697), .A2(n18677), .B1(n18676), .B2(n18694), .ZN(
        n18680) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18700), .B1(
        n18678), .B2(n18698), .ZN(n18679) );
  OAI211_X1 U21778 ( .C1(n18704), .C2(n18681), .A(n18680), .B(n18679), .ZN(
        P3_U2992) );
  AOI22_X1 U21779 ( .A1(n18697), .A2(n18683), .B1(n18682), .B2(n18694), .ZN(
        n18686) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18700), .B1(
        n18684), .B2(n18698), .ZN(n18685) );
  OAI211_X1 U21781 ( .C1(n18704), .C2(n18687), .A(n18686), .B(n18685), .ZN(
        P3_U2993) );
  AOI22_X1 U21782 ( .A1(n18689), .A2(n18698), .B1(n18688), .B2(n18694), .ZN(
        n18692) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18700), .B1(
        n18697), .B2(n18690), .ZN(n18691) );
  OAI211_X1 U21784 ( .C1(n18704), .C2(n18693), .A(n18692), .B(n18691), .ZN(
        P3_U2994) );
  AOI22_X1 U21785 ( .A1(n18697), .A2(n18696), .B1(n18695), .B2(n18694), .ZN(
        n18702) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18700), .B1(
        n18699), .B2(n18698), .ZN(n18701) );
  OAI211_X1 U21787 ( .C1(n18704), .C2(n18703), .A(n18702), .B(n18701), .ZN(
        P3_U2995) );
  INV_X1 U21788 ( .A(n18705), .ZN(n18711) );
  NOR2_X1 U21789 ( .A1(n18717), .A2(n18706), .ZN(n18708) );
  OAI222_X1 U21790 ( .A1(n18712), .A2(n18711), .B1(n18710), .B2(n18709), .C1(
        n18708), .C2(n18707), .ZN(n18918) );
  OAI21_X1 U21791 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18713), .ZN(n18715) );
  OAI211_X1 U21792 ( .C1(n18742), .C2(n18716), .A(n18715), .B(n18714), .ZN(
        n18764) );
  INV_X1 U21793 ( .A(n18742), .ZN(n18753) );
  NOR2_X1 U21794 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18726), .ZN(
        n18746) );
  INV_X1 U21795 ( .A(n18746), .ZN(n18718) );
  NAND2_X1 U21796 ( .A1(n18892), .A2(n18740), .ZN(n18723) );
  AOI22_X1 U21797 ( .A1(n18719), .A2(n18718), .B1(n18717), .B2(n18723), .ZN(
        n18875) );
  NOR2_X1 U21798 ( .A1(n18753), .A2(n18875), .ZN(n18728) );
  AOI21_X1 U21799 ( .B1(n18722), .B2(n18721), .A(n18720), .ZN(n18730) );
  OAI21_X1 U21800 ( .B1(n18730), .B2(n18724), .A(n18723), .ZN(n18725) );
  AOI21_X1 U21801 ( .B1(n18734), .B2(n18726), .A(n18725), .ZN(n18878) );
  NAND2_X1 U21802 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18878), .ZN(
        n18727) );
  OAI22_X1 U21803 ( .A1(n18728), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18753), .B2(n18727), .ZN(n18762) );
  NOR2_X1 U21804 ( .A1(n9588), .A2(n18905), .ZN(n18733) );
  OAI211_X1 U21805 ( .C1(n18733), .C2(n18732), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18892), .ZN(n18737) );
  OAI211_X1 U21806 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18735), .B(n18734), .ZN(
        n18736) );
  OAI211_X1 U21807 ( .C1(n18888), .C2(n18738), .A(n18737), .B(n18736), .ZN(
        n18739) );
  AOI21_X1 U21808 ( .B1(n18741), .B2(n18740), .A(n18739), .ZN(n18883) );
  AOI22_X1 U21809 ( .A1(n18753), .A2(n18892), .B1(n18883), .B2(n18742), .ZN(
        n18757) );
  NOR2_X1 U21810 ( .A1(n18744), .A2(n18743), .ZN(n18747) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18745), .B1(
        n18747), .B2(n18905), .ZN(n18901) );
  OAI22_X1 U21812 ( .A1(n18747), .A2(n18893), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18746), .ZN(n18897) );
  OR3_X1 U21813 ( .A1(n18901), .A2(n18750), .A3(n18748), .ZN(n18749) );
  AOI22_X1 U21814 ( .A1(n18901), .A2(n18750), .B1(n18897), .B2(n18749), .ZN(
        n18752) );
  OAI21_X1 U21815 ( .B1(n18753), .B2(n18752), .A(n18751), .ZN(n18756) );
  AND2_X1 U21816 ( .A1(n18757), .A2(n18756), .ZN(n18754) );
  OAI221_X1 U21817 ( .B1(n18757), .B2(n18756), .C1(n18755), .C2(n18754), .A(
        n18759), .ZN(n18761) );
  AOI21_X1 U21818 ( .B1(n18759), .B2(n18758), .A(n18757), .ZN(n18760) );
  AOI222_X1 U21819 ( .A1(n18762), .A2(n18761), .B1(n18762), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18761), .C2(n18760), .ZN(
        n18763) );
  NOR4_X1 U21820 ( .A1(n18765), .A2(n18918), .A3(n18764), .A4(n18763), .ZN(
        n18774) );
  NAND2_X1 U21821 ( .A1(n18926), .A2(n18938), .ZN(n18775) );
  NAND2_X1 U21822 ( .A1(n18775), .A2(n18766), .ZN(n18770) );
  OAI211_X1 U21823 ( .C1(n18768), .C2(n18767), .A(n18923), .B(n18774), .ZN(
        n18777) );
  NAND2_X1 U21824 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18777), .ZN(n18870) );
  NAND2_X1 U21825 ( .A1(n18885), .A2(n18938), .ZN(n18784) );
  INV_X1 U21826 ( .A(n18784), .ZN(n18931) );
  AOI22_X1 U21827 ( .A1(n18900), .A2(n18931), .B1(n18926), .B2(n18920), .ZN(
        n18769) );
  OAI21_X1 U21828 ( .B1(n18770), .B2(n18870), .A(n18769), .ZN(n18771) );
  OAI211_X1 U21829 ( .C1(n18774), .C2(n18773), .A(n18772), .B(n18771), .ZN(
        P3_U2996) );
  NAND2_X1 U21830 ( .A1(n18926), .A2(n18920), .ZN(n18780) );
  OR3_X1 U21831 ( .A1(n18885), .A2(n18928), .A3(n18775), .ZN(n18782) );
  NAND4_X1 U21832 ( .A1(n18778), .A2(n18777), .A3(n18776), .A4(n18775), .ZN(
        n18779) );
  NAND4_X1 U21833 ( .A1(n18781), .A2(n18780), .A3(n18782), .A4(n18779), .ZN(
        P3_U2997) );
  AND4_X1 U21834 ( .A1(n18784), .A2(n18783), .A3(n18871), .A4(n18782), .ZN(
        P3_U2998) );
  NOR2_X1 U21835 ( .A1(n18869), .A2(n20859), .ZN(P3_U2999) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18785), .ZN(
        P3_U3000) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18785), .ZN(
        P3_U3001) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18785), .ZN(
        P3_U3002) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18785), .ZN(
        P3_U3003) );
  NOR2_X1 U21840 ( .A1(n18869), .A2(n20809), .ZN(P3_U3004) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18785), .ZN(
        P3_U3005) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18785), .ZN(
        P3_U3006) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18785), .ZN(
        P3_U3007) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18785), .ZN(
        P3_U3008) );
  AND2_X1 U21845 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18785), .ZN(
        P3_U3009) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18785), .ZN(
        P3_U3010) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18785), .ZN(
        P3_U3011) );
  AND2_X1 U21848 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18785), .ZN(
        P3_U3012) );
  AND2_X1 U21849 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18785), .ZN(
        P3_U3013) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18785), .ZN(
        P3_U3014) );
  AND2_X1 U21851 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18785), .ZN(
        P3_U3015) );
  AND2_X1 U21852 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18785), .ZN(
        P3_U3016) );
  AND2_X1 U21853 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18785), .ZN(
        P3_U3017) );
  AND2_X1 U21854 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18785), .ZN(
        P3_U3018) );
  AND2_X1 U21855 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18785), .ZN(
        P3_U3019) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18785), .ZN(
        P3_U3020) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18785), .ZN(P3_U3021) );
  AND2_X1 U21858 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18785), .ZN(P3_U3022) );
  AND2_X1 U21859 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18785), .ZN(P3_U3023) );
  AND2_X1 U21860 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18785), .ZN(P3_U3024) );
  AND2_X1 U21861 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18785), .ZN(P3_U3025) );
  AND2_X1 U21862 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18785), .ZN(P3_U3026) );
  AND2_X1 U21863 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18785), .ZN(P3_U3027) );
  AND2_X1 U21864 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18785), .ZN(P3_U3028) );
  INV_X1 U21865 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18933) );
  INV_X1 U21866 ( .A(NA), .ZN(n20664) );
  OAI22_X1 U21867 ( .A1(n18786), .A2(n19731), .B1(P3_STATE_REG_0__SCAN_IN), 
        .B2(n20664), .ZN(n18787) );
  NOR2_X1 U21868 ( .A1(n18933), .A2(n18787), .ZN(n18789) );
  NAND2_X1 U21869 ( .A1(n18926), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18794) );
  NAND2_X1 U21870 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18794), .ZN(n18797) );
  INV_X1 U21871 ( .A(n18797), .ZN(n18788) );
  OAI22_X1 U21872 ( .A1(n18935), .A2(n18789), .B1(P3_STATE_REG_2__SCAN_IN), 
        .B2(n18788), .ZN(P3_U3029) );
  NOR2_X1 U21873 ( .A1(n18801), .A2(n19731), .ZN(n18796) );
  OAI22_X1 U21874 ( .A1(n18796), .A2(n18933), .B1(n19731), .B2(n18790), .ZN(
        n18791) );
  NAND2_X1 U21875 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18791), .ZN(n18793) );
  NAND3_X1 U21876 ( .A1(n18793), .A2(n18794), .A3(n18792), .ZN(P3_U3030) );
  OAI22_X1 U21877 ( .A1(NA), .A2(n18794), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18795) );
  OAI22_X1 U21878 ( .A1(n18796), .A2(n18795), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18800) );
  OAI211_X1 U21879 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n20664), .A(
        P3_STATE_REG_2__SCAN_IN), .B(n18797), .ZN(n18798) );
  OAI21_X1 U21880 ( .B1(n18800), .B2(n18799), .A(n18798), .ZN(P3_U3031) );
  OAI222_X1 U21881 ( .A1(n18907), .A2(n18861), .B1(n18802), .B2(n18935), .C1(
        n18803), .C2(n18857), .ZN(P3_U3032) );
  OAI222_X1 U21882 ( .A1(n18857), .A2(n18805), .B1(n18804), .B2(n18935), .C1(
        n18803), .C2(n18861), .ZN(P3_U3033) );
  OAI222_X1 U21883 ( .A1(n18857), .A2(n18807), .B1(n18806), .B2(n18935), .C1(
        n18805), .C2(n18861), .ZN(P3_U3034) );
  OAI222_X1 U21884 ( .A1(n18857), .A2(n18809), .B1(n18808), .B2(n18935), .C1(
        n18807), .C2(n18861), .ZN(P3_U3035) );
  OAI222_X1 U21885 ( .A1(n18857), .A2(n18811), .B1(n18810), .B2(n18935), .C1(
        n18809), .C2(n18861), .ZN(P3_U3036) );
  OAI222_X1 U21886 ( .A1(n18857), .A2(n18813), .B1(n18812), .B2(n18935), .C1(
        n18811), .C2(n18861), .ZN(P3_U3037) );
  OAI222_X1 U21887 ( .A1(n18857), .A2(n18816), .B1(n18814), .B2(n18935), .C1(
        n18813), .C2(n18861), .ZN(P3_U3038) );
  OAI222_X1 U21888 ( .A1(n18816), .A2(n18861), .B1(n18815), .B2(n18935), .C1(
        n18817), .C2(n18857), .ZN(P3_U3039) );
  OAI222_X1 U21889 ( .A1(n18857), .A2(n18819), .B1(n18818), .B2(n18935), .C1(
        n18817), .C2(n18861), .ZN(P3_U3040) );
  INV_X1 U21890 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18821) );
  OAI222_X1 U21891 ( .A1(n18857), .A2(n18821), .B1(n18820), .B2(n18935), .C1(
        n18819), .C2(n18861), .ZN(P3_U3041) );
  OAI222_X1 U21892 ( .A1(n18857), .A2(n18823), .B1(n18822), .B2(n18935), .C1(
        n18821), .C2(n18861), .ZN(P3_U3042) );
  INV_X1 U21893 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20777) );
  OAI222_X1 U21894 ( .A1(n18857), .A2(n20777), .B1(n18824), .B2(n18935), .C1(
        n18823), .C2(n18861), .ZN(P3_U3043) );
  OAI222_X1 U21895 ( .A1(n18857), .A2(n18827), .B1(n18825), .B2(n18935), .C1(
        n20777), .C2(n18861), .ZN(P3_U3044) );
  OAI222_X1 U21896 ( .A1(n18827), .A2(n18861), .B1(n18826), .B2(n18935), .C1(
        n18828), .C2(n18857), .ZN(P3_U3045) );
  OAI222_X1 U21897 ( .A1(n18857), .A2(n18830), .B1(n18829), .B2(n18935), .C1(
        n18828), .C2(n18861), .ZN(P3_U3046) );
  OAI222_X1 U21898 ( .A1(n18857), .A2(n18833), .B1(n18831), .B2(n18935), .C1(
        n18830), .C2(n18861), .ZN(P3_U3047) );
  OAI222_X1 U21899 ( .A1(n18833), .A2(n18861), .B1(n18832), .B2(n18935), .C1(
        n18834), .C2(n18857), .ZN(P3_U3048) );
  OAI222_X1 U21900 ( .A1(n18857), .A2(n18836), .B1(n18835), .B2(n18935), .C1(
        n18834), .C2(n18861), .ZN(P3_U3049) );
  OAI222_X1 U21901 ( .A1(n18857), .A2(n18838), .B1(n18837), .B2(n18935), .C1(
        n18836), .C2(n18861), .ZN(P3_U3050) );
  OAI222_X1 U21902 ( .A1(n18857), .A2(n20827), .B1(n18839), .B2(n18935), .C1(
        n18838), .C2(n18861), .ZN(P3_U3051) );
  OAI222_X1 U21903 ( .A1(n20827), .A2(n18861), .B1(n18840), .B2(n18935), .C1(
        n18841), .C2(n18857), .ZN(P3_U3052) );
  OAI222_X1 U21904 ( .A1(n18857), .A2(n18844), .B1(n18842), .B2(n18935), .C1(
        n18841), .C2(n18861), .ZN(P3_U3053) );
  OAI222_X1 U21905 ( .A1(n18844), .A2(n18861), .B1(n18843), .B2(n18935), .C1(
        n18845), .C2(n18857), .ZN(P3_U3054) );
  OAI222_X1 U21906 ( .A1(n18857), .A2(n18847), .B1(n18846), .B2(n18935), .C1(
        n18845), .C2(n18861), .ZN(P3_U3055) );
  OAI222_X1 U21907 ( .A1(n18857), .A2(n18849), .B1(n18848), .B2(n18935), .C1(
        n18847), .C2(n18861), .ZN(P3_U3056) );
  OAI222_X1 U21908 ( .A1(n18857), .A2(n18851), .B1(n18850), .B2(n18935), .C1(
        n18849), .C2(n18861), .ZN(P3_U3057) );
  INV_X1 U21909 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18854) );
  OAI222_X1 U21910 ( .A1(n18857), .A2(n18854), .B1(n18852), .B2(n18935), .C1(
        n18851), .C2(n18861), .ZN(P3_U3058) );
  OAI222_X1 U21911 ( .A1(n18854), .A2(n18861), .B1(n18853), .B2(n18935), .C1(
        n18855), .C2(n18857), .ZN(P3_U3059) );
  OAI222_X1 U21912 ( .A1(n18857), .A2(n18860), .B1(n18856), .B2(n18935), .C1(
        n18855), .C2(n18861), .ZN(P3_U3060) );
  OAI222_X1 U21913 ( .A1(n18861), .A2(n18860), .B1(n18859), .B2(n18935), .C1(
        n18858), .C2(n18857), .ZN(P3_U3061) );
  OAI22_X1 U21914 ( .A1(n18936), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18935), .ZN(n18862) );
  INV_X1 U21915 ( .A(n18862), .ZN(P3_U3274) );
  OAI22_X1 U21916 ( .A1(n18936), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18935), .ZN(n18863) );
  INV_X1 U21917 ( .A(n18863), .ZN(P3_U3275) );
  OAI22_X1 U21918 ( .A1(n18936), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18935), .ZN(n18864) );
  INV_X1 U21919 ( .A(n18864), .ZN(P3_U3276) );
  OAI22_X1 U21920 ( .A1(n18936), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18935), .ZN(n18865) );
  INV_X1 U21921 ( .A(n18865), .ZN(P3_U3277) );
  OAI21_X1 U21922 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n18869), .A(n18867), 
        .ZN(n18866) );
  INV_X1 U21923 ( .A(n18866), .ZN(P3_U3280) );
  OAI21_X1 U21924 ( .B1(n18869), .B2(n18868), .A(n18867), .ZN(P3_U3281) );
  INV_X1 U21925 ( .A(n18870), .ZN(n18873) );
  OAI21_X1 U21926 ( .B1(n18873), .B2(n18872), .A(n18871), .ZN(P3_U3282) );
  INV_X1 U21927 ( .A(n18874), .ZN(n18877) );
  NOR3_X1 U21928 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18875), .A3(
        n18884), .ZN(n18876) );
  AOI21_X1 U21929 ( .B1(n18877), .B2(n18900), .A(n18876), .ZN(n18882) );
  INV_X1 U21930 ( .A(n18906), .ZN(n18903) );
  OAI21_X1 U21931 ( .B1(n18884), .B2(n18878), .A(n18903), .ZN(n18879) );
  INV_X1 U21932 ( .A(n18879), .ZN(n18881) );
  OAI22_X1 U21933 ( .A1(n18906), .A2(n18882), .B1(n18881), .B2(n18880), .ZN(
        P3_U3285) );
  INV_X1 U21934 ( .A(n18883), .ZN(n18890) );
  INV_X1 U21935 ( .A(n18884), .ZN(n18939) );
  NOR2_X1 U21936 ( .A1(n18885), .A2(n18902), .ZN(n18894) );
  OAI22_X1 U21937 ( .A1(n18887), .A2(n18886), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18895) );
  INV_X1 U21938 ( .A(n18895), .ZN(n18889) );
  AOI222_X1 U21939 ( .A1(n18890), .A2(n18939), .B1(n18894), .B2(n18889), .C1(
        n18900), .C2(n18888), .ZN(n18891) );
  AOI22_X1 U21940 ( .A1(n18906), .A2(n18892), .B1(n18891), .B2(n18903), .ZN(
        P3_U3288) );
  INV_X1 U21941 ( .A(n18893), .ZN(n18896) );
  AOI222_X1 U21942 ( .A1(n18897), .A2(n18939), .B1(n18900), .B2(n18896), .C1(
        n18895), .C2(n18894), .ZN(n18898) );
  AOI22_X1 U21943 ( .A1(n18906), .A2(n18899), .B1(n18898), .B2(n18903), .ZN(
        P3_U3289) );
  AOI222_X1 U21944 ( .A1(n18902), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18939), 
        .B2(n18901), .C1(n18905), .C2(n18900), .ZN(n18904) );
  AOI22_X1 U21945 ( .A1(n18906), .A2(n18905), .B1(n18904), .B2(n18903), .ZN(
        P3_U3290) );
  AOI21_X1 U21946 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18908) );
  AOI22_X1 U21947 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18908), .B2(n18907), .ZN(n18910) );
  INV_X1 U21948 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18909) );
  AOI22_X1 U21949 ( .A1(n18911), .A2(n18910), .B1(n18909), .B2(n18914), .ZN(
        P3_U3292) );
  INV_X1 U21950 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18915) );
  NOR2_X1 U21951 ( .A1(n18914), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18912) );
  AOI22_X1 U21952 ( .A1(n18915), .A2(n18914), .B1(n18913), .B2(n18912), .ZN(
        P3_U3293) );
  INV_X1 U21953 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18942) );
  OAI22_X1 U21954 ( .A1(n18936), .A2(n18942), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18935), .ZN(n18916) );
  INV_X1 U21955 ( .A(n18916), .ZN(P3_U3294) );
  MUX2_X1 U21956 ( .A(P3_MORE_REG_SCAN_IN), .B(n18918), .S(n18917), .Z(
        P3_U3295) );
  AOI21_X1 U21957 ( .B1(n18920), .B2(n18919), .A(n18941), .ZN(n18921) );
  OAI21_X1 U21958 ( .B1(n18923), .B2(n18922), .A(n18921), .ZN(n18934) );
  OAI21_X1 U21959 ( .B1(n18925), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n18924), 
        .ZN(n18927) );
  AOI211_X1 U21960 ( .C1(n18940), .C2(n18927), .A(n18926), .B(n18938), .ZN(
        n18929) );
  NOR2_X1 U21961 ( .A1(n18929), .A2(n18928), .ZN(n18930) );
  OAI21_X1 U21962 ( .B1(n18931), .B2(n18930), .A(n18934), .ZN(n18932) );
  OAI21_X1 U21963 ( .B1(n18934), .B2(n18933), .A(n18932), .ZN(P3_U3296) );
  OAI22_X1 U21964 ( .A1(n18936), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18935), .ZN(n18937) );
  INV_X1 U21965 ( .A(n18937), .ZN(P3_U3297) );
  AOI21_X1 U21966 ( .B1(n18939), .B2(n18938), .A(n18941), .ZN(n18945) );
  AOI22_X1 U21967 ( .A1(n18945), .A2(n18942), .B1(n18941), .B2(n18940), .ZN(
        P3_U3298) );
  INV_X1 U21968 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18944) );
  AOI21_X1 U21969 ( .B1(n18945), .B2(n18944), .A(n18943), .ZN(P3_U3299) );
  AOI21_X1 U21970 ( .B1(n18947), .B2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n18946), 
        .ZN(n18948) );
  OAI21_X1 U21971 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n19552), .A(n18948), 
        .ZN(P2_U2814) );
  INV_X1 U21972 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18955) );
  NAND2_X1 U21973 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20815), .ZN(n19730) );
  NAND2_X1 U21974 ( .A1(n18955), .A2(n18949), .ZN(n19727) );
  OAI21_X1 U21975 ( .B1(n18955), .B2(n19730), .A(n19727), .ZN(n19796) );
  AOI21_X1 U21976 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19796), .ZN(n18950) );
  INV_X1 U21977 ( .A(n18950), .ZN(P2_U2815) );
  INV_X1 U21978 ( .A(n18951), .ZN(n18953) );
  AOI22_X1 U21979 ( .A1(n18953), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18952), 
        .B2(n19715), .ZN(n18954) );
  INV_X1 U21980 ( .A(n18954), .ZN(P2_U2816) );
  NAND2_X1 U21981 ( .A1(n18955), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19847) );
  INV_X2 U21982 ( .A(n19847), .ZN(n19783) );
  INV_X1 U21983 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n20875) );
  OAI21_X1 U21984 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n20815), .A(n18955), 
        .ZN(n18956) );
  AOI22_X1 U21985 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n19783), .B1(n20875), 
        .B2(n18956), .ZN(P2_U2817) );
  OAI21_X1 U21986 ( .B1(n19721), .B2(BS16), .A(n19796), .ZN(n19794) );
  OAI21_X1 U21987 ( .B1(n19796), .B2(n18957), .A(n19794), .ZN(P2_U2818) );
  NOR4_X1 U21988 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18961) );
  NOR4_X1 U21989 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18960) );
  NOR4_X1 U21990 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18959) );
  NOR4_X1 U21991 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18958) );
  NAND4_X1 U21992 ( .A1(n18961), .A2(n18960), .A3(n18959), .A4(n18958), .ZN(
        n18967) );
  NOR4_X1 U21993 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18965) );
  AOI211_X1 U21994 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_17__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18964) );
  NOR4_X1 U21995 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18963) );
  NOR4_X1 U21996 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18962) );
  NAND4_X1 U21997 ( .A1(n18965), .A2(n18964), .A3(n18963), .A4(n18962), .ZN(
        n18966) );
  NOR2_X1 U21998 ( .A1(n18967), .A2(n18966), .ZN(n18977) );
  INV_X1 U21999 ( .A(n18977), .ZN(n18975) );
  NOR2_X1 U22000 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18975), .ZN(n18970) );
  INV_X1 U22001 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18968) );
  AOI22_X1 U22002 ( .A1(n18970), .A2(n12092), .B1(n18975), .B2(n18968), .ZN(
        P2_U2820) );
  OR3_X1 U22003 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18974) );
  INV_X1 U22004 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18969) );
  AOI22_X1 U22005 ( .A1(n18970), .A2(n18974), .B1(n18975), .B2(n18969), .ZN(
        P2_U2821) );
  INV_X1 U22006 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19795) );
  NAND2_X1 U22007 ( .A1(n18970), .A2(n19795), .ZN(n18973) );
  OAI21_X1 U22008 ( .B1(n12092), .B2(n12076), .A(n18977), .ZN(n18971) );
  OAI21_X1 U22009 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18977), .A(n18971), 
        .ZN(n18972) );
  OAI221_X1 U22010 ( .B1(n18973), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18973), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18972), .ZN(P2_U2822) );
  INV_X1 U22011 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18976) );
  OAI221_X1 U22012 ( .B1(n18977), .B2(n18976), .C1(n18975), .C2(n18974), .A(
        n18973), .ZN(P2_U2823) );
  NAND2_X1 U22013 ( .A1(n9591), .A2(n18978), .ZN(n18979) );
  XOR2_X1 U22014 ( .A(n18980), .B(n18979), .Z(n18989) );
  INV_X1 U22015 ( .A(n18981), .ZN(n18983) );
  AOI22_X1 U22016 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19103), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19087), .ZN(n18982) );
  OAI21_X1 U22017 ( .B1(n18983), .B2(n19075), .A(n18982), .ZN(n18984) );
  AOI211_X1 U22018 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19112), .A(n19111), 
        .B(n18984), .ZN(n18988) );
  AOI22_X1 U22019 ( .A1(n18986), .A2(n19115), .B1(n18985), .B2(n19070), .ZN(
        n18987) );
  OAI211_X1 U22020 ( .C1(n19717), .C2(n18989), .A(n18988), .B(n18987), .ZN(
        P2_U2836) );
  OAI21_X1 U22021 ( .B1(n19764), .B2(n19091), .A(n11795), .ZN(n18992) );
  OAI22_X1 U22022 ( .A1(n18990), .A2(n19075), .B1(n13497), .B2(n19109), .ZN(
        n18991) );
  AOI211_X1 U22023 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19103), .A(
        n18992), .B(n18991), .ZN(n18999) );
  NOR2_X1 U22024 ( .A1(n19094), .A2(n18993), .ZN(n18995) );
  XNOR2_X1 U22025 ( .A(n18995), .B(n18994), .ZN(n18997) );
  AOI22_X1 U22026 ( .A1(n18997), .A2(n19098), .B1(n18996), .B2(n19115), .ZN(
        n18998) );
  OAI211_X1 U22027 ( .C1(n19000), .C2(n19107), .A(n18999), .B(n18998), .ZN(
        P2_U2837) );
  NAND2_X1 U22028 ( .A1(n9591), .A2(n19001), .ZN(n19002) );
  XOR2_X1 U22029 ( .A(n19003), .B(n19002), .Z(n19013) );
  INV_X1 U22030 ( .A(n19004), .ZN(n19006) );
  AOI22_X1 U22031 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19103), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19087), .ZN(n19005) );
  OAI21_X1 U22032 ( .B1(n19006), .B2(n19075), .A(n19005), .ZN(n19007) );
  AOI211_X1 U22033 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19112), .A(n19111), 
        .B(n19007), .ZN(n19012) );
  INV_X1 U22034 ( .A(n19008), .ZN(n19010) );
  AOI22_X1 U22035 ( .A1(n19010), .A2(n19115), .B1(n19070), .B2(n19009), .ZN(
        n19011) );
  OAI211_X1 U22036 ( .C1(n19717), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        P2_U2838) );
  NOR2_X1 U22037 ( .A1(n19094), .A2(n19014), .ZN(n19015) );
  XOR2_X1 U22038 ( .A(n19016), .B(n19015), .Z(n19026) );
  AOI22_X1 U22039 ( .A1(n19017), .A2(n19104), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19087), .ZN(n19018) );
  OAI211_X1 U22040 ( .C1(n19761), .C2(n19091), .A(n19018), .B(n19089), .ZN(
        n19024) );
  INV_X1 U22041 ( .A(n19019), .ZN(n19022) );
  OAI22_X1 U22042 ( .A1(n19022), .A2(n19021), .B1(n19107), .B2(n19020), .ZN(
        n19023) );
  AOI211_X1 U22043 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19103), .A(
        n19024), .B(n19023), .ZN(n19025) );
  OAI21_X1 U22044 ( .B1(n19717), .B2(n19026), .A(n19025), .ZN(P2_U2839) );
  OAI21_X1 U22045 ( .B1(n19759), .B2(n19091), .A(n11795), .ZN(n19029) );
  OAI22_X1 U22046 ( .A1(n19027), .A2(n19075), .B1(n14832), .B2(n19109), .ZN(
        n19028) );
  AOI211_X1 U22047 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19103), .A(
        n19029), .B(n19028), .ZN(n19036) );
  NAND2_X1 U22048 ( .A1(n9591), .A2(n19030), .ZN(n19032) );
  XNOR2_X1 U22049 ( .A(n19032), .B(n19031), .ZN(n19034) );
  AOI22_X1 U22050 ( .A1(n19034), .A2(n19098), .B1(n19115), .B2(n19033), .ZN(
        n19035) );
  OAI211_X1 U22051 ( .C1(n19037), .C2(n19107), .A(n19036), .B(n19035), .ZN(
        P2_U2840) );
  INV_X1 U22052 ( .A(n19038), .ZN(n19040) );
  AOI22_X1 U22053 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19103), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19087), .ZN(n19039) );
  OAI21_X1 U22054 ( .B1(n19040), .B2(n19075), .A(n19039), .ZN(n19041) );
  AOI211_X1 U22055 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19112), .A(n19111), 
        .B(n19041), .ZN(n19048) );
  NOR2_X1 U22056 ( .A1(n19094), .A2(n19042), .ZN(n19044) );
  XNOR2_X1 U22057 ( .A(n19044), .B(n19043), .ZN(n19046) );
  AOI22_X1 U22058 ( .A1(n19046), .A2(n19098), .B1(n19115), .B2(n19045), .ZN(
        n19047) );
  OAI211_X1 U22059 ( .C1(n19049), .C2(n19107), .A(n19048), .B(n19047), .ZN(
        P2_U2841) );
  OAI22_X1 U22060 ( .A1(n19050), .A2(n19075), .B1(n19109), .B2(n12713), .ZN(
        n19051) );
  INV_X1 U22061 ( .A(n19051), .ZN(n19052) );
  OAI211_X1 U22062 ( .C1(n19755), .C2(n19091), .A(n19052), .B(n19089), .ZN(
        n19053) );
  AOI21_X1 U22063 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19103), .A(
        n19053), .ZN(n19060) );
  NOR2_X1 U22064 ( .A1(n19094), .A2(n19054), .ZN(n19056) );
  XNOR2_X1 U22065 ( .A(n19056), .B(n19055), .ZN(n19058) );
  AOI22_X1 U22066 ( .A1(n19058), .A2(n19098), .B1(n19115), .B2(n19057), .ZN(
        n19059) );
  OAI211_X1 U22067 ( .C1(n19061), .C2(n19107), .A(n19060), .B(n19059), .ZN(
        P2_U2843) );
  NAND2_X1 U22068 ( .A1(n9591), .A2(n19062), .ZN(n19063) );
  XOR2_X1 U22069 ( .A(n19064), .B(n19063), .Z(n19074) );
  INV_X1 U22070 ( .A(n19065), .ZN(n19066) );
  AOI22_X1 U22071 ( .A1(n19066), .A2(n19104), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19103), .ZN(n19067) );
  OAI21_X1 U22072 ( .B1(n19109), .B2(n19068), .A(n19067), .ZN(n19069) );
  AOI211_X1 U22073 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19112), .A(n19111), 
        .B(n19069), .ZN(n19073) );
  AOI22_X1 U22074 ( .A1(n19071), .A2(n19115), .B1(n19070), .B2(n19141), .ZN(
        n19072) );
  OAI211_X1 U22075 ( .C1(n19717), .C2(n19074), .A(n19073), .B(n19072), .ZN(
        P2_U2844) );
  OAI21_X1 U22076 ( .B1(n12675), .B2(n19091), .A(n11795), .ZN(n19078) );
  OAI22_X1 U22077 ( .A1(n19076), .A2(n19075), .B1(n19109), .B2(n20801), .ZN(
        n19077) );
  AOI211_X1 U22078 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19103), .A(
        n19078), .B(n19077), .ZN(n19085) );
  NOR2_X1 U22079 ( .A1(n19094), .A2(n19079), .ZN(n19081) );
  XNOR2_X1 U22080 ( .A(n19081), .B(n19080), .ZN(n19083) );
  AOI22_X1 U22081 ( .A1(n19083), .A2(n19098), .B1(n19115), .B2(n19082), .ZN(
        n19084) );
  OAI211_X1 U22082 ( .C1(n19086), .C2(n19107), .A(n19085), .B(n19084), .ZN(
        P2_U2845) );
  AOI22_X1 U22083 ( .A1(n19088), .A2(n19104), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19087), .ZN(n19090) );
  OAI211_X1 U22084 ( .C1(n15413), .C2(n19091), .A(n19090), .B(n19089), .ZN(
        n19092) );
  AOI21_X1 U22085 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19103), .A(
        n19092), .ZN(n19101) );
  NOR2_X1 U22086 ( .A1(n19094), .A2(n19093), .ZN(n19096) );
  XNOR2_X1 U22087 ( .A(n19096), .B(n19095), .ZN(n19099) );
  AOI22_X1 U22088 ( .A1(n19099), .A2(n19098), .B1(n19115), .B2(n19097), .ZN(
        n19100) );
  OAI211_X1 U22089 ( .C1(n19102), .C2(n19107), .A(n19101), .B(n19100), .ZN(
        P2_U2847) );
  AOI22_X1 U22090 ( .A1(n19105), .A2(n19104), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19103), .ZN(n19126) );
  OAI22_X1 U22091 ( .A1(n19109), .A2(n19108), .B1(n19107), .B2(n19106), .ZN(
        n19110) );
  AOI211_X1 U22092 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19112), .A(n19111), .B(
        n19110), .ZN(n19125) );
  INV_X1 U22093 ( .A(n19113), .ZN(n19114) );
  AOI22_X1 U22094 ( .A1(n19117), .A2(n19116), .B1(n19115), .B2(n19114), .ZN(
        n19124) );
  INV_X1 U22095 ( .A(n19118), .ZN(n19122) );
  NOR2_X1 U22096 ( .A1(n19094), .A2(n19119), .ZN(n19121) );
  AOI21_X1 U22097 ( .B1(n19122), .B2(n19121), .A(n19717), .ZN(n19120) );
  OAI21_X1 U22098 ( .B1(n19122), .B2(n19121), .A(n19120), .ZN(n19123) );
  NAND4_X1 U22099 ( .A1(n19126), .A2(n19125), .A3(n19124), .A4(n19123), .ZN(
        P2_U2851) );
  INV_X1 U22100 ( .A(n19127), .ZN(n19128) );
  AOI22_X1 U22101 ( .A1(n19130), .A2(BUF2_REG_31__SCAN_IN), .B1(n19129), .B2(
        n19128), .ZN(n19134) );
  AOI22_X1 U22102 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19132), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19131), .ZN(n19133) );
  NAND2_X1 U22103 ( .A1(n19134), .A2(n19133), .ZN(P2_U2888) );
  INV_X1 U22104 ( .A(n19135), .ZN(n19142) );
  AOI22_X1 U22105 ( .A1(n19142), .A2(n19137), .B1(n19140), .B2(n19136), .ZN(
        n19138) );
  OAI21_X1 U22106 ( .B1(n19144), .B2(n20783), .A(n19138), .ZN(P2_U2906) );
  AOI22_X1 U22107 ( .A1(n19142), .A2(n19141), .B1(n19140), .B2(n19139), .ZN(
        n19143) );
  OAI21_X1 U22108 ( .B1(n19144), .B2(n19189), .A(n19143), .ZN(P2_U2908) );
  OAI21_X1 U22109 ( .B1(n19147), .B2(n19146), .A(n19145), .ZN(n19148) );
  AND2_X1 U22110 ( .A1(n19148), .A2(n19726), .ZN(n19180) );
  AND2_X1 U22111 ( .A1(n19197), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NAND2_X1 U22112 ( .A1(n19180), .A2(n19149), .ZN(n19178) );
  AOI22_X1 U22113 ( .A1(n19190), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22114 ( .B1(n19151), .B2(n19178), .A(n19150), .ZN(P2_U2921) );
  AOI22_X1 U22115 ( .A1(n19190), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19152) );
  OAI21_X1 U22116 ( .B1(n19153), .B2(n19178), .A(n19152), .ZN(P2_U2922) );
  INV_X1 U22117 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19155) );
  AOI22_X1 U22118 ( .A1(n19190), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19154) );
  OAI21_X1 U22119 ( .B1(n19155), .B2(n19178), .A(n19154), .ZN(P2_U2923) );
  AOI22_X1 U22120 ( .A1(n19190), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19156) );
  OAI21_X1 U22121 ( .B1(n19157), .B2(n19178), .A(n19156), .ZN(P2_U2924) );
  AOI22_X1 U22122 ( .A1(n19190), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22123 ( .B1(n20893), .B2(n19178), .A(n19158), .ZN(P2_U2925) );
  AOI22_X1 U22124 ( .A1(n19190), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U22125 ( .B1(n19160), .B2(n19178), .A(n19159), .ZN(P2_U2926) );
  AOI22_X1 U22126 ( .A1(n19190), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19161) );
  OAI21_X1 U22127 ( .B1(n19162), .B2(n19178), .A(n19161), .ZN(P2_U2927) );
  INV_X1 U22128 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22129 ( .A1(n19190), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U22130 ( .B1(n19164), .B2(n19178), .A(n19163), .ZN(P2_U2928) );
  INV_X1 U22131 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19166) );
  AOI22_X1 U22132 ( .A1(n19190), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19165) );
  OAI21_X1 U22133 ( .B1(n19166), .B2(n19178), .A(n19165), .ZN(P2_U2929) );
  INV_X1 U22134 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19168) );
  AOI22_X1 U22135 ( .A1(n19190), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19167) );
  OAI21_X1 U22136 ( .B1(n19168), .B2(n19178), .A(n19167), .ZN(P2_U2930) );
  INV_X1 U22137 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19170) );
  AOI22_X1 U22138 ( .A1(n19190), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19169) );
  OAI21_X1 U22139 ( .B1(n19170), .B2(n19178), .A(n19169), .ZN(P2_U2931) );
  INV_X1 U22140 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19172) );
  AOI22_X1 U22141 ( .A1(n19190), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22142 ( .B1(n19172), .B2(n19178), .A(n19171), .ZN(P2_U2932) );
  INV_X1 U22143 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19174) );
  AOI22_X1 U22144 ( .A1(n19190), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19173) );
  OAI21_X1 U22145 ( .B1(n19174), .B2(n19178), .A(n19173), .ZN(P2_U2933) );
  INV_X1 U22146 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19176) );
  AOI22_X1 U22147 ( .A1(n19190), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19175) );
  OAI21_X1 U22148 ( .B1(n19176), .B2(n19178), .A(n19175), .ZN(P2_U2934) );
  INV_X1 U22149 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19179) );
  AOI22_X1 U22150 ( .A1(n19190), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19177) );
  OAI21_X1 U22151 ( .B1(n19179), .B2(n19178), .A(n19177), .ZN(P2_U2935) );
  AOI22_X1 U22152 ( .A1(n19190), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22153 ( .B1(n19182), .B2(n19212), .A(n19181), .ZN(P2_U2936) );
  AOI22_X1 U22154 ( .A1(n19190), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U22155 ( .B1(n19184), .B2(n19212), .A(n19183), .ZN(P2_U2937) );
  AOI22_X1 U22156 ( .A1(n19190), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U22157 ( .B1(n20783), .B2(n19212), .A(n19185), .ZN(P2_U2938) );
  AOI22_X1 U22158 ( .A1(n19190), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U22159 ( .B1(n19187), .B2(n19212), .A(n19186), .ZN(P2_U2939) );
  AOI22_X1 U22160 ( .A1(n19190), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22161 ( .B1(n19189), .B2(n19212), .A(n19188), .ZN(P2_U2940) );
  AOI22_X1 U22162 ( .A1(n19190), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22163 ( .B1(n19192), .B2(n19212), .A(n19191), .ZN(P2_U2941) );
  INV_X1 U22164 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19194) );
  AOI22_X1 U22165 ( .A1(n19210), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22166 ( .B1(n19194), .B2(n19212), .A(n19193), .ZN(P2_U2942) );
  AOI22_X1 U22167 ( .A1(n19210), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U22168 ( .B1(n20780), .B2(n19212), .A(n19195), .ZN(P2_U2943) );
  AOI22_X1 U22169 ( .A1(n19210), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22170 ( .B1(n12334), .B2(n19212), .A(n19196), .ZN(P2_U2944) );
  AOI22_X1 U22171 ( .A1(n19210), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19197), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22172 ( .B1(n12085), .B2(n19212), .A(n19198), .ZN(P2_U2945) );
  INV_X1 U22173 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22174 ( .A1(n19210), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22175 ( .B1(n19200), .B2(n19212), .A(n19199), .ZN(P2_U2946) );
  AOI22_X1 U22176 ( .A1(n19210), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22177 ( .B1(n19202), .B2(n19212), .A(n19201), .ZN(P2_U2947) );
  INV_X1 U22178 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19204) );
  AOI22_X1 U22179 ( .A1(n19210), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U22180 ( .B1(n19204), .B2(n19212), .A(n19203), .ZN(P2_U2948) );
  INV_X1 U22181 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19206) );
  AOI22_X1 U22182 ( .A1(n19210), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22183 ( .B1(n19206), .B2(n19212), .A(n19205), .ZN(P2_U2949) );
  INV_X1 U22184 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19208) );
  AOI22_X1 U22185 ( .A1(n19210), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22186 ( .B1(n19208), .B2(n19212), .A(n19207), .ZN(P2_U2950) );
  AOI22_X1 U22187 ( .A1(n19210), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19209), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22188 ( .B1(n19213), .B2(n19212), .A(n19211), .ZN(P2_U2951) );
  INV_X1 U22189 ( .A(n19214), .ZN(n19217) );
  AOI22_X1 U22190 ( .A1(n19217), .A2(n19216), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19215), .ZN(n19229) );
  NOR3_X1 U22191 ( .A1(n19220), .A2(n19219), .A3(n19218), .ZN(n19226) );
  INV_X1 U22192 ( .A(n19221), .ZN(n19222) );
  OAI21_X1 U22193 ( .B1(n19224), .B2(n19223), .A(n19222), .ZN(n19225) );
  AOI211_X1 U22194 ( .C1(n9592), .C2(n19227), .A(n19226), .B(n19225), .ZN(
        n19228) );
  NAND2_X1 U22195 ( .A1(n19229), .A2(n19228), .ZN(P2_U3012) );
  AOI22_X1 U22196 ( .A1(n19615), .A2(n19707), .B1(n19246), .B2(n19666), .ZN(
        n19232) );
  AOI22_X1 U22197 ( .A1(n19667), .A2(n19247), .B1(n19252), .B2(n19668), .ZN(
        n19231) );
  OAI211_X1 U22198 ( .C1(n19251), .C2(n11361), .A(n19232), .B(n19231), .ZN(
        P2_U3049) );
  AOI22_X1 U22199 ( .A1(n19619), .A2(n19707), .B1(n19246), .B2(n19672), .ZN(
        n19235) );
  AOI22_X1 U22200 ( .A1(n19673), .A2(n19247), .B1(n19252), .B2(n19674), .ZN(
        n19234) );
  OAI211_X1 U22201 ( .C1(n19251), .C2(n12191), .A(n19235), .B(n19234), .ZN(
        P2_U3050) );
  AOI22_X1 U22202 ( .A1(n19623), .A2(n19707), .B1(n19246), .B2(n19678), .ZN(
        n19238) );
  AOI22_X1 U22203 ( .A1(n19679), .A2(n19247), .B1(n19252), .B2(n19680), .ZN(
        n19237) );
  OAI211_X1 U22204 ( .C1(n19251), .C2(n20842), .A(n19238), .B(n19237), .ZN(
        P2_U3051) );
  AOI22_X1 U22205 ( .A1(n19627), .A2(n19707), .B1(n19246), .B2(n19684), .ZN(
        n19241) );
  AOI22_X1 U22206 ( .A1(n19685), .A2(n19247), .B1(n19252), .B2(n19686), .ZN(
        n19240) );
  OAI211_X1 U22207 ( .C1(n19251), .C2(n12466), .A(n19241), .B(n19240), .ZN(
        P2_U3052) );
  AOI22_X1 U22208 ( .A1(n19631), .A2(n19707), .B1(n19246), .B2(n19690), .ZN(
        n19244) );
  AOI22_X1 U22209 ( .A1(n19691), .A2(n19247), .B1(n19252), .B2(n19692), .ZN(
        n19243) );
  OAI211_X1 U22210 ( .C1(n19251), .C2(n12490), .A(n19244), .B(n19243), .ZN(
        P2_U3053) );
  INV_X1 U22211 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19250) );
  AOI22_X1 U22212 ( .A1(n19641), .A2(n19707), .B1(n19246), .B2(n19703), .ZN(
        n19249) );
  AOI22_X1 U22213 ( .A1(n19704), .A2(n19247), .B1(n19252), .B2(n19706), .ZN(
        n19248) );
  OAI211_X1 U22214 ( .C1(n19251), .C2(n19250), .A(n19249), .B(n19248), .ZN(
        P2_U3055) );
  INV_X1 U22215 ( .A(n19258), .ZN(n19254) );
  NOR2_X1 U22216 ( .A1(n19461), .A2(n19253), .ZN(n19275) );
  OAI21_X1 U22217 ( .B1(n19254), .B2(n19275), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19255) );
  OAI21_X1 U22218 ( .B1(n19256), .B2(n19552), .A(n19255), .ZN(n19276) );
  AOI22_X1 U22219 ( .A1(n19276), .A2(n19653), .B1(n19652), .B2(n19275), .ZN(
        n19262) );
  OAI21_X1 U22220 ( .B1(n19399), .B2(n19469), .A(n19256), .ZN(n19260) );
  INV_X1 U22221 ( .A(n19275), .ZN(n19257) );
  OAI211_X1 U22222 ( .C1(n19258), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19257), 
        .B(n19552), .ZN(n19259) );
  NAND3_X1 U22223 ( .A1(n19260), .A2(n19655), .A3(n19259), .ZN(n19277) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19662), .ZN(n19261) );
  OAI211_X1 U22225 ( .C1(n19665), .C2(n19280), .A(n19262), .B(n19261), .ZN(
        P2_U3056) );
  AOI22_X1 U22226 ( .A1(n19276), .A2(n19667), .B1(n19666), .B2(n19275), .ZN(
        n19264) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19668), .ZN(n19263) );
  OAI211_X1 U22228 ( .C1(n19671), .C2(n19280), .A(n19264), .B(n19263), .ZN(
        P2_U3057) );
  AOI22_X1 U22229 ( .A1(n19276), .A2(n19673), .B1(n19672), .B2(n19275), .ZN(
        n19266) );
  AOI22_X1 U22230 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19674), .ZN(n19265) );
  OAI211_X1 U22231 ( .C1(n19677), .C2(n19280), .A(n19266), .B(n19265), .ZN(
        P2_U3058) );
  AOI22_X1 U22232 ( .A1(n19276), .A2(n19679), .B1(n19678), .B2(n19275), .ZN(
        n19268) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19680), .ZN(n19267) );
  OAI211_X1 U22234 ( .C1(n19683), .C2(n19280), .A(n19268), .B(n19267), .ZN(
        P2_U3059) );
  AOI22_X1 U22235 ( .A1(n19276), .A2(n19685), .B1(n19684), .B2(n19275), .ZN(
        n19270) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19686), .ZN(n19269) );
  OAI211_X1 U22237 ( .C1(n19689), .C2(n19280), .A(n19270), .B(n19269), .ZN(
        P2_U3060) );
  AOI22_X1 U22238 ( .A1(n19276), .A2(n19691), .B1(n19690), .B2(n19275), .ZN(
        n19272) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19692), .ZN(n19271) );
  OAI211_X1 U22240 ( .C1(n19695), .C2(n19280), .A(n19272), .B(n19271), .ZN(
        P2_U3061) );
  AOI22_X1 U22241 ( .A1(n19276), .A2(n19697), .B1(n19696), .B2(n19275), .ZN(
        n19274) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19698), .ZN(n19273) );
  OAI211_X1 U22243 ( .C1(n19701), .C2(n19280), .A(n19274), .B(n19273), .ZN(
        P2_U3062) );
  AOI22_X1 U22244 ( .A1(n19276), .A2(n19704), .B1(n19703), .B2(n19275), .ZN(
        n19279) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19277), .B1(
        n19298), .B2(n19706), .ZN(n19278) );
  OAI211_X1 U22246 ( .C1(n19712), .C2(n19280), .A(n19279), .B(n19278), .ZN(
        P2_U3063) );
  INV_X1 U22247 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19283) );
  AOI22_X1 U22248 ( .A1(n19297), .A2(n19667), .B1(n19296), .B2(n19666), .ZN(
        n19282) );
  AOI22_X1 U22249 ( .A1(n19299), .A2(n19668), .B1(n19298), .B2(n19615), .ZN(
        n19281) );
  OAI211_X1 U22250 ( .C1(n19303), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P2_U3065) );
  INV_X1 U22251 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19286) );
  AOI22_X1 U22252 ( .A1(n19297), .A2(n19673), .B1(n19296), .B2(n19672), .ZN(
        n19285) );
  AOI22_X1 U22253 ( .A1(n19299), .A2(n19674), .B1(n19298), .B2(n19619), .ZN(
        n19284) );
  OAI211_X1 U22254 ( .C1(n19303), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        P2_U3066) );
  AOI22_X1 U22255 ( .A1(n19297), .A2(n19679), .B1(n19296), .B2(n19678), .ZN(
        n19288) );
  AOI22_X1 U22256 ( .A1(n19299), .A2(n19680), .B1(n19298), .B2(n19623), .ZN(
        n19287) );
  OAI211_X1 U22257 ( .C1(n19303), .C2(n11433), .A(n19288), .B(n19287), .ZN(
        P2_U3067) );
  INV_X1 U22258 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19291) );
  AOI22_X1 U22259 ( .A1(n19297), .A2(n19685), .B1(n19296), .B2(n19684), .ZN(
        n19290) );
  AOI22_X1 U22260 ( .A1(n19299), .A2(n19686), .B1(n19298), .B2(n19627), .ZN(
        n19289) );
  OAI211_X1 U22261 ( .C1(n19303), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P2_U3068) );
  AOI22_X1 U22262 ( .A1(n19297), .A2(n19691), .B1(n19296), .B2(n19690), .ZN(
        n19293) );
  AOI22_X1 U22263 ( .A1(n19299), .A2(n19692), .B1(n19298), .B2(n19631), .ZN(
        n19292) );
  OAI211_X1 U22264 ( .C1(n19303), .C2(n11482), .A(n19293), .B(n19292), .ZN(
        P2_U3069) );
  AOI22_X1 U22265 ( .A1(n19297), .A2(n19697), .B1(n19296), .B2(n19696), .ZN(
        n19295) );
  AOI22_X1 U22266 ( .A1(n19299), .A2(n19698), .B1(n19298), .B2(n19635), .ZN(
        n19294) );
  OAI211_X1 U22267 ( .C1(n19303), .C2(n11522), .A(n19295), .B(n19294), .ZN(
        P2_U3070) );
  INV_X1 U22268 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19302) );
  AOI22_X1 U22269 ( .A1(n19297), .A2(n19704), .B1(n19296), .B2(n19703), .ZN(
        n19301) );
  AOI22_X1 U22270 ( .A1(n19299), .A2(n19706), .B1(n19298), .B2(n19641), .ZN(
        n19300) );
  OAI211_X1 U22271 ( .C1(n19303), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P2_U3071) );
  INV_X1 U22272 ( .A(n19304), .ZN(n19306) );
  INV_X1 U22273 ( .A(n19371), .ZN(n19305) );
  NAND2_X1 U22274 ( .A1(n19306), .A2(n19305), .ZN(n19551) );
  OR2_X1 U22275 ( .A1(n19551), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19312) );
  OAI21_X1 U22276 ( .B1(n19330), .B2(n19360), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19309) );
  INV_X1 U22277 ( .A(n19307), .ZN(n19310) );
  NOR3_X2 U22278 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19367), .ZN(n19328) );
  AOI211_X1 U22279 ( .C1(n19310), .C2(n12070), .A(n19328), .B(n19799), .ZN(
        n19308) );
  OAI21_X1 U22280 ( .B1(n19310), .B2(n19328), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19311) );
  OAI21_X1 U22281 ( .B1(n19312), .B2(n19552), .A(n19311), .ZN(n19329) );
  AOI22_X1 U22282 ( .A1(n19329), .A2(n19653), .B1(n19652), .B2(n19328), .ZN(
        n19314) );
  AOI22_X1 U22283 ( .A1(n19360), .A2(n19662), .B1(n19330), .B2(n19605), .ZN(
        n19313) );
  OAI211_X1 U22284 ( .C1(n19334), .C2(n19315), .A(n19314), .B(n19313), .ZN(
        P2_U3080) );
  AOI22_X1 U22285 ( .A1(n19329), .A2(n19667), .B1(n19666), .B2(n19328), .ZN(
        n19317) );
  AOI22_X1 U22286 ( .A1(n19360), .A2(n19668), .B1(n19330), .B2(n19615), .ZN(
        n19316) );
  OAI211_X1 U22287 ( .C1(n19334), .C2(n13270), .A(n19317), .B(n19316), .ZN(
        P2_U3081) );
  AOI22_X1 U22288 ( .A1(n19329), .A2(n19673), .B1(n19672), .B2(n19328), .ZN(
        n19319) );
  AOI22_X1 U22289 ( .A1(n19360), .A2(n19674), .B1(n19330), .B2(n19619), .ZN(
        n19318) );
  OAI211_X1 U22290 ( .C1(n19334), .C2(n13293), .A(n19319), .B(n19318), .ZN(
        P2_U3082) );
  AOI22_X1 U22291 ( .A1(n19329), .A2(n19679), .B1(n19678), .B2(n19328), .ZN(
        n19321) );
  AOI22_X1 U22292 ( .A1(n19360), .A2(n19680), .B1(n19330), .B2(n19623), .ZN(
        n19320) );
  OAI211_X1 U22293 ( .C1(n19334), .C2(n13320), .A(n19321), .B(n19320), .ZN(
        P2_U3083) );
  AOI22_X1 U22294 ( .A1(n19329), .A2(n19685), .B1(n19684), .B2(n19328), .ZN(
        n19323) );
  AOI22_X1 U22295 ( .A1(n19360), .A2(n19686), .B1(n19330), .B2(n19627), .ZN(
        n19322) );
  OAI211_X1 U22296 ( .C1(n19334), .C2(n13346), .A(n19323), .B(n19322), .ZN(
        P2_U3084) );
  AOI22_X1 U22297 ( .A1(n19329), .A2(n19691), .B1(n19690), .B2(n19328), .ZN(
        n19325) );
  AOI22_X1 U22298 ( .A1(n19360), .A2(n19692), .B1(n19330), .B2(n19631), .ZN(
        n19324) );
  OAI211_X1 U22299 ( .C1(n19334), .C2(n13369), .A(n19325), .B(n19324), .ZN(
        P2_U3085) );
  AOI22_X1 U22300 ( .A1(n19329), .A2(n19697), .B1(n19696), .B2(n19328), .ZN(
        n19327) );
  AOI22_X1 U22301 ( .A1(n19360), .A2(n19698), .B1(n19330), .B2(n19635), .ZN(
        n19326) );
  OAI211_X1 U22302 ( .C1(n19334), .C2(n11512), .A(n19327), .B(n19326), .ZN(
        P2_U3086) );
  AOI22_X1 U22303 ( .A1(n19329), .A2(n19704), .B1(n19703), .B2(n19328), .ZN(
        n19332) );
  AOI22_X1 U22304 ( .A1(n19360), .A2(n19706), .B1(n19330), .B2(n19641), .ZN(
        n19331) );
  OAI211_X1 U22305 ( .C1(n19334), .C2(n19333), .A(n19332), .B(n19331), .ZN(
        P2_U3087) );
  INV_X1 U22306 ( .A(n19399), .ZN(n19336) );
  INV_X1 U22307 ( .A(n19338), .ZN(n19335) );
  AOI21_X1 U22308 ( .B1(n19336), .B2(n19335), .A(n19552), .ZN(n19339) );
  NOR2_X1 U22309 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19367), .ZN(
        n19343) );
  NOR2_X1 U22310 ( .A1(n19367), .A2(n19461), .ZN(n19359) );
  INV_X1 U22311 ( .A(n19359), .ZN(n19340) );
  AOI21_X1 U22312 ( .B1(n19341), .B2(n19340), .A(n16425), .ZN(n19337) );
  AOI22_X1 U22313 ( .A1(n19662), .A2(n19369), .B1(n19652), .B2(n19359), .ZN(
        n19346) );
  INV_X1 U22314 ( .A(n19339), .ZN(n19344) );
  OAI211_X1 U22315 ( .C1(n19341), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19340), 
        .B(n19552), .ZN(n19342) );
  OAI211_X1 U22316 ( .C1(n19344), .C2(n19343), .A(n19655), .B(n19342), .ZN(
        n19361) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19605), .ZN(n19345) );
  OAI211_X1 U22318 ( .C1(n19364), .C2(n19614), .A(n19346), .B(n19345), .ZN(
        P2_U3088) );
  AOI22_X1 U22319 ( .A1(n19615), .A2(n19360), .B1(n19666), .B2(n19359), .ZN(
        n19348) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19361), .B1(
        n19369), .B2(n19668), .ZN(n19347) );
  OAI211_X1 U22321 ( .C1(n19364), .C2(n19618), .A(n19348), .B(n19347), .ZN(
        P2_U3089) );
  AOI22_X1 U22322 ( .A1(n19619), .A2(n19360), .B1(n19672), .B2(n19359), .ZN(
        n19350) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19361), .B1(
        n19369), .B2(n19674), .ZN(n19349) );
  OAI211_X1 U22324 ( .C1(n19364), .C2(n19622), .A(n19350), .B(n19349), .ZN(
        P2_U3090) );
  AOI22_X1 U22325 ( .A1(n19680), .A2(n19369), .B1(n19678), .B2(n19359), .ZN(
        n19352) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19623), .ZN(n19351) );
  OAI211_X1 U22327 ( .C1(n19364), .C2(n19626), .A(n19352), .B(n19351), .ZN(
        P2_U3091) );
  AOI22_X1 U22328 ( .A1(n19627), .A2(n19360), .B1(n19684), .B2(n19359), .ZN(
        n19354) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19361), .B1(
        n19369), .B2(n19686), .ZN(n19353) );
  OAI211_X1 U22330 ( .C1(n19364), .C2(n19630), .A(n19354), .B(n19353), .ZN(
        P2_U3092) );
  AOI22_X1 U22331 ( .A1(n19631), .A2(n19360), .B1(n19690), .B2(n19359), .ZN(
        n19356) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19361), .B1(
        n19369), .B2(n19692), .ZN(n19355) );
  OAI211_X1 U22333 ( .C1(n19364), .C2(n19634), .A(n19356), .B(n19355), .ZN(
        P2_U3093) );
  AOI22_X1 U22334 ( .A1(n19698), .A2(n19369), .B1(n19696), .B2(n19359), .ZN(
        n19358) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19635), .ZN(n19357) );
  OAI211_X1 U22336 ( .C1(n19364), .C2(n19638), .A(n19358), .B(n19357), .ZN(
        P2_U3094) );
  AOI22_X1 U22337 ( .A1(n19641), .A2(n19360), .B1(n19703), .B2(n19359), .ZN(
        n19363) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19361), .B1(
        n19369), .B2(n19706), .ZN(n19362) );
  OAI211_X1 U22339 ( .C1(n19364), .C2(n19646), .A(n19363), .B(n19362), .ZN(
        P2_U3095) );
  INV_X1 U22340 ( .A(n19365), .ZN(n19366) );
  NOR2_X1 U22341 ( .A1(n19367), .A2(n19494), .ZN(n19390) );
  NOR2_X1 U22342 ( .A1(n19366), .A2(n19390), .ZN(n19372) );
  OAI22_X1 U22343 ( .A1(n19372), .A2(n16425), .B1(n19367), .B2(n19497), .ZN(
        n19391) );
  AOI22_X1 U22344 ( .A1(n19391), .A2(n19653), .B1(n19652), .B2(n19390), .ZN(
        n19377) );
  OAI21_X1 U22345 ( .B1(n19369), .B2(n19396), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19374) );
  NAND2_X1 U22346 ( .A1(n19371), .A2(n19370), .ZN(n19373) );
  AOI22_X1 U22347 ( .A1(n19374), .A2(n19373), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19372), .ZN(n19375) );
  OAI211_X1 U22348 ( .C1(n19390), .C2(n12070), .A(n19375), .B(n19655), .ZN(
        n19392) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19662), .ZN(n19376) );
  OAI211_X1 U22350 ( .C1(n19665), .C2(n19395), .A(n19377), .B(n19376), .ZN(
        P2_U3096) );
  AOI22_X1 U22351 ( .A1(n19391), .A2(n19667), .B1(n19666), .B2(n19390), .ZN(
        n19379) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19668), .ZN(n19378) );
  OAI211_X1 U22353 ( .C1(n19671), .C2(n19395), .A(n19379), .B(n19378), .ZN(
        P2_U3097) );
  AOI22_X1 U22354 ( .A1(n19391), .A2(n19673), .B1(n19672), .B2(n19390), .ZN(
        n19381) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19674), .ZN(n19380) );
  OAI211_X1 U22356 ( .C1(n19677), .C2(n19395), .A(n19381), .B(n19380), .ZN(
        P2_U3098) );
  AOI22_X1 U22357 ( .A1(n19391), .A2(n19679), .B1(n19678), .B2(n19390), .ZN(
        n19383) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19680), .ZN(n19382) );
  OAI211_X1 U22359 ( .C1(n19683), .C2(n19395), .A(n19383), .B(n19382), .ZN(
        P2_U3099) );
  AOI22_X1 U22360 ( .A1(n19391), .A2(n19685), .B1(n19684), .B2(n19390), .ZN(
        n19385) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19686), .ZN(n19384) );
  OAI211_X1 U22362 ( .C1(n19689), .C2(n19395), .A(n19385), .B(n19384), .ZN(
        P2_U3100) );
  AOI22_X1 U22363 ( .A1(n19391), .A2(n19691), .B1(n19690), .B2(n19390), .ZN(
        n19387) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19692), .ZN(n19386) );
  OAI211_X1 U22365 ( .C1(n19695), .C2(n19395), .A(n19387), .B(n19386), .ZN(
        P2_U3101) );
  AOI22_X1 U22366 ( .A1(n19391), .A2(n19697), .B1(n19696), .B2(n19390), .ZN(
        n19389) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19698), .ZN(n19388) );
  OAI211_X1 U22368 ( .C1(n19701), .C2(n19395), .A(n19389), .B(n19388), .ZN(
        P2_U3102) );
  AOI22_X1 U22369 ( .A1(n19391), .A2(n19704), .B1(n19703), .B2(n19390), .ZN(
        n19394) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19392), .B1(
        n19396), .B2(n19706), .ZN(n19393) );
  OAI211_X1 U22371 ( .C1(n19712), .C2(n19395), .A(n19394), .B(n19393), .ZN(
        P2_U3103) );
  NOR2_X1 U22372 ( .A1(n19817), .A2(n19827), .ZN(n19602) );
  NAND2_X1 U22373 ( .A1(n19602), .A2(n19809), .ZN(n19400) );
  OR2_X1 U22374 ( .A1(n19400), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19398) );
  AOI21_X1 U22375 ( .B1(n16425), .B2(n19398), .A(n19403), .ZN(n19421) );
  INV_X1 U22376 ( .A(n19431), .ZN(n19434) );
  AOI22_X1 U22377 ( .A1(n19421), .A2(n19653), .B1(n19434), .B2(n19652), .ZN(
        n19408) );
  NOR2_X1 U22378 ( .A1(n19399), .A2(n19659), .ZN(n19798) );
  INV_X1 U22379 ( .A(n19400), .ZN(n19405) );
  AND2_X1 U22380 ( .A1(n19431), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19401) );
  OR2_X1 U22381 ( .A1(n19463), .A2(n19401), .ZN(n19402) );
  NOR2_X1 U22382 ( .A1(n19403), .A2(n19402), .ZN(n19404) );
  OAI21_X1 U22383 ( .B1(n19798), .B2(n19405), .A(n19404), .ZN(n19422) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19662), .ZN(n19407) );
  OAI211_X1 U22385 ( .C1(n19665), .C2(n19425), .A(n19408), .B(n19407), .ZN(
        P2_U3104) );
  AOI22_X1 U22386 ( .A1(n19421), .A2(n19667), .B1(n19434), .B2(n19666), .ZN(
        n19410) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19668), .ZN(n19409) );
  OAI211_X1 U22388 ( .C1(n19671), .C2(n19425), .A(n19410), .B(n19409), .ZN(
        P2_U3105) );
  AOI22_X1 U22389 ( .A1(n19421), .A2(n19673), .B1(n19434), .B2(n19672), .ZN(
        n19412) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19674), .ZN(n19411) );
  OAI211_X1 U22391 ( .C1(n19677), .C2(n19425), .A(n19412), .B(n19411), .ZN(
        P2_U3106) );
  AOI22_X1 U22392 ( .A1(n19421), .A2(n19679), .B1(n19434), .B2(n19678), .ZN(
        n19414) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19680), .ZN(n19413) );
  OAI211_X1 U22394 ( .C1(n19683), .C2(n19425), .A(n19414), .B(n19413), .ZN(
        P2_U3107) );
  AOI22_X1 U22395 ( .A1(n19421), .A2(n19685), .B1(n19434), .B2(n19684), .ZN(
        n19416) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19686), .ZN(n19415) );
  OAI211_X1 U22397 ( .C1(n19689), .C2(n19425), .A(n19416), .B(n19415), .ZN(
        P2_U3108) );
  AOI22_X1 U22398 ( .A1(n19421), .A2(n19691), .B1(n19434), .B2(n19690), .ZN(
        n19418) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19692), .ZN(n19417) );
  OAI211_X1 U22400 ( .C1(n19695), .C2(n19425), .A(n19418), .B(n19417), .ZN(
        P2_U3109) );
  AOI22_X1 U22401 ( .A1(n19421), .A2(n19697), .B1(n19434), .B2(n19696), .ZN(
        n19420) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19698), .ZN(n19419) );
  OAI211_X1 U22403 ( .C1(n19701), .C2(n19425), .A(n19420), .B(n19419), .ZN(
        P2_U3110) );
  AOI22_X1 U22404 ( .A1(n19421), .A2(n19704), .B1(n19434), .B2(n19703), .ZN(
        n19424) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19422), .B1(
        n19426), .B2(n19706), .ZN(n19423) );
  OAI211_X1 U22406 ( .C1(n19712), .C2(n19425), .A(n19424), .B(n19423), .ZN(
        P2_U3111) );
  NAND2_X1 U22407 ( .A1(n19427), .A2(n19827), .ZN(n19467) );
  NOR2_X1 U22408 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19467), .ZN(
        n19452) );
  AOI22_X1 U22409 ( .A1(n19662), .A2(n19489), .B1(n19652), .B2(n19452), .ZN(
        n19439) );
  NAND2_X1 U22410 ( .A1(n19799), .A2(n19457), .ZN(n19429) );
  INV_X1 U22411 ( .A(n19428), .ZN(n19600) );
  OAI21_X1 U22412 ( .B1(n19489), .B2(n19429), .A(n19600), .ZN(n19433) );
  INV_X1 U22413 ( .A(n11478), .ZN(n19435) );
  AOI21_X1 U22414 ( .B1(n19435), .B2(n12070), .A(n19799), .ZN(n19430) );
  AOI21_X1 U22415 ( .B1(n19433), .B2(n19431), .A(n19430), .ZN(n19432) );
  OAI21_X1 U22416 ( .B1(n19434), .B2(n19452), .A(n19433), .ZN(n19437) );
  OAI21_X1 U22417 ( .B1(n19435), .B2(n19452), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19436) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19454), .B1(
        n19653), .B2(n19453), .ZN(n19438) );
  OAI211_X1 U22419 ( .C1(n19665), .C2(n19457), .A(n19439), .B(n19438), .ZN(
        P2_U3112) );
  AOI22_X1 U22420 ( .A1(n19668), .A2(n19489), .B1(n19666), .B2(n19452), .ZN(
        n19441) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19454), .B1(
        n19667), .B2(n19453), .ZN(n19440) );
  OAI211_X1 U22422 ( .C1(n19671), .C2(n19457), .A(n19441), .B(n19440), .ZN(
        P2_U3113) );
  AOI22_X1 U22423 ( .A1(n19674), .A2(n19489), .B1(n19672), .B2(n19452), .ZN(
        n19443) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19454), .B1(
        n19673), .B2(n19453), .ZN(n19442) );
  OAI211_X1 U22425 ( .C1(n19677), .C2(n19457), .A(n19443), .B(n19442), .ZN(
        P2_U3114) );
  AOI22_X1 U22426 ( .A1(n19680), .A2(n19489), .B1(n19678), .B2(n19452), .ZN(
        n19445) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19454), .B1(
        n19679), .B2(n19453), .ZN(n19444) );
  OAI211_X1 U22428 ( .C1(n19683), .C2(n19457), .A(n19445), .B(n19444), .ZN(
        P2_U3115) );
  AOI22_X1 U22429 ( .A1(n19686), .A2(n19489), .B1(n19684), .B2(n19452), .ZN(
        n19447) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19454), .B1(
        n19685), .B2(n19453), .ZN(n19446) );
  OAI211_X1 U22431 ( .C1(n19689), .C2(n19457), .A(n19447), .B(n19446), .ZN(
        P2_U3116) );
  AOI22_X1 U22432 ( .A1(n19692), .A2(n19489), .B1(n19690), .B2(n19452), .ZN(
        n19449) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19454), .B1(
        n19691), .B2(n19453), .ZN(n19448) );
  OAI211_X1 U22434 ( .C1(n19695), .C2(n19457), .A(n19449), .B(n19448), .ZN(
        P2_U3117) );
  AOI22_X1 U22435 ( .A1(n19698), .A2(n19489), .B1(n19696), .B2(n19452), .ZN(
        n19451) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19454), .B1(
        n19697), .B2(n19453), .ZN(n19450) );
  OAI211_X1 U22437 ( .C1(n19701), .C2(n19457), .A(n19451), .B(n19450), .ZN(
        P2_U3118) );
  AOI22_X1 U22438 ( .A1(n19706), .A2(n19489), .B1(n19703), .B2(n19452), .ZN(
        n19456) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19454), .B1(
        n19704), .B2(n19453), .ZN(n19455) );
  OAI211_X1 U22440 ( .C1(n19712), .C2(n19457), .A(n19456), .B(n19455), .ZN(
        P2_U3119) );
  INV_X1 U22441 ( .A(n19469), .ZN(n19458) );
  AOI21_X1 U22442 ( .B1(n19459), .B2(n19458), .A(n19552), .ZN(n19464) );
  INV_X1 U22443 ( .A(n19460), .ZN(n19465) );
  NOR2_X1 U22444 ( .A1(n19461), .A2(n19498), .ZN(n19499) );
  AOI211_X1 U22445 ( .C1(n19465), .C2(n12070), .A(n19499), .B(n19799), .ZN(
        n19462) );
  INV_X1 U22446 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19473) );
  AOI22_X1 U22447 ( .A1(n19605), .A2(n19489), .B1(n19652), .B2(n19499), .ZN(
        n19472) );
  INV_X1 U22448 ( .A(n19464), .ZN(n19468) );
  OAI21_X1 U22449 ( .B1(n19465), .B2(n19499), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19466) );
  AOI22_X1 U22450 ( .A1(n19653), .A2(n19488), .B1(n19500), .B2(n19662), .ZN(
        n19471) );
  OAI211_X1 U22451 ( .C1(n19493), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P2_U3120) );
  AOI22_X1 U22452 ( .A1(n19668), .A2(n19500), .B1(n19666), .B2(n19499), .ZN(
        n19475) );
  AOI22_X1 U22453 ( .A1(n19489), .A2(n19615), .B1(n19667), .B2(n19488), .ZN(
        n19474) );
  OAI211_X1 U22454 ( .C1(n19493), .C2(n12343), .A(n19475), .B(n19474), .ZN(
        P2_U3121) );
  INV_X1 U22455 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n19478) );
  AOI22_X1 U22456 ( .A1(n19674), .A2(n19500), .B1(n19672), .B2(n19499), .ZN(
        n19477) );
  AOI22_X1 U22457 ( .A1(n19489), .A2(n19619), .B1(n19673), .B2(n19488), .ZN(
        n19476) );
  OAI211_X1 U22458 ( .C1(n19493), .C2(n19478), .A(n19477), .B(n19476), .ZN(
        P2_U3122) );
  AOI22_X1 U22459 ( .A1(n19623), .A2(n19489), .B1(n19678), .B2(n19499), .ZN(
        n19480) );
  AOI22_X1 U22460 ( .A1(n19679), .A2(n19488), .B1(n19500), .B2(n19680), .ZN(
        n19479) );
  OAI211_X1 U22461 ( .C1(n19493), .C2(n13158), .A(n19480), .B(n19479), .ZN(
        P2_U3123) );
  AOI22_X1 U22462 ( .A1(n19627), .A2(n19489), .B1(n19684), .B2(n19499), .ZN(
        n19482) );
  AOI22_X1 U22463 ( .A1(n19685), .A2(n19488), .B1(n19500), .B2(n19686), .ZN(
        n19481) );
  OAI211_X1 U22464 ( .C1(n19493), .C2(n19483), .A(n19482), .B(n19481), .ZN(
        P2_U3124) );
  AOI22_X1 U22465 ( .A1(n19631), .A2(n19489), .B1(n19690), .B2(n19499), .ZN(
        n19485) );
  AOI22_X1 U22466 ( .A1(n19691), .A2(n19488), .B1(n19500), .B2(n19692), .ZN(
        n19484) );
  OAI211_X1 U22467 ( .C1(n19493), .C2(n12739), .A(n19485), .B(n19484), .ZN(
        P2_U3125) );
  AOI22_X1 U22468 ( .A1(n19698), .A2(n19500), .B1(n19696), .B2(n19499), .ZN(
        n19487) );
  AOI22_X1 U22469 ( .A1(n19489), .A2(n19635), .B1(n19697), .B2(n19488), .ZN(
        n19486) );
  OAI211_X1 U22470 ( .C1(n19493), .C2(n11519), .A(n19487), .B(n19486), .ZN(
        P2_U3126) );
  AOI22_X1 U22471 ( .A1(n19706), .A2(n19500), .B1(n19703), .B2(n19499), .ZN(
        n19491) );
  AOI22_X1 U22472 ( .A1(n19489), .A2(n19641), .B1(n19704), .B2(n19488), .ZN(
        n19490) );
  OAI211_X1 U22473 ( .C1(n19493), .C2(n19492), .A(n19491), .B(n19490), .ZN(
        P2_U3127) );
  INV_X1 U22474 ( .A(n19502), .ZN(n19495) );
  NOR2_X1 U22475 ( .A1(n19494), .A2(n19498), .ZN(n19518) );
  OAI21_X1 U22476 ( .B1(n19495), .B2(n19518), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19496) );
  OAI21_X1 U22477 ( .B1(n19498), .B2(n19497), .A(n19496), .ZN(n19519) );
  AOI22_X1 U22478 ( .A1(n19519), .A2(n19653), .B1(n19652), .B2(n19518), .ZN(
        n19505) );
  AOI221_X1 U22479 ( .B1(n19500), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19539), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19499), .ZN(n19501) );
  AOI211_X1 U22480 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19502), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19501), .ZN(n19503) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19662), .ZN(n19504) );
  OAI211_X1 U22482 ( .C1(n19665), .C2(n19523), .A(n19505), .B(n19504), .ZN(
        P2_U3128) );
  AOI22_X1 U22483 ( .A1(n19519), .A2(n19667), .B1(n19666), .B2(n19518), .ZN(
        n19507) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19668), .ZN(n19506) );
  OAI211_X1 U22485 ( .C1(n19671), .C2(n19523), .A(n19507), .B(n19506), .ZN(
        P2_U3129) );
  AOI22_X1 U22486 ( .A1(n19519), .A2(n19673), .B1(n19672), .B2(n19518), .ZN(
        n19509) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19674), .ZN(n19508) );
  OAI211_X1 U22488 ( .C1(n19677), .C2(n19523), .A(n19509), .B(n19508), .ZN(
        P2_U3130) );
  AOI22_X1 U22489 ( .A1(n19519), .A2(n19679), .B1(n19678), .B2(n19518), .ZN(
        n19511) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19680), .ZN(n19510) );
  OAI211_X1 U22491 ( .C1(n19683), .C2(n19523), .A(n19511), .B(n19510), .ZN(
        P2_U3131) );
  AOI22_X1 U22492 ( .A1(n19519), .A2(n19685), .B1(n19684), .B2(n19518), .ZN(
        n19513) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19686), .ZN(n19512) );
  OAI211_X1 U22494 ( .C1(n19689), .C2(n19523), .A(n19513), .B(n19512), .ZN(
        P2_U3132) );
  AOI22_X1 U22495 ( .A1(n19519), .A2(n19691), .B1(n19690), .B2(n19518), .ZN(
        n19515) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19692), .ZN(n19514) );
  OAI211_X1 U22497 ( .C1(n19695), .C2(n19523), .A(n19515), .B(n19514), .ZN(
        P2_U3133) );
  AOI22_X1 U22498 ( .A1(n19519), .A2(n19697), .B1(n19696), .B2(n19518), .ZN(
        n19517) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19698), .ZN(n19516) );
  OAI211_X1 U22500 ( .C1(n19701), .C2(n19523), .A(n19517), .B(n19516), .ZN(
        P2_U3134) );
  AOI22_X1 U22501 ( .A1(n19519), .A2(n19704), .B1(n19703), .B2(n19518), .ZN(
        n19522) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19520), .B1(
        n19539), .B2(n19706), .ZN(n19521) );
  OAI211_X1 U22503 ( .C1(n19712), .C2(n19523), .A(n19522), .B(n19521), .ZN(
        P2_U3135) );
  AOI22_X1 U22504 ( .A1(n19538), .A2(n19667), .B1(n19537), .B2(n19666), .ZN(
        n19525) );
  AOI22_X1 U22505 ( .A1(n19549), .A2(n19668), .B1(n19539), .B2(n19615), .ZN(
        n19524) );
  OAI211_X1 U22506 ( .C1(n19543), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        P2_U3137) );
  AOI22_X1 U22507 ( .A1(n19538), .A2(n19673), .B1(n19537), .B2(n19672), .ZN(
        n19528) );
  AOI22_X1 U22508 ( .A1(n19549), .A2(n19674), .B1(n19539), .B2(n19619), .ZN(
        n19527) );
  OAI211_X1 U22509 ( .C1(n19543), .C2(n20775), .A(n19528), .B(n19527), .ZN(
        P2_U3138) );
  AOI22_X1 U22510 ( .A1(n19538), .A2(n19679), .B1(n19537), .B2(n19678), .ZN(
        n19530) );
  AOI22_X1 U22511 ( .A1(n19549), .A2(n19680), .B1(n19539), .B2(n19623), .ZN(
        n19529) );
  OAI211_X1 U22512 ( .C1(n19543), .C2(n13327), .A(n19530), .B(n19529), .ZN(
        P2_U3139) );
  AOI22_X1 U22513 ( .A1(n19538), .A2(n19685), .B1(n19537), .B2(n19684), .ZN(
        n19532) );
  AOI22_X1 U22514 ( .A1(n19549), .A2(n19686), .B1(n19539), .B2(n19627), .ZN(
        n19531) );
  OAI211_X1 U22515 ( .C1(n19543), .C2(n13353), .A(n19532), .B(n19531), .ZN(
        P2_U3140) );
  AOI22_X1 U22516 ( .A1(n19538), .A2(n19691), .B1(n19537), .B2(n19690), .ZN(
        n19534) );
  AOI22_X1 U22517 ( .A1(n19549), .A2(n19692), .B1(n19539), .B2(n19631), .ZN(
        n19533) );
  OAI211_X1 U22518 ( .C1(n19543), .C2(n13376), .A(n19534), .B(n19533), .ZN(
        P2_U3141) );
  AOI22_X1 U22519 ( .A1(n19538), .A2(n19697), .B1(n19537), .B2(n19696), .ZN(
        n19536) );
  AOI22_X1 U22520 ( .A1(n19549), .A2(n19698), .B1(n19539), .B2(n19635), .ZN(
        n19535) );
  OAI211_X1 U22521 ( .C1(n19543), .C2(n13399), .A(n19536), .B(n19535), .ZN(
        P2_U3142) );
  AOI22_X1 U22522 ( .A1(n19538), .A2(n19704), .B1(n19537), .B2(n19703), .ZN(
        n19541) );
  AOI22_X1 U22523 ( .A1(n19549), .A2(n19706), .B1(n19539), .B2(n19641), .ZN(
        n19540) );
  OAI211_X1 U22524 ( .C1(n19543), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        P2_U3143) );
  INV_X1 U22525 ( .A(n19544), .ZN(n19548) );
  INV_X1 U22526 ( .A(n19554), .ZN(n19546) );
  NOR2_X1 U22527 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19545), .ZN(
        n19571) );
  OAI21_X1 U22528 ( .B1(n19546), .B2(n19571), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19547) );
  OAI21_X1 U22529 ( .B1(n19551), .B2(n19548), .A(n19547), .ZN(n19572) );
  AOI22_X1 U22530 ( .A1(n19572), .A2(n19653), .B1(n19652), .B2(n19571), .ZN(
        n19558) );
  OAI21_X1 U22531 ( .B1(n19549), .B2(n19593), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19550) );
  OAI21_X1 U22532 ( .B1(n19551), .B2(n19809), .A(n19550), .ZN(n19556) );
  INV_X1 U22533 ( .A(n19571), .ZN(n19553) );
  OAI211_X1 U22534 ( .C1(n19554), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19553), 
        .B(n19552), .ZN(n19555) );
  NAND3_X1 U22535 ( .A1(n19556), .A2(n19655), .A3(n19555), .ZN(n19573) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19662), .ZN(n19557) );
  OAI211_X1 U22537 ( .C1(n19665), .C2(n19576), .A(n19558), .B(n19557), .ZN(
        P2_U3144) );
  AOI22_X1 U22538 ( .A1(n19572), .A2(n19667), .B1(n19666), .B2(n19571), .ZN(
        n19560) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19668), .ZN(n19559) );
  OAI211_X1 U22540 ( .C1(n19671), .C2(n19576), .A(n19560), .B(n19559), .ZN(
        P2_U3145) );
  AOI22_X1 U22541 ( .A1(n19572), .A2(n19673), .B1(n19672), .B2(n19571), .ZN(
        n19562) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19674), .ZN(n19561) );
  OAI211_X1 U22543 ( .C1(n19677), .C2(n19576), .A(n19562), .B(n19561), .ZN(
        P2_U3146) );
  AOI22_X1 U22544 ( .A1(n19572), .A2(n19679), .B1(n19678), .B2(n19571), .ZN(
        n19564) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19680), .ZN(n19563) );
  OAI211_X1 U22546 ( .C1(n19683), .C2(n19576), .A(n19564), .B(n19563), .ZN(
        P2_U3147) );
  AOI22_X1 U22547 ( .A1(n19572), .A2(n19685), .B1(n19684), .B2(n19571), .ZN(
        n19566) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19686), .ZN(n19565) );
  OAI211_X1 U22549 ( .C1(n19689), .C2(n19576), .A(n19566), .B(n19565), .ZN(
        P2_U3148) );
  AOI22_X1 U22550 ( .A1(n19572), .A2(n19691), .B1(n19690), .B2(n19571), .ZN(
        n19568) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19692), .ZN(n19567) );
  OAI211_X1 U22552 ( .C1(n19695), .C2(n19576), .A(n19568), .B(n19567), .ZN(
        P2_U3149) );
  AOI22_X1 U22553 ( .A1(n19572), .A2(n19697), .B1(n19696), .B2(n19571), .ZN(
        n19570) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19698), .ZN(n19569) );
  OAI211_X1 U22555 ( .C1(n19701), .C2(n19576), .A(n19570), .B(n19569), .ZN(
        P2_U3150) );
  AOI22_X1 U22556 ( .A1(n19572), .A2(n19704), .B1(n19703), .B2(n19571), .ZN(
        n19575) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19573), .B1(
        n19593), .B2(n19706), .ZN(n19574) );
  OAI211_X1 U22558 ( .C1(n19712), .C2(n19576), .A(n19575), .B(n19574), .ZN(
        P2_U3151) );
  AOI22_X1 U22559 ( .A1(n19592), .A2(n19667), .B1(n19591), .B2(n19666), .ZN(
        n19578) );
  AOI22_X1 U22560 ( .A1(n19642), .A2(n19668), .B1(n19593), .B2(n19615), .ZN(
        n19577) );
  OAI211_X1 U22561 ( .C1(n19597), .C2(n11367), .A(n19578), .B(n19577), .ZN(
        P2_U3153) );
  INV_X1 U22562 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19581) );
  AOI22_X1 U22563 ( .A1(n19592), .A2(n19673), .B1(n19591), .B2(n19672), .ZN(
        n19580) );
  AOI22_X1 U22564 ( .A1(n19642), .A2(n19674), .B1(n19593), .B2(n19619), .ZN(
        n19579) );
  OAI211_X1 U22565 ( .C1(n19597), .C2(n19581), .A(n19580), .B(n19579), .ZN(
        P2_U3154) );
  AOI22_X1 U22566 ( .A1(n19592), .A2(n19679), .B1(n19591), .B2(n19678), .ZN(
        n19583) );
  AOI22_X1 U22567 ( .A1(n19642), .A2(n19680), .B1(n19593), .B2(n19623), .ZN(
        n19582) );
  OAI211_X1 U22568 ( .C1(n19597), .C2(n12601), .A(n19583), .B(n19582), .ZN(
        P2_U3155) );
  AOI22_X1 U22569 ( .A1(n19592), .A2(n19685), .B1(n19591), .B2(n19684), .ZN(
        n19585) );
  AOI22_X1 U22570 ( .A1(n19642), .A2(n19686), .B1(n19593), .B2(n19627), .ZN(
        n19584) );
  OAI211_X1 U22571 ( .C1(n19597), .C2(n13178), .A(n19585), .B(n19584), .ZN(
        P2_U3156) );
  INV_X1 U22572 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n19588) );
  AOI22_X1 U22573 ( .A1(n19592), .A2(n19691), .B1(n19591), .B2(n19690), .ZN(
        n19587) );
  AOI22_X1 U22574 ( .A1(n19642), .A2(n19692), .B1(n19593), .B2(n19631), .ZN(
        n19586) );
  OAI211_X1 U22575 ( .C1(n19597), .C2(n19588), .A(n19587), .B(n19586), .ZN(
        P2_U3157) );
  AOI22_X1 U22576 ( .A1(n19592), .A2(n19697), .B1(n19591), .B2(n19696), .ZN(
        n19590) );
  AOI22_X1 U22577 ( .A1(n19642), .A2(n19698), .B1(n19593), .B2(n19635), .ZN(
        n19589) );
  OAI211_X1 U22578 ( .C1(n19597), .C2(n11511), .A(n19590), .B(n19589), .ZN(
        P2_U3158) );
  INV_X1 U22579 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U22580 ( .A1(n19592), .A2(n19704), .B1(n19591), .B2(n19703), .ZN(
        n19595) );
  AOI22_X1 U22581 ( .A1(n19642), .A2(n19706), .B1(n19593), .B2(n19641), .ZN(
        n19594) );
  OAI211_X1 U22582 ( .C1(n19597), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3159) );
  NAND3_X1 U22583 ( .A1(n19711), .A2(n19599), .A3(n19799), .ZN(n19601) );
  NAND2_X1 U22584 ( .A1(n19601), .A2(n19600), .ZN(n19607) );
  NAND2_X1 U22585 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19602), .ZN(
        n19660) );
  NOR2_X1 U22586 ( .A1(n19660), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19639) );
  INV_X1 U22587 ( .A(n19639), .ZN(n19608) );
  NAND2_X1 U22588 ( .A1(n19608), .A2(n19606), .ZN(n19604) );
  AOI21_X1 U22589 ( .B1(n19609), .B2(n19608), .A(n16425), .ZN(n19603) );
  AOI22_X1 U22590 ( .A1(n19605), .A2(n19642), .B1(n19652), .B2(n19639), .ZN(
        n19613) );
  OAI221_X1 U22591 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19607), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19606), .A(n19608), .ZN(n19611) );
  NAND3_X1 U22592 ( .A1(n19609), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19608), 
        .ZN(n19610) );
  NAND3_X1 U22593 ( .A1(n19611), .A2(n19655), .A3(n19610), .ZN(n19643) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19643), .B1(
        n19640), .B2(n19662), .ZN(n19612) );
  OAI211_X1 U22595 ( .C1(n19647), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P2_U3160) );
  AOI22_X1 U22596 ( .A1(n19615), .A2(n19642), .B1(n19666), .B2(n19639), .ZN(
        n19617) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19643), .B1(
        n19640), .B2(n19668), .ZN(n19616) );
  OAI211_X1 U22598 ( .C1(n19647), .C2(n19618), .A(n19617), .B(n19616), .ZN(
        P2_U3161) );
  AOI22_X1 U22599 ( .A1(n19674), .A2(n19640), .B1(n19672), .B2(n19639), .ZN(
        n19621) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19643), .B1(
        n19642), .B2(n19619), .ZN(n19620) );
  OAI211_X1 U22601 ( .C1(n19647), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P2_U3162) );
  AOI22_X1 U22602 ( .A1(n19623), .A2(n19642), .B1(n19678), .B2(n19639), .ZN(
        n19625) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19643), .B1(
        n19640), .B2(n19680), .ZN(n19624) );
  OAI211_X1 U22604 ( .C1(n19647), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3163) );
  AOI22_X1 U22605 ( .A1(n19627), .A2(n19642), .B1(n19684), .B2(n19639), .ZN(
        n19629) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19643), .B1(
        n19640), .B2(n19686), .ZN(n19628) );
  OAI211_X1 U22607 ( .C1(n19647), .C2(n19630), .A(n19629), .B(n19628), .ZN(
        P2_U3164) );
  AOI22_X1 U22608 ( .A1(n19692), .A2(n19640), .B1(n19690), .B2(n19639), .ZN(
        n19633) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19643), .B1(
        n19642), .B2(n19631), .ZN(n19632) );
  OAI211_X1 U22610 ( .C1(n19647), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P2_U3165) );
  AOI22_X1 U22611 ( .A1(n19698), .A2(n19640), .B1(n19696), .B2(n19639), .ZN(
        n19637) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19643), .B1(
        n19642), .B2(n19635), .ZN(n19636) );
  OAI211_X1 U22613 ( .C1(n19647), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3166) );
  AOI22_X1 U22614 ( .A1(n19706), .A2(n19640), .B1(n19703), .B2(n19639), .ZN(
        n19645) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19643), .B1(
        n19642), .B2(n19641), .ZN(n19644) );
  OAI211_X1 U22616 ( .C1(n19647), .C2(n19646), .A(n19645), .B(n19644), .ZN(
        P2_U3167) );
  INV_X1 U22617 ( .A(n19648), .ZN(n19649) );
  NOR3_X1 U22618 ( .A1(n19649), .A2(n19702), .A3(n16425), .ZN(n19654) );
  INV_X1 U22619 ( .A(n19660), .ZN(n19650) );
  AOI21_X1 U22620 ( .B1(n19650), .B2(n12070), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19651) );
  NOR2_X1 U22621 ( .A1(n19654), .A2(n19651), .ZN(n19705) );
  AOI22_X1 U22622 ( .A1(n19705), .A2(n19653), .B1(n19652), .B2(n19702), .ZN(
        n19664) );
  INV_X1 U22623 ( .A(n19654), .ZN(n19656) );
  OAI211_X1 U22624 ( .C1(n19702), .C2(n12070), .A(n19656), .B(n19655), .ZN(
        n19657) );
  AOI221_X1 U22625 ( .B1(n19660), .B2(n19659), .C1(n19660), .C2(n19658), .A(
        n19657), .ZN(n19661) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19662), .ZN(n19663) );
  OAI211_X1 U22627 ( .C1(n19665), .C2(n19711), .A(n19664), .B(n19663), .ZN(
        P2_U3168) );
  AOI22_X1 U22628 ( .A1(n19705), .A2(n19667), .B1(n19666), .B2(n19702), .ZN(
        n19670) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19668), .ZN(n19669) );
  OAI211_X1 U22630 ( .C1(n19671), .C2(n19711), .A(n19670), .B(n19669), .ZN(
        P2_U3169) );
  AOI22_X1 U22631 ( .A1(n19705), .A2(n19673), .B1(n19672), .B2(n19702), .ZN(
        n19676) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19674), .ZN(n19675) );
  OAI211_X1 U22633 ( .C1(n19677), .C2(n19711), .A(n19676), .B(n19675), .ZN(
        P2_U3170) );
  AOI22_X1 U22634 ( .A1(n19705), .A2(n19679), .B1(n19678), .B2(n19702), .ZN(
        n19682) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19680), .ZN(n19681) );
  OAI211_X1 U22636 ( .C1(n19683), .C2(n19711), .A(n19682), .B(n19681), .ZN(
        P2_U3171) );
  AOI22_X1 U22637 ( .A1(n19705), .A2(n19685), .B1(n19684), .B2(n19702), .ZN(
        n19688) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19686), .ZN(n19687) );
  OAI211_X1 U22639 ( .C1(n19689), .C2(n19711), .A(n19688), .B(n19687), .ZN(
        P2_U3172) );
  AOI22_X1 U22640 ( .A1(n19705), .A2(n19691), .B1(n19690), .B2(n19702), .ZN(
        n19694) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19692), .ZN(n19693) );
  OAI211_X1 U22642 ( .C1(n19695), .C2(n19711), .A(n19694), .B(n19693), .ZN(
        P2_U3173) );
  AOI22_X1 U22643 ( .A1(n19705), .A2(n19697), .B1(n19696), .B2(n19702), .ZN(
        n19700) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19698), .ZN(n19699) );
  OAI211_X1 U22645 ( .C1(n19701), .C2(n19711), .A(n19700), .B(n19699), .ZN(
        P2_U3174) );
  AOI22_X1 U22646 ( .A1(n19705), .A2(n19704), .B1(n19703), .B2(n19702), .ZN(
        n19710) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19708), .B1(
        n19707), .B2(n19706), .ZN(n19709) );
  OAI211_X1 U22648 ( .C1(n19712), .C2(n19711), .A(n19710), .B(n19709), .ZN(
        P2_U3175) );
  OAI221_X1 U22649 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n12070), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n19714), .A(n19713), .ZN(n19718) );
  OAI211_X1 U22650 ( .C1(n19719), .C2(n19715), .A(n19733), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19716) );
  OAI211_X1 U22651 ( .C1(n19719), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3177) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19720), .ZN(
        P2_U3179) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19720), .ZN(
        P2_U3180) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19720), .ZN(
        P2_U3181) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19720), .ZN(
        P2_U3182) );
  AND2_X1 U22656 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19720), .ZN(
        P2_U3183) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19720), .ZN(
        P2_U3184) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19720), .ZN(
        P2_U3185) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19720), .ZN(
        P2_U3186) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19720), .ZN(
        P2_U3187) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19720), .ZN(
        P2_U3188) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19720), .ZN(
        P2_U3189) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19720), .ZN(
        P2_U3190) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19720), .ZN(
        P2_U3191) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19720), .ZN(
        P2_U3192) );
  INV_X1 U22666 ( .A(P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20856) );
  NOR2_X1 U22667 ( .A1(n20856), .A2(n19796), .ZN(P2_U3193) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19720), .ZN(
        P2_U3194) );
  AND2_X1 U22669 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19720), .ZN(
        P2_U3195) );
  AND2_X1 U22670 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19720), .ZN(
        P2_U3196) );
  AND2_X1 U22671 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19720), .ZN(
        P2_U3197) );
  AND2_X1 U22672 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19720), .ZN(
        P2_U3198) );
  AND2_X1 U22673 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19720), .ZN(
        P2_U3199) );
  AND2_X1 U22674 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19720), .ZN(
        P2_U3200) );
  AND2_X1 U22675 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19720), .ZN(P2_U3201) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19720), .ZN(P2_U3202) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19720), .ZN(P2_U3203) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19720), .ZN(P2_U3204) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19720), .ZN(P2_U3205) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19720), .ZN(P2_U3206) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19720), .ZN(P2_U3207) );
  AND2_X1 U22682 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19720), .ZN(P2_U3208) );
  INV_X1 U22683 ( .A(n19721), .ZN(n19736) );
  NAND2_X1 U22684 ( .A1(n19736), .A2(n19847), .ZN(n19724) );
  NAND2_X1 U22685 ( .A1(n19733), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19735) );
  NAND3_X1 U22686 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19735), .ZN(n19722) );
  NOR2_X1 U22687 ( .A1(n20664), .A2(n19727), .ZN(n19740) );
  AOI21_X1 U22688 ( .B1(n20815), .B2(n19722), .A(n19740), .ZN(n19723) );
  OAI221_X1 U22689 ( .B1(n19724), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19724), .C2(n19731), .A(n19723), .ZN(P2_U3209) );
  INV_X1 U22690 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19725) );
  AOI21_X1 U22691 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19731), .A(n20815), 
        .ZN(n19732) );
  NOR2_X1 U22692 ( .A1(n19725), .A2(n19732), .ZN(n19728) );
  AOI21_X1 U22693 ( .B1(n19728), .B2(n19727), .A(n19726), .ZN(n19729) );
  OAI211_X1 U22694 ( .C1(n19731), .C2(n19730), .A(n19729), .B(n19735), .ZN(
        P2_U3210) );
  AOI21_X1 U22695 ( .B1(n19734), .B2(n19733), .A(n19732), .ZN(n19739) );
  OAI22_X1 U22696 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19736), .B1(NA), 
        .B2(n19735), .ZN(n19737) );
  OAI211_X1 U22697 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19737), .ZN(n19738) );
  OAI21_X1 U22698 ( .B1(n19740), .B2(n19739), .A(n19738), .ZN(P2_U3211) );
  NAND2_X1 U22699 ( .A1(n19783), .A2(n20815), .ZN(n19789) );
  CLKBUF_X1 U22700 ( .A(n19789), .Z(n19786) );
  OAI222_X1 U22701 ( .A1(n19786), .A2(n19743), .B1(n19741), .B2(n19783), .C1(
        n12076), .C2(n19787), .ZN(P2_U3212) );
  OAI222_X1 U22702 ( .A1(n19787), .A2(n19743), .B1(n19742), .B2(n19783), .C1(
        n19745), .C2(n19786), .ZN(P2_U3213) );
  OAI222_X1 U22703 ( .A1(n19787), .A2(n19745), .B1(n19744), .B2(n19783), .C1(
        n19746), .C2(n19786), .ZN(P2_U3214) );
  OAI222_X1 U22704 ( .A1(n19789), .A2(n14531), .B1(n19747), .B2(n19783), .C1(
        n19746), .C2(n19787), .ZN(P2_U3215) );
  OAI222_X1 U22705 ( .A1(n19789), .A2(n11792), .B1(n19748), .B2(n19783), .C1(
        n14531), .C2(n19787), .ZN(P2_U3216) );
  OAI222_X1 U22706 ( .A1(n19789), .A2(n14518), .B1(n19749), .B2(n19783), .C1(
        n11792), .C2(n19787), .ZN(P2_U3217) );
  OAI222_X1 U22707 ( .A1(n19789), .A2(n15413), .B1(n19750), .B2(n19783), .C1(
        n14518), .C2(n19787), .ZN(P2_U3218) );
  OAI222_X1 U22708 ( .A1(n19789), .A2(n12551), .B1(n19751), .B2(n19783), .C1(
        n15413), .C2(n19787), .ZN(P2_U3219) );
  OAI222_X1 U22709 ( .A1(n19786), .A2(n12675), .B1(n19752), .B2(n19783), .C1(
        n12551), .C2(n19787), .ZN(P2_U3220) );
  OAI222_X1 U22710 ( .A1(n19786), .A2(n12678), .B1(n19753), .B2(n19783), .C1(
        n12675), .C2(n19787), .ZN(P2_U3221) );
  OAI222_X1 U22711 ( .A1(n19786), .A2(n19755), .B1(n19754), .B2(n19783), .C1(
        n12678), .C2(n19787), .ZN(P2_U3222) );
  OAI222_X1 U22712 ( .A1(n19786), .A2(n14499), .B1(n19756), .B2(n19783), .C1(
        n19755), .C2(n19787), .ZN(P2_U3223) );
  OAI222_X1 U22713 ( .A1(n19786), .A2(n12920), .B1(n19757), .B2(n19783), .C1(
        n14499), .C2(n19787), .ZN(P2_U3224) );
  OAI222_X1 U22714 ( .A1(n19786), .A2(n19759), .B1(n19758), .B2(n19783), .C1(
        n12920), .C2(n19787), .ZN(P2_U3225) );
  OAI222_X1 U22715 ( .A1(n19789), .A2(n19761), .B1(n19760), .B2(n19783), .C1(
        n19759), .C2(n19787), .ZN(P2_U3226) );
  OAI222_X1 U22716 ( .A1(n19789), .A2(n13444), .B1(n19762), .B2(n19783), .C1(
        n19761), .C2(n19787), .ZN(P2_U3227) );
  OAI222_X1 U22717 ( .A1(n19789), .A2(n19764), .B1(n19763), .B2(n19783), .C1(
        n13444), .C2(n19787), .ZN(P2_U3228) );
  OAI222_X1 U22718 ( .A1(n19789), .A2(n19766), .B1(n19765), .B2(n19783), .C1(
        n19764), .C2(n19787), .ZN(P2_U3229) );
  OAI222_X1 U22719 ( .A1(n19789), .A2(n19768), .B1(n19767), .B2(n19783), .C1(
        n19766), .C2(n19787), .ZN(P2_U3230) );
  OAI222_X1 U22720 ( .A1(n19789), .A2(n19770), .B1(n19769), .B2(n19783), .C1(
        n19768), .C2(n19787), .ZN(P2_U3231) );
  OAI222_X1 U22721 ( .A1(n19786), .A2(n19772), .B1(n19771), .B2(n19783), .C1(
        n19770), .C2(n19787), .ZN(P2_U3232) );
  OAI222_X1 U22722 ( .A1(n19786), .A2(n19773), .B1(n20846), .B2(n19783), .C1(
        n19772), .C2(n19787), .ZN(P2_U3233) );
  OAI222_X1 U22723 ( .A1(n19786), .A2(n19775), .B1(n19774), .B2(n19783), .C1(
        n19773), .C2(n19787), .ZN(P2_U3234) );
  OAI222_X1 U22724 ( .A1(n19786), .A2(n19777), .B1(n19776), .B2(n19783), .C1(
        n19775), .C2(n19787), .ZN(P2_U3235) );
  OAI222_X1 U22725 ( .A1(n19786), .A2(n19779), .B1(n19778), .B2(n19783), .C1(
        n19777), .C2(n19787), .ZN(P2_U3236) );
  OAI222_X1 U22726 ( .A1(n19786), .A2(n14961), .B1(n19780), .B2(n19783), .C1(
        n19779), .C2(n19787), .ZN(P2_U3237) );
  OAI222_X1 U22727 ( .A1(n19787), .A2(n14961), .B1(n19781), .B2(n19783), .C1(
        n19782), .C2(n19786), .ZN(P2_U3238) );
  OAI222_X1 U22728 ( .A1(n19786), .A2(n14940), .B1(n19784), .B2(n19783), .C1(
        n19782), .C2(n19787), .ZN(P2_U3239) );
  OAI222_X1 U22729 ( .A1(n19786), .A2(n13539), .B1(n19785), .B2(n19783), .C1(
        n14940), .C2(n19787), .ZN(P2_U3240) );
  OAI222_X1 U22730 ( .A1(n19789), .A2(n14917), .B1(n19788), .B2(n19783), .C1(
        n13539), .C2(n19787), .ZN(P2_U3241) );
  OAI22_X1 U22731 ( .A1(n19847), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19783), .ZN(n19790) );
  INV_X1 U22732 ( .A(n19790), .ZN(P2_U3585) );
  MUX2_X1 U22733 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19847), .Z(P2_U3586) );
  OAI22_X1 U22734 ( .A1(n19847), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19783), .ZN(n19791) );
  INV_X1 U22735 ( .A(n19791), .ZN(P2_U3587) );
  OAI22_X1 U22736 ( .A1(n19847), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19783), .ZN(n19792) );
  INV_X1 U22737 ( .A(n19792), .ZN(P2_U3588) );
  OAI21_X1 U22738 ( .B1(n19796), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19794), 
        .ZN(n19793) );
  INV_X1 U22739 ( .A(n19793), .ZN(P2_U3591) );
  OAI21_X1 U22740 ( .B1(n19796), .B2(n19795), .A(n19794), .ZN(P2_U3592) );
  INV_X1 U22741 ( .A(n19797), .ZN(n19806) );
  NAND2_X1 U22742 ( .A1(n19798), .A2(n19799), .ZN(n19805) );
  NAND2_X1 U22743 ( .A1(n19799), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19822) );
  NOR2_X1 U22744 ( .A1(n19800), .A2(n19822), .ZN(n19810) );
  NAND3_X1 U22745 ( .A1(n19823), .A2(n19801), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19802) );
  AND2_X1 U22746 ( .A1(n19802), .A2(n19818), .ZN(n19811) );
  OAI21_X1 U22747 ( .B1(n19810), .B2(n19811), .A(n19803), .ZN(n19804) );
  OAI211_X1 U22748 ( .C1(n19806), .C2(n12070), .A(n19805), .B(n19804), .ZN(
        n19807) );
  INV_X1 U22749 ( .A(n19807), .ZN(n19808) );
  AOI22_X1 U22750 ( .A1(n19834), .A2(n19809), .B1(n19808), .B2(n19835), .ZN(
        P2_U3602) );
  AOI21_X1 U22751 ( .B1(n19812), .B2(n19811), .A(n19810), .ZN(n19813) );
  INV_X1 U22752 ( .A(n19813), .ZN(n19814) );
  AOI21_X1 U22753 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19815), .A(n19814), 
        .ZN(n19816) );
  AOI22_X1 U22754 ( .A1(n19834), .A2(n19817), .B1(n19816), .B2(n19835), .ZN(
        P2_U3603) );
  INV_X1 U22755 ( .A(n19818), .ZN(n19830) );
  AND2_X1 U22756 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19819) );
  OR3_X1 U22757 ( .A1(n19820), .A2(n19830), .A3(n19819), .ZN(n19821) );
  OAI21_X1 U22758 ( .B1(n19823), .B2(n19822), .A(n19821), .ZN(n19824) );
  AOI21_X1 U22759 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19825), .A(n19824), 
        .ZN(n19826) );
  AOI22_X1 U22760 ( .A1(n19834), .A2(n19827), .B1(n19826), .B2(n19835), .ZN(
        P2_U3604) );
  NAND3_X1 U22761 ( .A1(n19828), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19829) );
  OAI21_X1 U22762 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(n19832) );
  AOI21_X1 U22763 ( .B1(n19836), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19832), 
        .ZN(n19833) );
  OAI22_X1 U22764 ( .A1(n19836), .A2(n19835), .B1(n19834), .B2(n19833), .ZN(
        P2_U3605) );
  INV_X1 U22765 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19837) );
  AOI22_X1 U22766 ( .A1(n19783), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19837), 
        .B2(n19847), .ZN(P2_U3608) );
  INV_X1 U22767 ( .A(n19838), .ZN(n19842) );
  NAND2_X1 U22768 ( .A1(n19840), .A2(n19839), .ZN(n19841) );
  OAI211_X1 U22769 ( .C1(n19844), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        n19846) );
  MUX2_X1 U22770 ( .A(P2_MORE_REG_SCAN_IN), .B(n19846), .S(n19845), .Z(
        P2_U3609) );
  MUX2_X1 U22771 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .B(P2_M_IO_N_REG_SCAN_IN), 
        .S(n19847), .Z(P2_U3611) );
  AOI21_X1 U22772 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20670), .A(n20668), 
        .ZN(n19854) );
  INV_X1 U22773 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19848) );
  NAND2_X1 U22774 ( .A1(n20668), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20736) );
  AOI21_X1 U22775 ( .B1(n19854), .B2(n19848), .A(n20738), .ZN(P1_U2802) );
  OAI21_X1 U22776 ( .B1(n19850), .B2(n19849), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19851) );
  OAI21_X1 U22777 ( .B1(n19852), .B2(n20650), .A(n19851), .ZN(P1_U2803) );
  NAND2_X1 U22778 ( .A1(n20670), .A2(n20668), .ZN(n20658) );
  INV_X1 U22779 ( .A(n20658), .ZN(n19855) );
  INV_X1 U22780 ( .A(n20738), .ZN(n20750) );
  OAI21_X1 U22781 ( .B1(n19855), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20750), .ZN(
        n19853) );
  OAI21_X1 U22782 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20736), .A(n19853), 
        .ZN(P1_U2804) );
  NOR2_X1 U22783 ( .A1(n20738), .A2(n19854), .ZN(n20721) );
  OAI21_X1 U22784 ( .B1(BS16), .B2(n19855), .A(n20721), .ZN(n20719) );
  OAI21_X1 U22785 ( .B1(n20721), .B2(n20542), .A(n20719), .ZN(P1_U2805) );
  AOI21_X1 U22786 ( .B1(n19856), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20029), .ZN(
        n19857) );
  INV_X1 U22787 ( .A(n19857), .ZN(P1_U2806) );
  NOR4_X1 U22788 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19861) );
  NOR4_X1 U22789 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19860) );
  NOR4_X1 U22790 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n19859) );
  NOR4_X1 U22791 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19858) );
  NAND4_X1 U22792 ( .A1(n19861), .A2(n19860), .A3(n19859), .A4(n19858), .ZN(
        n19867) );
  NOR4_X1 U22793 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19865) );
  AOI211_X1 U22794 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_16__SCAN_IN), .B(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19864) );
  NOR4_X1 U22795 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19863) );
  NOR4_X1 U22796 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19862) );
  NAND4_X1 U22797 ( .A1(n19865), .A2(n19864), .A3(n19863), .A4(n19862), .ZN(
        n19866) );
  NOR2_X1 U22798 ( .A1(n19867), .A2(n19866), .ZN(n20731) );
  INV_X1 U22799 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19869) );
  NOR3_X1 U22800 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19870) );
  OAI21_X1 U22801 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19870), .A(n20731), .ZN(
        n19868) );
  OAI21_X1 U22802 ( .B1(n20731), .B2(n19869), .A(n19868), .ZN(P1_U2807) );
  INV_X1 U22803 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20720) );
  AOI21_X1 U22804 ( .B1(n12396), .B2(n20720), .A(n19870), .ZN(n19872) );
  INV_X1 U22805 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19871) );
  INV_X1 U22806 ( .A(n20731), .ZN(n20734) );
  AOI22_X1 U22807 ( .A1(n20731), .A2(n19872), .B1(n19871), .B2(n20734), .ZN(
        P1_U2808) );
  AND2_X1 U22808 ( .A1(n19874), .A2(n19873), .ZN(n19883) );
  OAI22_X1 U22809 ( .A1(n19876), .A2(n19926), .B1(n19939), .B2(n19875), .ZN(
        n19877) );
  AOI211_X1 U22810 ( .C1(n19934), .C2(P1_EBX_REG_9__SCAN_IN), .A(n20021), .B(
        n19877), .ZN(n19882) );
  AOI22_X1 U22811 ( .A1(n19880), .A2(n19904), .B1(n19879), .B2(n19878), .ZN(
        n19881) );
  OAI211_X1 U22812 ( .C1(n19884), .C2(n19883), .A(n19882), .B(n19881), .ZN(
        P1_U2831) );
  NAND4_X1 U22813 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n19917), .A4(n19893), .ZN(n19885) );
  OAI211_X1 U22814 ( .C1(n19926), .C2(n19886), .A(n20068), .B(n19885), .ZN(
        n19887) );
  AOI21_X1 U22815 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n19934), .A(n19887), .ZN(
        n19899) );
  NAND2_X1 U22816 ( .A1(n19888), .A2(n19904), .ZN(n19895) );
  NAND2_X1 U22817 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19892) );
  OAI21_X1 U22818 ( .B1(n19891), .B2(n19890), .A(n19889), .ZN(n19943) );
  AOI21_X1 U22819 ( .B1(n19923), .B2(n19892), .A(n19943), .ZN(n19903) );
  OR2_X1 U22820 ( .A1(n19903), .A2(n19893), .ZN(n19894) );
  OAI211_X1 U22821 ( .C1(n19948), .C2(n19896), .A(n19895), .B(n19894), .ZN(
        n19897) );
  INV_X1 U22822 ( .A(n19897), .ZN(n19898) );
  OAI211_X1 U22823 ( .C1(n19939), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        P1_U2833) );
  AOI21_X1 U22824 ( .B1(n19901), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20021), .ZN(n19912) );
  INV_X1 U22825 ( .A(n19902), .ZN(n19949) );
  AOI22_X1 U22826 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n19934), .B1(n19914), .B2(
        n19949), .ZN(n19911) );
  OR2_X1 U22827 ( .A1(n19903), .A2(n16152), .ZN(n19906) );
  NAND2_X1 U22828 ( .A1(n19951), .A2(n19904), .ZN(n19905) );
  OAI211_X1 U22829 ( .C1(n19948), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        n19908) );
  INV_X1 U22830 ( .A(n19908), .ZN(n19910) );
  NAND3_X1 U22831 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19917), .A3(n16152), 
        .ZN(n19909) );
  NAND4_X1 U22832 ( .A1(n19912), .A2(n19911), .A3(n19910), .A4(n19909), .ZN(
        P1_U2834) );
  AOI22_X1 U22833 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19934), .B1(n19914), .B2(
        n19913), .ZN(n19915) );
  OAI211_X1 U22834 ( .C1(n19926), .C2(n20862), .A(n19915), .B(n20068), .ZN(
        n19916) );
  AOI221_X1 U22835 ( .B1(n19917), .B2(n16161), .C1(n19943), .C2(
        P1_REIP_REG_5__SCAN_IN), .A(n19916), .ZN(n19920) );
  NAND2_X1 U22836 ( .A1(n19918), .A2(n19942), .ZN(n19919) );
  OAI211_X1 U22837 ( .C1(n19948), .C2(n19921), .A(n19920), .B(n19919), .ZN(
        P1_U2835) );
  NAND2_X1 U22838 ( .A1(n19923), .A2(n19922), .ZN(n19924) );
  OAI22_X1 U22839 ( .A1(n19927), .A2(n19926), .B1(n19925), .B2(n19924), .ZN(
        n19941) );
  INV_X1 U22840 ( .A(n19928), .ZN(n19929) );
  OAI21_X1 U22841 ( .B1(n19931), .B2(n19930), .A(n19929), .ZN(n19933) );
  NAND2_X1 U22842 ( .A1(n19933), .A2(n19932), .ZN(n20034) );
  NAND2_X1 U22843 ( .A1(n19934), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n19938) );
  AOI21_X1 U22844 ( .B1(n19936), .B2(n19935), .A(n20021), .ZN(n19937) );
  OAI211_X1 U22845 ( .C1(n19939), .C2(n20034), .A(n19938), .B(n19937), .ZN(
        n19940) );
  NOR2_X1 U22846 ( .A1(n19941), .A2(n19940), .ZN(n19946) );
  NAND2_X1 U22847 ( .A1(n20027), .A2(n19942), .ZN(n19945) );
  NAND2_X1 U22848 ( .A1(n19943), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n19944) );
  AND3_X1 U22849 ( .A1(n19946), .A2(n19945), .A3(n19944), .ZN(n19947) );
  OAI21_X1 U22850 ( .B1(n20032), .B2(n19948), .A(n19947), .ZN(P1_U2836) );
  AOI22_X1 U22851 ( .A1(n19951), .A2(n19956), .B1(n19950), .B2(n19949), .ZN(
        n19952) );
  OAI21_X1 U22852 ( .B1(n13839), .B2(n19953), .A(n19952), .ZN(P1_U2866) );
  NOR2_X1 U22853 ( .A1(n19954), .A2(n20034), .ZN(n19955) );
  AOI21_X1 U22854 ( .B1(n20027), .B2(n19956), .A(n19955), .ZN(n19957) );
  OAI21_X1 U22855 ( .B1(n13839), .B2(n19958), .A(n19957), .ZN(P1_U2868) );
  AOI22_X1 U22856 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19960) );
  OAI21_X1 U22857 ( .B1(n12262), .B2(n19989), .A(n19960), .ZN(P1_U2921) );
  INV_X1 U22858 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19962) );
  AOI22_X1 U22859 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19961) );
  OAI21_X1 U22860 ( .B1(n19962), .B2(n19989), .A(n19961), .ZN(P1_U2922) );
  AOI22_X1 U22861 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U22862 ( .B1(n13918), .B2(n19989), .A(n19963), .ZN(P1_U2923) );
  INV_X1 U22863 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U22864 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19964) );
  OAI21_X1 U22865 ( .B1(n19965), .B2(n19989), .A(n19964), .ZN(P1_U2924) );
  INV_X1 U22866 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U22867 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19966) );
  OAI21_X1 U22868 ( .B1(n19967), .B2(n19989), .A(n19966), .ZN(P1_U2925) );
  INV_X1 U22869 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U22870 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19968) );
  OAI21_X1 U22871 ( .B1(n19969), .B2(n19989), .A(n19968), .ZN(P1_U2926) );
  INV_X1 U22872 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U22873 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19970) );
  OAI21_X1 U22874 ( .B1(n19971), .B2(n19989), .A(n19970), .ZN(P1_U2927) );
  INV_X1 U22875 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U22876 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20742), .B1(n19986), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19972) );
  OAI21_X1 U22877 ( .B1(n19973), .B2(n19989), .A(n19972), .ZN(P1_U2928) );
  INV_X1 U22878 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U22879 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19974) );
  OAI21_X1 U22880 ( .B1(n19975), .B2(n19989), .A(n19974), .ZN(P1_U2929) );
  AOI22_X1 U22881 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19976) );
  OAI21_X1 U22882 ( .B1(n10730), .B2(n19989), .A(n19976), .ZN(P1_U2930) );
  AOI22_X1 U22883 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22884 ( .B1(n10720), .B2(n19989), .A(n19977), .ZN(P1_U2931) );
  AOI22_X1 U22885 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19978) );
  OAI21_X1 U22886 ( .B1(n19979), .B2(n19989), .A(n19978), .ZN(P1_U2932) );
  AOI22_X1 U22887 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22888 ( .B1(n19981), .B2(n19989), .A(n19980), .ZN(P1_U2933) );
  AOI22_X1 U22889 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22890 ( .B1(n19983), .B2(n19989), .A(n19982), .ZN(P1_U2934) );
  AOI22_X1 U22891 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U22892 ( .B1(n19985), .B2(n19989), .A(n19984), .ZN(P1_U2935) );
  AOI22_X1 U22893 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19987), .B1(n19986), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19988) );
  OAI21_X1 U22894 ( .B1(n20848), .B2(n19989), .A(n19988), .ZN(P1_U2936) );
  AOI22_X1 U22895 ( .A1(n20018), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20017), .ZN(n19991) );
  NAND2_X1 U22896 ( .A1(n20003), .A2(n19990), .ZN(n20005) );
  NAND2_X1 U22897 ( .A1(n19991), .A2(n20005), .ZN(P1_U2945) );
  AOI22_X1 U22898 ( .A1(n20018), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n19993) );
  NAND2_X1 U22899 ( .A1(n20003), .A2(n19992), .ZN(n20007) );
  NAND2_X1 U22900 ( .A1(n19993), .A2(n20007), .ZN(P1_U2946) );
  AOI22_X1 U22901 ( .A1(n20018), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n19995) );
  NAND2_X1 U22902 ( .A1(n20003), .A2(n19994), .ZN(n20009) );
  NAND2_X1 U22903 ( .A1(n19995), .A2(n20009), .ZN(P1_U2947) );
  AOI22_X1 U22904 ( .A1(n20018), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n19997) );
  NAND2_X1 U22905 ( .A1(n20003), .A2(n19996), .ZN(n20011) );
  NAND2_X1 U22906 ( .A1(n19997), .A2(n20011), .ZN(P1_U2948) );
  AOI22_X1 U22907 ( .A1(n20018), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n19999) );
  NAND2_X1 U22908 ( .A1(n20003), .A2(n19998), .ZN(n20013) );
  NAND2_X1 U22909 ( .A1(n19999), .A2(n20013), .ZN(P1_U2949) );
  AOI22_X1 U22910 ( .A1(n20018), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U22911 ( .A1(n20003), .A2(n20000), .ZN(n20015) );
  NAND2_X1 U22912 ( .A1(n20001), .A2(n20015), .ZN(P1_U2950) );
  AOI22_X1 U22913 ( .A1(n20018), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20017), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20004) );
  NAND2_X1 U22914 ( .A1(n20003), .A2(n20002), .ZN(n20019) );
  NAND2_X1 U22915 ( .A1(n20004), .A2(n20019), .ZN(P1_U2951) );
  AOI22_X1 U22916 ( .A1(n20018), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20006) );
  NAND2_X1 U22917 ( .A1(n20006), .A2(n20005), .ZN(P1_U2960) );
  AOI22_X1 U22918 ( .A1(n20018), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20017), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20008) );
  NAND2_X1 U22919 ( .A1(n20008), .A2(n20007), .ZN(P1_U2961) );
  AOI22_X1 U22920 ( .A1(n20018), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20017), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20010) );
  NAND2_X1 U22921 ( .A1(n20010), .A2(n20009), .ZN(P1_U2962) );
  AOI22_X1 U22922 ( .A1(n20018), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20017), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U22923 ( .A1(n20012), .A2(n20011), .ZN(P1_U2963) );
  AOI22_X1 U22924 ( .A1(n20018), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20017), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20014) );
  NAND2_X1 U22925 ( .A1(n20014), .A2(n20013), .ZN(P1_U2964) );
  AOI22_X1 U22926 ( .A1(n20018), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20017), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20016) );
  NAND2_X1 U22927 ( .A1(n20016), .A2(n20015), .ZN(P1_U2965) );
  AOI22_X1 U22928 ( .A1(n20018), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20017), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20020) );
  NAND2_X1 U22929 ( .A1(n20020), .A2(n20019), .ZN(P1_U2966) );
  AOI22_X1 U22930 ( .A1(n20022), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20021), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U22931 ( .B1(n20025), .B2(n20024), .A(n20023), .ZN(n20026) );
  INV_X1 U22932 ( .A(n20026), .ZN(n20037) );
  AOI22_X1 U22933 ( .A1(n20037), .A2(n20029), .B1(n20028), .B2(n20027), .ZN(
        n20030) );
  OAI211_X1 U22934 ( .C1(n20033), .C2(n20032), .A(n20031), .B(n20030), .ZN(
        P1_U2995) );
  OAI22_X1 U22935 ( .A1(n20083), .A2(n20034), .B1(n20068), .B2(n20673), .ZN(
        n20035) );
  INV_X1 U22936 ( .A(n20035), .ZN(n20042) );
  OAI21_X1 U22937 ( .B1(n20050), .B2(n20073), .A(n20036), .ZN(n20046) );
  AOI22_X1 U22938 ( .A1(n20037), .A2(n20075), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20046), .ZN(n20041) );
  OAI211_X1 U22939 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20039), .B(n20038), .ZN(n20040) );
  NAND3_X1 U22940 ( .A1(n20042), .A2(n20041), .A3(n20040), .ZN(P1_U3027) );
  AOI21_X1 U22941 ( .B1(n20071), .B2(n20044), .A(n20043), .ZN(n20048) );
  AOI22_X1 U22942 ( .A1(n20046), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20045), .B2(n20075), .ZN(n20047) );
  OAI211_X1 U22943 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20049), .A(
        n20048), .B(n20047), .ZN(P1_U3028) );
  OAI21_X1 U22944 ( .B1(n20052), .B2(n20051), .A(n20050), .ZN(n20054) );
  AOI22_X1 U22945 ( .A1(n20055), .A2(n20054), .B1(n20071), .B2(n20053), .ZN(
        n20066) );
  NOR2_X1 U22946 ( .A1(n20078), .A2(n20056), .ZN(n20061) );
  AOI21_X1 U22947 ( .B1(n20078), .B2(n20058), .A(n20057), .ZN(n20059) );
  INV_X1 U22948 ( .A(n20059), .ZN(n20060) );
  MUX2_X1 U22949 ( .A(n20061), .B(n20060), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n20064) );
  AND3_X1 U22950 ( .A1(n12486), .A2(n20062), .A3(n20075), .ZN(n20063) );
  NOR2_X1 U22951 ( .A1(n20064), .A2(n20063), .ZN(n20065) );
  OAI211_X1 U22952 ( .C1(n20068), .C2(n20067), .A(n20066), .B(n20065), .ZN(
        P1_U3029) );
  AOI21_X1 U22953 ( .B1(n20071), .B2(n20070), .A(n20069), .ZN(n20081) );
  OAI21_X1 U22954 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20073), .A(
        n20072), .ZN(n20088) );
  AOI22_X1 U22955 ( .A1(n20088), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20075), .B2(n20074), .ZN(n20080) );
  NAND3_X1 U22956 ( .A1(n20078), .A2(n20077), .A3(n20076), .ZN(n20079) );
  NAND3_X1 U22957 ( .A1(n20081), .A2(n20080), .A3(n20079), .ZN(P1_U3030) );
  OAI22_X1 U22958 ( .A1(n20085), .A2(n20084), .B1(n20083), .B2(n20082), .ZN(
        n20086) );
  INV_X1 U22959 ( .A(n20086), .ZN(n20092) );
  OAI22_X1 U22960 ( .A1(n20089), .A2(n20088), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20087), .ZN(n20090) );
  NAND3_X1 U22961 ( .A1(n20092), .A2(n20091), .A3(n20090), .ZN(P1_U3031) );
  NOR2_X1 U22962 ( .A1(n20094), .A2(n20093), .ZN(P1_U3032) );
  NOR2_X2 U22963 ( .A1(n20098), .A2(n20097), .ZN(n20138) );
  AOI22_X1 U22964 ( .A1(DATAI_16_), .A2(n20096), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20138), .ZN(n20602) );
  NOR2_X2 U22965 ( .A1(n20137), .A2(n20101), .ZN(n20591) );
  NOR3_X1 U22966 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20151) );
  INV_X1 U22967 ( .A(n20151), .ZN(n20147) );
  NOR2_X1 U22968 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20147), .ZN(
        n20140) );
  NAND2_X1 U22969 ( .A1(n9587), .A2(n20507), .ZN(n20450) );
  AOI22_X1 U22970 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20138), .B1(DATAI_24_), 
        .B2(n20096), .ZN(n20554) );
  INV_X1 U22971 ( .A(n20554), .ZN(n20599) );
  AOI22_X1 U22972 ( .A1(n20591), .A2(n20140), .B1(n20139), .B2(n20599), .ZN(
        n20113) );
  OR2_X1 U22973 ( .A1(n20109), .A2(n10675), .ZN(n20538) );
  AND2_X1 U22974 ( .A1(n20538), .A2(n20239), .ZN(n20408) );
  NAND2_X1 U22975 ( .A1(n20167), .A2(n20647), .ZN(n20102) );
  AOI21_X1 U22976 ( .B1(n20102), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20587), 
        .ZN(n20108) );
  NAND2_X1 U22977 ( .A1(n20104), .A2(n20540), .ZN(n20110) );
  INV_X1 U22978 ( .A(n20350), .ZN(n20105) );
  NAND2_X1 U22979 ( .A1(n20105), .A2(n20406), .ZN(n20236) );
  AOI22_X1 U22980 ( .A1(n20108), .A2(n20110), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20236), .ZN(n20106) );
  OAI211_X1 U22981 ( .C1(n20140), .C2(n20355), .A(n20408), .B(n20106), .ZN(
        n20143) );
  NOR2_X2 U22982 ( .A1(n20107), .A2(n20148), .ZN(n20592) );
  INV_X1 U22983 ( .A(n20108), .ZN(n20111) );
  NAND2_X1 U22984 ( .A1(n20109), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20410) );
  AOI22_X1 U22985 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20143), .B1(
        n20592), .B2(n20142), .ZN(n20112) );
  OAI211_X1 U22986 ( .C1(n20602), .C2(n20167), .A(n20113), .B(n20112), .ZN(
        P1_U3033) );
  AOI22_X1 U22987 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20138), .B1(DATAI_17_), 
        .B2(n20096), .ZN(n20608) );
  NOR2_X2 U22988 ( .A1(n20137), .A2(n10345), .ZN(n20603) );
  AOI22_X1 U22989 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20138), .B1(DATAI_25_), 
        .B2(n20096), .ZN(n20558) );
  INV_X1 U22990 ( .A(n20558), .ZN(n20605) );
  AOI22_X1 U22991 ( .A1(n20603), .A2(n20140), .B1(n20139), .B2(n20605), .ZN(
        n20116) );
  NOR2_X2 U22992 ( .A1(n20114), .A2(n20148), .ZN(n20604) );
  AOI22_X1 U22993 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20143), .B1(
        n20604), .B2(n20142), .ZN(n20115) );
  OAI211_X1 U22994 ( .C1(n20608), .C2(n20167), .A(n20116), .B(n20115), .ZN(
        P1_U3034) );
  AOI22_X1 U22995 ( .A1(DATAI_18_), .A2(n20096), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20138), .ZN(n20614) );
  AOI22_X1 U22996 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20138), .B1(DATAI_26_), 
        .B2(n20096), .ZN(n20562) );
  INV_X1 U22997 ( .A(n20562), .ZN(n20611) );
  AOI22_X1 U22998 ( .A1(n9726), .A2(n20140), .B1(n20139), .B2(n20611), .ZN(
        n20119) );
  NOR2_X2 U22999 ( .A1(n20117), .A2(n20148), .ZN(n20610) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20143), .B1(
        n20610), .B2(n20142), .ZN(n20118) );
  OAI211_X1 U23001 ( .C1(n20614), .C2(n20167), .A(n20119), .B(n20118), .ZN(
        P1_U3035) );
  AOI22_X1 U23002 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20138), .B1(DATAI_19_), 
        .B2(n20096), .ZN(n20620) );
  NOR2_X2 U23003 ( .A1(n20137), .A2(n20120), .ZN(n20615) );
  AOI22_X1 U23004 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20138), .B1(DATAI_27_), 
        .B2(n20096), .ZN(n20566) );
  INV_X1 U23005 ( .A(n20566), .ZN(n20617) );
  AOI22_X1 U23006 ( .A1(n20615), .A2(n20140), .B1(n20139), .B2(n20617), .ZN(
        n20123) );
  NOR2_X2 U23007 ( .A1(n20121), .A2(n20148), .ZN(n20616) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20143), .B1(
        n20616), .B2(n20142), .ZN(n20122) );
  OAI211_X1 U23009 ( .C1(n20620), .C2(n20167), .A(n20123), .B(n20122), .ZN(
        P1_U3036) );
  AOI22_X1 U23010 ( .A1(DATAI_20_), .A2(n20096), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20138), .ZN(n20626) );
  NOR2_X2 U23011 ( .A1(n20137), .A2(n20124), .ZN(n20621) );
  AOI22_X1 U23012 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20138), .B1(DATAI_28_), 
        .B2(n20096), .ZN(n20570) );
  INV_X1 U23013 ( .A(n20570), .ZN(n20623) );
  AOI22_X1 U23014 ( .A1(n20621), .A2(n20140), .B1(n20139), .B2(n20623), .ZN(
        n20127) );
  NOR2_X2 U23015 ( .A1(n20125), .A2(n20148), .ZN(n20622) );
  AOI22_X1 U23016 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20143), .B1(
        n20622), .B2(n20142), .ZN(n20126) );
  OAI211_X1 U23017 ( .C1(n20626), .C2(n20167), .A(n20127), .B(n20126), .ZN(
        P1_U3037) );
  AOI22_X1 U23018 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20138), .B1(DATAI_21_), 
        .B2(n20096), .ZN(n20632) );
  NOR2_X2 U23019 ( .A1(n20137), .A2(n20128), .ZN(n20627) );
  AOI22_X1 U23020 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20138), .B1(DATAI_29_), 
        .B2(n20096), .ZN(n20574) );
  INV_X1 U23021 ( .A(n20574), .ZN(n20629) );
  AOI22_X1 U23022 ( .A1(n20627), .A2(n20140), .B1(n20139), .B2(n20629), .ZN(
        n20131) );
  NOR2_X2 U23023 ( .A1(n20129), .A2(n20148), .ZN(n20628) );
  AOI22_X1 U23024 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20143), .B1(
        n20628), .B2(n20142), .ZN(n20130) );
  OAI211_X1 U23025 ( .C1(n20632), .C2(n20167), .A(n20131), .B(n20130), .ZN(
        P1_U3038) );
  AOI22_X1 U23026 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20138), .B1(DATAI_22_), 
        .B2(n20096), .ZN(n20637) );
  AOI22_X1 U23027 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20138), .B1(DATAI_30_), 
        .B2(n20096), .ZN(n20578) );
  INV_X1 U23028 ( .A(n20578), .ZN(n20634) );
  AOI22_X1 U23029 ( .A1(n9684), .A2(n20140), .B1(n20139), .B2(n20634), .ZN(
        n20135) );
  NOR2_X2 U23030 ( .A1(n20133), .A2(n20148), .ZN(n20633) );
  AOI22_X1 U23031 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20143), .B1(
        n20633), .B2(n20142), .ZN(n20134) );
  OAI211_X1 U23032 ( .C1(n20637), .C2(n20167), .A(n20135), .B(n20134), .ZN(
        P1_U3039) );
  NOR2_X2 U23033 ( .A1(n20137), .A2(n20136), .ZN(n20638) );
  AOI22_X1 U23034 ( .A1(DATAI_31_), .A2(n20096), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20138), .ZN(n20586) );
  INV_X1 U23035 ( .A(n20586), .ZN(n20642) );
  AOI22_X1 U23036 ( .A1(n20638), .A2(n20140), .B1(n20139), .B2(n20642), .ZN(
        n20145) );
  NOR2_X2 U23037 ( .A1(n20141), .A2(n20148), .ZN(n20641) );
  AOI22_X1 U23038 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20143), .B1(
        n20641), .B2(n20142), .ZN(n20144) );
  OAI211_X1 U23039 ( .C1(n20648), .C2(n20167), .A(n20145), .B(n20144), .ZN(
        P1_U3040) );
  INV_X1 U23040 ( .A(n20511), .ZN(n20376) );
  NOR2_X1 U23041 ( .A1(n20509), .A2(n20147), .ZN(n20168) );
  AOI21_X1 U23042 ( .B1(n20104), .B2(n20376), .A(n20168), .ZN(n20149) );
  OAI22_X1 U23043 ( .A1(n20149), .A2(n20587), .B1(n20147), .B2(n10675), .ZN(
        n20169) );
  AOI22_X1 U23044 ( .A1(n20592), .A2(n20169), .B1(n20591), .B2(n20168), .ZN(
        n20153) );
  OAI211_X1 U23045 ( .C1(n20208), .C2(n20542), .A(n20510), .B(n20149), .ZN(
        n20150) );
  OAI211_X1 U23046 ( .C1(n20510), .C2(n20151), .A(n20597), .B(n20150), .ZN(
        n20171) );
  INV_X1 U23047 ( .A(n20167), .ZN(n20170) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20171), .B1(
        n20170), .B2(n20599), .ZN(n20152) );
  OAI211_X1 U23049 ( .C1(n20602), .C2(n20198), .A(n20153), .B(n20152), .ZN(
        P1_U3041) );
  AOI22_X1 U23050 ( .A1(n20604), .A2(n20169), .B1(n20603), .B2(n20168), .ZN(
        n20155) );
  INV_X1 U23051 ( .A(n20198), .ZN(n20164) );
  INV_X1 U23052 ( .A(n20608), .ZN(n20555) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20555), .ZN(n20154) );
  OAI211_X1 U23054 ( .C1(n20558), .C2(n20167), .A(n20155), .B(n20154), .ZN(
        P1_U3042) );
  AOI22_X1 U23055 ( .A1(n20610), .A2(n20169), .B1(n9726), .B2(n20168), .ZN(
        n20157) );
  INV_X1 U23056 ( .A(n20614), .ZN(n20559) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20559), .ZN(n20156) );
  OAI211_X1 U23058 ( .C1(n20562), .C2(n20167), .A(n20157), .B(n20156), .ZN(
        P1_U3043) );
  AOI22_X1 U23059 ( .A1(n20616), .A2(n20169), .B1(n20615), .B2(n20168), .ZN(
        n20159) );
  INV_X1 U23060 ( .A(n20620), .ZN(n20563) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20563), .ZN(n20158) );
  OAI211_X1 U23062 ( .C1(n20566), .C2(n20167), .A(n20159), .B(n20158), .ZN(
        P1_U3044) );
  AOI22_X1 U23063 ( .A1(n20622), .A2(n20169), .B1(n20621), .B2(n20168), .ZN(
        n20161) );
  INV_X1 U23064 ( .A(n20626), .ZN(n20567) );
  AOI22_X1 U23065 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20567), .ZN(n20160) );
  OAI211_X1 U23066 ( .C1(n20570), .C2(n20167), .A(n20161), .B(n20160), .ZN(
        P1_U3045) );
  AOI22_X1 U23067 ( .A1(n20628), .A2(n20169), .B1(n20627), .B2(n20168), .ZN(
        n20163) );
  INV_X1 U23068 ( .A(n20632), .ZN(n20571) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20571), .ZN(n20162) );
  OAI211_X1 U23070 ( .C1(n20574), .C2(n20167), .A(n20163), .B(n20162), .ZN(
        P1_U3046) );
  AOI22_X1 U23071 ( .A1(n20633), .A2(n20169), .B1(n9684), .B2(n20168), .ZN(
        n20166) );
  INV_X1 U23072 ( .A(n20637), .ZN(n20575) );
  AOI22_X1 U23073 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20171), .B1(
        n20164), .B2(n20575), .ZN(n20165) );
  OAI211_X1 U23074 ( .C1(n20578), .C2(n20167), .A(n20166), .B(n20165), .ZN(
        P1_U3047) );
  AOI22_X1 U23075 ( .A1(n20641), .A2(n20169), .B1(n20638), .B2(n20168), .ZN(
        n20173) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20171), .B1(
        n20170), .B2(n20642), .ZN(n20172) );
  OAI211_X1 U23077 ( .C1(n20648), .C2(n20198), .A(n20173), .B(n20172), .ZN(
        P1_U3048) );
  NAND2_X1 U23078 ( .A1(n9587), .A2(n10688), .ZN(n20541) );
  INV_X1 U23079 ( .A(n20541), .ZN(n20174) );
  INV_X1 U23080 ( .A(n20591), .ZN(n20403) );
  NAND3_X1 U23081 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20474), .A3(
        n10625), .ZN(n20211) );
  NOR2_X1 U23082 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20211), .ZN(
        n20194) );
  INV_X1 U23083 ( .A(n20194), .ZN(n20197) );
  OAI22_X1 U23084 ( .A1(n20198), .A2(n20554), .B1(n20403), .B2(n20197), .ZN(
        n20175) );
  INV_X1 U23085 ( .A(n20175), .ZN(n20183) );
  NAND3_X1 U23086 ( .A1(n20198), .A2(n20510), .A3(n20228), .ZN(n20176) );
  NAND2_X1 U23087 ( .A1(n20176), .A2(n20476), .ZN(n20178) );
  NAND2_X1 U23088 ( .A1(n20104), .A2(n20544), .ZN(n20180) );
  AOI22_X1 U23089 ( .A1(n20178), .A2(n20180), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20197), .ZN(n20177) );
  OAI21_X1 U23090 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20406), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20290) );
  NAND3_X1 U23091 ( .A1(n20408), .A2(n20177), .A3(n20290), .ZN(n20201) );
  INV_X1 U23092 ( .A(n20178), .ZN(n20181) );
  INV_X1 U23093 ( .A(n20406), .ZN(n20179) );
  NAND2_X1 U23094 ( .A1(n20179), .A2(n20474), .ZN(n20293) );
  OAI22_X1 U23095 ( .A1(n20181), .A2(n20180), .B1(n20410), .B2(n20293), .ZN(
        n20200) );
  AOI22_X1 U23096 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20201), .B1(
        n20592), .B2(n20200), .ZN(n20182) );
  OAI211_X1 U23097 ( .C1(n20602), .C2(n20228), .A(n20183), .B(n20182), .ZN(
        P1_U3049) );
  AOI22_X1 U23098 ( .A1(n20229), .A2(n20555), .B1(n20603), .B2(n20194), .ZN(
        n20185) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20201), .B1(
        n20604), .B2(n20200), .ZN(n20184) );
  OAI211_X1 U23100 ( .C1(n20558), .C2(n20198), .A(n20185), .B(n20184), .ZN(
        P1_U3050) );
  AOI22_X1 U23101 ( .A1(n20229), .A2(n20559), .B1(n9726), .B2(n20194), .ZN(
        n20187) );
  AOI22_X1 U23102 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20201), .B1(
        n20610), .B2(n20200), .ZN(n20186) );
  OAI211_X1 U23103 ( .C1(n20562), .C2(n20198), .A(n20187), .B(n20186), .ZN(
        P1_U3051) );
  AOI22_X1 U23104 ( .A1(n20229), .A2(n20563), .B1(n20194), .B2(n20615), .ZN(
        n20189) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20201), .B1(
        n20616), .B2(n20200), .ZN(n20188) );
  OAI211_X1 U23106 ( .C1(n20566), .C2(n20198), .A(n20189), .B(n20188), .ZN(
        P1_U3052) );
  AOI22_X1 U23107 ( .A1(n20229), .A2(n20567), .B1(n20194), .B2(n20621), .ZN(
        n20191) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20201), .B1(
        n20622), .B2(n20200), .ZN(n20190) );
  OAI211_X1 U23109 ( .C1(n20570), .C2(n20198), .A(n20191), .B(n20190), .ZN(
        P1_U3053) );
  AOI22_X1 U23110 ( .A1(n20229), .A2(n20571), .B1(n20194), .B2(n20627), .ZN(
        n20193) );
  AOI22_X1 U23111 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20201), .B1(
        n20628), .B2(n20200), .ZN(n20192) );
  OAI211_X1 U23112 ( .C1(n20574), .C2(n20198), .A(n20193), .B(n20192), .ZN(
        P1_U3054) );
  AOI22_X1 U23113 ( .A1(n20229), .A2(n20575), .B1(n20194), .B2(n9684), .ZN(
        n20196) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20201), .B1(
        n20633), .B2(n20200), .ZN(n20195) );
  OAI211_X1 U23115 ( .C1(n20578), .C2(n20198), .A(n20196), .B(n20195), .ZN(
        P1_U3055) );
  INV_X1 U23116 ( .A(n20638), .ZN(n20433) );
  OAI22_X1 U23117 ( .A1(n20198), .A2(n20586), .B1(n20433), .B2(n20197), .ZN(
        n20199) );
  INV_X1 U23118 ( .A(n20199), .ZN(n20203) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20201), .B1(
        n20641), .B2(n20200), .ZN(n20202) );
  OAI211_X1 U23120 ( .C1(n20648), .C2(n20228), .A(n20203), .B(n20202), .ZN(
        P1_U3056) );
  INV_X1 U23121 ( .A(n20450), .ZN(n20204) );
  AOI22_X1 U23122 ( .A1(n20229), .A2(n20599), .B1(n20591), .B2(n10228), .ZN(
        n20215) );
  NAND2_X1 U23123 ( .A1(n20207), .A2(n20206), .ZN(n20588) );
  INV_X1 U23124 ( .A(n20588), .ZN(n20441) );
  AOI21_X1 U23125 ( .B1(n20104), .B2(n20441), .A(n10228), .ZN(n20213) );
  AOI21_X1 U23126 ( .B1(n20208), .B2(n20510), .A(n20446), .ZN(n20212) );
  INV_X1 U23127 ( .A(n20212), .ZN(n20209) );
  AOI22_X1 U23128 ( .A1(n20213), .A2(n20209), .B1(n20587), .B2(n20211), .ZN(
        n20210) );
  NAND2_X1 U23129 ( .A1(n20597), .A2(n20210), .ZN(n20231) );
  OAI22_X1 U23130 ( .A1(n20213), .A2(n20212), .B1(n10675), .B2(n20211), .ZN(
        n20230) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20231), .B1(
        n20592), .B2(n20230), .ZN(n20214) );
  OAI211_X1 U23132 ( .C1(n20602), .C2(n20255), .A(n20215), .B(n20214), .ZN(
        P1_U3057) );
  INV_X1 U23133 ( .A(n20255), .ZN(n20258) );
  AOI22_X1 U23134 ( .A1(n20258), .A2(n20555), .B1(n20603), .B2(n10228), .ZN(
        n20217) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20231), .B1(
        n20604), .B2(n20230), .ZN(n20216) );
  OAI211_X1 U23136 ( .C1(n20558), .C2(n20228), .A(n20217), .B(n20216), .ZN(
        P1_U3058) );
  AOI22_X1 U23137 ( .A1(n20229), .A2(n20611), .B1(n9726), .B2(n10228), .ZN(
        n20219) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20231), .B1(
        n20610), .B2(n20230), .ZN(n20218) );
  OAI211_X1 U23139 ( .C1(n20614), .C2(n20255), .A(n20219), .B(n20218), .ZN(
        P1_U3059) );
  AOI22_X1 U23140 ( .A1(n20229), .A2(n20617), .B1(n20615), .B2(n10228), .ZN(
        n20221) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20231), .B1(
        n20616), .B2(n20230), .ZN(n20220) );
  OAI211_X1 U23142 ( .C1(n20620), .C2(n20255), .A(n20221), .B(n20220), .ZN(
        P1_U3060) );
  AOI22_X1 U23143 ( .A1(n20258), .A2(n20567), .B1(n20621), .B2(n10228), .ZN(
        n20223) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20231), .B1(
        n20622), .B2(n20230), .ZN(n20222) );
  OAI211_X1 U23145 ( .C1(n20570), .C2(n20228), .A(n20223), .B(n20222), .ZN(
        P1_U3061) );
  AOI22_X1 U23146 ( .A1(n20258), .A2(n20571), .B1(n20627), .B2(n10228), .ZN(
        n20225) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20231), .B1(
        n20628), .B2(n20230), .ZN(n20224) );
  OAI211_X1 U23148 ( .C1(n20574), .C2(n20228), .A(n20225), .B(n20224), .ZN(
        P1_U3062) );
  AOI22_X1 U23149 ( .A1(n20258), .A2(n20575), .B1(n9684), .B2(n10228), .ZN(
        n20227) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20231), .B1(
        n20633), .B2(n20230), .ZN(n20226) );
  OAI211_X1 U23151 ( .C1(n20578), .C2(n20228), .A(n20227), .B(n20226), .ZN(
        P1_U3063) );
  AOI22_X1 U23152 ( .A1(n20229), .A2(n20642), .B1(n20638), .B2(n10228), .ZN(
        n20233) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20231), .B1(
        n20641), .B2(n20230), .ZN(n20232) );
  OAI211_X1 U23154 ( .C1(n20648), .C2(n20255), .A(n20233), .B(n20232), .ZN(
        P1_U3064) );
  NOR2_X1 U23155 ( .A1(n20479), .A2(n20234), .ZN(n20318) );
  NAND3_X1 U23156 ( .A1(n20318), .A2(n20510), .A3(n20540), .ZN(n20235) );
  OAI21_X1 U23157 ( .B1(n20538), .B2(n20236), .A(n20235), .ZN(n20257) );
  NOR3_X1 U23158 ( .A1(n10625), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20266) );
  INV_X1 U23159 ( .A(n20266), .ZN(n20263) );
  NOR2_X1 U23160 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20263), .ZN(
        n20256) );
  AOI22_X1 U23161 ( .A1(n20592), .A2(n20257), .B1(n20591), .B2(n20256), .ZN(
        n20242) );
  AOI21_X1 U23162 ( .B1(n20255), .B2(n20287), .A(n20542), .ZN(n20237) );
  AOI21_X1 U23163 ( .B1(n20318), .B2(n20540), .A(n20237), .ZN(n20238) );
  NOR2_X1 U23164 ( .A1(n20238), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20240) );
  AND2_X1 U23165 ( .A1(n20410), .A2(n20239), .ZN(n20548) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20259), .B1(
        n20258), .B2(n20599), .ZN(n20241) );
  OAI211_X1 U23167 ( .C1(n20602), .C2(n20287), .A(n20242), .B(n20241), .ZN(
        P1_U3065) );
  AOI22_X1 U23168 ( .A1(n20604), .A2(n20257), .B1(n20603), .B2(n20256), .ZN(
        n20244) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20555), .ZN(n20243) );
  OAI211_X1 U23170 ( .C1(n20558), .C2(n20255), .A(n20244), .B(n20243), .ZN(
        P1_U3066) );
  AOI22_X1 U23171 ( .A1(n20610), .A2(n20257), .B1(n9726), .B2(n20256), .ZN(
        n20246) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20559), .ZN(n20245) );
  OAI211_X1 U23173 ( .C1(n20562), .C2(n20255), .A(n20246), .B(n20245), .ZN(
        P1_U3067) );
  AOI22_X1 U23174 ( .A1(n20616), .A2(n20257), .B1(n20615), .B2(n20256), .ZN(
        n20248) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20563), .ZN(n20247) );
  OAI211_X1 U23176 ( .C1(n20566), .C2(n20255), .A(n20248), .B(n20247), .ZN(
        P1_U3068) );
  AOI22_X1 U23177 ( .A1(n20622), .A2(n20257), .B1(n20621), .B2(n20256), .ZN(
        n20250) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20567), .ZN(n20249) );
  OAI211_X1 U23179 ( .C1(n20570), .C2(n20255), .A(n20250), .B(n20249), .ZN(
        P1_U3069) );
  AOI22_X1 U23180 ( .A1(n20628), .A2(n20257), .B1(n20627), .B2(n20256), .ZN(
        n20252) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20571), .ZN(n20251) );
  OAI211_X1 U23182 ( .C1(n20574), .C2(n20255), .A(n20252), .B(n20251), .ZN(
        P1_U3070) );
  AOI22_X1 U23183 ( .A1(n20633), .A2(n20257), .B1(n9684), .B2(n20256), .ZN(
        n20254) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20259), .B1(
        n20279), .B2(n20575), .ZN(n20253) );
  OAI211_X1 U23185 ( .C1(n20578), .C2(n20255), .A(n20254), .B(n20253), .ZN(
        P1_U3071) );
  AOI22_X1 U23186 ( .A1(n20641), .A2(n20257), .B1(n20638), .B2(n20256), .ZN(
        n20261) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20259), .B1(
        n20258), .B2(n20642), .ZN(n20260) );
  OAI211_X1 U23188 ( .C1(n20648), .C2(n20287), .A(n20261), .B(n20260), .ZN(
        P1_U3072) );
  NOR2_X1 U23189 ( .A1(n20509), .A2(n20263), .ZN(n20282) );
  AOI21_X1 U23190 ( .B1(n20318), .B2(n20376), .A(n20282), .ZN(n20264) );
  OAI22_X1 U23191 ( .A1(n20264), .A2(n20587), .B1(n20263), .B2(n10675), .ZN(
        n20283) );
  AOI22_X1 U23192 ( .A1(n20592), .A2(n20283), .B1(n20591), .B2(n20282), .ZN(
        n20268) );
  OAI211_X1 U23193 ( .C1(n20325), .C2(n20542), .A(n20510), .B(n20264), .ZN(
        n20265) );
  OAI211_X1 U23194 ( .C1(n20510), .C2(n20266), .A(n20597), .B(n20265), .ZN(
        n20284) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20284), .B1(
        n20279), .B2(n20599), .ZN(n20267) );
  OAI211_X1 U23196 ( .C1(n20602), .C2(n20298), .A(n20268), .B(n20267), .ZN(
        P1_U3073) );
  AOI22_X1 U23197 ( .A1(n20604), .A2(n20283), .B1(n20603), .B2(n20282), .ZN(
        n20270) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20555), .ZN(n20269) );
  OAI211_X1 U23199 ( .C1(n20558), .C2(n20287), .A(n20270), .B(n20269), .ZN(
        P1_U3074) );
  AOI22_X1 U23200 ( .A1(n20610), .A2(n20283), .B1(n9726), .B2(n20282), .ZN(
        n20272) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20559), .ZN(n20271) );
  OAI211_X1 U23202 ( .C1(n20562), .C2(n20287), .A(n20272), .B(n20271), .ZN(
        P1_U3075) );
  AOI22_X1 U23203 ( .A1(n20616), .A2(n20283), .B1(n20615), .B2(n20282), .ZN(
        n20274) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20563), .ZN(n20273) );
  OAI211_X1 U23205 ( .C1(n20566), .C2(n20287), .A(n20274), .B(n20273), .ZN(
        P1_U3076) );
  AOI22_X1 U23206 ( .A1(n20622), .A2(n20283), .B1(n20621), .B2(n20282), .ZN(
        n20276) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20284), .B1(
        n20279), .B2(n20623), .ZN(n20275) );
  OAI211_X1 U23208 ( .C1(n20626), .C2(n20298), .A(n20276), .B(n20275), .ZN(
        P1_U3077) );
  AOI22_X1 U23209 ( .A1(n20628), .A2(n20283), .B1(n20627), .B2(n20282), .ZN(
        n20278) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20284), .B1(
        n20279), .B2(n20629), .ZN(n20277) );
  OAI211_X1 U23211 ( .C1(n20632), .C2(n20298), .A(n20278), .B(n20277), .ZN(
        P1_U3078) );
  AOI22_X1 U23212 ( .A1(n20633), .A2(n20283), .B1(n9684), .B2(n20282), .ZN(
        n20281) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20284), .B1(
        n20279), .B2(n20634), .ZN(n20280) );
  OAI211_X1 U23214 ( .C1(n20637), .C2(n20298), .A(n20281), .B(n20280), .ZN(
        P1_U3079) );
  AOI22_X1 U23215 ( .A1(n20641), .A2(n20283), .B1(n20638), .B2(n20282), .ZN(
        n20286) );
  INV_X1 U23216 ( .A(n20648), .ZN(n20581) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20581), .ZN(n20285) );
  OAI211_X1 U23218 ( .C1(n20586), .C2(n20287), .A(n20286), .B(n20285), .ZN(
        P1_U3080) );
  NAND2_X1 U23219 ( .A1(n20509), .A2(n20324), .ZN(n20289) );
  INV_X1 U23220 ( .A(n20289), .ZN(n20311) );
  INV_X1 U23221 ( .A(n20336), .ZN(n20343) );
  INV_X1 U23222 ( .A(n20602), .ZN(n20551) );
  AOI22_X1 U23223 ( .A1(n20591), .A2(n20311), .B1(n20343), .B2(n20551), .ZN(
        n20297) );
  NAND2_X1 U23224 ( .A1(n20298), .A2(n20336), .ZN(n20288) );
  AOI21_X1 U23225 ( .B1(n20288), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20587), 
        .ZN(n20292) );
  NAND2_X1 U23226 ( .A1(n20318), .A2(n20544), .ZN(n20294) );
  AOI22_X1 U23227 ( .A1(n20292), .A2(n20294), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20289), .ZN(n20291) );
  NAND3_X1 U23228 ( .A1(n20548), .A2(n20291), .A3(n20290), .ZN(n20314) );
  INV_X1 U23229 ( .A(n20292), .ZN(n20295) );
  OAI22_X1 U23230 ( .A1(n20295), .A2(n20294), .B1(n20293), .B2(n20538), .ZN(
        n20313) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20314), .B1(
        n20592), .B2(n20313), .ZN(n20296) );
  OAI211_X1 U23232 ( .C1(n20554), .C2(n20298), .A(n20297), .B(n20296), .ZN(
        P1_U3081) );
  AOI22_X1 U23233 ( .A1(n20312), .A2(n20605), .B1(n20603), .B2(n20311), .ZN(
        n20300) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20314), .B1(
        n20604), .B2(n20313), .ZN(n20299) );
  OAI211_X1 U23235 ( .C1(n20608), .C2(n20336), .A(n20300), .B(n20299), .ZN(
        P1_U3082) );
  AOI22_X1 U23236 ( .A1(n20312), .A2(n20611), .B1(n9726), .B2(n20311), .ZN(
        n20302) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20314), .B1(
        n20610), .B2(n20313), .ZN(n20301) );
  OAI211_X1 U23238 ( .C1(n20614), .C2(n20336), .A(n20302), .B(n20301), .ZN(
        P1_U3083) );
  AOI22_X1 U23239 ( .A1(n20312), .A2(n20617), .B1(n20615), .B2(n20311), .ZN(
        n20304) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20314), .B1(
        n20616), .B2(n20313), .ZN(n20303) );
  OAI211_X1 U23241 ( .C1(n20620), .C2(n20336), .A(n20304), .B(n20303), .ZN(
        P1_U3084) );
  AOI22_X1 U23242 ( .A1(n20312), .A2(n20623), .B1(n20621), .B2(n20311), .ZN(
        n20306) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20314), .B1(
        n20622), .B2(n20313), .ZN(n20305) );
  OAI211_X1 U23244 ( .C1(n20626), .C2(n20336), .A(n20306), .B(n20305), .ZN(
        P1_U3085) );
  AOI22_X1 U23245 ( .A1(n20312), .A2(n20629), .B1(n20627), .B2(n20311), .ZN(
        n20308) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20314), .B1(
        n20628), .B2(n20313), .ZN(n20307) );
  OAI211_X1 U23247 ( .C1(n20632), .C2(n20336), .A(n20308), .B(n20307), .ZN(
        P1_U3086) );
  AOI22_X1 U23248 ( .A1(n20312), .A2(n20634), .B1(n9684), .B2(n20311), .ZN(
        n20310) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20314), .B1(
        n20633), .B2(n20313), .ZN(n20309) );
  OAI211_X1 U23250 ( .C1(n20637), .C2(n20336), .A(n20310), .B(n20309), .ZN(
        P1_U3087) );
  AOI22_X1 U23251 ( .A1(n20312), .A2(n20642), .B1(n20638), .B2(n20311), .ZN(
        n20316) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20314), .B1(
        n20641), .B2(n20313), .ZN(n20315) );
  OAI211_X1 U23253 ( .C1(n20648), .C2(n20336), .A(n20316), .B(n20315), .ZN(
        P1_U3088) );
  INV_X1 U23254 ( .A(n20317), .ZN(n20341) );
  AOI21_X1 U23255 ( .B1(n20318), .B2(n20441), .A(n20341), .ZN(n20321) );
  OAI22_X1 U23256 ( .A1(n20321), .A2(n20587), .B1(n20319), .B2(n10675), .ZN(
        n20342) );
  AOI22_X1 U23257 ( .A1(n20592), .A2(n20342), .B1(n20341), .B2(n20591), .ZN(
        n20327) );
  INV_X1 U23258 ( .A(n20325), .ZN(n20320) );
  NOR2_X1 U23259 ( .A1(n20320), .A2(n20587), .ZN(n20322) );
  OAI21_X1 U23260 ( .B1(n20322), .B2(n20446), .A(n20321), .ZN(n20323) );
  OAI211_X1 U23261 ( .C1(n20324), .C2(n20510), .A(n20597), .B(n20323), .ZN(
        n20344) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20344), .B1(
        n20372), .B2(n20551), .ZN(n20326) );
  OAI211_X1 U23263 ( .C1(n20554), .C2(n20336), .A(n20327), .B(n20326), .ZN(
        P1_U3089) );
  AOI22_X1 U23264 ( .A1(n20604), .A2(n20342), .B1(n20341), .B2(n20603), .ZN(
        n20329) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20344), .B1(
        n20343), .B2(n20605), .ZN(n20328) );
  OAI211_X1 U23266 ( .C1(n20608), .C2(n20347), .A(n20329), .B(n20328), .ZN(
        P1_U3090) );
  AOI22_X1 U23267 ( .A1(n20610), .A2(n20342), .B1(n20341), .B2(n9726), .ZN(
        n20331) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20344), .B1(
        n20372), .B2(n20559), .ZN(n20330) );
  OAI211_X1 U23269 ( .C1(n20562), .C2(n20336), .A(n20331), .B(n20330), .ZN(
        P1_U3091) );
  AOI22_X1 U23270 ( .A1(n20616), .A2(n20342), .B1(n20341), .B2(n20615), .ZN(
        n20333) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20344), .B1(
        n20372), .B2(n20563), .ZN(n20332) );
  OAI211_X1 U23272 ( .C1(n20566), .C2(n20336), .A(n20333), .B(n20332), .ZN(
        P1_U3092) );
  AOI22_X1 U23273 ( .A1(n20622), .A2(n20342), .B1(n20341), .B2(n20621), .ZN(
        n20335) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20344), .B1(
        n20372), .B2(n20567), .ZN(n20334) );
  OAI211_X1 U23275 ( .C1(n20570), .C2(n20336), .A(n20335), .B(n20334), .ZN(
        P1_U3093) );
  AOI22_X1 U23276 ( .A1(n20628), .A2(n20342), .B1(n20341), .B2(n20627), .ZN(
        n20338) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20344), .B1(
        n20343), .B2(n20629), .ZN(n20337) );
  OAI211_X1 U23278 ( .C1(n20632), .C2(n20347), .A(n20338), .B(n20337), .ZN(
        P1_U3094) );
  AOI22_X1 U23279 ( .A1(n20633), .A2(n20342), .B1(n20341), .B2(n9684), .ZN(
        n20340) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20344), .B1(
        n20343), .B2(n20634), .ZN(n20339) );
  OAI211_X1 U23281 ( .C1(n20637), .C2(n20347), .A(n20340), .B(n20339), .ZN(
        P1_U3095) );
  AOI22_X1 U23282 ( .A1(n20641), .A2(n20342), .B1(n20341), .B2(n20638), .ZN(
        n20346) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20344), .B1(
        n20343), .B2(n20642), .ZN(n20345) );
  OAI211_X1 U23284 ( .C1(n20648), .C2(n20347), .A(n20346), .B(n20345), .ZN(
        P1_U3096) );
  NOR3_X1 U23285 ( .A1(n20474), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20380) );
  INV_X1 U23286 ( .A(n20380), .ZN(n20377) );
  NOR2_X1 U23287 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20377), .ZN(
        n20370) );
  AOI21_X1 U23288 ( .B1(n20442), .B2(n20540), .A(n20370), .ZN(n20352) );
  NAND2_X1 U23289 ( .A1(n20350), .A2(n20406), .ZN(n20484) );
  OAI22_X1 U23290 ( .A1(n20352), .A2(n20587), .B1(n20410), .B2(n20484), .ZN(
        n20371) );
  AOI22_X1 U23291 ( .A1(n20592), .A2(n20371), .B1(n20591), .B2(n20370), .ZN(
        n20357) );
  INV_X1 U23292 ( .A(n20402), .ZN(n20351) );
  OAI21_X1 U23293 ( .B1(n20351), .B2(n20372), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20353) );
  NAND2_X1 U23294 ( .A1(n20353), .A2(n20352), .ZN(n20354) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20599), .ZN(n20356) );
  OAI211_X1 U23296 ( .C1(n20602), .C2(n20402), .A(n20357), .B(n20356), .ZN(
        P1_U3097) );
  AOI22_X1 U23297 ( .A1(n20604), .A2(n20371), .B1(n20603), .B2(n20370), .ZN(
        n20359) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20605), .ZN(n20358) );
  OAI211_X1 U23299 ( .C1(n20608), .C2(n20402), .A(n20359), .B(n20358), .ZN(
        P1_U3098) );
  AOI22_X1 U23300 ( .A1(n20610), .A2(n20371), .B1(n9726), .B2(n20370), .ZN(
        n20361) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20611), .ZN(n20360) );
  OAI211_X1 U23302 ( .C1(n20614), .C2(n20402), .A(n20361), .B(n20360), .ZN(
        P1_U3099) );
  AOI22_X1 U23303 ( .A1(n20616), .A2(n20371), .B1(n20615), .B2(n20370), .ZN(
        n20363) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20617), .ZN(n20362) );
  OAI211_X1 U23305 ( .C1(n20620), .C2(n20402), .A(n20363), .B(n20362), .ZN(
        P1_U3100) );
  AOI22_X1 U23306 ( .A1(n20622), .A2(n20371), .B1(n20621), .B2(n20370), .ZN(
        n20365) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20623), .ZN(n20364) );
  OAI211_X1 U23308 ( .C1(n20626), .C2(n20402), .A(n20365), .B(n20364), .ZN(
        P1_U3101) );
  AOI22_X1 U23309 ( .A1(n20628), .A2(n20371), .B1(n20627), .B2(n20370), .ZN(
        n20367) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20629), .ZN(n20366) );
  OAI211_X1 U23311 ( .C1(n20632), .C2(n20402), .A(n20367), .B(n20366), .ZN(
        P1_U3102) );
  AOI22_X1 U23312 ( .A1(n20633), .A2(n20371), .B1(n9684), .B2(n20370), .ZN(
        n20369) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20634), .ZN(n20368) );
  OAI211_X1 U23314 ( .C1(n20637), .C2(n20402), .A(n20369), .B(n20368), .ZN(
        P1_U3103) );
  AOI22_X1 U23315 ( .A1(n20641), .A2(n20371), .B1(n20638), .B2(n20370), .ZN(
        n20375) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20373), .B1(
        n20372), .B2(n20642), .ZN(n20374) );
  OAI211_X1 U23317 ( .C1(n20648), .C2(n20402), .A(n20375), .B(n20374), .ZN(
        P1_U3104) );
  NOR2_X1 U23318 ( .A1(n20509), .A2(n20377), .ZN(n20396) );
  AOI21_X1 U23319 ( .B1(n20442), .B2(n20376), .A(n20396), .ZN(n20378) );
  OAI22_X1 U23320 ( .A1(n20378), .A2(n20587), .B1(n20377), .B2(n10675), .ZN(
        n20397) );
  AOI22_X1 U23321 ( .A1(n20592), .A2(n20397), .B1(n20591), .B2(n20396), .ZN(
        n20383) );
  OAI211_X1 U23322 ( .C1(n20451), .C2(n20542), .A(n20510), .B(n20378), .ZN(
        n20379) );
  OAI211_X1 U23323 ( .C1(n20510), .C2(n20380), .A(n20597), .B(n20379), .ZN(
        n20399) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20551), .ZN(n20382) );
  OAI211_X1 U23325 ( .C1(n20554), .C2(n20402), .A(n20383), .B(n20382), .ZN(
        P1_U3105) );
  AOI22_X1 U23326 ( .A1(n20604), .A2(n20397), .B1(n20603), .B2(n20396), .ZN(
        n20385) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20555), .ZN(n20384) );
  OAI211_X1 U23328 ( .C1(n20558), .C2(n20402), .A(n20385), .B(n20384), .ZN(
        P1_U3106) );
  AOI22_X1 U23329 ( .A1(n20610), .A2(n20397), .B1(n9726), .B2(n20396), .ZN(
        n20387) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20559), .ZN(n20386) );
  OAI211_X1 U23331 ( .C1(n20562), .C2(n20402), .A(n20387), .B(n20386), .ZN(
        P1_U3107) );
  AOI22_X1 U23332 ( .A1(n20616), .A2(n20397), .B1(n20615), .B2(n20396), .ZN(
        n20389) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20563), .ZN(n20388) );
  OAI211_X1 U23334 ( .C1(n20566), .C2(n20402), .A(n20389), .B(n20388), .ZN(
        P1_U3108) );
  AOI22_X1 U23335 ( .A1(n20622), .A2(n20397), .B1(n20621), .B2(n20396), .ZN(
        n20391) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20567), .ZN(n20390) );
  OAI211_X1 U23337 ( .C1(n20570), .C2(n20402), .A(n20391), .B(n20390), .ZN(
        P1_U3109) );
  AOI22_X1 U23338 ( .A1(n20628), .A2(n20397), .B1(n20627), .B2(n20396), .ZN(
        n20393) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20571), .ZN(n20392) );
  OAI211_X1 U23340 ( .C1(n20574), .C2(n20402), .A(n20393), .B(n20392), .ZN(
        P1_U3110) );
  AOI22_X1 U23341 ( .A1(n20633), .A2(n20397), .B1(n9684), .B2(n20396), .ZN(
        n20395) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20575), .ZN(n20394) );
  OAI211_X1 U23343 ( .C1(n20578), .C2(n20402), .A(n20395), .B(n20394), .ZN(
        P1_U3111) );
  AOI22_X1 U23344 ( .A1(n20641), .A2(n20397), .B1(n20638), .B2(n20396), .ZN(
        n20401) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20399), .B1(
        n20398), .B2(n20581), .ZN(n20400) );
  OAI211_X1 U23346 ( .C1(n20586), .C2(n20402), .A(n20401), .B(n20400), .ZN(
        P1_U3112) );
  NOR3_X1 U23347 ( .A1(n20474), .A2(n10622), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20449) );
  NAND2_X1 U23348 ( .A1(n20509), .A2(n20449), .ZN(n20432) );
  OAI22_X1 U23349 ( .A1(n20434), .A2(n20554), .B1(n20403), .B2(n20432), .ZN(
        n20404) );
  INV_X1 U23350 ( .A(n20404), .ZN(n20414) );
  NAND2_X1 U23351 ( .A1(n20434), .A2(n20473), .ZN(n20405) );
  AOI21_X1 U23352 ( .B1(n20405), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20587), 
        .ZN(n20409) );
  NAND2_X1 U23353 ( .A1(n20442), .A2(n20544), .ZN(n20411) );
  AOI22_X1 U23354 ( .A1(n20409), .A2(n20411), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20432), .ZN(n20407) );
  OR2_X1 U23355 ( .A1(n20406), .A2(n20474), .ZN(n20539) );
  NAND2_X1 U23356 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20539), .ZN(n20547) );
  NAND3_X1 U23357 ( .A1(n20408), .A2(n20407), .A3(n20547), .ZN(n20437) );
  INV_X1 U23358 ( .A(n20409), .ZN(n20412) );
  OAI22_X1 U23359 ( .A1(n20412), .A2(n20411), .B1(n20410), .B2(n20539), .ZN(
        n20436) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20437), .B1(
        n20592), .B2(n20436), .ZN(n20413) );
  OAI211_X1 U23361 ( .C1(n20602), .C2(n20473), .A(n20414), .B(n20413), .ZN(
        P1_U3113) );
  INV_X1 U23362 ( .A(n20603), .ZN(n20415) );
  OAI22_X1 U23363 ( .A1(n20434), .A2(n20558), .B1(n20415), .B2(n20432), .ZN(
        n20416) );
  INV_X1 U23364 ( .A(n20416), .ZN(n20418) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20437), .B1(
        n20604), .B2(n20436), .ZN(n20417) );
  OAI211_X1 U23366 ( .C1(n20608), .C2(n20473), .A(n20418), .B(n20417), .ZN(
        P1_U3114) );
  INV_X1 U23367 ( .A(n9726), .ZN(n20419) );
  OAI22_X1 U23368 ( .A1(n20434), .A2(n20562), .B1(n20419), .B2(n20432), .ZN(
        n20420) );
  INV_X1 U23369 ( .A(n20420), .ZN(n20422) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20437), .B1(
        n20610), .B2(n20436), .ZN(n20421) );
  OAI211_X1 U23371 ( .C1(n20614), .C2(n20473), .A(n20422), .B(n20421), .ZN(
        P1_U3115) );
  INV_X1 U23372 ( .A(n20432), .ZN(n20429) );
  AOI22_X1 U23373 ( .A1(n20462), .A2(n20563), .B1(n20615), .B2(n20429), .ZN(
        n20424) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20437), .B1(
        n20616), .B2(n20436), .ZN(n20423) );
  OAI211_X1 U23375 ( .C1(n20566), .C2(n20434), .A(n20424), .B(n20423), .ZN(
        P1_U3116) );
  AOI22_X1 U23376 ( .A1(n20462), .A2(n20567), .B1(n20621), .B2(n20429), .ZN(
        n20426) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20437), .B1(
        n20622), .B2(n20436), .ZN(n20425) );
  OAI211_X1 U23378 ( .C1(n20570), .C2(n20434), .A(n20426), .B(n20425), .ZN(
        P1_U3117) );
  AOI22_X1 U23379 ( .A1(n20462), .A2(n20571), .B1(n20627), .B2(n20429), .ZN(
        n20428) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20437), .B1(
        n20628), .B2(n20436), .ZN(n20427) );
  OAI211_X1 U23381 ( .C1(n20574), .C2(n20434), .A(n20428), .B(n20427), .ZN(
        P1_U3118) );
  AOI22_X1 U23382 ( .A1(n20462), .A2(n20575), .B1(n9684), .B2(n20429), .ZN(
        n20431) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20437), .B1(
        n20633), .B2(n20436), .ZN(n20430) );
  OAI211_X1 U23384 ( .C1(n20578), .C2(n20434), .A(n20431), .B(n20430), .ZN(
        P1_U3119) );
  OAI22_X1 U23385 ( .A1(n20434), .A2(n20586), .B1(n20433), .B2(n20432), .ZN(
        n20435) );
  INV_X1 U23386 ( .A(n20435), .ZN(n20439) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20437), .B1(
        n20641), .B2(n20436), .ZN(n20438) );
  OAI211_X1 U23388 ( .C1(n20648), .C2(n20473), .A(n20439), .B(n20438), .ZN(
        P1_U3120) );
  NOR2_X1 U23389 ( .A1(n20440), .A2(n20474), .ZN(n20467) );
  AOI21_X1 U23390 ( .B1(n20442), .B2(n20441), .A(n20467), .ZN(n20445) );
  INV_X1 U23391 ( .A(n20449), .ZN(n20443) );
  OAI22_X1 U23392 ( .A1(n20445), .A2(n20587), .B1(n20443), .B2(n10675), .ZN(
        n20468) );
  AOI22_X1 U23393 ( .A1(n20592), .A2(n20468), .B1(n20591), .B2(n20467), .ZN(
        n20453) );
  INV_X1 U23394 ( .A(n20451), .ZN(n20444) );
  NOR2_X1 U23395 ( .A1(n20444), .A2(n20587), .ZN(n20447) );
  OAI21_X1 U23396 ( .B1(n20447), .B2(n20446), .A(n20445), .ZN(n20448) );
  OAI211_X1 U23397 ( .C1(n20510), .C2(n20449), .A(n20597), .B(n20448), .ZN(
        n20470) );
  INV_X1 U23398 ( .A(n20506), .ZN(n20469) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20470), .B1(
        n20469), .B2(n20551), .ZN(n20452) );
  OAI211_X1 U23400 ( .C1(n20554), .C2(n20473), .A(n20453), .B(n20452), .ZN(
        P1_U3121) );
  AOI22_X1 U23401 ( .A1(n20604), .A2(n20468), .B1(n20603), .B2(n20467), .ZN(
        n20455) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20470), .B1(
        n20469), .B2(n20555), .ZN(n20454) );
  OAI211_X1 U23403 ( .C1(n20558), .C2(n20473), .A(n20455), .B(n20454), .ZN(
        P1_U3122) );
  AOI22_X1 U23404 ( .A1(n20610), .A2(n20468), .B1(n9726), .B2(n20467), .ZN(
        n20457) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20470), .B1(
        n20462), .B2(n20611), .ZN(n20456) );
  OAI211_X1 U23406 ( .C1(n20614), .C2(n20506), .A(n20457), .B(n20456), .ZN(
        P1_U3123) );
  AOI22_X1 U23407 ( .A1(n20616), .A2(n20468), .B1(n20615), .B2(n20467), .ZN(
        n20459) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20470), .B1(
        n20462), .B2(n20617), .ZN(n20458) );
  OAI211_X1 U23409 ( .C1(n20620), .C2(n20506), .A(n20459), .B(n20458), .ZN(
        P1_U3124) );
  AOI22_X1 U23410 ( .A1(n20622), .A2(n20468), .B1(n20621), .B2(n20467), .ZN(
        n20461) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20470), .B1(
        n20469), .B2(n20567), .ZN(n20460) );
  OAI211_X1 U23412 ( .C1(n20570), .C2(n20473), .A(n20461), .B(n20460), .ZN(
        P1_U3125) );
  AOI22_X1 U23413 ( .A1(n20628), .A2(n20468), .B1(n20627), .B2(n20467), .ZN(
        n20464) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20470), .B1(
        n20462), .B2(n20629), .ZN(n20463) );
  OAI211_X1 U23415 ( .C1(n20632), .C2(n20506), .A(n20464), .B(n20463), .ZN(
        P1_U3126) );
  AOI22_X1 U23416 ( .A1(n20633), .A2(n20468), .B1(n9684), .B2(n20467), .ZN(
        n20466) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20470), .B1(
        n20469), .B2(n20575), .ZN(n20465) );
  OAI211_X1 U23418 ( .C1(n20578), .C2(n20473), .A(n20466), .B(n20465), .ZN(
        P1_U3127) );
  AOI22_X1 U23419 ( .A1(n20641), .A2(n20468), .B1(n20638), .B2(n20467), .ZN(
        n20472) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20470), .B1(
        n20469), .B2(n20581), .ZN(n20471) );
  OAI211_X1 U23421 ( .C1(n20586), .C2(n20473), .A(n20472), .B(n20471), .ZN(
        P1_U3128) );
  NOR3_X1 U23422 ( .A1(n10625), .A2(n20474), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20517) );
  NAND2_X1 U23423 ( .A1(n20509), .A2(n20517), .ZN(n20480) );
  INV_X1 U23424 ( .A(n20480), .ZN(n20501) );
  AOI22_X1 U23425 ( .A1(n20534), .A2(n20551), .B1(n20591), .B2(n20501), .ZN(
        n20488) );
  INV_X1 U23426 ( .A(n20484), .ZN(n20482) );
  NAND3_X1 U23427 ( .A1(n20475), .A2(n20506), .A3(n20510), .ZN(n20477) );
  NAND2_X1 U23428 ( .A1(n20477), .A2(n20476), .ZN(n20483) );
  NOR2_X1 U23429 ( .A1(n20479), .A2(n20478), .ZN(n20545) );
  NAND2_X1 U23430 ( .A1(n20545), .A2(n20540), .ZN(n20485) );
  AOI22_X1 U23431 ( .A1(n20483), .A2(n20485), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20480), .ZN(n20481) );
  OAI211_X1 U23432 ( .C1(n20482), .C2(n10675), .A(n20548), .B(n20481), .ZN(
        n20503) );
  INV_X1 U23433 ( .A(n20483), .ZN(n20486) );
  OAI22_X1 U23434 ( .A1(n20486), .A2(n20485), .B1(n20538), .B2(n20484), .ZN(
        n20502) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20503), .B1(
        n20592), .B2(n20502), .ZN(n20487) );
  OAI211_X1 U23436 ( .C1(n20554), .C2(n20506), .A(n20488), .B(n20487), .ZN(
        P1_U3129) );
  AOI22_X1 U23437 ( .A1(n20534), .A2(n20555), .B1(n20603), .B2(n20501), .ZN(
        n20490) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20503), .B1(
        n20604), .B2(n20502), .ZN(n20489) );
  OAI211_X1 U23439 ( .C1(n20558), .C2(n20506), .A(n20490), .B(n20489), .ZN(
        P1_U3130) );
  AOI22_X1 U23440 ( .A1(n20534), .A2(n20559), .B1(n9726), .B2(n20501), .ZN(
        n20492) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20503), .B1(
        n20610), .B2(n20502), .ZN(n20491) );
  OAI211_X1 U23442 ( .C1(n20562), .C2(n20506), .A(n20492), .B(n20491), .ZN(
        P1_U3131) );
  AOI22_X1 U23443 ( .A1(n20534), .A2(n20563), .B1(n20615), .B2(n20501), .ZN(
        n20494) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20503), .B1(
        n20616), .B2(n20502), .ZN(n20493) );
  OAI211_X1 U23445 ( .C1(n20566), .C2(n20506), .A(n20494), .B(n20493), .ZN(
        P1_U3132) );
  AOI22_X1 U23446 ( .A1(n20534), .A2(n20567), .B1(n20621), .B2(n20501), .ZN(
        n20496) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20503), .B1(
        n20622), .B2(n20502), .ZN(n20495) );
  OAI211_X1 U23448 ( .C1(n20570), .C2(n20506), .A(n20496), .B(n20495), .ZN(
        P1_U3133) );
  AOI22_X1 U23449 ( .A1(n20534), .A2(n20571), .B1(n20627), .B2(n20501), .ZN(
        n20498) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20503), .B1(
        n20628), .B2(n20502), .ZN(n20497) );
  OAI211_X1 U23451 ( .C1(n20574), .C2(n20506), .A(n20498), .B(n20497), .ZN(
        P1_U3134) );
  AOI22_X1 U23452 ( .A1(n20534), .A2(n20575), .B1(n9684), .B2(n20501), .ZN(
        n20500) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20503), .B1(
        n20633), .B2(n20502), .ZN(n20499) );
  OAI211_X1 U23454 ( .C1(n20578), .C2(n20506), .A(n20500), .B(n20499), .ZN(
        P1_U3135) );
  AOI22_X1 U23455 ( .A1(n20534), .A2(n20581), .B1(n20638), .B2(n20501), .ZN(
        n20505) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20503), .B1(
        n20641), .B2(n20502), .ZN(n20504) );
  OAI211_X1 U23457 ( .C1(n20586), .C2(n20506), .A(n20505), .B(n20504), .ZN(
        P1_U3136) );
  INV_X1 U23458 ( .A(n20515), .ZN(n20508) );
  INV_X1 U23459 ( .A(n20517), .ZN(n20512) );
  NOR2_X1 U23460 ( .A1(n20509), .A2(n20512), .ZN(n20532) );
  INV_X1 U23461 ( .A(n20532), .ZN(n20513) );
  NAND2_X1 U23462 ( .A1(n20545), .A2(n20510), .ZN(n20589) );
  OAI222_X1 U23463 ( .A1(n20513), .A2(n20587), .B1(n10675), .B2(n20512), .C1(
        n20511), .C2(n20589), .ZN(n20533) );
  AOI22_X1 U23464 ( .A1(n20592), .A2(n20533), .B1(n20591), .B2(n20532), .ZN(
        n20519) );
  NOR2_X1 U23465 ( .A1(n20515), .A2(n20514), .ZN(n20516) );
  OAI21_X1 U23466 ( .B1(n20517), .B2(n20516), .A(n20597), .ZN(n20535) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20599), .ZN(n20518) );
  OAI211_X1 U23468 ( .C1(n20602), .C2(n20585), .A(n20519), .B(n20518), .ZN(
        P1_U3137) );
  AOI22_X1 U23469 ( .A1(n20604), .A2(n20533), .B1(n20603), .B2(n20532), .ZN(
        n20521) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20605), .ZN(n20520) );
  OAI211_X1 U23471 ( .C1(n20608), .C2(n20585), .A(n20521), .B(n20520), .ZN(
        P1_U3138) );
  AOI22_X1 U23472 ( .A1(n20610), .A2(n20533), .B1(n9726), .B2(n20532), .ZN(
        n20523) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20611), .ZN(n20522) );
  OAI211_X1 U23474 ( .C1(n20614), .C2(n20585), .A(n20523), .B(n20522), .ZN(
        P1_U3139) );
  AOI22_X1 U23475 ( .A1(n20616), .A2(n20533), .B1(n20615), .B2(n20532), .ZN(
        n20525) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20617), .ZN(n20524) );
  OAI211_X1 U23477 ( .C1(n20620), .C2(n20585), .A(n20525), .B(n20524), .ZN(
        P1_U3140) );
  AOI22_X1 U23478 ( .A1(n20622), .A2(n20533), .B1(n20621), .B2(n20532), .ZN(
        n20527) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20623), .ZN(n20526) );
  OAI211_X1 U23480 ( .C1(n20626), .C2(n20585), .A(n20527), .B(n20526), .ZN(
        P1_U3141) );
  AOI22_X1 U23481 ( .A1(n20628), .A2(n20533), .B1(n20627), .B2(n20532), .ZN(
        n20529) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20629), .ZN(n20528) );
  OAI211_X1 U23483 ( .C1(n20632), .C2(n20585), .A(n20529), .B(n20528), .ZN(
        P1_U3142) );
  AOI22_X1 U23484 ( .A1(n20633), .A2(n20533), .B1(n9684), .B2(n20532), .ZN(
        n20531) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20634), .ZN(n20530) );
  OAI211_X1 U23486 ( .C1(n20637), .C2(n20585), .A(n20531), .B(n20530), .ZN(
        P1_U3143) );
  AOI22_X1 U23487 ( .A1(n20641), .A2(n20533), .B1(n20638), .B2(n20532), .ZN(
        n20537) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20535), .B1(
        n20534), .B2(n20642), .ZN(n20536) );
  OAI211_X1 U23489 ( .C1(n20648), .C2(n20585), .A(n20537), .B(n20536), .ZN(
        P1_U3144) );
  OAI22_X1 U23490 ( .A1(n20589), .A2(n20540), .B1(n20539), .B2(n20538), .ZN(
        n20580) );
  NOR2_X1 U23491 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20594), .ZN(
        n20579) );
  AOI22_X1 U23492 ( .A1(n20592), .A2(n20580), .B1(n20591), .B2(n20579), .ZN(
        n20553) );
  OR2_X1 U23493 ( .A1(n20595), .A2(n20541), .ZN(n20550) );
  AOI21_X1 U23494 ( .B1(n20585), .B2(n20550), .A(n20542), .ZN(n20543) );
  AOI21_X1 U23495 ( .B1(n20545), .B2(n20544), .A(n20543), .ZN(n20546) );
  NOR2_X1 U23496 ( .A1(n20546), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20551), .ZN(n20552) );
  OAI211_X1 U23498 ( .C1(n20554), .C2(n20585), .A(n20553), .B(n20552), .ZN(
        P1_U3145) );
  AOI22_X1 U23499 ( .A1(n20604), .A2(n20580), .B1(n20603), .B2(n20579), .ZN(
        n20557) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20555), .ZN(n20556) );
  OAI211_X1 U23501 ( .C1(n20558), .C2(n20585), .A(n20557), .B(n20556), .ZN(
        P1_U3146) );
  AOI22_X1 U23502 ( .A1(n20610), .A2(n20580), .B1(n9726), .B2(n20579), .ZN(
        n20561) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20559), .ZN(n20560) );
  OAI211_X1 U23504 ( .C1(n20562), .C2(n20585), .A(n20561), .B(n20560), .ZN(
        P1_U3147) );
  AOI22_X1 U23505 ( .A1(n20616), .A2(n20580), .B1(n20615), .B2(n20579), .ZN(
        n20565) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20563), .ZN(n20564) );
  OAI211_X1 U23507 ( .C1(n20566), .C2(n20585), .A(n20565), .B(n20564), .ZN(
        P1_U3148) );
  AOI22_X1 U23508 ( .A1(n20622), .A2(n20580), .B1(n20621), .B2(n20579), .ZN(
        n20569) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20567), .ZN(n20568) );
  OAI211_X1 U23510 ( .C1(n20570), .C2(n20585), .A(n20569), .B(n20568), .ZN(
        P1_U3149) );
  AOI22_X1 U23511 ( .A1(n20628), .A2(n20580), .B1(n20627), .B2(n20579), .ZN(
        n20573) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20571), .ZN(n20572) );
  OAI211_X1 U23513 ( .C1(n20574), .C2(n20585), .A(n20573), .B(n20572), .ZN(
        P1_U3150) );
  AOI22_X1 U23514 ( .A1(n20633), .A2(n20580), .B1(n9684), .B2(n20579), .ZN(
        n20577) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20575), .ZN(n20576) );
  OAI211_X1 U23516 ( .C1(n20578), .C2(n20585), .A(n20577), .B(n20576), .ZN(
        P1_U3151) );
  AOI22_X1 U23517 ( .A1(n20641), .A2(n20580), .B1(n20638), .B2(n20579), .ZN(
        n20584) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20582), .B1(
        n20643), .B2(n20581), .ZN(n20583) );
  OAI211_X1 U23519 ( .C1(n20586), .C2(n20585), .A(n20584), .B(n20583), .ZN(
        P1_U3152) );
  OAI222_X1 U23520 ( .A1(n20589), .A2(n20588), .B1(n10675), .B2(n20594), .C1(
        n20587), .C2(n20590), .ZN(n20640) );
  INV_X1 U23521 ( .A(n20590), .ZN(n20639) );
  AOI22_X1 U23522 ( .A1(n20592), .A2(n20640), .B1(n20639), .B2(n20591), .ZN(
        n20601) );
  INV_X1 U23523 ( .A(n20593), .ZN(n20596) );
  OAI21_X1 U23524 ( .B1(n20596), .B2(n20595), .A(n20594), .ZN(n20598) );
  NAND2_X1 U23525 ( .A1(n20598), .A2(n20597), .ZN(n20644) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20599), .ZN(n20600) );
  OAI211_X1 U23527 ( .C1(n20602), .C2(n20647), .A(n20601), .B(n20600), .ZN(
        P1_U3153) );
  AOI22_X1 U23528 ( .A1(n20604), .A2(n20640), .B1(n20639), .B2(n20603), .ZN(
        n20607) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20605), .ZN(n20606) );
  OAI211_X1 U23530 ( .C1(n20608), .C2(n20647), .A(n20607), .B(n20606), .ZN(
        P1_U3154) );
  AOI22_X1 U23531 ( .A1(n20610), .A2(n20640), .B1(n20639), .B2(n9726), .ZN(
        n20613) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20611), .ZN(n20612) );
  OAI211_X1 U23533 ( .C1(n20614), .C2(n20647), .A(n20613), .B(n20612), .ZN(
        P1_U3155) );
  AOI22_X1 U23534 ( .A1(n20616), .A2(n20640), .B1(n20639), .B2(n20615), .ZN(
        n20619) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20617), .ZN(n20618) );
  OAI211_X1 U23536 ( .C1(n20620), .C2(n20647), .A(n20619), .B(n20618), .ZN(
        P1_U3156) );
  AOI22_X1 U23537 ( .A1(n20622), .A2(n20640), .B1(n20639), .B2(n20621), .ZN(
        n20625) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20623), .ZN(n20624) );
  OAI211_X1 U23539 ( .C1(n20626), .C2(n20647), .A(n20625), .B(n20624), .ZN(
        P1_U3157) );
  AOI22_X1 U23540 ( .A1(n20628), .A2(n20640), .B1(n20639), .B2(n20627), .ZN(
        n20631) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20629), .ZN(n20630) );
  OAI211_X1 U23542 ( .C1(n20632), .C2(n20647), .A(n20631), .B(n20630), .ZN(
        P1_U3158) );
  AOI22_X1 U23543 ( .A1(n20633), .A2(n20640), .B1(n20639), .B2(n9684), .ZN(
        n20636) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20634), .ZN(n20635) );
  OAI211_X1 U23545 ( .C1(n20637), .C2(n20647), .A(n20636), .B(n20635), .ZN(
        P1_U3159) );
  AOI22_X1 U23546 ( .A1(n20641), .A2(n20640), .B1(n20639), .B2(n20638), .ZN(
        n20646) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20642), .ZN(n20645) );
  OAI211_X1 U23548 ( .C1(n20648), .C2(n20647), .A(n20646), .B(n20645), .ZN(
        P1_U3160) );
  NOR2_X1 U23549 ( .A1(n20650), .A2(n20649), .ZN(n20653) );
  OAI21_X1 U23550 ( .B1(n20653), .B2(n10675), .A(n20651), .ZN(P1_U3163) );
  INV_X1 U23551 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20840) );
  NOR2_X1 U23552 ( .A1(n20721), .A2(n20840), .ZN(P1_U3164) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20654), .ZN(
        P1_U3165) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20654), .ZN(
        P1_U3166) );
  AND2_X1 U23555 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20654), .ZN(
        P1_U3167) );
  AND2_X1 U23556 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20654), .ZN(
        P1_U3168) );
  AND2_X1 U23557 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20654), .ZN(
        P1_U3169) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20654), .ZN(
        P1_U3170) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20654), .ZN(
        P1_U3171) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20654), .ZN(
        P1_U3172) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20654), .ZN(
        P1_U3173) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20654), .ZN(
        P1_U3174) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20654), .ZN(
        P1_U3175) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20654), .ZN(
        P1_U3176) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20654), .ZN(
        P1_U3177) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20654), .ZN(
        P1_U3178) );
  INV_X1 U23567 ( .A(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20781) );
  NOR2_X1 U23568 ( .A1(n20721), .A2(n20781), .ZN(P1_U3179) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20654), .ZN(
        P1_U3180) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20654), .ZN(
        P1_U3181) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20654), .ZN(
        P1_U3182) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20654), .ZN(
        P1_U3183) );
  INV_X1 U23573 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20895) );
  NOR2_X1 U23574 ( .A1(n20721), .A2(n20895), .ZN(P1_U3184) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20654), .ZN(
        P1_U3185) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20654), .ZN(P1_U3186) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20654), .ZN(P1_U3187) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20654), .ZN(P1_U3188) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20654), .ZN(P1_U3189) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20654), .ZN(P1_U3190) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20654), .ZN(P1_U3191) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20654), .ZN(P1_U3192) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20654), .ZN(P1_U3193) );
  NAND2_X1 U23584 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n20655) );
  OAI211_X1 U23585 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n20664), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n20655), .ZN(n20656) );
  OAI21_X1 U23586 ( .B1(n20657), .B2(n20656), .A(n20750), .ZN(n20659) );
  OAI211_X1 U23587 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20662), .A(n20659), 
        .B(n20658), .ZN(P1_U3194) );
  OAI21_X1 U23588 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20664), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20669) );
  OAI211_X1 U23589 ( .C1(NA), .C2(n20741), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20670), .ZN(n20660) );
  OAI211_X1 U23590 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20661), .A(HOLD), .B(
        n20660), .ZN(n20667) );
  INV_X1 U23591 ( .A(n20662), .ZN(n20663) );
  OAI221_X1 U23592 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20665), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n20664), .A(n20663), .ZN(n20666) );
  OAI221_X1 U23593 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20669), .C1(n20668), 
        .C2(n20667), .A(n20666), .ZN(P1_U3196) );
  OR2_X1 U23594 ( .A1(n20736), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20707) );
  INV_X1 U23595 ( .A(n20707), .ZN(n20711) );
  OR2_X1 U23596 ( .A1(n20670), .A2(n20750), .ZN(n20709) );
  INV_X1 U23597 ( .A(n20709), .ZN(n20712) );
  AOI222_X1 U23598 ( .A1(n20711), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20750), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20712), .ZN(n20671) );
  INV_X1 U23599 ( .A(n20671), .ZN(P1_U3197) );
  AOI222_X1 U23600 ( .A1(n20712), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20750), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20711), .ZN(n20672) );
  INV_X1 U23601 ( .A(n20672), .ZN(P1_U3198) );
  OAI222_X1 U23602 ( .A1(n20709), .A2(n20675), .B1(n20674), .B2(n20738), .C1(
        n20673), .C2(n20707), .ZN(P1_U3199) );
  AOI222_X1 U23603 ( .A1(n20711), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20712), .ZN(n20676) );
  INV_X1 U23604 ( .A(n20676), .ZN(P1_U3200) );
  AOI222_X1 U23605 ( .A1(n20712), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20750), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20711), .ZN(n20677) );
  INV_X1 U23606 ( .A(n20677), .ZN(P1_U3201) );
  AOI222_X1 U23607 ( .A1(n20712), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20711), .ZN(n20678) );
  INV_X1 U23608 ( .A(n20678), .ZN(P1_U3202) );
  AOI222_X1 U23609 ( .A1(n20712), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20711), .ZN(n20679) );
  INV_X1 U23610 ( .A(n20679), .ZN(P1_U3203) );
  AOI222_X1 U23611 ( .A1(n20711), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20712), .ZN(n20680) );
  INV_X1 U23612 ( .A(n20680), .ZN(P1_U3204) );
  AOI222_X1 U23613 ( .A1(n20712), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20711), .ZN(n20681) );
  INV_X1 U23614 ( .A(n20681), .ZN(P1_U3205) );
  AOI222_X1 U23615 ( .A1(n20711), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20712), .ZN(n20682) );
  INV_X1 U23616 ( .A(n20682), .ZN(P1_U3206) );
  AOI222_X1 U23617 ( .A1(n20712), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20711), .ZN(n20683) );
  INV_X1 U23618 ( .A(n20683), .ZN(P1_U3207) );
  AOI222_X1 U23619 ( .A1(n20711), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20712), .ZN(n20684) );
  INV_X1 U23620 ( .A(n20684), .ZN(P1_U3208) );
  INV_X1 U23621 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20865) );
  OAI222_X1 U23622 ( .A1(n20709), .A2(n20686), .B1(n20865), .B2(n20738), .C1(
        n20685), .C2(n20707), .ZN(P1_U3209) );
  AOI222_X1 U23623 ( .A1(n20711), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20712), .ZN(n20687) );
  INV_X1 U23624 ( .A(n20687), .ZN(P1_U3210) );
  AOI222_X1 U23625 ( .A1(n20712), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20711), .ZN(n20688) );
  INV_X1 U23626 ( .A(n20688), .ZN(P1_U3211) );
  AOI222_X1 U23627 ( .A1(n20712), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20711), .ZN(n20689) );
  INV_X1 U23628 ( .A(n20689), .ZN(P1_U3212) );
  AOI22_X1 U23629 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20711), .ZN(n20690) );
  OAI21_X1 U23630 ( .B1(n20691), .B2(n20709), .A(n20690), .ZN(P1_U3213) );
  AOI22_X1 U23631 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20712), .ZN(n20692) );
  OAI21_X1 U23632 ( .B1(n20693), .B2(n20707), .A(n20692), .ZN(P1_U3214) );
  AOI222_X1 U23633 ( .A1(n20711), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20712), .ZN(n20694) );
  INV_X1 U23634 ( .A(n20694), .ZN(P1_U3215) );
  AOI222_X1 U23635 ( .A1(n20712), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20711), .ZN(n20695) );
  INV_X1 U23636 ( .A(n20695), .ZN(P1_U3216) );
  AOI222_X1 U23637 ( .A1(n20712), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20711), .ZN(n20696) );
  INV_X1 U23638 ( .A(n20696), .ZN(P1_U3217) );
  AOI22_X1 U23639 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20711), .ZN(n20697) );
  OAI21_X1 U23640 ( .B1(n20698), .B2(n20709), .A(n20697), .ZN(P1_U3218) );
  AOI22_X1 U23641 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20712), .ZN(n20699) );
  OAI21_X1 U23642 ( .B1(n20701), .B2(n20707), .A(n20699), .ZN(P1_U3219) );
  AOI22_X1 U23643 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n20711), .ZN(n20700) );
  OAI21_X1 U23644 ( .B1(n20701), .B2(n20709), .A(n20700), .ZN(P1_U3220) );
  AOI22_X1 U23645 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n20750), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n20712), .ZN(n20702) );
  OAI21_X1 U23646 ( .B1(n20703), .B2(n20707), .A(n20702), .ZN(P1_U3221) );
  AOI222_X1 U23647 ( .A1(n20712), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20711), .ZN(n20704) );
  INV_X1 U23648 ( .A(n20704), .ZN(P1_U3222) );
  AOI22_X1 U23649 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20711), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20736), .ZN(n20705) );
  OAI21_X1 U23650 ( .B1(n20821), .B2(n20709), .A(n20705), .ZN(P1_U3223) );
  AOI22_X1 U23651 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20712), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20736), .ZN(n20706) );
  OAI21_X1 U23652 ( .B1(n20710), .B2(n20707), .A(n20706), .ZN(P1_U3224) );
  AOI22_X1 U23653 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20711), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20736), .ZN(n20708) );
  OAI21_X1 U23654 ( .B1(n20710), .B2(n20709), .A(n20708), .ZN(P1_U3225) );
  AOI222_X1 U23655 ( .A1(n20712), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20711), .ZN(n20713) );
  INV_X1 U23656 ( .A(n20713), .ZN(P1_U3226) );
  OAI22_X1 U23657 ( .A1(n20750), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20738), .ZN(n20714) );
  INV_X1 U23658 ( .A(n20714), .ZN(P1_U3458) );
  OAI22_X1 U23659 ( .A1(n20750), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20738), .ZN(n20715) );
  INV_X1 U23660 ( .A(n20715), .ZN(P1_U3459) );
  OAI22_X1 U23661 ( .A1(n20750), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20738), .ZN(n20716) );
  INV_X1 U23662 ( .A(n20716), .ZN(P1_U3460) );
  OAI22_X1 U23663 ( .A1(n20750), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20738), .ZN(n20717) );
  INV_X1 U23664 ( .A(n20717), .ZN(P1_U3461) );
  OAI21_X1 U23665 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20721), .A(n20719), 
        .ZN(n20718) );
  INV_X1 U23666 ( .A(n20718), .ZN(P1_U3464) );
  OAI21_X1 U23667 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(P1_U3465) );
  OAI22_X1 U23668 ( .A1(n20725), .A2(n20724), .B1(n20723), .B2(n20722), .ZN(
        n20727) );
  MUX2_X1 U23669 ( .A(n20727), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20726), .Z(P1_U3469) );
  AOI21_X1 U23670 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20728) );
  AOI22_X1 U23671 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20728), .B2(n12396), .ZN(n20730) );
  INV_X1 U23672 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20729) );
  AOI22_X1 U23673 ( .A1(n20731), .A2(n20730), .B1(n20729), .B2(n20734), .ZN(
        P1_U3481) );
  INV_X1 U23674 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20735) );
  NOR2_X1 U23675 ( .A1(n20734), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20732) );
  AOI22_X1 U23676 ( .A1(n20735), .A2(n20734), .B1(n20733), .B2(n20732), .ZN(
        P1_U3482) );
  AOI22_X1 U23677 ( .A1(n20738), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20737), 
        .B2(n20736), .ZN(P1_U3483) );
  AOI211_X1 U23678 ( .C1(n20742), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        n20749) );
  OAI211_X1 U23679 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20744), .A(n20743), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20746) );
  AOI21_X1 U23680 ( .B1(n20746), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20745), 
        .ZN(n20748) );
  NAND2_X1 U23681 ( .A1(n20749), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20747) );
  OAI21_X1 U23682 ( .B1(n20749), .B2(n20748), .A(n20747), .ZN(P1_U3485) );
  MUX2_X1 U23683 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20750), .Z(P1_U3486) );
  NOR4_X1 U23684 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__3__SCAN_IN), .A3(P3_INSTQUEUE_REG_6__3__SCAN_IN), 
        .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n20754) );
  NOR4_X1 U23685 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P3_EBX_REG_23__SCAN_IN), .A3(P3_EBX_REG_7__SCAN_IN), .A4(
        P3_REIP_REG_13__SCAN_IN), .ZN(n20753) );
  NOR4_X1 U23686 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(BUF1_REG_21__SCAN_IN), .A4(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n20752) );
  NOR4_X1 U23687 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A4(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20751) );
  NAND4_X1 U23688 ( .A1(n20754), .A2(n20753), .A3(n20752), .A4(n20751), .ZN(
        n20771) );
  NAND4_X1 U23689 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_13__3__SCAN_IN), .A3(P1_REIP_REG_10__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n20770) );
  NOR4_X1 U23690 ( .A1(n20824), .A2(n20780), .A3(n20797), .A4(n20825), .ZN(
        n20757) );
  NOR4_X1 U23691 ( .A1(n11360), .A2(n11786), .A3(n20821), .A4(n20822), .ZN(
        n20756) );
  NOR3_X1 U23692 ( .A1(n20811), .A2(n20814), .A3(n20827), .ZN(n20755) );
  NAND4_X1 U23693 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20757), .A3(n20756), 
        .A4(n20755), .ZN(n20769) );
  NOR4_X1 U23694 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(
        P1_ADDRESS_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20767) );
  NOR4_X1 U23695 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(READY2), .ZN(n20766) );
  INV_X1 U23696 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n20864) );
  NAND4_X1 U23697 ( .A1(n20783), .A2(n20815), .A3(n20887), .A4(n20864), .ZN(
        n20758) );
  NOR4_X1 U23698 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(n20759), .A4(n20758), .ZN(n20765)
         );
  INV_X1 U23699 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20871) );
  NAND4_X1 U23700 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20871), .A3(n20829), .A4(
        n20792), .ZN(n20763) );
  NAND4_X1 U23701 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(P3_LWORD_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20762) );
  NAND4_X1 U23702 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P1_LWORD_REG_1__SCAN_IN), .A4(
        P2_UWORD_REG_6__SCAN_IN), .ZN(n20761) );
  NAND4_X1 U23703 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(P2_EAX_REG_26__SCAN_IN), 
        .A3(P2_DATAO_REG_15__SCAN_IN), .A4(P2_D_C_N_REG_SCAN_IN), .ZN(n20760)
         );
  NOR4_X1 U23704 ( .A1(n20763), .A2(n20762), .A3(n20761), .A4(n20760), .ZN(
        n20764) );
  NAND4_X1 U23705 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20768) );
  NOR4_X1 U23706 ( .A1(n20771), .A2(n20770), .A3(n20769), .A4(n20768), .ZN(
        n20910) );
  AOI22_X1 U23707 ( .A1(n20772), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(U215), .ZN(n20908) );
  AOI22_X1 U23708 ( .A1(n20775), .A2(keyinput16), .B1(keyinput1), .B2(n20774), 
        .ZN(n20773) );
  OAI221_X1 U23709 ( .B1(n20775), .B2(keyinput16), .C1(n20774), .C2(keyinput1), 
        .A(n20773), .ZN(n20788) );
  INV_X1 U23710 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23711 ( .A1(n20778), .A2(keyinput51), .B1(keyinput3), .B2(n20777), 
        .ZN(n20776) );
  OAI221_X1 U23712 ( .B1(n20778), .B2(keyinput51), .C1(n20777), .C2(keyinput3), 
        .A(n20776), .ZN(n20787) );
  AOI22_X1 U23713 ( .A1(n20781), .A2(keyinput43), .B1(n20780), .B2(keyinput21), 
        .ZN(n20779) );
  OAI221_X1 U23714 ( .B1(n20781), .B2(keyinput43), .C1(n20780), .C2(keyinput21), .A(n20779), .ZN(n20786) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U23716 ( .A1(n20784), .A2(keyinput0), .B1(n20783), .B2(keyinput17), 
        .ZN(n20782) );
  OAI221_X1 U23717 ( .B1(n20784), .B2(keyinput0), .C1(n20783), .C2(keyinput17), 
        .A(n20782), .ZN(n20785) );
  NOR4_X1 U23718 ( .A1(n20788), .A2(n20787), .A3(n20786), .A4(n20785), .ZN(
        n20837) );
  AOI22_X1 U23719 ( .A1(n20791), .A2(keyinput47), .B1(n20790), .B2(keyinput55), 
        .ZN(n20789) );
  OAI221_X1 U23720 ( .B1(n20791), .B2(keyinput47), .C1(n20790), .C2(keyinput55), .A(n20789), .ZN(n20795) );
  XOR2_X1 U23721 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B(keyinput14), .Z(
        n20794) );
  XNOR2_X1 U23722 ( .A(n20792), .B(keyinput6), .ZN(n20793) );
  OR3_X1 U23723 ( .A1(n20795), .A2(n20794), .A3(n20793), .ZN(n20804) );
  AOI22_X1 U23724 ( .A1(n20798), .A2(keyinput46), .B1(n20797), .B2(keyinput57), 
        .ZN(n20796) );
  OAI221_X1 U23725 ( .B1(n20798), .B2(keyinput46), .C1(n20797), .C2(keyinput57), .A(n20796), .ZN(n20803) );
  INV_X1 U23726 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n20800) );
  AOI22_X1 U23727 ( .A1(n20801), .A2(keyinput48), .B1(keyinput53), .B2(n20800), 
        .ZN(n20799) );
  OAI221_X1 U23728 ( .B1(n20801), .B2(keyinput48), .C1(n20800), .C2(keyinput53), .A(n20799), .ZN(n20802) );
  NOR3_X1 U23729 ( .A1(n20804), .A2(n20803), .A3(n20802), .ZN(n20836) );
  AOI22_X1 U23730 ( .A1(n20806), .A2(keyinput7), .B1(n12920), .B2(keyinput26), 
        .ZN(n20805) );
  OAI221_X1 U23731 ( .B1(n20806), .B2(keyinput7), .C1(n12920), .C2(keyinput26), 
        .A(n20805), .ZN(n20819) );
  AOI22_X1 U23732 ( .A1(n20809), .A2(keyinput4), .B1(n20808), .B2(keyinput44), 
        .ZN(n20807) );
  OAI221_X1 U23733 ( .B1(n20809), .B2(keyinput4), .C1(n20808), .C2(keyinput44), 
        .A(n20807), .ZN(n20818) );
  AOI22_X1 U23734 ( .A1(n20812), .A2(keyinput42), .B1(n20811), .B2(keyinput60), 
        .ZN(n20810) );
  OAI221_X1 U23735 ( .B1(n20812), .B2(keyinput42), .C1(n20811), .C2(keyinput60), .A(n20810), .ZN(n20817) );
  AOI22_X1 U23736 ( .A1(n20815), .A2(keyinput23), .B1(keyinput36), .B2(n20814), 
        .ZN(n20813) );
  OAI221_X1 U23737 ( .B1(n20815), .B2(keyinput23), .C1(n20814), .C2(keyinput36), .A(n20813), .ZN(n20816) );
  NOR4_X1 U23738 ( .A1(n20819), .A2(n20818), .A3(n20817), .A4(n20816), .ZN(
        n20835) );
  AOI22_X1 U23739 ( .A1(n20822), .A2(keyinput52), .B1(n20821), .B2(keyinput2), 
        .ZN(n20820) );
  OAI221_X1 U23740 ( .B1(n20822), .B2(keyinput52), .C1(n20821), .C2(keyinput2), 
        .A(n20820), .ZN(n20833) );
  AOI22_X1 U23741 ( .A1(n20825), .A2(keyinput35), .B1(n20824), .B2(keyinput33), 
        .ZN(n20823) );
  OAI221_X1 U23742 ( .B1(n20825), .B2(keyinput35), .C1(n20824), .C2(keyinput33), .A(n20823), .ZN(n20832) );
  AOI22_X1 U23743 ( .A1(n11786), .A2(keyinput31), .B1(keyinput54), .B2(n20827), 
        .ZN(n20826) );
  OAI221_X1 U23744 ( .B1(n11786), .B2(keyinput31), .C1(n20827), .C2(keyinput54), .A(n20826), .ZN(n20831) );
  AOI22_X1 U23745 ( .A1(n11360), .A2(keyinput39), .B1(keyinput29), .B2(n20829), 
        .ZN(n20828) );
  OAI221_X1 U23746 ( .B1(n11360), .B2(keyinput39), .C1(n20829), .C2(keyinput29), .A(n20828), .ZN(n20830) );
  NOR4_X1 U23747 ( .A1(n20833), .A2(n20832), .A3(n20831), .A4(n20830), .ZN(
        n20834) );
  NAND4_X1 U23748 ( .A1(n20837), .A2(n20836), .A3(n20835), .A4(n20834), .ZN(
        n20906) );
  INV_X1 U23749 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n20839) );
  AOI22_X1 U23750 ( .A1(n20840), .A2(keyinput41), .B1(n20839), .B2(keyinput27), 
        .ZN(n20838) );
  OAI221_X1 U23751 ( .B1(n20840), .B2(keyinput41), .C1(n20839), .C2(keyinput27), .A(n20838), .ZN(n20853) );
  INV_X1 U23752 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n20843) );
  AOI22_X1 U23753 ( .A1(n20843), .A2(keyinput56), .B1(n20842), .B2(keyinput32), 
        .ZN(n20841) );
  OAI221_X1 U23754 ( .B1(n20843), .B2(keyinput56), .C1(n20842), .C2(keyinput32), .A(n20841), .ZN(n20852) );
  AOI22_X1 U23755 ( .A1(n20846), .A2(keyinput15), .B1(n20845), .B2(keyinput8), 
        .ZN(n20844) );
  OAI221_X1 U23756 ( .B1(n20846), .B2(keyinput15), .C1(n20845), .C2(keyinput8), 
        .A(n20844), .ZN(n20851) );
  INV_X1 U23757 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n20849) );
  AOI22_X1 U23758 ( .A1(n20849), .A2(keyinput25), .B1(n20848), .B2(keyinput49), 
        .ZN(n20847) );
  OAI221_X1 U23759 ( .B1(n20849), .B2(keyinput25), .C1(n20848), .C2(keyinput49), .A(n20847), .ZN(n20850) );
  NOR4_X1 U23760 ( .A1(n20853), .A2(n20852), .A3(n20851), .A4(n20850), .ZN(
        n20904) );
  INV_X1 U23761 ( .A(READY2), .ZN(n20855) );
  AOI22_X1 U23762 ( .A1(n20856), .A2(keyinput18), .B1(n20855), .B2(keyinput58), 
        .ZN(n20854) );
  OAI221_X1 U23763 ( .B1(n20856), .B2(keyinput18), .C1(n20855), .C2(keyinput58), .A(n20854), .ZN(n20869) );
  AOI22_X1 U23764 ( .A1(n20859), .A2(keyinput13), .B1(n20858), .B2(keyinput12), 
        .ZN(n20857) );
  OAI221_X1 U23765 ( .B1(n20859), .B2(keyinput13), .C1(n20858), .C2(keyinput12), .A(n20857), .ZN(n20868) );
  AOI22_X1 U23766 ( .A1(n20862), .A2(keyinput38), .B1(n20861), .B2(keyinput40), 
        .ZN(n20860) );
  OAI221_X1 U23767 ( .B1(n20862), .B2(keyinput38), .C1(n20861), .C2(keyinput40), .A(n20860), .ZN(n20867) );
  AOI22_X1 U23768 ( .A1(n20865), .A2(keyinput30), .B1(keyinput63), .B2(n20864), 
        .ZN(n20863) );
  OAI221_X1 U23769 ( .B1(n20865), .B2(keyinput30), .C1(n20864), .C2(keyinput63), .A(n20863), .ZN(n20866) );
  NOR4_X1 U23770 ( .A1(n20869), .A2(n20868), .A3(n20867), .A4(n20866), .ZN(
        n20903) );
  INV_X1 U23771 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U23772 ( .A1(n20872), .A2(keyinput10), .B1(n20871), .B2(keyinput5), 
        .ZN(n20870) );
  OAI221_X1 U23773 ( .B1(n20872), .B2(keyinput10), .C1(n20871), .C2(keyinput5), 
        .A(n20870), .ZN(n20885) );
  AOI22_X1 U23774 ( .A1(n20875), .A2(keyinput59), .B1(n20874), .B2(keyinput61), 
        .ZN(n20873) );
  OAI221_X1 U23775 ( .B1(n20875), .B2(keyinput59), .C1(n20874), .C2(keyinput61), .A(n20873), .ZN(n20884) );
  AOI22_X1 U23776 ( .A1(n20878), .A2(keyinput24), .B1(n20877), .B2(keyinput20), 
        .ZN(n20876) );
  OAI221_X1 U23777 ( .B1(n20878), .B2(keyinput24), .C1(n20877), .C2(keyinput20), .A(n20876), .ZN(n20883) );
  INV_X1 U23778 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20881) );
  INV_X1 U23779 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U23780 ( .A1(n20881), .A2(keyinput45), .B1(n20880), .B2(keyinput9), 
        .ZN(n20879) );
  OAI221_X1 U23781 ( .B1(n20881), .B2(keyinput45), .C1(n20880), .C2(keyinput9), 
        .A(n20879), .ZN(n20882) );
  NOR4_X1 U23782 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n20902) );
  AOI22_X1 U23783 ( .A1(n20887), .A2(keyinput34), .B1(n14499), .B2(keyinput62), 
        .ZN(n20886) );
  OAI221_X1 U23784 ( .B1(n20887), .B2(keyinput34), .C1(n14499), .C2(keyinput62), .A(n20886), .ZN(n20900) );
  INV_X1 U23785 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23786 ( .A1(n20890), .A2(keyinput28), .B1(keyinput22), .B2(n20889), 
        .ZN(n20888) );
  OAI221_X1 U23787 ( .B1(n20890), .B2(keyinput28), .C1(n20889), .C2(keyinput22), .A(n20888), .ZN(n20899) );
  AOI22_X1 U23788 ( .A1(n20893), .A2(keyinput19), .B1(keyinput50), .B2(n20892), 
        .ZN(n20891) );
  OAI221_X1 U23789 ( .B1(n20893), .B2(keyinput19), .C1(n20892), .C2(keyinput50), .A(n20891), .ZN(n20898) );
  INV_X1 U23790 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U23791 ( .A1(n20896), .A2(keyinput37), .B1(keyinput11), .B2(n20895), 
        .ZN(n20894) );
  OAI221_X1 U23792 ( .B1(n20896), .B2(keyinput37), .C1(n20895), .C2(keyinput11), .A(n20894), .ZN(n20897) );
  NOR4_X1 U23793 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20901) );
  NAND4_X1 U23794 ( .A1(n20904), .A2(n20903), .A3(n20902), .A4(n20901), .ZN(
        n20905) );
  NOR2_X1 U23795 ( .A1(n20906), .A2(n20905), .ZN(n20907) );
  XOR2_X1 U23796 ( .A(n20908), .B(n20907), .Z(n20909) );
  XNOR2_X1 U23797 ( .A(n20910), .B(n20909), .ZN(U274) );
  AND2_X1 U11723 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10245) );
  XOR2_X1 U11109 ( .A(n13598), .B(n13597), .Z(n14065) );
  CLKBUF_X1 U11086 ( .A(n10816), .Z(n11084) );
  CLKBUF_X1 U11095 ( .A(n12658), .Z(n13579) );
  NAND2_X2 U11100 ( .A1(n12501), .A2(n13585), .ZN(n13590) );
  CLKBUF_X1 U11104 ( .A(n11556), .Z(n11646) );
  CLKBUF_X1 U11140 ( .A(n12446), .Z(n9587) );
  CLKBUF_X1 U11354 ( .A(n18731), .Z(n9588) );
  XNOR2_X1 U11387 ( .A(n13652), .B(n13630), .ZN(n13927) );
  CLKBUF_X1 U11404 ( .A(n19210), .Z(n19190) );
  CLKBUF_X1 U12177 ( .A(n11942), .Z(n11990) );
  CLKBUF_X1 U12485 ( .A(n17924), .Z(n9589) );
endmodule

