

module b14_C_gen_AntiSAT_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744;

  OR2_X1 U2281 ( .A1(n3907), .A2(n2149), .ZN(n2733) );
  INV_X2 U2282 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X2 U2283 ( .A(n3462), .ZN(n3505) );
  INV_X2 U2284 ( .A(n2302), .ZN(n3636) );
  NAND2_X1 U2285 ( .A1(n2627), .A2(n3795), .ZN(n2836) );
  INV_X1 U2286 ( .A(n2872), .ZN(n4198) );
  AND2_X1 U2287 ( .A1(n2046), .A2(n2292), .ZN(n2725) );
  NOR2_X1 U2288 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2267)
         );
  INV_X1 U2289 ( .A(n3503), .ZN(n3461) );
  INV_X1 U2290 ( .A(n3504), .ZN(n2887) );
  AND2_X1 U2291 ( .A1(n2836), .A2(n2847), .ZN(n3451) );
  OR2_X1 U2292 ( .A1(n3934), .A2(n2584), .ZN(n2252) );
  MUX2_X1 U2294 ( .A(DATAI_3_), .B(n3832), .S(n2040), .Z(n3045) );
  OAI21_X1 U2295 ( .B1(n2040), .B2(n2157), .A(n2156), .ZN(n2872) );
  NAND3_X1 U2296 ( .A1(n2690), .A2(n4409), .A3(n2741), .ZN(n2835) );
  AND2_X1 U2297 ( .A1(n2287), .A2(n2286), .ZN(n2039) );
  OAI21_X2 U2298 ( .B1(n3066), .B2(n2351), .A(n2350), .ZN(n3077) );
  OAI21_X1 U2301 ( .B1(n2733), .B2(n4551), .A(n2259), .ZN(n2732) );
  AOI21_X1 U2302 ( .B1(n4347), .B2(n4346), .A(n4345), .ZN(n4348) );
  AOI21_X1 U2303 ( .B1(n4221), .B2(n4347), .A(n4220), .ZN(n4222) );
  AOI21_X1 U2304 ( .B1(n3481), .B2(n3448), .A(n3447), .ZN(n3562) );
  NAND2_X1 U2305 ( .A1(n4216), .A2(n2715), .ZN(n2716) );
  OAI22_X1 U2306 ( .A1(n3205), .A2(n4515), .B1(n3219), .B2(n2079), .ZN(n4432)
         );
  NAND2_X1 U2307 ( .A1(n2854), .A2(n2855), .ZN(n2896) );
  AND2_X2 U2308 ( .A1(n3013), .A2(n4513), .ZN(n4525) );
  INV_X1 U2309 ( .A(n3818), .ZN(n3108) );
  NAND4_X2 U2311 ( .A1(n2318), .A2(n2317), .A3(n2316), .A4(n2315), .ZN(n4183)
         );
  INV_X1 U2312 ( .A(n2977), .ZN(n2888) );
  INV_X2 U2313 ( .A(n3451), .ZN(n3508) );
  NAND2_X1 U2314 ( .A1(n2109), .A2(n2835), .ZN(n3504) );
  CLKBUF_X3 U2315 ( .A(n2303), .Z(n3639) );
  INV_X1 U2316 ( .A(n3045), .ZN(n2942) );
  NAND2_X1 U2318 ( .A1(n2749), .A2(IR_REG_31__SCAN_IN), .ZN(n2283) );
  XNOR2_X1 U2319 ( .A(n2280), .B(IR_REG_29__SCAN_IN), .ZN(n2746) );
  OR2_X1 U2320 ( .A1(n2282), .A2(n2748), .ZN(n2280) );
  AND2_X1 U2321 ( .A1(n2620), .A2(n2254), .ZN(n2282) );
  AND2_X1 U2322 ( .A1(n2442), .A2(n2276), .ZN(n2620) );
  AND2_X1 U2323 ( .A1(n2133), .A2(n2278), .ZN(n2132) );
  AND4_X1 U2324 ( .A1(n2275), .A2(n2274), .A3(n2273), .A4(n2272), .ZN(n2276)
         );
  AND3_X1 U2325 ( .A1(n2265), .A2(n2319), .A3(n2266), .ZN(n2075) );
  AND3_X1 U2326 ( .A1(n2669), .A2(n2277), .A3(n2623), .ZN(n2278) );
  NOR2_X2 U2327 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2308)
         );
  INV_X1 U2328 ( .A(IR_REG_3__SCAN_IN), .ZN(n2319) );
  NOR2_X1 U2329 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2669)
         );
  NOR2_X1 U2330 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2277)
         );
  INV_X1 U2331 ( .A(IR_REG_15__SCAN_IN), .ZN(n2481) );
  NOR2_X1 U2332 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2272)
         );
  NOR2_X1 U2333 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2273)
         );
  OAI21_X2 U2334 ( .B1(n3176), .B2(n2240), .A(n2239), .ZN(n3191) );
  OAI21_X2 U2335 ( .B1(n3947), .B2(n2574), .A(n2573), .ZN(n3934) );
  NAND2_X2 U2336 ( .A1(n2563), .A2(n2562), .ZN(n3947) );
  NOR2_X2 U2337 ( .A1(n3974), .A2(n4236), .ZN(n3952) );
  OR2_X2 U2338 ( .A1(n3993), .A2(n2703), .ZN(n3974) );
  NAND2_X2 U2339 ( .A1(n2294), .A2(n2293), .ZN(n2040) );
  NAND2_X2 U2340 ( .A1(n2294), .A2(n2293), .ZN(n2041) );
  NAND2_X1 U2341 ( .A1(n2294), .A2(n2293), .ZN(n2560) );
  NOR2_X1 U2342 ( .A1(n3172), .A2(n3124), .ZN(n2360) );
  NOR2_X1 U2343 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2274)
         );
  INV_X1 U2344 ( .A(IR_REG_13__SCAN_IN), .ZN(n2444) );
  AOI21_X1 U2345 ( .B1(n2236), .B2(n2238), .A(n2061), .ZN(n2235) );
  AOI21_X1 U2346 ( .B1(n2188), .B2(n2191), .A(n2187), .ZN(n2186) );
  INV_X1 U2347 ( .A(n3235), .ZN(n2187) );
  INV_X1 U2348 ( .A(n2188), .ZN(n2107) );
  NOR2_X1 U2349 ( .A1(n2540), .A2(n2233), .ZN(n2232) );
  INV_X1 U2350 ( .A(n2533), .ZN(n2233) );
  NAND2_X1 U2351 ( .A1(n4303), .A2(n3379), .ZN(n2227) );
  INV_X1 U2352 ( .A(IR_REG_26__SCAN_IN), .ZN(n2256) );
  INV_X1 U2353 ( .A(IR_REG_27__SCAN_IN), .ZN(n2279) );
  INV_X1 U2354 ( .A(n2271), .ZN(n2133) );
  INV_X1 U2355 ( .A(n2945), .ZN(n2172) );
  OR2_X1 U2356 ( .A1(n2585), .A2(n3615), .ZN(n2596) );
  INV_X1 U2357 ( .A(n2488), .ZN(n3635) );
  XNOR2_X1 U2358 ( .A(n3207), .B(n4534), .ZN(n4443) );
  NAND2_X1 U2359 ( .A1(n4452), .A2(n4453), .ZN(n4451) );
  NAND2_X1 U2360 ( .A1(n4494), .A2(n2470), .ZN(n4493) );
  NOR2_X1 U2361 ( .A1(n2592), .A2(n2251), .ZN(n2250) );
  INV_X1 U2362 ( .A(n2583), .ZN(n2251) );
  AOI21_X1 U2363 ( .B1(n3914), .B2(n2660), .A(n2659), .ZN(n3370) );
  NAND2_X1 U2364 ( .A1(n2216), .A2(n2215), .ZN(n4110) );
  AOI21_X1 U2365 ( .B1(n2218), .B2(n2222), .A(n2060), .ZN(n2215) );
  NOR2_X1 U2366 ( .A1(n3191), .A2(n2264), .ZN(n2397) );
  NAND2_X1 U2367 ( .A1(n2726), .A2(n2255), .ZN(n2294) );
  NOR2_X1 U2368 ( .A1(n2271), .A2(IR_REG_21__SCAN_IN), .ZN(n2074) );
  OAI21_X1 U2369 ( .B1(n2518), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2520) );
  AND2_X1 U2370 ( .A1(n2492), .A2(n2444), .ZN(n2201) );
  INV_X1 U2371 ( .A(n3416), .ZN(n3419) );
  INV_X1 U2372 ( .A(n3417), .ZN(n3418) );
  OR2_X1 U2373 ( .A1(n3493), .A2(n2184), .ZN(n2183) );
  INV_X1 U2374 ( .A(n3602), .ZN(n2184) );
  NAND2_X1 U2375 ( .A1(n2073), .A2(n3472), .ZN(n3392) );
  INV_X1 U2376 ( .A(n3473), .ZN(n2071) );
  OR2_X1 U2377 ( .A1(n2881), .A2(n2081), .ZN(n2080) );
  AND2_X1 U2378 ( .A1(n4414), .A2(REG2_REG_7__SCAN_IN), .ZN(n2081) );
  NAND2_X1 U2379 ( .A1(n4454), .A2(n3209), .ZN(n3210) );
  INV_X1 U2380 ( .A(n3857), .ZN(n2089) );
  AND2_X1 U2381 ( .A1(n3773), .A2(n3772), .ZN(n2144) );
  NAND2_X1 U2382 ( .A1(n2144), .A2(n2044), .ZN(n2143) );
  AND2_X1 U2383 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
  INV_X1 U2384 ( .A(n3693), .ZN(n2146) );
  INV_X1 U2385 ( .A(n4074), .ZN(n2148) );
  INV_X1 U2386 ( .A(n3670), .ZN(n2140) );
  INV_X1 U2387 ( .A(n3668), .ZN(n2137) );
  INV_X1 U2388 ( .A(n2746), .ZN(n2214) );
  NAND2_X1 U2389 ( .A1(n3651), .A2(n2637), .ZN(n2636) );
  NAND2_X1 U2390 ( .A1(n2594), .A2(REG3_REG_27__SCAN_IN), .ZN(n2608) );
  NOR2_X1 U2391 ( .A1(n3609), .A2(n2102), .ZN(n2101) );
  INV_X1 U2392 ( .A(n3532), .ZN(n2102) );
  NAND2_X1 U2393 ( .A1(n2175), .A2(n2173), .ZN(n2072) );
  NOR2_X1 U2394 ( .A1(n3585), .A2(n2174), .ZN(n2173) );
  NAND2_X1 U2395 ( .A1(n2197), .A2(n2058), .ZN(n2195) );
  AOI21_X1 U2396 ( .B1(n2186), .B2(n2107), .A(n2052), .ZN(n2106) );
  INV_X1 U2397 ( .A(n2186), .ZN(n2108) );
  XNOR2_X1 U2398 ( .A(n2941), .B(n3508), .ZN(n2988) );
  NAND2_X1 U2399 ( .A1(n2100), .A2(n3610), .ZN(n2099) );
  NAND2_X1 U2400 ( .A1(n2101), .A2(n3531), .ZN(n2100) );
  AOI21_X1 U2401 ( .B1(n2834), .B2(n2887), .A(n2837), .ZN(n2851) );
  AND2_X1 U2402 ( .A1(n3330), .A2(n3329), .ZN(n3376) );
  NAND2_X1 U2403 ( .A1(n3399), .A2(n3398), .ZN(n3400) );
  INV_X1 U2404 ( .A(n4183), .ZN(n2998) );
  INV_X1 U2405 ( .A(n3142), .ZN(n2192) );
  NAND2_X1 U2406 ( .A1(n2839), .A2(n2069), .ZN(n2168) );
  AOI21_X1 U2407 ( .B1(n2887), .B2(n3058), .A(n2070), .ZN(n2069) );
  AND2_X1 U2408 ( .A1(n2947), .A2(IR_REG_0__SCAN_IN), .ZN(n2070) );
  NAND2_X1 U2409 ( .A1(n2168), .A2(n2840), .ZN(n2853) );
  AND2_X1 U2410 ( .A1(n3594), .A2(n3433), .ZN(n2197) );
  INV_X1 U2411 ( .A(n2901), .ZN(n2899) );
  OR2_X1 U2412 ( .A1(n2846), .A2(n3506), .ZN(n2850) );
  AND2_X1 U2413 ( .A1(n2336), .A2(REG3_REG_5__SCAN_IN), .ZN(n2352) );
  OR2_X1 U2414 ( .A1(n4412), .A2(n2824), .ZN(n2847) );
  AND2_X1 U2415 ( .A1(n2572), .A2(n2571), .ZN(n3486) );
  NOR2_X1 U2416 ( .A1(n2302), .A2(n2328), .ZN(n2329) );
  INV_X1 U2417 ( .A(n2086), .ZN(n2083) );
  OAI21_X1 U2418 ( .B1(n2926), .B2(n2083), .A(n2082), .ZN(n2085) );
  AOI21_X1 U2419 ( .B1(n2086), .B2(n2324), .A(n2771), .ZN(n2082) );
  NOR2_X1 U2420 ( .A1(n2810), .A2(n2809), .ZN(n2881) );
  XNOR2_X1 U2421 ( .A(n2080), .B(n4413), .ZN(n3205) );
  OAI21_X1 U2422 ( .B1(n2877), .B2(n2212), .A(n2211), .ZN(n2879) );
  NAND2_X1 U2423 ( .A1(n4414), .A2(REG1_REG_7__SCAN_IN), .ZN(n2211) );
  NOR2_X1 U2424 ( .A1(n4414), .A2(REG1_REG_7__SCAN_IN), .ZN(n2212) );
  NAND2_X1 U2425 ( .A1(n4430), .A2(n3206), .ZN(n3207) );
  NAND2_X1 U2426 ( .A1(n4443), .A2(REG2_REG_10__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U2427 ( .A1(n4447), .A2(n3224), .ZN(n4452) );
  XNOR2_X1 U2428 ( .A(n3210), .B(n2167), .ZN(n4465) );
  NAND2_X1 U2429 ( .A1(n4465), .A2(REG2_REG_12__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U2430 ( .A1(n4469), .A2(n3227), .ZN(n3229) );
  NAND2_X1 U2431 ( .A1(n3229), .A2(n3228), .ZN(n3843) );
  XNOR2_X1 U2432 ( .A(n3859), .B(n4531), .ZN(n4475) );
  NAND2_X1 U2433 ( .A1(n4493), .A2(n3865), .ZN(n2091) );
  NAND2_X1 U2434 ( .A1(n2091), .A2(n3866), .ZN(n3875) );
  NAND2_X1 U2435 ( .A1(n3875), .A2(n2165), .ZN(n2164) );
  NAND2_X1 U2436 ( .A1(n3872), .A2(n2166), .ZN(n2165) );
  INV_X1 U2437 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2166) );
  NAND2_X1 U2438 ( .A1(n2207), .A2(n2210), .ZN(n2208) );
  INV_X1 U2439 ( .A(n2246), .ZN(n2245) );
  NAND2_X1 U2440 ( .A1(n2053), .A2(n2253), .ZN(n2243) );
  OAI21_X1 U2441 ( .B1(n2606), .B2(n2247), .A(n2605), .ZN(n2246) );
  NAND2_X1 U2442 ( .A1(n3370), .A2(n3787), .ZN(n3369) );
  OR2_X1 U2443 ( .A1(n3950), .A2(n3720), .ZN(n3930) );
  OR2_X1 U2444 ( .A1(n2543), .A2(n2542), .ZN(n2553) );
  NAND2_X1 U2445 ( .A1(n2525), .A2(REG3_REG_20__SCAN_IN), .ZN(n2543) );
  AOI21_X1 U2446 ( .B1(n2232), .B2(n2045), .A(n2059), .ZN(n2231) );
  NAND2_X1 U2447 ( .A1(n4016), .A2(n2232), .ZN(n2230) );
  INV_X1 U2448 ( .A(n4069), .ZN(n2506) );
  AND2_X1 U2449 ( .A1(n4041), .A2(n4042), .ZN(n4069) );
  NAND2_X1 U2450 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  AOI21_X1 U2451 ( .B1(n2221), .B2(n2220), .A(n2219), .ZN(n2218) );
  INV_X1 U2452 ( .A(n2224), .ZN(n2220) );
  INV_X1 U2453 ( .A(n2227), .ZN(n2223) );
  AND2_X1 U2454 ( .A1(n2227), .A2(n2434), .ZN(n2224) );
  OAI21_X1 U2455 ( .B1(n3193), .B2(n3192), .A(n3671), .ZN(n3262) );
  INV_X1 U2456 ( .A(n2241), .ZN(n2240) );
  AOI21_X1 U2457 ( .B1(n2241), .B2(n2262), .A(n2051), .ZN(n2239) );
  AOI21_X1 U2458 ( .B1(n3731), .B2(n2242), .A(n2382), .ZN(n2241) );
  NAND2_X1 U2459 ( .A1(n2372), .A2(REG3_REG_8__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U2460 ( .A1(n2352), .A2(REG3_REG_6__SCAN_IN), .ZN(n2363) );
  AND2_X1 U2461 ( .A1(n2642), .A2(n3668), .ZN(n3731) );
  NAND2_X1 U2462 ( .A1(n2640), .A2(n3663), .ZN(n3068) );
  NAND2_X1 U2463 ( .A1(n2975), .A2(n2114), .ZN(n2640) );
  NOR2_X1 U2464 ( .A1(n2639), .A2(n2115), .ZN(n2114) );
  INV_X1 U2465 ( .A(n3809), .ZN(n4240) );
  NOR2_X2 U2466 ( .A1(n4078), .A2(n4274), .ZN(n4079) );
  NOR2_X1 U2467 ( .A1(n3176), .A2(n3731), .ZN(n4547) );
  INV_X1 U2468 ( .A(n4306), .ZN(n4098) );
  AND4_X1 U2469 ( .A1(n2345), .A2(n2344), .A3(n2343), .A4(n2342), .ZN(n3125)
         );
  INV_X1 U2470 ( .A(n4537), .ZN(n4543) );
  AND2_X1 U2471 ( .A1(n2627), .A2(n3057), .ZN(n4285) );
  AND2_X1 U2472 ( .A1(n2692), .A2(n4409), .ZN(n2751) );
  AND2_X1 U2473 ( .A1(n2835), .A2(n4527), .ZN(n2831) );
  AND2_X1 U2474 ( .A1(n2278), .A2(n2055), .ZN(n2131) );
  INV_X1 U2475 ( .A(n2620), .ZN(n2621) );
  INV_X1 U2476 ( .A(IR_REG_19__SCAN_IN), .ZN(n2519) );
  AND2_X1 U2477 ( .A1(n2201), .A2(n2200), .ZN(n2199) );
  INV_X1 U2478 ( .A(IR_REG_17__SCAN_IN), .ZN(n2200) );
  INV_X1 U2479 ( .A(n2308), .ZN(n2204) );
  NAND2_X1 U2480 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2078)
         );
  AND2_X1 U2481 ( .A1(n2526), .A2(n2512), .ZN(n4052) );
  OAI21_X1 U2482 ( .B1(n3530), .B2(n2098), .A(n2094), .ZN(n3513) );
  OR2_X1 U2483 ( .A1(n2099), .A2(n3501), .ZN(n2098) );
  AOI21_X1 U2484 ( .B1(n2097), .B2(n2096), .A(n2095), .ZN(n2094) );
  NOR2_X1 U2485 ( .A1(n3499), .A2(n3500), .ZN(n2095) );
  NAND2_X1 U2486 ( .A1(n3030), .A2(n3029), .ZN(n3035) );
  INV_X1 U2487 ( .A(n3984), .ZN(n4024) );
  AND2_X1 U2488 ( .A1(n2596), .A2(n2586), .ZN(n3924) );
  INV_X1 U2489 ( .A(n4084), .ZN(n4292) );
  NAND4_X1 U2490 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n4141)
         );
  OR2_X1 U2491 ( .A1(n2610), .A2(n3343), .ZN(n2426) );
  INV_X1 U2492 ( .A(n3279), .ZN(n3815) );
  INV_X1 U2493 ( .A(IR_REG_5__SCAN_IN), .ZN(n2347) );
  NOR2_X1 U2494 ( .A1(n2802), .A2(n2213), .ZN(n2877) );
  AND2_X1 U2495 ( .A1(n2803), .A2(n4415), .ZN(n2213) );
  NAND2_X1 U2496 ( .A1(n4455), .A2(n4456), .ZN(n4454) );
  INV_X1 U2497 ( .A(n2208), .ZN(n3880) );
  NAND2_X1 U2498 ( .A1(n2163), .A2(n4464), .ZN(n2162) );
  NAND2_X1 U2499 ( .A1(n2164), .A2(n4503), .ZN(n2163) );
  AOI21_X1 U2500 ( .B1(n4505), .B2(ADDR_REG_18__SCAN_IN), .A(n4504), .ZN(n2161) );
  NOR2_X1 U2501 ( .A1(n2164), .A2(n4503), .ZN(n4502) );
  NOR2_X1 U2502 ( .A1(n3880), .A2(n3881), .ZN(n4508) );
  NAND2_X1 U2503 ( .A1(n2208), .A2(n2209), .ZN(n4506) );
  INV_X1 U2504 ( .A(n4412), .ZN(n3887) );
  OAI21_X1 U2505 ( .B1(n2207), .B2(n2206), .A(n2205), .ZN(n3884) );
  AOI21_X1 U2506 ( .B1(n2209), .B2(n3852), .A(n2068), .ZN(n2205) );
  AND2_X1 U2507 ( .A1(n4426), .A2(n2785), .ZN(n4507) );
  OR2_X1 U2508 ( .A1(n3370), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2509 ( .A1(n2244), .A2(n2593), .ZN(n3364) );
  NAND2_X1 U2510 ( .A1(n2252), .A2(n2250), .ZN(n2244) );
  AND2_X1 U2511 ( .A1(n2616), .A2(n2615), .ZN(n3507) );
  NAND2_X1 U2512 ( .A1(n2252), .A2(n2583), .ZN(n3911) );
  INV_X1 U2513 ( .A(n3705), .ZN(n2130) );
  INV_X1 U2514 ( .A(IR_REG_14__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U2515 ( .A1(n3376), .A2(n3375), .ZN(n2180) );
  NOR2_X1 U2516 ( .A1(n2399), .A2(n4704), .ZN(n2409) );
  NOR2_X1 U2517 ( .A1(n2457), .A2(n3627), .ZN(n2474) );
  NOR2_X1 U2518 ( .A1(n4482), .A2(n2159), .ZN(n3864) );
  AND2_X1 U2519 ( .A1(n3862), .A2(REG2_REG_15__SCAN_IN), .ZN(n2159) );
  AOI21_X1 U2520 ( .B1(n2127), .B2(n2130), .A(n2126), .ZN(n2125) );
  INV_X1 U2521 ( .A(n3706), .ZN(n2126) );
  NOR2_X1 U2522 ( .A1(n2129), .A2(n2128), .ZN(n2127) );
  INV_X1 U2523 ( .A(n3642), .ZN(n2129) );
  NOR2_X1 U2524 ( .A1(n2130), .A2(n3787), .ZN(n2128) );
  OR2_X1 U2525 ( .A1(n2248), .A2(n2250), .ZN(n2247) );
  INV_X1 U2526 ( .A(n2593), .ZN(n2248) );
  INV_X1 U2527 ( .A(n2606), .ZN(n2249) );
  INV_X1 U2528 ( .A(n3930), .ZN(n3914) );
  AND2_X1 U2529 ( .A1(n2509), .A2(REG3_REG_19__SCAN_IN), .ZN(n2525) );
  INV_X1 U2530 ( .A(n2237), .ZN(n2236) );
  OAI21_X1 U2531 ( .B1(n4091), .B2(n2238), .A(n2499), .ZN(n2237) );
  NAND2_X1 U2532 ( .A1(n2498), .A2(n2497), .ZN(n2499) );
  INV_X1 U2533 ( .A(n2485), .ZN(n2238) );
  NOR2_X1 U2534 ( .A1(n2500), .A2(n3605), .ZN(n2509) );
  AND2_X1 U2535 ( .A1(n4137), .A2(n3727), .ZN(n3685) );
  NAND2_X1 U2536 ( .A1(n3067), .A2(n3648), .ZN(n2112) );
  AND2_X1 U2537 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2336) );
  NAND2_X1 U2538 ( .A1(n2148), .A2(n2147), .ZN(n4040) );
  OR2_X1 U2539 ( .A1(n4111), .A2(n4281), .ZN(n4078) );
  NAND2_X1 U2540 ( .A1(n3264), .A2(n3294), .ZN(n3265) );
  NAND2_X1 U2541 ( .A1(n2464), .A2(n2481), .ZN(n2491) );
  OR3_X1 U2542 ( .A1(n2391), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2394) );
  NOR2_X1 U2543 ( .A1(n2394), .A2(IR_REG_9__SCAN_IN), .ZN(n2418) );
  OAI21_X1 U2544 ( .B1(n3377), .B2(n2179), .A(n2177), .ZN(n2181) );
  INV_X1 U2545 ( .A(n2178), .ZN(n2177) );
  OAI21_X1 U2546 ( .B1(n2179), .B2(n3375), .A(n3584), .ZN(n2178) );
  NAND2_X1 U2547 ( .A1(n3585), .A2(n2180), .ZN(n2179) );
  INV_X1 U2548 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4704) );
  INV_X1 U2549 ( .A(n2099), .ZN(n2096) );
  NOR2_X1 U2550 ( .A1(n3501), .A2(n2101), .ZN(n2097) );
  INV_X1 U2551 ( .A(n2836), .ZN(n2109) );
  NAND2_X1 U2552 ( .A1(n2564), .A2(REG3_REG_24__SCAN_IN), .ZN(n2575) );
  INV_X1 U2553 ( .A(n2566), .ZN(n2564) );
  INV_X1 U2554 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2383) );
  AOI21_X1 U2555 ( .B1(n2190), .B2(n2189), .A(n2067), .ZN(n2188) );
  INV_X1 U2556 ( .A(n3160), .ZN(n2189) );
  OAI21_X1 U2557 ( .B1(n3406), .B2(n2185), .A(n2062), .ZN(n3571) );
  OR2_X1 U2558 ( .A1(n2066), .A2(n3493), .ZN(n2185) );
  NAND2_X1 U2559 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  INV_X1 U2560 ( .A(n3376), .ZN(n2176) );
  OR2_X1 U2561 ( .A1(n3521), .A2(n2058), .ZN(n2198) );
  OR2_X1 U2562 ( .A1(n2448), .A2(n2447), .ZN(n2457) );
  INV_X1 U2563 ( .A(n2828), .ZN(n2858) );
  INV_X1 U2564 ( .A(n3393), .ZN(n2104) );
  INV_X1 U2565 ( .A(n3392), .ZN(n2105) );
  INV_X1 U2566 ( .A(IR_REG_6__SCAN_IN), .ZN(n2370) );
  AND2_X1 U2567 ( .A1(n2085), .A2(n2084), .ZN(n2806) );
  NAND2_X1 U2568 ( .A1(n4416), .A2(REG2_REG_5__SCAN_IN), .ZN(n2084) );
  INV_X1 U2569 ( .A(n2080), .ZN(n2079) );
  NAND2_X1 U2570 ( .A1(n4451), .A2(n3225), .ZN(n3226) );
  AND2_X1 U2571 ( .A1(n2442), .A2(n2444), .ZN(n2493) );
  NAND2_X1 U2572 ( .A1(n3843), .A2(n3844), .ZN(n3845) );
  NAND2_X1 U2573 ( .A1(n2088), .A2(n2087), .ZN(n3859) );
  OR2_X1 U2574 ( .A1(n3856), .A2(REG2_REG_13__SCAN_IN), .ZN(n2087) );
  NAND2_X1 U2575 ( .A1(n4463), .A2(n2050), .ZN(n2088) );
  NOR2_X1 U2576 ( .A1(n4475), .A2(n2451), .ZN(n4474) );
  XNOR2_X1 U2577 ( .A(n3864), .B(n3863), .ZN(n4494) );
  AND2_X1 U2578 ( .A1(n4509), .A2(n3850), .ZN(n2209) );
  INV_X1 U2579 ( .A(n2209), .ZN(n2206) );
  NAND2_X1 U2580 ( .A1(n2125), .A2(n2718), .ZN(n2124) );
  INV_X1 U2581 ( .A(n2119), .ZN(n2118) );
  OAI22_X1 U2582 ( .A1(n2121), .A2(n2120), .B1(n3717), .B2(n2125), .ZN(n2119)
         );
  NOR2_X1 U2583 ( .A1(n2127), .A2(n3717), .ZN(n2120) );
  INV_X1 U2584 ( .A(n2125), .ZN(n2121) );
  AND2_X1 U2585 ( .A1(n2127), .A2(n3717), .ZN(n2122) );
  AND2_X1 U2586 ( .A1(n2143), .A2(n3774), .ZN(n2142) );
  AND2_X1 U2587 ( .A1(n2559), .A2(n2558), .ZN(n3987) );
  OR2_X1 U2588 ( .A1(n3485), .A2(n2610), .ZN(n2559) );
  OAI21_X1 U2589 ( .B1(n4074), .B2(n2044), .A(n3772), .ZN(n4001) );
  NAND2_X1 U2590 ( .A1(n2148), .A2(n2145), .ZN(n4019) );
  OR2_X1 U2591 ( .A1(n2486), .A2(n4681), .ZN(n2500) );
  NAND2_X1 U2592 ( .A1(n2421), .A2(REG3_REG_12__SCAN_IN), .ZN(n2436) );
  AOI21_X1 U2593 ( .B1(n2139), .B2(n2137), .A(n2136), .ZN(n2135) );
  INV_X1 U2594 ( .A(n2139), .ZN(n2138) );
  INV_X1 U2595 ( .A(n3667), .ZN(n2136) );
  AND2_X1 U2596 ( .A1(n3125), .A2(n3036), .ZN(n2351) );
  AND4_X1 U2597 ( .A1(n2369), .A2(n2368), .A3(n2367), .A4(n2366), .ZN(n3279)
         );
  INV_X1 U2598 ( .A(n3015), .ZN(n3020) );
  NAND2_X1 U2599 ( .A1(n2960), .A2(n3654), .ZN(n2976) );
  NAND2_X1 U2600 ( .A1(n2976), .A2(n3735), .ZN(n2975) );
  AND2_X1 U2601 ( .A1(n3658), .A2(n3656), .ZN(n3735) );
  NAND2_X1 U2602 ( .A1(n2867), .A2(n2637), .ZN(n2961) );
  NAND3_X1 U2603 ( .A1(n2110), .A2(n2637), .A3(n3651), .ZN(n2867) );
  NAND2_X1 U2604 ( .A1(n3936), .A2(n3923), .ZN(n3922) );
  AND2_X1 U2605 ( .A1(n3952), .A2(n3937), .ZN(n3936) );
  NAND2_X1 U2606 ( .A1(n4005), .A2(n3994), .ZN(n3993) );
  AND2_X1 U2607 ( .A1(n4031), .A2(n4009), .ZN(n4005) );
  NOR2_X2 U2608 ( .A1(n4049), .A2(n4030), .ZN(n4031) );
  NOR2_X1 U2609 ( .A1(n2560), .A2(n4586), .ZN(n4030) );
  NAND2_X1 U2610 ( .A1(n4079), .A2(n4058), .ZN(n4057) );
  OR2_X1 U2611 ( .A1(n4126), .A2(n2467), .ZN(n4111) );
  NAND2_X1 U2612 ( .A1(n4148), .A2(n4300), .ZN(n4126) );
  INV_X1 U2613 ( .A(n4127), .ZN(n4300) );
  AND4_X1 U2614 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n4317)
         );
  OR2_X1 U2615 ( .A1(n2610), .A2(n4165), .ZN(n2414) );
  INV_X1 U2616 ( .A(n3124), .ZN(n3119) );
  INV_X1 U2617 ( .A(n4325), .ZN(n4546) );
  AND2_X1 U2618 ( .A1(n4419), .A2(n2759), .ZN(n4291) );
  INV_X1 U2619 ( .A(n4304), .ZN(n4329) );
  INV_X1 U2620 ( .A(n4291), .ZN(n4316) );
  AND2_X1 U2621 ( .A1(n2057), .A2(n2278), .ZN(n2254) );
  AND2_X1 U2622 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2292)
         );
  NAND2_X1 U2623 ( .A1(n2047), .A2(n2291), .ZN(n2726) );
  INV_X1 U2624 ( .A(IR_REG_20__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U2625 ( .A1(n2617), .A2(IR_REG_31__SCAN_IN), .ZN(n2619) );
  AND2_X1 U2626 ( .A1(n2333), .A2(n2321), .ZN(n3832) );
  AND4_X1 U2627 ( .A1(n2357), .A2(n2356), .A3(n2355), .A4(n2354), .ZN(n3172)
         );
  OR2_X1 U2628 ( .A1(n2610), .A2(n3130), .ZN(n2355) );
  AOI21_X1 U2629 ( .B1(n3530), .B2(n2101), .A(n2099), .ZN(n2093) );
  NAND2_X1 U2630 ( .A1(n2196), .A2(n2194), .ZN(n3481) );
  AND2_X1 U2631 ( .A1(n2195), .A2(n3440), .ZN(n2194) );
  AND2_X1 U2632 ( .A1(n3483), .A2(n3484), .ZN(n3440) );
  INV_X1 U2633 ( .A(n3244), .ZN(n3245) );
  NOR2_X1 U2634 ( .A1(n3406), .A2(n2066), .ZN(n2182) );
  NAND2_X1 U2635 ( .A1(n3159), .A2(n3160), .ZN(n2193) );
  INV_X1 U2636 ( .A(DATAI_1_), .ZN(n2157) );
  NAND2_X1 U2637 ( .A1(n2853), .A2(n2852), .ZN(n2855) );
  AND2_X1 U2638 ( .A1(n2549), .A2(n2548), .ZN(n4258) );
  AND3_X1 U2639 ( .A1(n2504), .A2(n2503), .A3(n2502), .ZN(n4277) );
  NAND3_X1 U2640 ( .A1(n2170), .A2(n2171), .A3(n2996), .ZN(n3030) );
  INV_X1 U2641 ( .A(n3251), .ZN(n3195) );
  AND2_X1 U2642 ( .A1(n2198), .A2(n3433), .ZN(n3593) );
  AND4_X1 U2643 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n4330)
         );
  NAND2_X1 U2644 ( .A1(n2898), .A2(n2899), .ZN(n2946) );
  INV_X1 U2645 ( .A(n4060), .ZN(n4058) );
  INV_X1 U2646 ( .A(n3634), .ZN(n3618) );
  AND4_X1 U2647 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n4295)
         );
  INV_X1 U2648 ( .A(n3617), .ZN(n3629) );
  INV_X1 U2649 ( .A(n3582), .ZN(n3625) );
  INV_X1 U2650 ( .A(n3578), .ZN(n3631) );
  NAND2_X1 U2651 ( .A1(n2603), .A2(n2602), .ZN(n3919) );
  NAND2_X1 U2652 ( .A1(n2581), .A2(n2580), .ZN(n3809) );
  INV_X1 U2653 ( .A(n3486), .ZN(n4228) );
  INV_X1 U2654 ( .A(n3987), .ZN(n4237) );
  INV_X1 U2655 ( .A(n4258), .ZN(n3810) );
  NAND2_X1 U2656 ( .A1(n2538), .A2(n2537), .ZN(n3984) );
  OR2_X1 U2657 ( .A1(n3576), .A2(n2610), .ZN(n2532) );
  NAND2_X1 U2658 ( .A1(n2517), .A2(n2516), .ZN(n4022) );
  INV_X1 U2659 ( .A(n4277), .ZN(n3811) );
  NAND4_X1 U2660 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .ZN(n3813)
         );
  OR2_X1 U2661 ( .A1(n2610), .A2(n3197), .ZN(n2389) );
  NAND4_X1 U2662 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3814)
         );
  NAND3_X1 U2663 ( .A1(n2332), .A2(n2331), .A3(n2330), .ZN(n3818) );
  OR2_X1 U2664 ( .A1(n2488), .A2(n2324), .ZN(n2332) );
  OR2_X1 U2665 ( .A1(n3639), .A2(n2982), .ZN(n2318) );
  NOR2_X1 U2666 ( .A1(n2914), .A2(n2913), .ZN(n2912) );
  AOI21_X1 U2667 ( .B1(n2926), .B2(REG2_REG_4__SCAN_IN), .A(n2083), .ZN(n2772)
         );
  XNOR2_X1 U2668 ( .A(n2806), .B(n4415), .ZN(n2808) );
  INV_X1 U2669 ( .A(n2879), .ZN(n3220) );
  NAND2_X1 U2670 ( .A1(n4442), .A2(n3208), .ZN(n4455) );
  XNOR2_X1 U2671 ( .A(n3226), .B(n2167), .ZN(n4470) );
  NAND2_X1 U2672 ( .A1(n4463), .A2(n3211), .ZN(n3858) );
  XNOR2_X1 U2673 ( .A(n3845), .B(n4531), .ZN(n4479) );
  NAND2_X1 U2674 ( .A1(n2090), .A2(n4464), .ZN(n3867) );
  NAND2_X1 U2675 ( .A1(n3369), .A2(n3705), .ZN(n2720) );
  AND2_X1 U2676 ( .A1(n2591), .A2(n2590), .ZN(n4231) );
  NOR2_X1 U2677 ( .A1(n3992), .A2(n2229), .ZN(n2228) );
  INV_X1 U2678 ( .A(n2231), .ZN(n2229) );
  NAND2_X1 U2679 ( .A1(n4090), .A2(n2485), .ZN(n4076) );
  OAI21_X1 U2680 ( .B1(n3338), .B2(n2222), .A(n2218), .ZN(n4123) );
  NAND2_X1 U2681 ( .A1(n2217), .A2(n2221), .ZN(n4125) );
  NAND2_X1 U2682 ( .A1(n3338), .A2(n2224), .ZN(n2217) );
  INV_X1 U2683 ( .A(n2433), .ZN(n2225) );
  NAND2_X1 U2684 ( .A1(n3338), .A2(n2434), .ZN(n2226) );
  INV_X1 U2685 ( .A(n3813), .ZN(n3272) );
  INV_X1 U2686 ( .A(n4196), .ZN(n4519) );
  NOR2_X1 U2687 ( .A1(n4547), .A2(n2262), .ZN(n3276) );
  OAI21_X1 U2688 ( .B1(n3068), .B2(n3067), .A(n3648), .ZN(n2113) );
  INV_X1 U2689 ( .A(n3036), .ZN(n3102) );
  INV_X1 U2690 ( .A(n3172), .ZN(n3816) );
  INV_X1 U2691 ( .A(n4105), .ZN(n4153) );
  AND2_X1 U2692 ( .A1(n4516), .A2(n4304), .ZN(n4190) );
  NAND2_X1 U2693 ( .A1(n4543), .A2(n2832), .ZN(n4513) );
  NAND2_X1 U2694 ( .A1(n2730), .A2(n2150), .ZN(n2149) );
  AOI21_X1 U2695 ( .B1(n4216), .B2(n4304), .A(n2729), .ZN(n2150) );
  OAI21_X1 U2696 ( .B1(n3365), .B2(n3515), .A(n2705), .ZN(n3353) );
  AND2_X1 U2697 ( .A1(n2674), .A2(n2673), .ZN(n2741) );
  NAND2_X1 U2698 ( .A1(n2680), .A2(IR_REG_31__SCAN_IN), .ZN(n2668) );
  AND2_X1 U2699 ( .A1(n2758), .A2(STATE_REG_SCAN_IN), .ZN(n4527) );
  AND2_X1 U2700 ( .A1(n2617), .A2(n2521), .ZN(n4412) );
  NAND2_X1 U2701 ( .A1(n2442), .A2(n2201), .ZN(n2495) );
  INV_X1 U2702 ( .A(n3862), .ZN(n4530) );
  NAND2_X1 U2703 ( .A1(n2203), .A2(n2202), .ZN(n2311) );
  NAND2_X1 U2704 ( .A1(n2748), .A2(n2265), .ZN(n2202) );
  INV_X1 U2705 ( .A(n2160), .ZN(n4511) );
  OAI21_X1 U2706 ( .B1(n4502), .B2(n2162), .A(n2161), .ZN(n2160) );
  NAND2_X1 U2707 ( .A1(n2153), .A2(n2152), .ZN(U3351) );
  NAND2_X1 U2708 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2152) );
  OR2_X1 U2709 ( .A1(U3149), .A2(n2154), .ZN(n2153) );
  INV_X1 U2710 ( .A(n2300), .ZN(n2846) );
  AND2_X1 U2711 ( .A1(n2290), .A2(n2289), .ZN(n2042) );
  INV_X1 U2712 ( .A(n2222), .ZN(n2221) );
  NOR2_X1 U2713 ( .A1(n2043), .A2(n2223), .ZN(n2222) );
  INV_X1 U2714 ( .A(n2262), .ZN(n2242) );
  NOR2_X1 U2715 ( .A1(n2433), .A2(n2065), .ZN(n2043) );
  INV_X1 U2716 ( .A(n4282), .ZN(n2498) );
  NAND2_X1 U2717 ( .A1(n2105), .A2(n2104), .ZN(n3540) );
  NAND2_X1 U2718 ( .A1(n2652), .A2(n2145), .ZN(n2044) );
  NAND2_X1 U2719 ( .A1(n2859), .A2(n3058), .ZN(n3055) );
  INV_X1 U2720 ( .A(n3055), .ZN(n2110) );
  NOR2_X1 U2721 ( .A1(n4255), .A2(n4030), .ZN(n2045) );
  NAND2_X1 U2722 ( .A1(n2076), .A2(n3245), .ZN(n3307) );
  INV_X1 U2723 ( .A(n3852), .ZN(n2210) );
  INV_X1 U2724 ( .A(n2560), .ZN(n2539) );
  XNOR2_X1 U2725 ( .A(n2078), .B(IR_REG_1__SCAN_IN), .ZN(n2158) );
  XNOR2_X1 U2726 ( .A(n2619), .B(n2618), .ZN(n2627) );
  NAND2_X1 U2727 ( .A1(n2308), .A2(n2265), .ZN(n2309) );
  OR2_X1 U2728 ( .A1(n4408), .A2(n2746), .ZN(n2302) );
  INV_X1 U2729 ( .A(n2191), .ZN(n2190) );
  OR2_X1 U2730 ( .A1(n3181), .A2(n2192), .ZN(n2191) );
  OR2_X1 U2731 ( .A1(n2673), .A2(IR_REG_26__SCAN_IN), .ZN(n2046) );
  NOR2_X1 U2732 ( .A1(n2182), .A2(n3602), .ZN(n3492) );
  NAND4_X1 U2733 ( .A1(n2134), .A2(n2133), .A3(n2276), .A4(n2131), .ZN(n2047)
         );
  OAI21_X1 U2734 ( .B1(n4016), .B2(n2045), .A(n2533), .ZN(n4003) );
  NAND2_X1 U2735 ( .A1(n2746), .A2(n2284), .ZN(n2303) );
  INV_X1 U2736 ( .A(n2093), .ZN(n3502) );
  AND2_X1 U2737 ( .A1(n2898), .A2(n2986), .ZN(n2048) );
  NAND2_X1 U2738 ( .A1(n2230), .A2(n2231), .ZN(n3991) );
  AND2_X1 U2739 ( .A1(n2990), .A2(n2989), .ZN(n2049) );
  AND2_X1 U2740 ( .A1(n3211), .A2(n2089), .ZN(n2050) );
  AND2_X1 U2741 ( .A1(n3814), .A2(n3287), .ZN(n2051) );
  AND2_X1 U2742 ( .A1(n3239), .A2(n3238), .ZN(n2052) );
  INV_X1 U2743 ( .A(IR_REG_21__SCAN_IN), .ZN(n2623) );
  AND2_X1 U2744 ( .A1(n2249), .A2(n2593), .ZN(n2053) );
  NAND2_X1 U2745 ( .A1(n2198), .A2(n2197), .ZN(n3482) );
  INV_X1 U2746 ( .A(IR_REG_28__SCAN_IN), .ZN(n2255) );
  AND2_X1 U2747 ( .A1(n2891), .A2(n2890), .ZN(n2054) );
  NAND2_X1 U2748 ( .A1(n2075), .A2(n2308), .ZN(n2346) );
  INV_X1 U2749 ( .A(n2346), .ZN(n2134) );
  AND2_X1 U2750 ( .A1(n2279), .A2(n2256), .ZN(n2055) );
  AND2_X1 U2751 ( .A1(n2112), .A2(n3661), .ZN(n2056) );
  AND2_X1 U2752 ( .A1(n2055), .A2(n2255), .ZN(n2057) );
  INV_X1 U2753 ( .A(IR_REG_31__SCAN_IN), .ZN(n2748) );
  XNOR2_X1 U2754 ( .A(n2668), .B(IR_REG_24__SCAN_IN), .ZN(n2690) );
  INV_X1 U2755 ( .A(n3717), .ZN(n2718) );
  XNOR2_X1 U2756 ( .A(n2406), .B(IR_REG_10__SCAN_IN), .ZN(n3222) );
  AND2_X1 U2757 ( .A1(n3523), .A2(n3522), .ZN(n2058) );
  NAND2_X1 U2758 ( .A1(n3321), .A2(n3320), .ZN(n3377) );
  NAND2_X1 U2759 ( .A1(n2072), .A2(n2181), .ZN(n3471) );
  NAND2_X1 U2760 ( .A1(n4092), .A2(n4091), .ZN(n4090) );
  NAND2_X1 U2761 ( .A1(n2300), .A2(n4198), .ZN(n3651) );
  AND2_X1 U2762 ( .A1(n4024), .A2(n4009), .ZN(n2059) );
  INV_X1 U2763 ( .A(n3726), .ZN(n2147) );
  NAND2_X1 U2764 ( .A1(n3683), .A2(n3646), .ZN(n4124) );
  INV_X1 U2765 ( .A(n4124), .ZN(n2219) );
  AND2_X1 U2766 ( .A1(n4295), .A2(n4300), .ZN(n2060) );
  AND2_X1 U2767 ( .A1(n4282), .A2(n4274), .ZN(n2061) );
  AND2_X1 U2768 ( .A1(n2183), .A2(n3420), .ZN(n2062) );
  AND2_X1 U2769 ( .A1(n3553), .A2(n3403), .ZN(n2063) );
  AND2_X1 U2770 ( .A1(n2226), .A2(n2225), .ZN(n2064) );
  AND2_X1 U2771 ( .A1(n4317), .A2(n4145), .ZN(n2065) );
  NAND2_X1 U2772 ( .A1(n2946), .A2(n2945), .ZN(n2987) );
  INV_X1 U2773 ( .A(n3375), .ZN(n2174) );
  NAND2_X1 U2774 ( .A1(n3135), .A2(n3134), .ZN(n3159) );
  OAI21_X1 U2775 ( .B1(n3159), .B2(n2191), .A(n2188), .ZN(n3236) );
  NAND2_X1 U2776 ( .A1(n2193), .A2(n3142), .ZN(n3182) );
  OAI21_X1 U2777 ( .B1(n3159), .B2(n2108), .A(n2106), .ZN(n3243) );
  AND2_X1 U2778 ( .A1(n3410), .A2(n3409), .ZN(n2066) );
  AND2_X1 U2779 ( .A1(n4426), .A2(n3801), .ZN(n4464) );
  AND2_X1 U2780 ( .A1(n3149), .A2(n3148), .ZN(n2067) );
  INV_X1 U2781 ( .A(n4462), .ZN(n2167) );
  NOR2_X1 U2782 ( .A1(n4528), .A2(n3882), .ZN(n2068) );
  OR2_X1 U2783 ( .A1(n3922), .A2(n4213), .ZN(n2704) );
  NAND2_X1 U2784 ( .A1(n2899), .A2(n2048), .ZN(n2170) );
  NAND3_X1 U2785 ( .A1(n2072), .A2(n2181), .A3(n2071), .ZN(n2073) );
  NAND2_X1 U2786 ( .A1(n2092), .A2(n2176), .ZN(n2175) );
  NAND3_X1 U2787 ( .A1(n2276), .A2(n2074), .A3(n2134), .ZN(n2665) );
  NOR2_X2 U2788 ( .A1(n2346), .A2(n2271), .ZN(n2442) );
  NAND4_X1 U2789 ( .A1(n2267), .A2(n2270), .A3(n2269), .A4(n2268), .ZN(n2271)
         );
  INV_X1 U2790 ( .A(n3243), .ZN(n2076) );
  OAI21_X1 U2791 ( .B1(n3530), .B2(n3531), .A(n3532), .ZN(n3613) );
  AOI21_X2 U2792 ( .B1(n3560), .B2(n3563), .A(n3562), .ZN(n3530) );
  OAI21_X1 U2793 ( .B1(n2158), .B2(REG2_REG_1__SCAN_IN), .A(n2077), .ZN(n2765)
         );
  NAND2_X1 U2794 ( .A1(n2158), .A2(REG2_REG_1__SCAN_IN), .ZN(n2077) );
  INV_X1 U2795 ( .A(n2085), .ZN(n2790) );
  NAND2_X1 U2796 ( .A1(n2768), .A2(n4417), .ZN(n2086) );
  OAI21_X1 U2797 ( .B1(n3866), .B2(n2091), .A(n3875), .ZN(n2090) );
  XNOR2_X1 U2798 ( .A(n2944), .B(n2054), .ZN(n2897) );
  XNOR2_X1 U2799 ( .A(n2889), .B(n3451), .ZN(n2944) );
  INV_X1 U2800 ( .A(n3377), .ZN(n2092) );
  NAND2_X1 U2801 ( .A1(n2103), .A2(n3400), .ZN(n3550) );
  NAND3_X1 U2802 ( .A1(n2169), .A2(n3395), .A3(n3540), .ZN(n2103) );
  NAND2_X1 U2803 ( .A1(n2171), .A2(n2170), .ZN(n2994) );
  INV_X1 U2804 ( .A(n2835), .ZN(n2947) );
  NAND2_X1 U2805 ( .A1(n3746), .A2(n2961), .ZN(n2960) );
  NAND2_X1 U2806 ( .A1(n3068), .A2(n3648), .ZN(n2111) );
  NAND2_X1 U2807 ( .A1(n2111), .A2(n2056), .ZN(n2641) );
  XNOR2_X1 U2808 ( .A(n2113), .B(n3733), .ZN(n3090) );
  NAND2_X1 U2809 ( .A1(n2975), .A2(n3658), .ZN(n2116) );
  INV_X1 U2810 ( .A(n3658), .ZN(n2115) );
  XNOR2_X1 U2811 ( .A(n2116), .B(n3745), .ZN(n3019) );
  NAND2_X1 U2812 ( .A1(n2123), .A2(n2117), .ZN(n2728) );
  AOI21_X1 U2813 ( .B1(n3370), .B2(n2122), .A(n2118), .ZN(n2117) );
  NAND3_X1 U2814 ( .A1(n2132), .A2(n2134), .A3(n2276), .ZN(n2673) );
  OAI21_X1 U2815 ( .B1(n3169), .B2(n2138), .A(n2135), .ZN(n3193) );
  OAI21_X1 U2816 ( .B1(n3169), .B2(n2643), .A(n3668), .ZN(n3277) );
  AOI21_X1 U2817 ( .B1(n2643), .B2(n3668), .A(n2140), .ZN(n2139) );
  NAND2_X1 U2818 ( .A1(n2141), .A2(n2142), .ZN(n2656) );
  NAND2_X1 U2819 ( .A1(n4074), .A2(n2144), .ZN(n2141) );
  NAND2_X1 U2820 ( .A1(n2647), .A2(n3683), .ZN(n4106) );
  NAND2_X1 U2821 ( .A1(n2649), .A2(n2648), .ZN(n4107) );
  NAND2_X1 U2822 ( .A1(n2641), .A2(n3665), .ZN(n3169) );
  NAND2_X1 U2823 ( .A1(n4101), .A2(n4100), .ZN(n4099) );
  NAND2_X1 U2824 ( .A1(n2646), .A2(n3681), .ZN(n3764) );
  NAND2_X1 U2825 ( .A1(n4107), .A2(n3647), .ZN(n4101) );
  NAND2_X1 U2826 ( .A1(n4099), .A2(n3767), .ZN(n4074) );
  CLKBUF_X1 U2827 ( .A(n2158), .Z(n2151) );
  NAND2_X1 U2828 ( .A1(n2151), .A2(REG1_REG_1__SCAN_IN), .ZN(n2778) );
  INV_X1 U2829 ( .A(n2151), .ZN(n2154) );
  XNOR2_X1 U2830 ( .A(n2158), .B(n2777), .ZN(n3822) );
  MUX2_X1 U2831 ( .A(REG2_REG_1__SCAN_IN), .B(n2763), .S(n2151), .Z(n3826) );
  NOR2_X1 U2832 ( .A1(n3824), .A2(n2155), .ZN(n2914) );
  AND2_X1 U2833 ( .A1(n2158), .A2(REG2_REG_1__SCAN_IN), .ZN(n2155) );
  NAND2_X1 U2834 ( .A1(n2041), .A2(n2151), .ZN(n2156) );
  NAND2_X1 U2835 ( .A1(n3833), .A2(n2151), .ZN(n3831) );
  OAI21_X1 U2836 ( .B1(n2840), .B2(n2168), .A(n2853), .ZN(n2909) );
  NAND2_X1 U2837 ( .A1(n3541), .A2(n3623), .ZN(n2169) );
  NAND2_X1 U2838 ( .A1(n3392), .A2(n3393), .ZN(n3541) );
  AOI21_X1 U2839 ( .B1(n2986), .B2(n2172), .A(n2049), .ZN(n2171) );
  NAND2_X1 U2840 ( .A1(n2175), .A2(n3375), .ZN(n3587) );
  INV_X1 U2841 ( .A(n3406), .ZN(n3601) );
  NAND2_X1 U2842 ( .A1(n3571), .A2(n3572), .ZN(n3570) );
  NAND2_X1 U2843 ( .A1(n3521), .A2(n2197), .ZN(n2196) );
  NAND2_X1 U2844 ( .A1(n2442), .A2(n2199), .ZN(n2518) );
  NAND3_X1 U2845 ( .A1(n2204), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2203) );
  INV_X1 U2846 ( .A(n3853), .ZN(n2207) );
  NAND2_X1 U2847 ( .A1(n4408), .A2(n2214), .ZN(n2314) );
  NAND3_X1 U2848 ( .A1(n2214), .A2(n4408), .A3(REG2_REG_1__SCAN_IN), .ZN(n2289) );
  XNOR2_X2 U2849 ( .A(n2283), .B(IR_REG_30__SCAN_IN), .ZN(n4408) );
  NAND2_X2 U2850 ( .A1(n2042), .A2(n2039), .ZN(n2300) );
  NAND3_X1 U2851 ( .A1(n2042), .A2(n2039), .A3(n2872), .ZN(n2637) );
  NAND2_X1 U2852 ( .A1(n3338), .A2(n2218), .ZN(n2216) );
  NAND2_X1 U2853 ( .A1(n2230), .A2(n2228), .ZN(n3990) );
  NAND2_X1 U2854 ( .A1(n2234), .A2(n2235), .ZN(n4066) );
  NAND2_X1 U2855 ( .A1(n4092), .A2(n2236), .ZN(n2234) );
  OAI21_X1 U2856 ( .B1(n3934), .B2(n2243), .A(n2245), .ZN(n2714) );
  INV_X1 U2857 ( .A(n2584), .ZN(n2253) );
  OR2_X1 U2858 ( .A1(n2314), .A2(n3062), .ZN(n2297) );
  AOI21_X2 U2859 ( .B1(n2974), .B2(n2323), .A(n2322), .ZN(n3004) );
  NAND2_X1 U2860 ( .A1(n2746), .A2(n4408), .ZN(n2450) );
  INV_X1 U2861 ( .A(n3814), .ZN(n3254) );
  OR2_X1 U2862 ( .A1(n4559), .A2(REG1_REG_29__SCAN_IN), .ZN(n2257) );
  INV_X1 U2863 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U2864 ( .A1(n3817), .A2(n3102), .ZN(n2350) );
  NOR2_X1 U2865 ( .A1(n2610), .A2(n3022), .ZN(n2258) );
  OR2_X1 U2866 ( .A1(n4553), .A2(REG0_REG_29__SCAN_IN), .ZN(n2259) );
  INV_X1 U2867 ( .A(n4318), .ZN(n3812) );
  AND4_X1 U2868 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n4318)
         );
  AND4_X1 U2869 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n4301)
         );
  INV_X1 U2870 ( .A(n4301), .ZN(n2468) );
  AND2_X1 U2871 ( .A1(n3272), .A2(n3195), .ZN(n2396) );
  INV_X1 U2872 ( .A(n3780), .ZN(n2660) );
  OR2_X1 U2873 ( .A1(n3905), .A2(n4336), .ZN(n2260) );
  OR2_X1 U2874 ( .A1(n3905), .A2(n4406), .ZN(n2261) );
  AND2_X1 U2875 ( .A1(n3815), .A2(n3170), .ZN(n2262) );
  AND2_X1 U2876 ( .A1(n4301), .A2(n4118), .ZN(n2263) );
  INV_X1 U2877 ( .A(n4109), .ZN(n2648) );
  INV_X1 U2878 ( .A(n4118), .ZN(n2467) );
  NAND2_X1 U2879 ( .A1(n2956), .A2(n2313), .ZN(n2974) );
  AND2_X1 U2880 ( .A1(n3813), .A2(n3251), .ZN(n2264) );
  AND2_X1 U2881 ( .A1(n3770), .A2(n3767), .ZN(n4100) );
  INV_X1 U2882 ( .A(IR_REG_4__SCAN_IN), .ZN(n2266) );
  INV_X1 U2883 ( .A(n3543), .ZN(n3395) );
  NAND2_X1 U2884 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  INV_X1 U2885 ( .A(n4274), .ZN(n2497) );
  NAND2_X1 U2886 ( .A1(n3404), .A2(n3552), .ZN(n3405) );
  INV_X1 U2887 ( .A(n3703), .ZN(n2659) );
  INV_X1 U2888 ( .A(IR_REG_2__SCAN_IN), .ZN(n2265) );
  INV_X1 U2889 ( .A(n2553), .ZN(n2552) );
  OR2_X1 U2890 ( .A1(n2859), .A2(n3506), .ZN(n2839) );
  INV_X1 U2891 ( .A(n2596), .ZN(n2594) );
  NAND2_X1 U2892 ( .A1(n2285), .A2(REG0_REG_1__SCAN_IN), .ZN(n2286) );
  INV_X1 U2893 ( .A(n3992), .ZN(n2550) );
  NAND2_X1 U2894 ( .A1(n3654), .A2(n3650), .ZN(n2638) );
  NAND2_X1 U2895 ( .A1(n2552), .A2(REG3_REG_23__SCAN_IN), .ZN(n2566) );
  INV_X1 U2896 ( .A(n3506), .ZN(n3464) );
  OR2_X1 U2897 ( .A1(n2575), .A2(n4684), .ZN(n2585) );
  NAND2_X1 U2898 ( .A1(n2474), .A2(REG3_REG_16__SCAN_IN), .ZN(n2486) );
  OR2_X1 U2899 ( .A1(n4237), .A2(n3975), .ZN(n3723) );
  NAND2_X1 U2900 ( .A1(n4318), .A2(n4168), .ZN(n2420) );
  NAND2_X1 U2901 ( .A1(n3818), .A2(n3020), .ZN(n3663) );
  INV_X1 U2902 ( .A(n2638), .ZN(n3746) );
  AND2_X1 U2903 ( .A1(n3151), .A2(n3150), .ZN(n3181) );
  INV_X1 U2904 ( .A(n3550), .ZN(n3551) );
  INV_X1 U2905 ( .A(n2995), .ZN(n2996) );
  INV_X1 U2906 ( .A(n4022), .ZN(n4062) );
  AND2_X1 U2907 ( .A1(n2409), .A2(REG3_REG_11__SCAN_IN), .ZN(n2421) );
  AND2_X1 U2908 ( .A1(n2833), .A2(n4513), .ZN(n3628) );
  OR2_X1 U2909 ( .A1(n3516), .A2(n2610), .ZN(n2616) );
  OR2_X1 U2910 ( .A1(n2610), .A2(n3175), .ZN(n2367) );
  INV_X1 U2911 ( .A(n4323), .ZN(n4290) );
  AND2_X1 U2912 ( .A1(n3968), .A2(n2654), .ZN(n3992) );
  NAND2_X1 U2913 ( .A1(n3659), .A2(n3663), .ZN(n3745) );
  AND2_X1 U2914 ( .A1(n2662), .A2(n2661), .ZN(n4306) );
  OR2_X1 U2915 ( .A1(n3056), .A2(n4410), .ZN(n4537) );
  NOR2_X1 U2916 ( .A1(n2395), .A2(n2418), .ZN(n3215) );
  NOR2_X1 U2917 ( .A1(n2363), .A2(n2362), .ZN(n2372) );
  OR2_X1 U2918 ( .A1(n2384), .A2(n2383), .ZN(n2399) );
  OR2_X1 U2919 ( .A1(n2436), .A2(n2435), .ZN(n2448) );
  NAND2_X1 U2920 ( .A1(n2896), .A2(n2895), .ZN(n2901) );
  AND2_X1 U2921 ( .A1(n2858), .A2(n2857), .ZN(n3617) );
  OR2_X1 U2922 ( .A1(n3939), .A2(n2610), .ZN(n2581) );
  AND3_X1 U2923 ( .A1(n2480), .A2(n2479), .A3(n2478), .ZN(n4084) );
  AND2_X1 U2924 ( .A1(n2770), .A2(n2769), .ZN(n4426) );
  NAND2_X1 U2925 ( .A1(n4028), .A2(n4537), .ZN(n4325) );
  AND3_X1 U2926 ( .A1(n2697), .A2(n2816), .A3(n2696), .ZN(n2708) );
  INV_X1 U2927 ( .A(n2830), .ZN(n3795) );
  XNOR2_X1 U2928 ( .A(n2432), .B(IR_REG_12__SCAN_IN), .ZN(n4462) );
  INV_X1 U2929 ( .A(n3832), .ZN(n2780) );
  AND2_X1 U2930 ( .A1(n2770), .A2(n2761), .ZN(n4505) );
  NAND2_X1 U2931 ( .A1(n2858), .A2(n2842), .ZN(n3582) );
  AND2_X1 U2932 ( .A1(n2951), .A2(n2950), .ZN(n3634) );
  INV_X1 U2933 ( .A(n3507), .ZN(n4216) );
  NAND2_X1 U2934 ( .A1(n2532), .A2(n2531), .ZN(n4255) );
  INV_X1 U2935 ( .A(n4317), .ZN(n4303) );
  INV_X1 U2936 ( .A(n3125), .ZN(n3817) );
  OR2_X1 U2937 ( .A1(n4336), .A2(n3353), .ZN(n2706) );
  NAND2_X1 U2938 ( .A1(n4559), .A2(n4285), .ZN(n4336) );
  NAND2_X1 U2939 ( .A1(n2708), .A2(n2818), .ZN(n4557) );
  OR2_X1 U2940 ( .A1(n3353), .A2(n4406), .ZN(n2711) );
  NAND2_X1 U2941 ( .A1(n4553), .A2(n4285), .ZN(n4406) );
  INV_X1 U2942 ( .A(n4553), .ZN(n4551) );
  INV_X1 U2943 ( .A(n3222), .ZN(n4534) );
  NOR2_X2 U2944 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2270)
         );
  NOR2_X2 U2945 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2269)
         );
  NOR2_X2 U2946 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2268)
         );
  INV_X1 U2947 ( .A(n2491), .ZN(n2275) );
  INV_X1 U2948 ( .A(IR_REG_29__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2949 ( .A1(n2282), .A2(n2281), .ZN(n2749) );
  INV_X1 U2950 ( .A(n4408), .ZN(n2284) );
  OR2_X1 U2951 ( .A1(n2303), .A2(n2777), .ZN(n2287) );
  INV_X1 U2952 ( .A(n2302), .ZN(n2285) );
  INV_X1 U2953 ( .A(n2450), .ZN(n2288) );
  NAND2_X1 U2954 ( .A1(n2288), .A2(REG3_REG_1__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2955 ( .A1(n2279), .A2(n2748), .ZN(n2291) );
  NAND2_X2 U2956 ( .A1(n2725), .A2(IR_REG_28__SCAN_IN), .ZN(n2293) );
  INV_X1 U2957 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3061) );
  OR2_X1 U2958 ( .A1(n2450), .A2(n3061), .ZN(n2299) );
  INV_X1 U2959 ( .A(n2303), .ZN(n2477) );
  NAND2_X1 U2960 ( .A1(n2477), .A2(REG1_REG_0__SCAN_IN), .ZN(n2298) );
  INV_X1 U2961 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3062) );
  INV_X1 U2962 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2295) );
  OR2_X1 U2963 ( .A1(n2302), .A2(n2295), .ZN(n2296) );
  NAND4_X1 U2964 ( .A1(n2299), .A2(n2298), .A3(n2297), .A4(n2296), .ZN(n2834)
         );
  INV_X1 U2965 ( .A(n2834), .ZN(n2859) );
  MUX2_X1 U2966 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2041), .Z(n3058) );
  INV_X2 U2967 ( .A(n3058), .ZN(n3054) );
  NOR2_X1 U2968 ( .A1(n2859), .A2(n3054), .ZN(n2864) );
  NAND2_X1 U2969 ( .A1(n2636), .A2(n2864), .ZN(n2866) );
  NAND2_X1 U2970 ( .A1(n2300), .A2(n2872), .ZN(n2301) );
  NAND2_X1 U2971 ( .A1(n2866), .A2(n2301), .ZN(n2957) );
  INV_X1 U2972 ( .A(n2957), .ZN(n2312) );
  NAND2_X1 U2973 ( .A1(n2285), .A2(REG0_REG_2__SCAN_IN), .ZN(n2307) );
  INV_X1 U2974 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2776) );
  OR2_X1 U2975 ( .A1(n2303), .A2(n2776), .ZN(n2306) );
  INV_X1 U2976 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2919) );
  OR2_X1 U2977 ( .A1(n2450), .A2(n2919), .ZN(n2305) );
  INV_X1 U2978 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4177) );
  OR2_X1 U2979 ( .A1(n2314), .A2(n4177), .ZN(n2304) );
  NAND4_X1 U2980 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n2977)
         );
  INV_X1 U2981 ( .A(n2309), .ZN(n2310) );
  NOR2_X2 U2982 ( .A1(n2311), .A2(n2310), .ZN(n4418) );
  MUX2_X1 U2983 ( .A(DATAI_2_), .B(n4418), .S(n2041), .Z(n4181) );
  NAND2_X1 U2984 ( .A1(n2888), .A2(n4181), .ZN(n3654) );
  INV_X2 U2985 ( .A(n4181), .ZN(n2967) );
  NAND2_X1 U2986 ( .A1(n2977), .A2(n2967), .ZN(n3650) );
  NAND2_X1 U2987 ( .A1(n2312), .A2(n2638), .ZN(n2956) );
  NAND2_X1 U2988 ( .A1(n2888), .A2(n2967), .ZN(n2313) );
  INV_X1 U2989 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2982) );
  OR2_X1 U2990 ( .A1(n2610), .A2(REG3_REG_3__SCAN_IN), .ZN(n2317) );
  NAND2_X1 U2991 ( .A1(n3636), .A2(REG0_REG_3__SCAN_IN), .ZN(n2316) );
  INV_X1 U2992 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2767) );
  OR2_X1 U2993 ( .A1(n2314), .A2(n2767), .ZN(n2315) );
  NAND2_X1 U2994 ( .A1(n2309), .A2(IR_REG_31__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2995 ( .A1(n2320), .A2(n2319), .ZN(n2333) );
  OR2_X1 U2996 ( .A1(n2320), .A2(n2319), .ZN(n2321) );
  NAND2_X1 U2997 ( .A1(n4183), .A2(n3045), .ZN(n2323) );
  NOR2_X1 U2998 ( .A1(n4183), .A2(n3045), .ZN(n2322) );
  INV_X1 U2999 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2324) );
  INV_X1 U3000 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2325) );
  OR2_X1 U3001 ( .A1(n3639), .A2(n2325), .ZN(n2331) );
  INV_X1 U3002 ( .A(n2336), .ZN(n2338) );
  INV_X1 U3003 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3046) );
  INV_X1 U3004 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U3005 ( .A1(n3046), .A2(n2326), .ZN(n2327) );
  NAND2_X1 U3006 ( .A1(n2338), .A2(n2327), .ZN(n3022) );
  INV_X1 U3007 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2328) );
  NOR2_X1 U3008 ( .A1(n2258), .A2(n2329), .ZN(n2330) );
  NAND2_X1 U3009 ( .A1(n2333), .A2(IR_REG_31__SCAN_IN), .ZN(n2334) );
  XNOR2_X1 U3010 ( .A(n2334), .B(IR_REG_4__SCAN_IN), .ZN(n4417) );
  MUX2_X1 U3011 ( .A(DATAI_4_), .B(n4417), .S(n2041), .Z(n3015) );
  NAND2_X1 U3012 ( .A1(n3108), .A2(n3015), .ZN(n3659) );
  NAND2_X1 U3013 ( .A1(n3004), .A2(n3745), .ZN(n3003) );
  NAND2_X1 U3014 ( .A1(n3818), .A2(n3015), .ZN(n2335) );
  NAND2_X1 U3015 ( .A1(n3636), .A2(REG0_REG_5__SCAN_IN), .ZN(n2345) );
  INV_X1 U3016 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2792) );
  OR2_X1 U3017 ( .A1(n3639), .A2(n2792), .ZN(n2344) );
  INV_X1 U3018 ( .A(n2352), .ZN(n2340) );
  INV_X1 U3019 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U3020 ( .A1(n2338), .A2(n2337), .ZN(n2339) );
  NAND2_X1 U3021 ( .A1(n2340), .A2(n2339), .ZN(n3103) );
  OR2_X1 U3022 ( .A1(n2610), .A2(n3103), .ZN(n2343) );
  INV_X1 U3023 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2341) );
  OR2_X1 U3024 ( .A1(n2488), .A2(n2341), .ZN(n2342) );
  INV_X1 U3025 ( .A(DATAI_5_), .ZN(n2349) );
  NAND2_X1 U3026 ( .A1(n2346), .A2(IR_REG_31__SCAN_IN), .ZN(n2348) );
  XNOR2_X1 U3027 ( .A(n2348), .B(n2347), .ZN(n2793) );
  MUX2_X1 U3028 ( .A(n2349), .B(n2793), .S(n2041), .Z(n3036) );
  NAND2_X1 U3029 ( .A1(n3636), .A2(REG0_REG_6__SCAN_IN), .ZN(n2357) );
  INV_X1 U3030 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3093) );
  OR2_X1 U3031 ( .A1(n2488), .A2(n3093), .ZN(n2356) );
  OAI21_X1 U3032 ( .B1(n2352), .B2(REG3_REG_6__SCAN_IN), .A(n2363), .ZN(n3130)
         );
  INV_X1 U3033 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2353) );
  OR2_X1 U3034 ( .A1(n3639), .A2(n2353), .ZN(n2354) );
  INV_X1 U3035 ( .A(DATAI_6_), .ZN(n2359) );
  NOR2_X1 U3036 ( .A1(n2346), .A2(IR_REG_5__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3037 ( .A1(n2371), .A2(n2748), .ZN(n2358) );
  XNOR2_X1 U3038 ( .A(n2358), .B(n2370), .ZN(n2797) );
  MUX2_X1 U3039 ( .A(n2359), .B(n2797), .S(n2040), .Z(n3124) );
  OAI22_X2 U3040 ( .A1(n3077), .A2(n2360), .B1(n3119), .B2(n3816), .ZN(n3176)
         );
  NAND2_X1 U3041 ( .A1(n3636), .A2(REG0_REG_7__SCAN_IN), .ZN(n2369) );
  INV_X1 U3042 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2361) );
  OR2_X1 U3043 ( .A1(n2488), .A2(n2361), .ZN(n2368) );
  AND2_X1 U3044 ( .A1(n2363), .A2(n2362), .ZN(n2364) );
  OR2_X1 U3045 ( .A1(n2364), .A2(n2372), .ZN(n3175) );
  INV_X1 U3046 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2365) );
  OR2_X1 U3047 ( .A1(n3639), .A2(n2365), .ZN(n2366) );
  NAND2_X1 U3048 ( .A1(n2371), .A2(n2370), .ZN(n2391) );
  NAND2_X1 U3049 ( .A1(n2391), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U3050 ( .A(n2379), .B(IR_REG_7__SCAN_IN), .ZN(n4414) );
  MUX2_X1 U3051 ( .A(DATAI_7_), .B(n4414), .S(n2041), .Z(n3170) );
  NAND2_X1 U3052 ( .A1(n3279), .A2(n3170), .ZN(n2642) );
  INV_X1 U3053 ( .A(n3170), .ZN(n3167) );
  NAND2_X1 U3054 ( .A1(n3815), .A2(n3167), .ZN(n3668) );
  NAND2_X1 U3055 ( .A1(n3636), .A2(REG0_REG_8__SCAN_IN), .ZN(n2377) );
  INV_X1 U3056 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3217) );
  OR2_X1 U3057 ( .A1(n3639), .A2(n3217), .ZN(n2376) );
  OR2_X1 U3058 ( .A1(n2372), .A2(REG3_REG_8__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3059 ( .A1(n2384), .A2(n2373), .ZN(n4514) );
  OR2_X1 U3060 ( .A1(n2610), .A2(n4514), .ZN(n2375) );
  INV_X1 U3061 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4515) );
  OR2_X1 U3062 ( .A1(n2488), .A2(n4515), .ZN(n2374) );
  INV_X1 U3063 ( .A(IR_REG_7__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3064 ( .A1(n2379), .A2(n2378), .ZN(n2380) );
  NAND2_X1 U3065 ( .A1(n2380), .A2(IR_REG_31__SCAN_IN), .ZN(n2381) );
  XNOR2_X1 U3066 ( .A(n2381), .B(IR_REG_8__SCAN_IN), .ZN(n4413) );
  MUX2_X1 U3067 ( .A(DATAI_8_), .B(n4413), .S(n2040), .Z(n3287) );
  NOR2_X1 U3068 ( .A1(n3814), .A2(n3287), .ZN(n2382) );
  INV_X1 U3069 ( .A(n3287), .ZN(n3278) );
  NAND2_X1 U3070 ( .A1(n3636), .A2(REG0_REG_9__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3071 ( .A1(n2384), .A2(n2383), .ZN(n2385) );
  NAND2_X1 U3072 ( .A1(n2399), .A2(n2385), .ZN(n3197) );
  INV_X1 U3073 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2386) );
  OR2_X1 U3074 ( .A1(n3639), .A2(n2386), .ZN(n2388) );
  INV_X1 U3075 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3076 ( .A1(n2488), .A2(n3204), .ZN(n2387) );
  NAND2_X1 U3077 ( .A1(n2394), .A2(IR_REG_31__SCAN_IN), .ZN(n2392) );
  MUX2_X1 U3078 ( .A(IR_REG_31__SCAN_IN), .B(n2392), .S(IR_REG_9__SCAN_IN), 
        .Z(n2393) );
  INV_X1 U3079 ( .A(n2393), .ZN(n2395) );
  MUX2_X1 U3080 ( .A(DATAI_9_), .B(n3215), .S(n2041), .Z(n3251) );
  NOR2_X1 U3081 ( .A1(n2397), .A2(n2396), .ZN(n3263) );
  NAND2_X1 U3082 ( .A1(n3636), .A2(REG0_REG_10__SCAN_IN), .ZN(n2405) );
  INV_X1 U3083 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3084 ( .A1(n3639), .A2(n2398), .ZN(n2404) );
  INV_X1 U3085 ( .A(n2409), .ZN(n2411) );
  NAND2_X1 U3086 ( .A1(n2399), .A2(n4704), .ZN(n2400) );
  NAND2_X1 U3087 ( .A1(n2411), .A2(n2400), .ZN(n3268) );
  OR2_X1 U3088 ( .A1(n2610), .A2(n3268), .ZN(n2403) );
  INV_X1 U3089 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2401) );
  OR2_X1 U3090 ( .A1(n2488), .A2(n2401), .ZN(n2402) );
  INV_X1 U3091 ( .A(DATAI_10_), .ZN(n4721) );
  OR2_X1 U3092 ( .A1(n2418), .A2(n2748), .ZN(n2406) );
  MUX2_X1 U3093 ( .A(n4721), .B(n4534), .S(n2040), .Z(n3294) );
  NAND2_X1 U3094 ( .A1(n4330), .A2(n3294), .ZN(n2408) );
  NOR2_X1 U3095 ( .A1(n4330), .A2(n3294), .ZN(n2407) );
  AOI21_X1 U3096 ( .B1(n3263), .B2(n2408), .A(n2407), .ZN(n4157) );
  NAND2_X1 U3097 ( .A1(n3636), .A2(REG0_REG_11__SCAN_IN), .ZN(n2416) );
  INV_X1 U3098 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4334) );
  OR2_X1 U3099 ( .A1(n3639), .A2(n4334), .ZN(n2415) );
  INV_X1 U3100 ( .A(n2421), .ZN(n2423) );
  INV_X1 U3101 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3102 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  NAND2_X1 U3103 ( .A1(n2423), .A2(n2412), .ZN(n4165) );
  INV_X1 U3104 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4166) );
  OR2_X1 U3105 ( .A1(n2488), .A2(n4166), .ZN(n2413) );
  INV_X1 U3106 ( .A(IR_REG_10__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3107 ( .A1(n2418), .A2(n2417), .ZN(n2419) );
  NAND2_X1 U3108 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2430) );
  XNOR2_X1 U3109 ( .A(n2430), .B(IR_REG_11__SCAN_IN), .ZN(n3214) );
  MUX2_X1 U3110 ( .A(DATAI_11_), .B(n3214), .S(n2040), .Z(n3309) );
  NAND2_X1 U3111 ( .A1(n4318), .A2(n3309), .ZN(n3680) );
  INV_X1 U3112 ( .A(n3309), .ZN(n4168) );
  NAND2_X1 U3113 ( .A1(n3812), .A2(n4168), .ZN(n3679) );
  NAND2_X1 U3114 ( .A1(n3680), .A2(n3679), .ZN(n4159) );
  NAND2_X1 U3115 ( .A1(n4157), .A2(n4159), .ZN(n4156) );
  NAND2_X1 U3116 ( .A1(n4156), .A2(n2420), .ZN(n3338) );
  NAND2_X1 U3117 ( .A1(n3636), .A2(REG0_REG_12__SCAN_IN), .ZN(n2428) );
  INV_X1 U3118 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3344) );
  OR2_X1 U3119 ( .A1(n2488), .A2(n3344), .ZN(n2427) );
  INV_X1 U3120 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3121 ( .A1(n2423), .A2(n2422), .ZN(n2424) );
  NAND2_X1 U3122 ( .A1(n2436), .A2(n2424), .ZN(n3343) );
  INV_X1 U3123 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4327) );
  OR2_X1 U3124 ( .A1(n3639), .A2(n4327), .ZN(n2425) );
  INV_X1 U3125 ( .A(IR_REG_11__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3126 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  NAND2_X1 U3127 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  MUX2_X1 U3128 ( .A(DATAI_12_), .B(n4462), .S(n2560), .Z(n3346) );
  NAND2_X1 U3129 ( .A1(n4141), .A2(n3346), .ZN(n2434) );
  NOR2_X1 U3130 ( .A1(n4141), .A2(n3346), .ZN(n2433) );
  NAND2_X1 U3131 ( .A1(n3636), .A2(REG0_REG_13__SCAN_IN), .ZN(n2441) );
  INV_X1 U3132 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4150) );
  OR2_X1 U3133 ( .A1(n2488), .A2(n4150), .ZN(n2440) );
  INV_X1 U3134 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3135 ( .A1(n2436), .A2(n2435), .ZN(n2437) );
  NAND2_X1 U3136 ( .A1(n2448), .A2(n2437), .ZN(n4149) );
  OR2_X1 U3137 ( .A1(n2450), .A2(n4149), .ZN(n2439) );
  INV_X1 U3138 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4314) );
  OR2_X1 U3139 ( .A1(n3639), .A2(n4314), .ZN(n2438) );
  INV_X1 U3140 ( .A(DATAI_13_), .ZN(n2446) );
  NOR2_X1 U3141 ( .A1(n2442), .A2(n2748), .ZN(n2443) );
  MUX2_X1 U3142 ( .A(n2748), .B(n2443), .S(IR_REG_13__SCAN_IN), .Z(n2445) );
  OR2_X1 U3143 ( .A1(n2445), .A2(n2493), .ZN(n3232) );
  MUX2_X1 U3144 ( .A(n2446), .B(n3232), .S(n2560), .Z(n4145) );
  INV_X1 U3145 ( .A(n4145), .ZN(n3379) );
  NAND2_X1 U3146 ( .A1(n3636), .A2(REG0_REG_14__SCAN_IN), .ZN(n2455) );
  INV_X1 U3147 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4310) );
  OR2_X1 U31480 ( .A1(n3639), .A2(n4310), .ZN(n2454) );
  INV_X1 U31490 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2447) );
  NAND2_X1 U3150 ( .A1(n2448), .A2(n2447), .ZN(n2449) );
  NAND2_X1 U3151 ( .A1(n2457), .A2(n2449), .ZN(n3476) );
  OR2_X1 U3152 ( .A1(n2450), .A2(n3476), .ZN(n2453) );
  INV_X1 U3153 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3154 ( .A1(n2488), .A2(n2451), .ZN(n2452) );
  OR2_X1 U3155 ( .A1(n2493), .A2(n2748), .ZN(n2456) );
  XNOR2_X1 U3156 ( .A(n2456), .B(IR_REG_14__SCAN_IN), .ZN(n3855) );
  MUX2_X1 U3157 ( .A(DATAI_14_), .B(n3855), .S(n2560), .Z(n4127) );
  NAND2_X1 U3158 ( .A1(n4295), .A2(n4127), .ZN(n3683) );
  INV_X1 U3159 ( .A(n4295), .ZN(n4113) );
  NAND2_X1 U3160 ( .A1(n4113), .A2(n4300), .ZN(n3646) );
  NAND2_X1 U3161 ( .A1(n3636), .A2(REG0_REG_15__SCAN_IN), .ZN(n2463) );
  INV_X1 U3162 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3627) );
  INV_X1 U3163 ( .A(n2474), .ZN(n2475) );
  NAND2_X1 U3164 ( .A1(n2457), .A2(n3627), .ZN(n2458) );
  NAND2_X1 U3165 ( .A1(n2475), .A2(n2458), .ZN(n4114) );
  OR2_X1 U3166 ( .A1(n4114), .A2(n2610), .ZN(n2462) );
  INV_X1 U3167 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2459) );
  OR2_X1 U3168 ( .A1(n2488), .A2(n2459), .ZN(n2461) );
  INV_X1 U3169 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4298) );
  OR2_X1 U3170 ( .A1(n3639), .A2(n4298), .ZN(n2460) );
  INV_X1 U3171 ( .A(DATAI_15_), .ZN(n2466) );
  NAND2_X1 U3172 ( .A1(n2493), .A2(n2464), .ZN(n2465) );
  NAND2_X1 U3173 ( .A1(n2465), .A2(IR_REG_31__SCAN_IN), .ZN(n2482) );
  XNOR2_X1 U3174 ( .A(n2482), .B(IR_REG_15__SCAN_IN), .ZN(n3862) );
  MUX2_X1 U3175 ( .A(n2466), .B(n4530), .S(n2560), .Z(n4118) );
  AOI21_X2 U3176 ( .B1(n4110), .B2(n2469), .A(n2263), .ZN(n4092) );
  INV_X1 U3177 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2470) );
  OR2_X1 U3178 ( .A1(n2488), .A2(n2470), .ZN(n2473) );
  INV_X1 U3179 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3180 ( .A1(n2302), .A2(n2471), .ZN(n2472) );
  AND2_X1 U3181 ( .A1(n2473), .A2(n2472), .ZN(n2480) );
  INV_X1 U3182 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U3183 ( .A1(n2475), .A2(n4718), .ZN(n2476) );
  NAND2_X1 U3184 ( .A1(n2486), .A2(n2476), .ZN(n3545) );
  OR2_X1 U3185 ( .A1(n3545), .A2(n2610), .ZN(n2479) );
  NAND2_X1 U3186 ( .A1(n2477), .A2(REG1_REG_16__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3187 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  NAND2_X1 U3188 ( .A1(n2483), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  XNOR2_X1 U3189 ( .A(n2484), .B(IR_REG_16__SCAN_IN), .ZN(n3863) );
  MUX2_X1 U3190 ( .A(DATAI_16_), .B(n3863), .S(n2560), .Z(n4281) );
  NAND2_X1 U3191 ( .A1(n4084), .A2(n4281), .ZN(n3770) );
  INV_X1 U3192 ( .A(n4281), .ZN(n4097) );
  NAND2_X1 U3193 ( .A1(n4292), .A2(n4097), .ZN(n3767) );
  NAND2_X1 U3194 ( .A1(n4292), .A2(n4281), .ZN(n2485) );
  INV_X1 U3195 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U3196 ( .A1(n2486), .A2(n4681), .ZN(n2487) );
  NAND2_X1 U3197 ( .A1(n2500), .A2(n2487), .ZN(n3555) );
  AOI22_X1 U3198 ( .A1(n2477), .A2(REG1_REG_17__SCAN_IN), .B1(n3636), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3199 ( .A1(n3635), .A2(REG2_REG_17__SCAN_IN), .ZN(n2489) );
  OAI211_X1 U3200 ( .C1(n3555), .C2(n2610), .A(n2490), .B(n2489), .ZN(n4282)
         );
  NOR2_X1 U3201 ( .A1(n2491), .A2(IR_REG_16__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3202 ( .A1(n2495), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  MUX2_X1 U3203 ( .A(IR_REG_31__SCAN_IN), .B(n2494), .S(IR_REG_17__SCAN_IN), 
        .Z(n2496) );
  AND2_X1 U3204 ( .A1(n2496), .A2(n2518), .ZN(n3876) );
  MUX2_X1 U3205 ( .A(DATAI_17_), .B(n3876), .S(n2560), .Z(n4274) );
  INV_X1 U3206 ( .A(n4066), .ZN(n2507) );
  INV_X1 U3207 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3605) );
  INV_X1 U3208 ( .A(n2509), .ZN(n2511) );
  NAND2_X1 U3209 ( .A1(n2500), .A2(n3605), .ZN(n2501) );
  NAND2_X1 U32100 ( .A1(n2511), .A2(n2501), .ZN(n4065) );
  OR2_X1 U32110 ( .A1(n4065), .A2(n2610), .ZN(n2504) );
  AOI22_X1 U32120 ( .A1(n2477), .A2(REG1_REG_18__SCAN_IN), .B1(n3636), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U32130 ( .A1(n3635), .A2(REG2_REG_18__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U32140 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2505) );
  XNOR2_X1 U32150 ( .A(n2505), .B(IR_REG_18__SCAN_IN), .ZN(n3879) );
  MUX2_X1 U32160 ( .A(DATAI_18_), .B(n3879), .S(n2560), .Z(n4060) );
  NAND2_X1 U32170 ( .A1(n4277), .A2(n4060), .ZN(n4041) );
  NAND2_X1 U32180 ( .A1(n3811), .A2(n4058), .ZN(n4042) );
  NAND2_X1 U32190 ( .A1(n2507), .A2(n2506), .ZN(n4067) );
  NAND2_X1 U32200 ( .A1(n4277), .A2(n4058), .ZN(n2508) );
  NAND2_X1 U32210 ( .A1(n4067), .A2(n2508), .ZN(n4038) );
  INV_X1 U32220 ( .A(n2525), .ZN(n2526) );
  INV_X1 U32230 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32240 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  NAND2_X1 U32250 ( .A1(n4052), .A2(n2288), .ZN(n2517) );
  INV_X1 U32260 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U32270 ( .A1(n3635), .A2(REG2_REG_19__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32280 ( .A1(n3636), .A2(REG0_REG_19__SCAN_IN), .ZN(n2513) );
  OAI211_X1 U32290 ( .C1(n4269), .C2(n3639), .A(n2514), .B(n2513), .ZN(n2515)
         );
  INV_X1 U32300 ( .A(n2515), .ZN(n2516) );
  NAND2_X1 U32310 ( .A1(n2520), .A2(n2519), .ZN(n2617) );
  OR2_X1 U32320 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  MUX2_X1 U32330 ( .A(DATAI_19_), .B(n4412), .S(n2560), .Z(n3494) );
  NAND2_X1 U32340 ( .A1(n4022), .A2(n3494), .ZN(n2522) );
  NAND2_X1 U32350 ( .A1(n4038), .A2(n2522), .ZN(n2524) );
  INV_X1 U32360 ( .A(n3494), .ZN(n4050) );
  NAND2_X1 U32370 ( .A1(n4062), .A2(n4050), .ZN(n2523) );
  NAND2_X1 U32380 ( .A1(n2524), .A2(n2523), .ZN(n4016) );
  INV_X1 U32390 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U32400 ( .A1(n2526), .A2(n4564), .ZN(n2527) );
  NAND2_X1 U32410 ( .A1(n2543), .A2(n2527), .ZN(n3576) );
  INV_X1 U32420 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U32430 ( .A1(n3635), .A2(REG2_REG_20__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32440 ( .A1(n3636), .A2(REG0_REG_20__SCAN_IN), .ZN(n2528) );
  OAI211_X1 U32450 ( .C1(n4265), .C2(n3639), .A(n2529), .B(n2528), .ZN(n2530)
         );
  INV_X1 U32460 ( .A(n2530), .ZN(n2531) );
  INV_X1 U32470 ( .A(DATAI_20_), .ZN(n4586) );
  NAND2_X1 U32480 ( .A1(n4255), .A2(n4030), .ZN(n2533) );
  XNOR2_X1 U32490 ( .A(n2543), .B(REG3_REG_21__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U32500 ( .A1(n4007), .A2(n2288), .ZN(n2538) );
  INV_X1 U32510 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U32520 ( .A1(n3636), .A2(REG0_REG_21__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32530 ( .A1(n3635), .A2(REG2_REG_21__SCAN_IN), .ZN(n2534) );
  OAI211_X1 U32540 ( .C1(n3639), .C2(n4261), .A(n2535), .B(n2534), .ZN(n2536)
         );
  INV_X1 U32550 ( .A(n2536), .ZN(n2537) );
  NAND2_X1 U32560 ( .A1(n2539), .A2(DATAI_21_), .ZN(n4009) );
  NOR2_X1 U32570 ( .A1(n4024), .A2(n4009), .ZN(n2540) );
  INV_X1 U32580 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3525) );
  INV_X1 U32590 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2541) );
  OAI21_X1 U32600 ( .B1(n2543), .B2(n3525), .A(n2541), .ZN(n2544) );
  NAND2_X1 U32610 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2542) );
  NAND2_X1 U32620 ( .A1(n2544), .A2(n2553), .ZN(n3996) );
  OR2_X1 U32630 ( .A1(n3996), .A2(n2610), .ZN(n2549) );
  INV_X1 U32640 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U32650 ( .A1(n3636), .A2(REG0_REG_22__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32660 ( .A1(n3635), .A2(REG2_REG_22__SCAN_IN), .ZN(n2545) );
  OAI211_X1 U32670 ( .C1(n3639), .C2(n4252), .A(n2546), .B(n2545), .ZN(n2547)
         );
  INV_X1 U32680 ( .A(n2547), .ZN(n2548) );
  INV_X1 U32690 ( .A(DATAI_22_), .ZN(n4595) );
  NOR2_X1 U32700 ( .A1(n2560), .A2(n4595), .ZN(n3983) );
  NAND2_X1 U32710 ( .A1(n4258), .A2(n3983), .ZN(n3968) );
  INV_X1 U32720 ( .A(n3983), .ZN(n3994) );
  NAND2_X1 U32730 ( .A1(n3810), .A2(n3994), .ZN(n2654) );
  NAND2_X1 U32740 ( .A1(n3810), .A2(n3983), .ZN(n2551) );
  NAND2_X1 U32750 ( .A1(n3990), .A2(n2551), .ZN(n3964) );
  INV_X1 U32760 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U32770 ( .A1(n2553), .A2(n4565), .ZN(n2554) );
  NAND2_X1 U32780 ( .A1(n2566), .A2(n2554), .ZN(n3485) );
  INV_X1 U32790 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4247) );
  NAND2_X1 U32800 ( .A1(n3635), .A2(REG2_REG_23__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U32810 ( .A1(n3636), .A2(REG0_REG_23__SCAN_IN), .ZN(n2555) );
  OAI211_X1 U32820 ( .C1(n4247), .C2(n3639), .A(n2556), .B(n2555), .ZN(n2557)
         );
  INV_X1 U32830 ( .A(n2557), .ZN(n2558) );
  NAND2_X1 U32840 ( .A1(n2539), .A2(DATAI_23_), .ZN(n3975) );
  NAND2_X1 U32850 ( .A1(n3987), .A2(n3975), .ZN(n2561) );
  NAND2_X1 U32860 ( .A1(n3964), .A2(n2561), .ZN(n2563) );
  INV_X1 U32870 ( .A(n3975), .ZN(n2703) );
  NAND2_X1 U32880 ( .A1(n4237), .A2(n2703), .ZN(n2562) );
  INV_X1 U32890 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U32900 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  NAND2_X1 U32910 ( .A1(n2575), .A2(n2567), .ZN(n3957) );
  OR2_X1 U32920 ( .A1(n3957), .A2(n2610), .ZN(n2572) );
  INV_X1 U32930 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4243) );
  NAND2_X1 U32940 ( .A1(n3635), .A2(REG2_REG_24__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32950 ( .A1(n3636), .A2(REG0_REG_24__SCAN_IN), .ZN(n2568) );
  OAI211_X1 U32960 ( .C1(n4243), .C2(n3639), .A(n2569), .B(n2568), .ZN(n2570)
         );
  INV_X1 U32970 ( .A(n2570), .ZN(n2571) );
  NAND2_X1 U32980 ( .A1(n2539), .A2(DATAI_24_), .ZN(n3954) );
  NOR2_X1 U32990 ( .A1(n3486), .A2(n3954), .ZN(n2574) );
  NAND2_X1 U33000 ( .A1(n3486), .A2(n3954), .ZN(n2573) );
  INV_X1 U33010 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U33020 ( .A1(n2575), .A2(n4684), .ZN(n2576) );
  NAND2_X1 U33030 ( .A1(n2585), .A2(n2576), .ZN(n3939) );
  INV_X1 U33040 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U33050 ( .A1(n3636), .A2(REG0_REG_25__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U33060 ( .A1(n3635), .A2(REG2_REG_25__SCAN_IN), .ZN(n2577) );
  OAI211_X1 U33070 ( .C1(n4234), .C2(n3639), .A(n2578), .B(n2577), .ZN(n2579)
         );
  INV_X1 U33080 ( .A(n2579), .ZN(n2580) );
  INV_X1 U33090 ( .A(DATAI_25_), .ZN(n2582) );
  NOR2_X1 U33100 ( .A1(n2560), .A2(n2582), .ZN(n4227) );
  NOR2_X1 U33110 ( .A1(n3809), .A2(n4227), .ZN(n2584) );
  NAND2_X1 U33120 ( .A1(n3809), .A2(n4227), .ZN(n2583) );
  INV_X1 U33130 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U33140 ( .A1(n2585), .A2(n3615), .ZN(n2586) );
  NAND2_X1 U33150 ( .A1(n3924), .A2(n2288), .ZN(n2591) );
  INV_X1 U33160 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4225) );
  NAND2_X1 U33170 ( .A1(n3635), .A2(REG2_REG_26__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U33180 ( .A1(n3636), .A2(REG0_REG_26__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U33190 ( .C1(n4225), .C2(n3639), .A(n2588), .B(n2587), .ZN(n2589)
         );
  INV_X1 U33200 ( .A(n2589), .ZN(n2590) );
  NAND2_X1 U33210 ( .A1(n2539), .A2(DATAI_26_), .ZN(n3923) );
  NOR2_X1 U33220 ( .A1(n4231), .A2(n3923), .ZN(n2592) );
  NAND2_X1 U33230 ( .A1(n4231), .A2(n3923), .ZN(n2593) );
  INV_X1 U33240 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33250 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  NAND2_X1 U33260 ( .A1(n2608), .A2(n2597), .ZN(n3467) );
  OR2_X1 U33270 ( .A1(n3467), .A2(n2610), .ZN(n2603) );
  INV_X1 U33280 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U33290 ( .A1(n3635), .A2(REG2_REG_27__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U33300 ( .A1(n3636), .A2(REG0_REG_27__SCAN_IN), .ZN(n2598) );
  OAI211_X1 U33310 ( .C1(n2600), .C2(n3639), .A(n2599), .B(n2598), .ZN(n2601)
         );
  INV_X1 U33320 ( .A(n2601), .ZN(n2602) );
  INV_X1 U33330 ( .A(DATAI_27_), .ZN(n2604) );
  NOR2_X1 U33340 ( .A1(n2560), .A2(n2604), .ZN(n4213) );
  NOR2_X1 U33350 ( .A1(n3919), .A2(n4213), .ZN(n2606) );
  NAND2_X1 U33360 ( .A1(n3919), .A2(n4213), .ZN(n2605) );
  INV_X1 U33370 ( .A(n2608), .ZN(n2607) );
  NAND2_X1 U33380 ( .A1(n2607), .A2(REG3_REG_28__SCAN_IN), .ZN(n3904) );
  INV_X1 U33390 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U33400 ( .A1(n2608), .A2(n3514), .ZN(n2609) );
  NAND2_X1 U33410 ( .A1(n3904), .A2(n2609), .ZN(n3516) );
  INV_X1 U33420 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33430 ( .A1(n3635), .A2(REG2_REG_28__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U33440 ( .A1(n3636), .A2(REG0_REG_28__SCAN_IN), .ZN(n2611) );
  OAI211_X1 U33450 ( .C1(n2613), .C2(n3639), .A(n2612), .B(n2611), .ZN(n2614)
         );
  INV_X1 U33460 ( .A(n2614), .ZN(n2615) );
  INV_X1 U33470 ( .A(DATAI_28_), .ZN(n4687) );
  NOR2_X1 U33480 ( .A1(n2560), .A2(n4687), .ZN(n2715) );
  NAND2_X1 U33490 ( .A1(n3507), .A2(n2715), .ZN(n3706) );
  INV_X1 U33500 ( .A(n2715), .ZN(n3515) );
  NAND2_X1 U33510 ( .A1(n4216), .A2(n3515), .ZN(n3642) );
  NAND2_X1 U33520 ( .A1(n3706), .A2(n3642), .ZN(n2713) );
  XNOR2_X1 U3353 ( .A(n2714), .B(n2713), .ZN(n3352) );
  NAND2_X1 U33540 ( .A1(n2621), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  MUX2_X1 U3355 ( .A(IR_REG_31__SCAN_IN), .B(n2622), .S(IR_REG_21__SCAN_IN), 
        .Z(n2624) );
  NAND2_X1 U3356 ( .A1(n2624), .A2(n2665), .ZN(n2830) );
  NAND2_X1 U3357 ( .A1(n2665), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  XNOR2_X1 U3358 ( .A(n2625), .B(IR_REG_22__SCAN_IN), .ZN(n4410) );
  XNOR2_X1 U3359 ( .A(n2836), .B(n4410), .ZN(n2626) );
  NAND2_X1 U3360 ( .A1(n2626), .A2(n3887), .ZN(n4028) );
  NAND2_X1 U3361 ( .A1(n2627), .A2(n4412), .ZN(n3056) );
  NAND2_X1 U3362 ( .A1(n2047), .A2(IR_REG_31__SCAN_IN), .ZN(n2628) );
  XNOR2_X1 U3363 ( .A(n2628), .B(n2255), .ZN(n4419) );
  AND2_X1 U3364 ( .A1(n3795), .A2(n4410), .ZN(n2759) );
  OR2_X1 U3365 ( .A1(n3904), .A2(n2610), .ZN(n2634) );
  INV_X1 U3366 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3367 ( .A1(n3635), .A2(REG2_REG_29__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3368 ( .A1(n3636), .A2(REG0_REG_29__SCAN_IN), .ZN(n2629) );
  OAI211_X1 U3369 ( .C1(n2631), .C2(n3639), .A(n2630), .B(n2629), .ZN(n2632)
         );
  INV_X1 U3370 ( .A(n2632), .ZN(n2633) );
  NAND2_X1 U3371 ( .A1(n2634), .A2(n2633), .ZN(n3807) );
  INV_X1 U3372 ( .A(n3919), .ZN(n3704) );
  INV_X1 U3373 ( .A(n2759), .ZN(n2820) );
  NOR2_X2 U3374 ( .A1(n4419), .A2(n2820), .ZN(n4304) );
  INV_X1 U3375 ( .A(n2627), .ZN(n4411) );
  INV_X1 U3376 ( .A(n4410), .ZN(n2824) );
  AND2_X1 U3377 ( .A1(n2824), .A2(n2830), .ZN(n3057) );
  NAND2_X1 U3378 ( .A1(n4411), .A2(n3057), .ZN(n4323) );
  OAI22_X1 U3379 ( .A1(n3704), .A2(n4329), .B1(n4323), .B2(n3515), .ZN(n2635)
         );
  AOI21_X1 U3380 ( .B1(n4291), .B2(n3807), .A(n2635), .ZN(n2664) );
  NAND2_X1 U3381 ( .A1(n2998), .A2(n3045), .ZN(n3658) );
  NAND2_X1 U3382 ( .A1(n4183), .A2(n2942), .ZN(n3656) );
  INV_X1 U3383 ( .A(n3659), .ZN(n2639) );
  AND2_X1 U3384 ( .A1(n3817), .A2(n3036), .ZN(n3067) );
  NAND2_X1 U3385 ( .A1(n3125), .A2(n3102), .ZN(n3648) );
  NAND2_X1 U3386 ( .A1(n3816), .A2(n3124), .ZN(n3661) );
  NAND2_X1 U3387 ( .A1(n3172), .A2(n3119), .ZN(n3665) );
  INV_X1 U3388 ( .A(n2642), .ZN(n2643) );
  NAND2_X1 U3389 ( .A1(n3254), .A2(n3287), .ZN(n3670) );
  NAND2_X1 U3390 ( .A1(n3814), .A2(n3278), .ZN(n3667) );
  AND2_X1 U3391 ( .A1(n3813), .A2(n3195), .ZN(n3192) );
  NAND2_X1 U3392 ( .A1(n3272), .A2(n3251), .ZN(n3671) );
  INV_X1 U3393 ( .A(n4330), .ZN(n4172) );
  NAND2_X1 U3394 ( .A1(n4172), .A2(n3294), .ZN(n3678) );
  NAND2_X1 U3395 ( .A1(n3262), .A2(n3678), .ZN(n2644) );
  INV_X1 U3396 ( .A(n3294), .ZN(n3267) );
  NAND2_X1 U3397 ( .A1(n4330), .A2(n3267), .ZN(n3645) );
  NAND2_X1 U3398 ( .A1(n2644), .A2(n3645), .ZN(n4158) );
  NAND2_X1 U3399 ( .A1(n4158), .A2(n3679), .ZN(n2645) );
  NAND2_X1 U3400 ( .A1(n2645), .A2(n3680), .ZN(n3339) );
  INV_X1 U3401 ( .A(n3346), .ZN(n4322) );
  NAND2_X1 U3402 ( .A1(n4141), .A2(n4322), .ZN(n4137) );
  NAND2_X1 U3403 ( .A1(n4303), .A2(n4145), .ZN(n3727) );
  NAND2_X1 U3404 ( .A1(n3339), .A2(n3685), .ZN(n2646) );
  NOR2_X1 U3405 ( .A1(n4141), .A2(n4322), .ZN(n4138) );
  NOR2_X1 U3406 ( .A1(n4303), .A2(n4145), .ZN(n3728) );
  AOI21_X1 U3407 ( .B1(n3685), .B2(n4138), .A(n3728), .ZN(n3681) );
  NAND2_X1 U3408 ( .A1(n3764), .A2(n2219), .ZN(n2647) );
  INV_X1 U3409 ( .A(n4106), .ZN(n2649) );
  NAND2_X1 U3410 ( .A1(n4301), .A2(n2467), .ZN(n3682) );
  NAND2_X1 U3411 ( .A1(n2468), .A2(n4118), .ZN(n3647) );
  NAND2_X1 U3412 ( .A1(n3682), .A2(n3647), .ZN(n4109) );
  AND2_X1 U3413 ( .A1(n4282), .A2(n2497), .ZN(n3726) );
  NAND2_X1 U3414 ( .A1(n4022), .A2(n4050), .ZN(n3724) );
  NAND2_X1 U3415 ( .A1(n3724), .A2(n4042), .ZN(n3693) );
  INV_X1 U3416 ( .A(n4030), .ZN(n3577) );
  NAND2_X1 U3417 ( .A1(n4255), .A2(n3577), .ZN(n2652) );
  INV_X1 U3418 ( .A(n2652), .ZN(n3694) );
  OR2_X1 U3419 ( .A1(n4282), .A2(n2497), .ZN(n4039) );
  AND2_X1 U3420 ( .A1(n4041), .A2(n4039), .ZN(n2650) );
  NAND2_X1 U3421 ( .A1(n4062), .A2(n3494), .ZN(n3725) );
  OAI21_X1 U3422 ( .B1(n3693), .B2(n2650), .A(n3725), .ZN(n4017) );
  NOR2_X1 U3423 ( .A1(n4255), .A2(n3577), .ZN(n2651) );
  OR2_X1 U3424 ( .A1(n4017), .A2(n2651), .ZN(n2653) );
  NAND2_X1 U3425 ( .A1(n2653), .A2(n2652), .ZN(n3772) );
  OR2_X1 U3426 ( .A1(n3984), .A2(n4009), .ZN(n3721) );
  AND2_X1 U3427 ( .A1(n3968), .A2(n3721), .ZN(n3773) );
  NAND2_X1 U3428 ( .A1(n4237), .A2(n3975), .ZN(n3722) );
  NAND2_X1 U3429 ( .A1(n3722), .A2(n2654), .ZN(n3700) );
  AND2_X1 U3430 ( .A1(n3984), .A2(n4009), .ZN(n3965) );
  AND2_X1 U3431 ( .A1(n3968), .A2(n3965), .ZN(n2655) );
  NOR2_X1 U3432 ( .A1(n3700), .A2(n2655), .ZN(n3774) );
  NAND2_X1 U3433 ( .A1(n2656), .A2(n3723), .ZN(n3950) );
  NOR2_X1 U3434 ( .A1(n4228), .A2(n3954), .ZN(n3720) );
  INV_X1 U3435 ( .A(n3923), .ZN(n2657) );
  NAND2_X1 U3436 ( .A1(n4231), .A2(n2657), .ZN(n2658) );
  NAND2_X1 U3437 ( .A1(n4240), .A2(n4227), .ZN(n3912) );
  NAND2_X1 U3438 ( .A1(n2658), .A2(n3912), .ZN(n3780) );
  INV_X1 U3439 ( .A(n4227), .ZN(n3937) );
  NAND2_X1 U3440 ( .A1(n3809), .A2(n3937), .ZN(n3759) );
  NAND2_X1 U3441 ( .A1(n4228), .A2(n3954), .ZN(n3929) );
  NAND2_X1 U3442 ( .A1(n3759), .A2(n3929), .ZN(n3913) );
  INV_X1 U3443 ( .A(n4231), .ZN(n3808) );
  AND2_X1 U3444 ( .A1(n3808), .A2(n3923), .ZN(n3783) );
  AOI21_X1 U3445 ( .B1(n2660), .B2(n3913), .A(n3783), .ZN(n3703) );
  XNOR2_X1 U3446 ( .A(n3919), .B(n4213), .ZN(n3787) );
  NAND2_X1 U3447 ( .A1(n3704), .A2(n4213), .ZN(n3705) );
  INV_X1 U3448 ( .A(n2713), .ZN(n3762) );
  XNOR2_X1 U3449 ( .A(n2720), .B(n3762), .ZN(n2663) );
  NAND2_X1 U3450 ( .A1(n4411), .A2(n3795), .ZN(n2662) );
  OR2_X1 U3451 ( .A1(n3887), .A2(n2824), .ZN(n2661) );
  NAND2_X1 U3452 ( .A1(n2663), .A2(n4098), .ZN(n3359) );
  OAI211_X1 U3453 ( .C1(n3352), .C2(n4546), .A(n2664), .B(n3359), .ZN(n2709)
         );
  INV_X1 U3454 ( .A(n2665), .ZN(n2667) );
  INV_X1 U3455 ( .A(IR_REG_22__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3456 ( .A1(n2667), .A2(n2666), .ZN(n2671) );
  NAND2_X1 U3457 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2678) );
  INV_X1 U34580 ( .A(IR_REG_23__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U34590 ( .A1(n2678), .A2(n2677), .ZN(n2680) );
  INV_X1 U3460 ( .A(n2669), .ZN(n2670) );
  OAI21_X1 U3461 ( .B1(n2671), .B2(n2670), .A(IR_REG_31__SCAN_IN), .ZN(n2672)
         );
  MUX2_X1 U3462 ( .A(IR_REG_31__SCAN_IN), .B(n2672), .S(IR_REG_25__SCAN_IN), 
        .Z(n2674) );
  NAND2_X1 U3463 ( .A1(n2673), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  MUX2_X1 U3464 ( .A(IR_REG_31__SCAN_IN), .B(n2675), .S(IR_REG_26__SCAN_IN), 
        .Z(n2676) );
  AND2_X1 U3465 ( .A1(n2676), .A2(n2046), .ZN(n4409) );
  OR2_X1 U3466 ( .A1(n2678), .A2(n2677), .ZN(n2679) );
  NAND2_X1 U34670 ( .A1(n2680), .A2(n2679), .ZN(n2758) );
  NAND2_X1 U3468 ( .A1(n2627), .A2(n3887), .ZN(n2819) );
  NAND2_X1 U34690 ( .A1(n2819), .A2(n2759), .ZN(n3010) );
  OAI211_X1 U3470 ( .C1(n4537), .C2(n3795), .A(n2831), .B(n3010), .ZN(n2681)
         );
  INV_X1 U34710 ( .A(n2681), .ZN(n2697) );
  NOR4_X1 U3472 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2685) );
  NOR4_X1 U34730 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2684) );
  NOR4_X1 U3474 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2683) );
  NOR4_X1 U34750 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2682) );
  NAND4_X1 U3476 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n2694)
         );
  NOR2_X1 U34770 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2689) );
  NOR4_X1 U3478 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U34790 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2687) );
  NOR4_X1 U3480 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2686) );
  NAND4_X1 U34810 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n2693)
         );
  INV_X1 U3482 ( .A(n2741), .ZN(n2695) );
  NAND2_X1 U34830 ( .A1(n2695), .A2(B_REG_SCAN_IN), .ZN(n2691) );
  MUX2_X1 U3484 ( .A(n2691), .B(B_REG_SCAN_IN), .S(n2690), .Z(n2692) );
  OAI21_X1 U34850 ( .B1(n2694), .B2(n2693), .A(n2751), .ZN(n2816) );
  INV_X1 U3486 ( .A(D_REG_1__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U34870 ( .A1(n2751), .A2(n3007), .ZN(n2817) );
  INV_X1 U3488 ( .A(n4409), .ZN(n2698) );
  NAND2_X1 U34890 ( .A1(n2695), .A2(n2698), .ZN(n2815) );
  NAND2_X1 U3490 ( .A1(n2817), .A2(n2815), .ZN(n2696) );
  INV_X1 U34910 ( .A(D_REG_0__SCAN_IN), .ZN(n2755) );
  INV_X1 U3492 ( .A(n2690), .ZN(n2699) );
  AND2_X1 U34930 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  AOI21_X1 U3494 ( .B1(n2751), .B2(n2755), .A(n2700), .ZN(n2818) );
  INV_X2 U34950 ( .A(n4557), .ZN(n4559) );
  MUX2_X1 U3496 ( .A(REG1_REG_28__SCAN_IN), .B(n2709), .S(n4559), .Z(n2701) );
  INV_X1 U34970 ( .A(n2701), .ZN(n2707) );
  NAND2_X1 U3498 ( .A1(n4198), .A2(n3054), .ZN(n2971) );
  NAND2_X1 U34990 ( .A1(n2967), .A2(n2942), .ZN(n2702) );
  NOR2_X2 U3500 ( .A1(n2971), .A2(n2702), .ZN(n3021) );
  NAND2_X1 U35010 ( .A1(n3021), .A2(n3020), .ZN(n3072) );
  NOR2_X2 U3502 ( .A1(n3072), .A2(n3102), .ZN(n3082) );
  NAND2_X1 U35030 ( .A1(n3082), .A2(n3124), .ZN(n3166) );
  OR2_X2 U3504 ( .A1(n3166), .A2(n3170), .ZN(n3286) );
  NOR2_X2 U35050 ( .A1(n3286), .A2(n3287), .ZN(n3285) );
  AND2_X2 U35060 ( .A1(n3285), .A2(n3195), .ZN(n3264) );
  OR2_X2 U35070 ( .A1(n3265), .A2(n3309), .ZN(n4167) );
  NOR2_X2 U35080 ( .A1(n4167), .A2(n3346), .ZN(n4146) );
  AND2_X2 U35090 ( .A1(n4146), .A2(n4145), .ZN(n4148) );
  OR2_X2 U35100 ( .A1(n4057), .A2(n3494), .ZN(n4049) );
  INV_X1 U35110 ( .A(n3954), .ZN(n4236) );
  INV_X1 U35120 ( .A(n2704), .ZN(n3365) );
  NOR2_X2 U35130 ( .A1(n2704), .A2(n2715), .ZN(n2731) );
  INV_X1 U35140 ( .A(n2731), .ZN(n2705) );
  NAND2_X1 U35150 ( .A1(n2707), .A2(n2706), .ZN(U3546) );
  INV_X1 U35160 ( .A(n2818), .ZN(n3012) );
  AND2_X2 U35170 ( .A1(n2708), .A2(n3012), .ZN(n4553) );
  MUX2_X1 U35180 ( .A(REG0_REG_28__SCAN_IN), .B(n2709), .S(n4553), .Z(n2710)
         );
  INV_X1 U35190 ( .A(n2710), .ZN(n2712) );
  NAND2_X1 U35200 ( .A1(n2712), .A2(n2711), .ZN(U3514) );
  NAND2_X1 U35210 ( .A1(n2714), .A2(n2713), .ZN(n2717) );
  NAND2_X1 U35220 ( .A1(n2717), .A2(n2716), .ZN(n2719) );
  NAND2_X1 U35230 ( .A1(n2539), .A2(DATAI_29_), .ZN(n3902) );
  XNOR2_X1 U35240 ( .A(n3807), .B(n3902), .ZN(n3717) );
  XNOR2_X1 U35250 ( .A(n2719), .B(n2718), .ZN(n3900) );
  NAND2_X1 U35260 ( .A1(n3900), .A2(n4325), .ZN(n2730) );
  NOR2_X1 U35270 ( .A1(n4323), .A2(n3902), .ZN(n2729) );
  NAND2_X1 U35280 ( .A1(n3635), .A2(REG2_REG_30__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U35290 ( .A1(n3636), .A2(REG0_REG_30__SCAN_IN), .ZN(n2723) );
  INV_X1 U35300 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2721) );
  OR2_X1 U35310 ( .A1(n3639), .A2(n2721), .ZN(n2722) );
  AND3_X1 U35320 ( .A1(n2724), .A2(n2723), .A3(n2722), .ZN(n3707) );
  NOR2_X1 U35330 ( .A1(n2726), .A2(n2725), .ZN(n4424) );
  NAND2_X1 U35340 ( .A1(n4424), .A2(B_REG_SCAN_IN), .ZN(n2727) );
  NAND2_X1 U35350 ( .A1(n4291), .A2(n2727), .ZN(n3893) );
  OAI22_X1 U35360 ( .A1(n2728), .A2(n4306), .B1(n3707), .B2(n3893), .ZN(n3907)
         );
  NAND2_X1 U35370 ( .A1(n2731), .A2(n3902), .ZN(n4208) );
  OAI21_X1 U35380 ( .B1(n2731), .B2(n3902), .A(n4208), .ZN(n3905) );
  NAND2_X1 U35390 ( .A1(n2732), .A2(n2261), .ZN(U3515) );
  OR2_X1 U35400 ( .A1(n2733), .A2(n4557), .ZN(n2734) );
  NAND2_X1 U35410 ( .A1(n2734), .A2(n2257), .ZN(n2735) );
  NAND2_X1 U35420 ( .A1(n2735), .A2(n2260), .ZN(U3547) );
  INV_X1 U35430 ( .A(n4527), .ZN(n2753) );
  OR2_X1 U35440 ( .A1(n2835), .A2(n2753), .ZN(n3819) );
  INV_X2 U35450 ( .A(n3819), .ZN(U4043) );
  INV_X1 U35460 ( .A(DATAI_3_), .ZN(n2736) );
  MUX2_X1 U35470 ( .A(n2780), .B(n2736), .S(U3149), .Z(n2737) );
  INV_X1 U35480 ( .A(n2737), .ZN(U3349) );
  INV_X1 U35490 ( .A(n3232), .ZN(n3856) );
  NAND2_X1 U35500 ( .A1(n3856), .A2(STATE_REG_SCAN_IN), .ZN(n2738) );
  OAI21_X1 U35510 ( .B1(STATE_REG_SCAN_IN), .B2(n2446), .A(n2738), .ZN(U3339)
         );
  INV_X1 U35520 ( .A(DATAI_17_), .ZN(n4598) );
  NAND2_X1 U35530 ( .A1(n3876), .A2(STATE_REG_SCAN_IN), .ZN(n2739) );
  OAI21_X1 U35540 ( .B1(STATE_REG_SCAN_IN), .B2(n4598), .A(n2739), .ZN(U3335)
         );
  INV_X1 U35550 ( .A(DATAI_21_), .ZN(n4720) );
  NAND2_X1 U35560 ( .A1(n3795), .A2(STATE_REG_SCAN_IN), .ZN(n2740) );
  OAI21_X1 U35570 ( .B1(STATE_REG_SCAN_IN), .B2(n4720), .A(n2740), .ZN(U3331)
         );
  NAND2_X1 U35580 ( .A1(n2741), .A2(STATE_REG_SCAN_IN), .ZN(n2742) );
  OAI21_X1 U35590 ( .B1(STATE_REG_SCAN_IN), .B2(n2582), .A(n2742), .ZN(U3327)
         );
  NAND2_X1 U35600 ( .A1(n4424), .A2(STATE_REG_SCAN_IN), .ZN(n2743) );
  OAI21_X1 U35610 ( .B1(STATE_REG_SCAN_IN), .B2(n2604), .A(n2743), .ZN(U3325)
         );
  INV_X1 U35620 ( .A(n3215), .ZN(n4438) );
  INV_X1 U35630 ( .A(DATAI_9_), .ZN(n2744) );
  MUX2_X1 U35640 ( .A(n4438), .B(n2744), .S(U3149), .Z(n2745) );
  INV_X1 U35650 ( .A(n2745), .ZN(U3343) );
  INV_X1 U35660 ( .A(DATAI_29_), .ZN(n4596) );
  NAND2_X1 U35670 ( .A1(n2746), .A2(STATE_REG_SCAN_IN), .ZN(n2747) );
  OAI21_X1 U35680 ( .B1(STATE_REG_SCAN_IN), .B2(n4596), .A(n2747), .ZN(U3323)
         );
  INV_X1 U35690 ( .A(DATAI_31_), .ZN(n4706) );
  OR4_X1 U35700 ( .A1(n2749), .A2(IR_REG_30__SCAN_IN), .A3(n2748), .A4(U3149), 
        .ZN(n2750) );
  OAI21_X1 U35710 ( .B1(STATE_REG_SCAN_IN), .B2(n4706), .A(n2750), .ZN(U3321)
         );
  INV_X1 U35720 ( .A(n2751), .ZN(n2752) );
  NAND2_X2 U35730 ( .A1(n2752), .A2(n2831), .ZN(n4526) );
  NOR3_X1 U35740 ( .A1(n2753), .A2(n2690), .A3(n4409), .ZN(n2754) );
  AOI21_X1 U35750 ( .B1(n4526), .B2(n2755), .A(n2754), .ZN(U3458) );
  INV_X1 U35760 ( .A(n2815), .ZN(n2756) );
  AOI22_X1 U35770 ( .A1(n4526), .A2(n3007), .B1(n2756), .B2(n4527), .ZN(U3459)
         );
  INV_X1 U35780 ( .A(n2831), .ZN(n3008) );
  INV_X1 U35790 ( .A(n2758), .ZN(n2757) );
  NAND2_X1 U35800 ( .A1(n2757), .A2(STATE_REG_SCAN_IN), .ZN(n3805) );
  NAND2_X1 U35810 ( .A1(n3008), .A2(n3805), .ZN(n2770) );
  AND2_X1 U3582 ( .A1(n2759), .A2(n2758), .ZN(n2760) );
  NOR2_X1 U3583 ( .A1(n2760), .A2(n2560), .ZN(n2769) );
  INV_X1 U3584 ( .A(n2769), .ZN(n2761) );
  NOR2_X1 U3585 ( .A1(n4505), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3586 ( .A1(n3819), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2762) );
  OAI21_X1 U3587 ( .B1(n3707), .B2(n3819), .A(n2762), .ZN(U3580) );
  INV_X1 U3588 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2763) );
  INV_X1 U3589 ( .A(IR_REG_0__SCAN_IN), .ZN(n2764) );
  NOR3_X1 U3590 ( .A1(n2765), .A2(n3062), .A3(n2764), .ZN(n3824) );
  MUX2_X1 U3591 ( .A(n4177), .B(REG2_REG_2__SCAN_IN), .S(n4418), .Z(n2913) );
  AOI21_X1 U3592 ( .B1(n4418), .B2(REG2_REG_2__SCAN_IN), .A(n2912), .ZN(n2766)
         );
  XNOR2_X1 U3593 ( .A(n2766), .B(n2780), .ZN(n3836) );
  OAI22_X1 U3594 ( .A1(n3836), .A2(n2767), .B1(n2766), .B2(n2780), .ZN(n2768)
         );
  INV_X1 U3595 ( .A(n4417), .ZN(n2931) );
  XNOR2_X1 U3596 ( .A(n2768), .B(n2931), .ZN(n2926) );
  MUX2_X1 U3597 ( .A(REG2_REG_5__SCAN_IN), .B(n2341), .S(n2793), .Z(n2771) );
  INV_X1 U3598 ( .A(n4419), .ZN(n2908) );
  AND2_X1 U3599 ( .A1(n2908), .A2(n4424), .ZN(n3801) );
  INV_X1 U3600 ( .A(n4464), .ZN(n4501) );
  AOI211_X1 U3601 ( .C1(n2772), .C2(n2771), .A(n4501), .B(n2790), .ZN(n2775)
         );
  NAND2_X1 U3602 ( .A1(n4426), .A2(n4419), .ZN(n4512) );
  AND2_X1 U3603 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3038) );
  AOI21_X1 U3604 ( .B1(n4505), .B2(ADDR_REG_5__SCAN_IN), .A(n3038), .ZN(n2773)
         );
  OAI21_X1 U3605 ( .B1(n4512), .B2(n2793), .A(n2773), .ZN(n2774) );
  NOR2_X1 U3606 ( .A1(n2775), .A2(n2774), .ZN(n2789) );
  XNOR2_X1 U3607 ( .A(n2793), .B(REG1_REG_5__SCAN_IN), .ZN(n2787) );
  XNOR2_X1 U3608 ( .A(n4418), .B(n2776), .ZN(n2917) );
  INV_X1 U3609 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2777) );
  AND2_X1 U3610 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3821)
         );
  NAND2_X1 U3611 ( .A1(n3822), .A2(n3821), .ZN(n3820) );
  NAND2_X1 U3612 ( .A1(n3820), .A2(n2778), .ZN(n2916) );
  NAND2_X1 U3613 ( .A1(n2917), .A2(n2916), .ZN(n2915) );
  NAND2_X1 U3614 ( .A1(n4418), .A2(REG1_REG_2__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U3615 ( .A1(n2915), .A2(n2779), .ZN(n2781) );
  XNOR2_X1 U3616 ( .A(n2781), .B(n2780), .ZN(n3835) );
  NAND2_X1 U3617 ( .A1(n3835), .A2(REG1_REG_3__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U3618 ( .A1(n2781), .A2(n3832), .ZN(n2782) );
  NAND2_X1 U3619 ( .A1(n3834), .A2(n2782), .ZN(n2783) );
  INV_X1 U3620 ( .A(n2783), .ZN(n2784) );
  XNOR2_X1 U3621 ( .A(n2783), .B(n2931), .ZN(n2928) );
  NAND2_X1 U3622 ( .A1(n2928), .A2(REG1_REG_4__SCAN_IN), .ZN(n2927) );
  OAI21_X1 U3623 ( .B1(n2784), .B2(n2931), .A(n2927), .ZN(n2786) );
  INV_X1 U3624 ( .A(n4424), .ZN(n2785) );
  NAND2_X1 U3625 ( .A1(n2786), .A2(n2787), .ZN(n2791) );
  OAI211_X1 U3626 ( .C1(n2787), .C2(n2786), .A(n4507), .B(n2791), .ZN(n2788)
         );
  NAND2_X1 U3627 ( .A1(n2789), .A2(n2788), .ZN(U3245) );
  INV_X1 U3628 ( .A(n2793), .ZN(n4416) );
  INV_X1 U3629 ( .A(n2797), .ZN(n4415) );
  XOR2_X1 U3630 ( .A(REG2_REG_6__SCAN_IN), .B(n2808), .Z(n2800) );
  OAI21_X1 U3631 ( .B1(n2793), .B2(n2792), .A(n2791), .ZN(n2803) );
  XOR2_X1 U3632 ( .A(n2797), .B(n2803), .Z(n2795) );
  INV_X1 U3633 ( .A(n4507), .ZN(n2794) );
  NOR2_X1 U3634 ( .A1(n2795), .A2(n2353), .ZN(n2802) );
  AOI211_X1 U3635 ( .C1(n2795), .C2(n2353), .A(n2794), .B(n2802), .ZN(n2799)
         );
  AND2_X1 U3636 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3127) );
  AOI21_X1 U3637 ( .B1(n4505), .B2(ADDR_REG_6__SCAN_IN), .A(n3127), .ZN(n2796)
         );
  OAI21_X1 U3638 ( .B1(n4512), .B2(n2797), .A(n2796), .ZN(n2798) );
  AOI211_X1 U3639 ( .C1(n2800), .C2(n4464), .A(n2799), .B(n2798), .ZN(n2801)
         );
  INV_X1 U3640 ( .A(n2801), .ZN(U3246) );
  MUX2_X1 U3641 ( .A(REG1_REG_7__SCAN_IN), .B(n2365), .S(n4414), .Z(n2804) );
  XNOR2_X1 U3642 ( .A(n2877), .B(n2804), .ZN(n2813) );
  INV_X1 U3643 ( .A(n4414), .ZN(n2878) );
  NOR2_X1 U3644 ( .A1(STATE_REG_SCAN_IN), .A2(n2362), .ZN(n3163) );
  AOI21_X1 U3645 ( .B1(n4505), .B2(ADDR_REG_7__SCAN_IN), .A(n3163), .ZN(n2805)
         );
  OAI21_X1 U3646 ( .B1(n4512), .B2(n2878), .A(n2805), .ZN(n2812) );
  INV_X1 U3647 ( .A(n2806), .ZN(n2807) );
  AOI22_X1 U3648 ( .A1(n2808), .A2(REG2_REG_6__SCAN_IN), .B1(n4415), .B2(n2807), .ZN(n2810) );
  MUX2_X1 U3649 ( .A(n2361), .B(REG2_REG_7__SCAN_IN), .S(n4414), .Z(n2809) );
  AOI211_X1 U3650 ( .C1(n2810), .C2(n2809), .A(n4501), .B(n2881), .ZN(n2811)
         );
  AOI211_X1 U3651 ( .C1(n4507), .C2(n2813), .A(n2812), .B(n2811), .ZN(n2814)
         );
  INV_X1 U3652 ( .A(n2814), .ZN(U3247) );
  AND2_X1 U3653 ( .A1(n2816), .A2(n2815), .ZN(n3011) );
  NAND3_X1 U3654 ( .A1(n3011), .A2(n2818), .A3(n2817), .ZN(n2828) );
  NAND2_X1 U3655 ( .A1(n2819), .A2(n3057), .ZN(n2821) );
  NAND2_X1 U3656 ( .A1(n2821), .A2(n2820), .ZN(n2841) );
  NAND2_X1 U3657 ( .A1(n2841), .A2(n4323), .ZN(n2822) );
  NAND2_X1 U3658 ( .A1(n2828), .A2(n2822), .ZN(n2823) );
  NAND2_X1 U3659 ( .A1(n2823), .A2(n3010), .ZN(n2948) );
  INV_X1 U3660 ( .A(n2948), .ZN(n2827) );
  INV_X1 U3661 ( .A(n2847), .ZN(n2825) );
  NAND2_X1 U3662 ( .A1(n2825), .A2(n4527), .ZN(n2826) );
  NOR2_X1 U3663 ( .A1(n3505), .A2(n2826), .ZN(n3802) );
  NAND2_X1 U3664 ( .A1(n2828), .A2(n3802), .ZN(n2949) );
  NAND3_X1 U3665 ( .A1(n2827), .A2(n2831), .A3(n2949), .ZN(n2904) );
  INV_X1 U3666 ( .A(n2904), .ZN(n2863) );
  AND2_X1 U3667 ( .A1(n4290), .A2(n2831), .ZN(n2829) );
  NAND2_X1 U3668 ( .A1(n2858), .A2(n2829), .ZN(n2833) );
  AND2_X1 U3669 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  INV_X1 U3670 ( .A(n3628), .ZN(n3595) );
  NOR2_X1 U3671 ( .A1(n3054), .A2(n3503), .ZN(n2837) );
  NAND2_X1 U3672 ( .A1(n2947), .A2(REG1_REG_0__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U3673 ( .A1(n2851), .A2(n2838), .ZN(n2840) );
  OR2_X4 U3674 ( .A1(n3503), .A2(n4285), .ZN(n3506) );
  NOR2_X1 U3675 ( .A1(n2841), .A2(n3008), .ZN(n2842) );
  AND2_X1 U3676 ( .A1(n3802), .A2(n4419), .ZN(n2843) );
  NAND2_X1 U3677 ( .A1(n2858), .A2(n2843), .ZN(n3578) );
  OAI22_X1 U3678 ( .A1(n2909), .A2(n3582), .B1(n2846), .B2(n3578), .ZN(n2844)
         );
  AOI21_X1 U3679 ( .B1(n3058), .B2(n3595), .A(n2844), .ZN(n2845) );
  OAI21_X1 U3680 ( .B1(n2863), .B2(n3061), .A(n2845), .ZN(U3229) );
  INV_X1 U3681 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4194) );
  OAI22_X1 U3682 ( .A1(n2846), .A2(n3504), .B1(n3503), .B2(n4198), .ZN(n2848)
         );
  XNOR2_X1 U3683 ( .A(n2848), .B(n3451), .ZN(n2892) );
  NAND2_X1 U3684 ( .A1(n2872), .A2(n2887), .ZN(n2849) );
  NAND2_X1 U3685 ( .A1(n2850), .A2(n2849), .ZN(n2893) );
  XNOR2_X1 U3686 ( .A(n2892), .B(n2893), .ZN(n2854) );
  NAND2_X1 U3687 ( .A1(n2851), .A2(n3451), .ZN(n2852) );
  OAI211_X1 U3688 ( .C1(n2854), .C2(n2855), .A(n2896), .B(n3625), .ZN(n2862)
         );
  INV_X1 U3689 ( .A(n3802), .ZN(n2856) );
  NOR2_X1 U3690 ( .A1(n2856), .A2(n4419), .ZN(n2857) );
  OAI22_X1 U3691 ( .A1(n3629), .A2(n2859), .B1(n2888), .B2(n3578), .ZN(n2860)
         );
  AOI21_X1 U3692 ( .B1(n2872), .B2(n3595), .A(n2860), .ZN(n2861) );
  OAI211_X1 U3693 ( .C1(n2863), .C2(n4194), .A(n2862), .B(n2861), .ZN(U3219)
         );
  OR2_X1 U3694 ( .A1(n2636), .A2(n2864), .ZN(n2865) );
  AND2_X1 U3695 ( .A1(n2866), .A2(n2865), .ZN(n4192) );
  INV_X1 U3696 ( .A(n4192), .ZN(n2871) );
  INV_X1 U3697 ( .A(n2636), .ZN(n3747) );
  OAI21_X1 U3698 ( .B1(n3747), .B2(n2110), .A(n2867), .ZN(n2868) );
  INV_X1 U3699 ( .A(n4028), .ZN(n4162) );
  AOI22_X1 U3700 ( .A1(n4098), .A2(n2868), .B1(n4192), .B2(n4162), .ZN(n4189)
         );
  OAI22_X1 U3701 ( .A1(n2888), .A2(n4316), .B1(n4323), .B2(n4198), .ZN(n2869)
         );
  AOI21_X1 U3702 ( .B1(n4304), .B2(n2834), .A(n2869), .ZN(n2870) );
  OAI211_X1 U3703 ( .C1(n4537), .C2(n2871), .A(n4189), .B(n2870), .ZN(n2937)
         );
  NAND2_X1 U3704 ( .A1(n2872), .A2(n3058), .ZN(n2873) );
  NAND2_X1 U3705 ( .A1(n2971), .A2(n2873), .ZN(n4195) );
  INV_X1 U3706 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2874) );
  OAI22_X1 U3707 ( .A1(n4406), .A2(n4195), .B1(n4553), .B2(n2874), .ZN(n2875)
         );
  AOI21_X1 U3708 ( .B1(n2937), .B2(n4553), .A(n2875), .ZN(n2876) );
  INV_X1 U3709 ( .A(n2876), .ZN(U3469) );
  INV_X1 U3710 ( .A(n4413), .ZN(n3219) );
  XNOR2_X1 U3711 ( .A(n2879), .B(n4413), .ZN(n3218) );
  XNOR2_X1 U3712 ( .A(n3218), .B(REG1_REG_8__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3713 ( .A1(n2880), .A2(n4507), .ZN(n2886) );
  XNOR2_X1 U3714 ( .A(REG2_REG_8__SCAN_IN), .B(n3205), .ZN(n2882) );
  NAND2_X1 U3715 ( .A1(n4464), .A2(n2882), .ZN(n2883) );
  NAND2_X1 U3716 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3153) );
  NAND2_X1 U3717 ( .A1(n2883), .A2(n3153), .ZN(n2884) );
  AOI21_X1 U3718 ( .B1(n4505), .B2(ADDR_REG_8__SCAN_IN), .A(n2884), .ZN(n2885)
         );
  OAI211_X1 U3719 ( .C1(n4512), .C2(n3219), .A(n2886), .B(n2885), .ZN(U3248)
         );
  OAI22_X1 U3720 ( .A1(n2888), .A2(n3504), .B1(n3503), .B2(n2967), .ZN(n2889)
         );
  OR2_X1 U3721 ( .A1(n2888), .A2(n3506), .ZN(n2891) );
  NAND2_X1 U3722 ( .A1(n4181), .A2(n2887), .ZN(n2890) );
  INV_X1 U3723 ( .A(n2892), .ZN(n2894) );
  NAND2_X1 U3724 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  INV_X1 U3725 ( .A(n2897), .ZN(n2898) );
  INV_X1 U3726 ( .A(n2946), .ZN(n2900) );
  AOI21_X1 U3727 ( .B1(n2897), .B2(n2901), .A(n2900), .ZN(n2906) );
  AOI22_X1 U3728 ( .A1(n3631), .A2(n4183), .B1(n3617), .B2(n2300), .ZN(n2902)
         );
  OAI21_X1 U3729 ( .B1(n3628), .B2(n2967), .A(n2902), .ZN(n2903) );
  AOI21_X1 U3730 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2904), .A(n2903), .ZN(n2905)
         );
  OAI21_X1 U3731 ( .B1(n2906), .B2(n3582), .A(n2905), .ZN(U3234) );
  NAND2_X1 U3732 ( .A1(n4424), .A2(n3062), .ZN(n2907) );
  NAND2_X1 U3733 ( .A1(n2908), .A2(n2907), .ZN(n4425) );
  NAND2_X1 U3734 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3823) );
  NOR2_X1 U3735 ( .A1(n2909), .A2(n4424), .ZN(n2910) );
  AOI211_X1 U3736 ( .C1(n4424), .C2(n3823), .A(n4419), .B(n2910), .ZN(n2911)
         );
  AOI211_X1 U3737 ( .C1(n2764), .C2(n4425), .A(n3819), .B(n2911), .ZN(n2932)
         );
  AOI211_X1 U3738 ( .C1(n2914), .C2(n2913), .A(n2912), .B(n4501), .ZN(n2925)
         );
  OAI211_X1 U3739 ( .C1(n2917), .C2(n2916), .A(n4507), .B(n2915), .ZN(n2918)
         );
  INV_X1 U3740 ( .A(n2918), .ZN(n2924) );
  INV_X1 U3741 ( .A(n4418), .ZN(n2922) );
  NOR2_X1 U3742 ( .A1(n2919), .A2(STATE_REG_SCAN_IN), .ZN(n2920) );
  AOI21_X1 U3743 ( .B1(n4505), .B2(ADDR_REG_2__SCAN_IN), .A(n2920), .ZN(n2921)
         );
  OAI21_X1 U3744 ( .B1(n4512), .B2(n2922), .A(n2921), .ZN(n2923) );
  OR4_X1 U3745 ( .A1(n2932), .A2(n2925), .A3(n2924), .A4(n2923), .ZN(U3242) );
  XOR2_X1 U3746 ( .A(REG2_REG_4__SCAN_IN), .B(n2926), .Z(n2934) );
  OAI211_X1 U3747 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2928), .A(n4507), .B(n2927), 
        .ZN(n2930) );
  AND2_X1 U3748 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3000) );
  AOI21_X1 U3749 ( .B1(n4505), .B2(ADDR_REG_4__SCAN_IN), .A(n3000), .ZN(n2929)
         );
  OAI211_X1 U3750 ( .C1(n4512), .C2(n2931), .A(n2930), .B(n2929), .ZN(n2933)
         );
  AOI211_X1 U3751 ( .C1(n4464), .C2(n2934), .A(n2933), .B(n2932), .ZN(n2935)
         );
  INV_X1 U3752 ( .A(n2935), .ZN(U3244) );
  OAI22_X1 U3753 ( .A1(n4336), .A2(n4195), .B1(n4559), .B2(n2777), .ZN(n2936)
         );
  AOI21_X1 U3754 ( .B1(n2937), .B2(n4559), .A(n2936), .ZN(n2938) );
  INV_X1 U3755 ( .A(n2938), .ZN(U3519) );
  NAND2_X1 U3756 ( .A1(n4183), .A2(n2887), .ZN(n2940) );
  NAND2_X1 U3757 ( .A1(n3045), .A2(n3461), .ZN(n2939) );
  NAND2_X1 U3758 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  NOR2_X1 U3759 ( .A1(n2942), .A2(n3504), .ZN(n2943) );
  AOI21_X1 U3760 ( .B1(n4183), .B2(n3464), .A(n2943), .ZN(n2989) );
  XNOR2_X1 U3761 ( .A(n2988), .B(n2989), .ZN(n2986) );
  NAND2_X1 U3762 ( .A1(n2944), .A2(n2054), .ZN(n2945) );
  XOR2_X1 U3763 ( .A(n2986), .B(n2987), .Z(n2955) );
  OAI22_X1 U3764 ( .A1(n3629), .A2(n2888), .B1(n3108), .B2(n3578), .ZN(n2953)
         );
  OAI21_X1 U3765 ( .B1(n2948), .B2(n2947), .A(STATE_REG_SCAN_IN), .ZN(n2951)
         );
  AND2_X1 U3766 ( .A1(n2949), .A2(n3805), .ZN(n2950) );
  MUX2_X1 U3767 ( .A(n3618), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2952) );
  AOI211_X1 U3768 ( .C1(n3045), .C2(n3595), .A(n2953), .B(n2952), .ZN(n2954)
         );
  OAI21_X1 U3769 ( .B1(n2955), .B2(n3582), .A(n2954), .ZN(U3215) );
  NAND2_X1 U3770 ( .A1(n2957), .A2(n3746), .ZN(n2958) );
  NAND2_X1 U3771 ( .A1(n2956), .A2(n2958), .ZN(n4179) );
  AOI22_X1 U3772 ( .A1(n4183), .A2(n4291), .B1(n4181), .B2(n4290), .ZN(n2959)
         );
  OAI21_X1 U3773 ( .B1(n2846), .B2(n4329), .A(n2959), .ZN(n2966) );
  NAND2_X1 U3774 ( .A1(n4179), .A2(n4162), .ZN(n2964) );
  OAI21_X1 U3775 ( .B1(n3746), .B2(n2961), .A(n2960), .ZN(n2962) );
  NAND2_X1 U3776 ( .A1(n2962), .A2(n4098), .ZN(n2963) );
  AND2_X1 U3777 ( .A1(n2964), .A2(n2963), .ZN(n4178) );
  INV_X1 U3778 ( .A(n4178), .ZN(n2965) );
  AOI211_X1 U3779 ( .C1(n4543), .C2(n4179), .A(n2966), .B(n2965), .ZN(n2970)
         );
  INV_X1 U3780 ( .A(n4406), .ZN(n4346) );
  XNOR2_X1 U3781 ( .A(n2971), .B(n2967), .ZN(n4184) );
  AOI22_X1 U3782 ( .A1(n4346), .A2(n4184), .B1(REG0_REG_2__SCAN_IN), .B2(n4551), .ZN(n2968) );
  OAI21_X1 U3783 ( .B1(n2970), .B2(n4551), .A(n2968), .ZN(U3471) );
  INV_X1 U3784 ( .A(n4336), .ZN(n4221) );
  AOI22_X1 U3785 ( .A1(n4221), .A2(n4184), .B1(REG1_REG_2__SCAN_IN), .B2(n4557), .ZN(n2969) );
  OAI21_X1 U3786 ( .B1(n2970), .B2(n4557), .A(n2969), .ZN(U3520) );
  INV_X1 U3787 ( .A(n3021), .ZN(n2973) );
  OAI21_X1 U3788 ( .B1(n2971), .B2(n4181), .A(n3045), .ZN(n2972) );
  NAND2_X1 U3789 ( .A1(n2973), .A2(n2972), .ZN(n3049) );
  XNOR2_X1 U3790 ( .A(n2974), .B(n3735), .ZN(n3053) );
  OAI21_X1 U3791 ( .B1(n3735), .B2(n2976), .A(n2975), .ZN(n2978) );
  AOI22_X1 U3792 ( .A1(n2978), .A2(n4098), .B1(n4304), .B2(n2977), .ZN(n3043)
         );
  AOI22_X1 U3793 ( .A1(n3818), .A2(n4291), .B1(n4290), .B2(n3045), .ZN(n2979)
         );
  OAI211_X1 U3794 ( .C1(n4546), .C2(n3053), .A(n3043), .B(n2979), .ZN(n2984)
         );
  NAND2_X1 U3795 ( .A1(n2984), .A2(n4553), .ZN(n2981) );
  NAND2_X1 U3796 ( .A1(n4551), .A2(REG0_REG_3__SCAN_IN), .ZN(n2980) );
  OAI211_X1 U3797 ( .C1(n3049), .C2(n4406), .A(n2981), .B(n2980), .ZN(U3473)
         );
  OAI22_X1 U3798 ( .A1(n4336), .A2(n3049), .B1(n4559), .B2(n2982), .ZN(n2983)
         );
  AOI21_X1 U3799 ( .B1(n2984), .B2(n4559), .A(n2983), .ZN(n2985) );
  INV_X1 U3800 ( .A(n2985), .ZN(U3521) );
  INV_X1 U3801 ( .A(n2988), .ZN(n2990) );
  OAI22_X1 U3802 ( .A1(n3108), .A2(n3504), .B1(n3503), .B2(n3020), .ZN(n2991)
         );
  XNOR2_X1 U3803 ( .A(n2991), .B(n3508), .ZN(n3028) );
  OR2_X1 U3804 ( .A1(n3108), .A2(n3506), .ZN(n2993) );
  NAND2_X1 U3805 ( .A1(n3015), .A2(n3462), .ZN(n2992) );
  NAND2_X1 U3806 ( .A1(n2993), .A2(n2992), .ZN(n3027) );
  XNOR2_X1 U3807 ( .A(n3028), .B(n3027), .ZN(n2995) );
  AOI21_X1 U3808 ( .B1(n2994), .B2(n2995), .A(n3582), .ZN(n2997) );
  NAND2_X1 U3809 ( .A1(n2997), .A2(n3030), .ZN(n3002) );
  OAI22_X1 U3810 ( .A1(n2998), .A2(n3629), .B1(n3628), .B2(n3020), .ZN(n2999)
         );
  AOI211_X1 U3811 ( .C1(n3631), .C2(n3817), .A(n3000), .B(n2999), .ZN(n3001)
         );
  OAI211_X1 U3812 ( .C1(n3634), .C2(n3022), .A(n3002), .B(n3001), .ZN(U3227)
         );
  INV_X1 U3813 ( .A(n3003), .ZN(n3006) );
  NOR2_X1 U3814 ( .A1(n3004), .A2(n3745), .ZN(n3005) );
  OR2_X1 U3815 ( .A1(n3006), .A2(n3005), .ZN(n3026) );
  OAI21_X1 U3816 ( .B1(n3008), .B2(n3007), .A(n4526), .ZN(n3009) );
  NAND4_X1 U3817 ( .A1(n3012), .A2(n3011), .A3(n3010), .A4(n3009), .ZN(n3013)
         );
  OR2_X1 U3818 ( .A1(n2836), .A2(n3887), .ZN(n3041) );
  INV_X1 U3819 ( .A(n3041), .ZN(n3014) );
  AND2_X1 U3820 ( .A1(n4516), .A2(n3014), .ZN(n4520) );
  INV_X1 U3821 ( .A(n4520), .ZN(n4175) );
  INV_X1 U3822 ( .A(n3026), .ZN(n4544) );
  AOI22_X1 U3823 ( .A1(n4183), .A2(n4304), .B1(n3015), .B2(n4290), .ZN(n3016)
         );
  OAI21_X1 U3824 ( .B1(n3125), .B2(n4316), .A(n3016), .ZN(n3017) );
  AOI21_X1 U3825 ( .B1(n4544), .B2(n4162), .A(n3017), .ZN(n3018) );
  OAI21_X1 U3826 ( .B1(n4306), .B2(n3019), .A(n3018), .ZN(n4541) );
  OAI211_X1 U3827 ( .C1(n3021), .C2(n3020), .A(n3072), .B(n4285), .ZN(n4540)
         );
  OAI22_X1 U3828 ( .A1(n4540), .A2(n4412), .B1(n4513), .B2(n3022), .ZN(n3023)
         );
  OAI21_X1 U3829 ( .B1(n4541), .B2(n3023), .A(n4516), .ZN(n3025) );
  NAND2_X1 U3830 ( .A1(n4525), .A2(REG2_REG_4__SCAN_IN), .ZN(n3024) );
  OAI211_X1 U3831 ( .C1(n3026), .C2(n4175), .A(n3025), .B(n3024), .ZN(U3286)
         );
  NAND2_X1 U3832 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  OAI22_X1 U3833 ( .A1(n3125), .A2(n3504), .B1(n3503), .B2(n3036), .ZN(n3031)
         );
  XNOR2_X1 U3834 ( .A(n3031), .B(n3451), .ZN(n3113) );
  OR2_X1 U3835 ( .A1(n3125), .A2(n3506), .ZN(n3033) );
  NAND2_X1 U3836 ( .A1(n3102), .A2(n3462), .ZN(n3032) );
  NAND2_X1 U3837 ( .A1(n3033), .A2(n3032), .ZN(n3114) );
  XNOR2_X1 U3838 ( .A(n3113), .B(n3114), .ZN(n3034) );
  NAND2_X1 U3839 ( .A1(n3035), .A2(n3034), .ZN(n3117) );
  OAI211_X1 U3840 ( .C1(n3035), .C2(n3034), .A(n3117), .B(n3625), .ZN(n3040)
         );
  OAI22_X1 U3841 ( .A1(n3108), .A2(n3629), .B1(n3628), .B2(n3036), .ZN(n3037)
         );
  AOI211_X1 U3842 ( .C1(n3631), .C2(n3816), .A(n3038), .B(n3037), .ZN(n3039)
         );
  OAI211_X1 U3843 ( .C1(n3634), .C2(n3103), .A(n3040), .B(n3039), .ZN(U3224)
         );
  NAND2_X1 U3844 ( .A1(n4028), .A2(n3041), .ZN(n3042) );
  NAND2_X1 U3845 ( .A1(n4516), .A2(n3042), .ZN(n4105) );
  INV_X1 U3846 ( .A(n3043), .ZN(n3051) );
  INV_X2 U3847 ( .A(n4525), .ZN(n4516) );
  AND2_X1 U3848 ( .A1(n4285), .A2(n3887), .ZN(n3044) );
  NAND2_X1 U3849 ( .A1(n4516), .A2(n3044), .ZN(n4196) );
  NAND2_X1 U3850 ( .A1(n4516), .A2(n4290), .ZN(n4197) );
  INV_X1 U3851 ( .A(n4197), .ZN(n4182) );
  NAND2_X1 U3852 ( .A1(n4516), .A2(n4291), .ZN(n4083) );
  INV_X1 U3853 ( .A(n4083), .ZN(n4191) );
  AOI22_X1 U3854 ( .A1(n4182), .A2(n3045), .B1(n4191), .B2(n3818), .ZN(n3048)
         );
  INV_X1 U3855 ( .A(n4513), .ZN(n4180) );
  AOI22_X1 U3856 ( .A1(n4525), .A2(REG2_REG_3__SCAN_IN), .B1(n4180), .B2(n3046), .ZN(n3047) );
  OAI211_X1 U3857 ( .C1(n4196), .C2(n3049), .A(n3048), .B(n3047), .ZN(n3050)
         );
  AOI21_X1 U3858 ( .B1(n3051), .B2(n4516), .A(n3050), .ZN(n3052) );
  OAI21_X1 U3859 ( .B1(n4105), .B2(n3053), .A(n3052), .ZN(U3287) );
  NAND2_X1 U3860 ( .A1(n2834), .A2(n3054), .ZN(n3652) );
  AND2_X1 U3861 ( .A1(n3055), .A2(n3652), .ZN(n4538) );
  INV_X1 U3862 ( .A(n3056), .ZN(n3060) );
  NAND2_X1 U3863 ( .A1(n3058), .A2(n3057), .ZN(n4535) );
  AOI21_X1 U3864 ( .B1(n4306), .B2(n4028), .A(n4538), .ZN(n3059) );
  AOI21_X1 U3865 ( .B1(n4291), .B2(n2300), .A(n3059), .ZN(n4536) );
  OAI21_X1 U3866 ( .B1(n3060), .B2(n4535), .A(n4536), .ZN(n3064) );
  OAI22_X1 U3867 ( .A1(n4516), .A2(n3062), .B1(n3061), .B2(n4513), .ZN(n3063)
         );
  AOI21_X1 U3868 ( .B1(n3064), .B2(n4516), .A(n3063), .ZN(n3065) );
  OAI21_X1 U3869 ( .B1(n4538), .B2(n4175), .A(n3065), .ZN(U3290) );
  INV_X1 U3870 ( .A(n3067), .ZN(n3662) );
  AND2_X1 U3871 ( .A1(n3662), .A2(n3648), .ZN(n3743) );
  XOR2_X1 U3872 ( .A(n3066), .B(n3743), .Z(n3110) );
  XOR2_X1 U3873 ( .A(n3743), .B(n3068), .Z(n3069) );
  NAND2_X1 U3874 ( .A1(n3069), .A2(n4098), .ZN(n3112) );
  AOI22_X1 U3875 ( .A1(n3816), .A2(n4291), .B1(n4290), .B2(n3102), .ZN(n3070)
         );
  OAI211_X1 U3876 ( .C1(n3108), .C2(n4329), .A(n3112), .B(n3070), .ZN(n3071)
         );
  AOI21_X1 U3877 ( .B1(n3110), .B2(n4325), .A(n3071), .ZN(n3076) );
  AND2_X1 U3878 ( .A1(n3072), .A2(n3102), .ZN(n3073) );
  NOR2_X1 U3879 ( .A1(n3082), .A2(n3073), .ZN(n3105) );
  AOI22_X1 U3880 ( .A1(n4221), .A2(n3105), .B1(REG1_REG_5__SCAN_IN), .B2(n4557), .ZN(n3074) );
  OAI21_X1 U3881 ( .B1(n3076), .B2(n4557), .A(n3074), .ZN(U3523) );
  AOI22_X1 U3882 ( .A1(n4346), .A2(n3105), .B1(REG0_REG_5__SCAN_IN), .B2(n4551), .ZN(n3075) );
  OAI21_X1 U3883 ( .B1(n3076), .B2(n4551), .A(n3075), .ZN(U3477) );
  INV_X1 U3884 ( .A(n3077), .ZN(n3078) );
  AND2_X1 U3885 ( .A1(n3665), .A2(n3661), .ZN(n3733) );
  XNOR2_X1 U3886 ( .A(n3078), .B(n3733), .ZN(n3091) );
  AOI22_X1 U3887 ( .A1(n3815), .A2(n4291), .B1(n3119), .B2(n4290), .ZN(n3079)
         );
  OAI21_X1 U3888 ( .B1(n3125), .B2(n4329), .A(n3079), .ZN(n3080) );
  AOI21_X1 U3889 ( .B1(n3090), .B2(n4098), .A(n3080), .ZN(n3081) );
  OAI21_X1 U3890 ( .B1(n3091), .B2(n4546), .A(n3081), .ZN(n3088) );
  OR2_X1 U3891 ( .A1(n3082), .A2(n3124), .ZN(n3083) );
  NAND2_X1 U3892 ( .A1(n3166), .A2(n3083), .ZN(n3092) );
  INV_X1 U3893 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3084) );
  OAI22_X1 U3894 ( .A1(n3092), .A2(n4406), .B1(n4553), .B2(n3084), .ZN(n3085)
         );
  AOI21_X1 U3895 ( .B1(n3088), .B2(n4553), .A(n3085), .ZN(n3086) );
  INV_X1 U3896 ( .A(n3086), .ZN(U3479) );
  OAI22_X1 U3897 ( .A1(n3092), .A2(n4336), .B1(n4559), .B2(n2353), .ZN(n3087)
         );
  AOI21_X1 U3898 ( .B1(n3088), .B2(n4559), .A(n3087), .ZN(n3089) );
  INV_X1 U3899 ( .A(n3089), .ZN(U3524) );
  NAND2_X1 U3900 ( .A1(n4516), .A2(n4098), .ZN(n4136) );
  INV_X1 U3901 ( .A(n3090), .ZN(n3101) );
  INV_X1 U3902 ( .A(n3091), .ZN(n3099) );
  INV_X1 U3903 ( .A(n3092), .ZN(n3095) );
  OAI22_X1 U3904 ( .A1(n4516), .A2(n3093), .B1(n3130), .B2(n4513), .ZN(n3094)
         );
  AOI21_X1 U3905 ( .B1(n3095), .B2(n4519), .A(n3094), .ZN(n3097) );
  AOI22_X1 U3906 ( .A1(n4182), .A2(n3119), .B1(n4190), .B2(n3817), .ZN(n3096)
         );
  OAI211_X1 U3907 ( .C1(n3279), .C2(n4083), .A(n3097), .B(n3096), .ZN(n3098)
         );
  AOI21_X1 U3908 ( .B1(n3099), .B2(n4153), .A(n3098), .ZN(n3100) );
  OAI21_X1 U3909 ( .B1(n4136), .B2(n3101), .A(n3100), .ZN(U3284) );
  INV_X1 U3910 ( .A(n4190), .ZN(n4131) );
  AOI22_X1 U3911 ( .A1(n4182), .A2(n3102), .B1(n4191), .B2(n3816), .ZN(n3107)
         );
  OAI22_X1 U3912 ( .A1(n4516), .A2(n2341), .B1(n3103), .B2(n4513), .ZN(n3104)
         );
  AOI21_X1 U3913 ( .B1(n4519), .B2(n3105), .A(n3104), .ZN(n3106) );
  OAI211_X1 U3914 ( .C1(n3108), .C2(n4131), .A(n3107), .B(n3106), .ZN(n3109)
         );
  AOI21_X1 U3915 ( .B1(n3110), .B2(n4153), .A(n3109), .ZN(n3111) );
  OAI21_X1 U3916 ( .B1(n4525), .B2(n3112), .A(n3111), .ZN(U3285) );
  INV_X1 U3917 ( .A(n3113), .ZN(n3115) );
  NAND2_X1 U3918 ( .A1(n3115), .A2(n3114), .ZN(n3116) );
  NAND2_X1 U3919 ( .A1(n3117), .A2(n3116), .ZN(n3133) );
  OAI22_X1 U3920 ( .A1(n3172), .A2(n3504), .B1(n3503), .B2(n3124), .ZN(n3118)
         );
  XNOR2_X1 U3921 ( .A(n3118), .B(n3508), .ZN(n3131) );
  OR2_X1 U3922 ( .A1(n3172), .A2(n3506), .ZN(n3121) );
  NAND2_X1 U3923 ( .A1(n3119), .A2(n3462), .ZN(n3120) );
  NAND2_X1 U3924 ( .A1(n3121), .A2(n3120), .ZN(n3132) );
  XNOR2_X1 U3925 ( .A(n3131), .B(n3132), .ZN(n3122) );
  XNOR2_X1 U3926 ( .A(n3133), .B(n3122), .ZN(n3123) );
  NAND2_X1 U3927 ( .A1(n3123), .A2(n3625), .ZN(n3129) );
  OAI22_X1 U3928 ( .A1(n3125), .A2(n3629), .B1(n3628), .B2(n3124), .ZN(n3126)
         );
  AOI211_X1 U3929 ( .C1(n3631), .C2(n3815), .A(n3127), .B(n3126), .ZN(n3128)
         );
  OAI211_X1 U3930 ( .C1(n3634), .C2(n3130), .A(n3129), .B(n3128), .ZN(U3236)
         );
  OAI21_X1 U3931 ( .B1(n3133), .B2(n3132), .A(n3131), .ZN(n3135) );
  NAND2_X1 U3932 ( .A1(n3133), .A2(n3132), .ZN(n3134) );
  OAI22_X1 U3933 ( .A1(n3279), .A2(n3504), .B1(n3503), .B2(n3167), .ZN(n3136)
         );
  XNOR2_X1 U3934 ( .A(n3136), .B(n3451), .ZN(n3139) );
  OR2_X1 U3935 ( .A1(n3279), .A2(n3506), .ZN(n3138) );
  NAND2_X1 U3936 ( .A1(n3170), .A2(n3462), .ZN(n3137) );
  NAND2_X1 U3937 ( .A1(n3138), .A2(n3137), .ZN(n3140) );
  XNOR2_X1 U3938 ( .A(n3139), .B(n3140), .ZN(n3160) );
  INV_X1 U3939 ( .A(n3139), .ZN(n3141) );
  NAND2_X1 U3940 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  NAND2_X1 U3941 ( .A1(n3814), .A2(n3462), .ZN(n3144) );
  NAND2_X1 U3942 ( .A1(n3287), .A2(n3461), .ZN(n3143) );
  NAND2_X1 U3943 ( .A1(n3144), .A2(n3143), .ZN(n3145) );
  XNOR2_X1 U3944 ( .A(n3145), .B(n3508), .ZN(n3151) );
  INV_X1 U3945 ( .A(n3151), .ZN(n3149) );
  NAND2_X1 U3946 ( .A1(n3814), .A2(n3464), .ZN(n3147) );
  NAND2_X1 U3947 ( .A1(n3287), .A2(n3462), .ZN(n3146) );
  NAND2_X1 U3948 ( .A1(n3147), .A2(n3146), .ZN(n3150) );
  INV_X1 U3949 ( .A(n3150), .ZN(n3148) );
  NOR2_X1 U3950 ( .A1(n2067), .A2(n3181), .ZN(n3152) );
  XNOR2_X1 U3951 ( .A(n3182), .B(n3152), .ZN(n3158) );
  INV_X1 U3952 ( .A(n4514), .ZN(n3156) );
  AOI22_X1 U3953 ( .A1(n3595), .A2(n3287), .B1(n3617), .B2(n3815), .ZN(n3154)
         );
  OAI211_X1 U3954 ( .C1(n3272), .C2(n3578), .A(n3154), .B(n3153), .ZN(n3155)
         );
  AOI21_X1 U3955 ( .B1(n3156), .B2(n3618), .A(n3155), .ZN(n3157) );
  OAI21_X1 U3956 ( .B1(n3158), .B2(n3582), .A(n3157), .ZN(U3218) );
  XOR2_X1 U3957 ( .A(n3159), .B(n3160), .Z(n3161) );
  NAND2_X1 U3958 ( .A1(n3161), .A2(n3625), .ZN(n3165) );
  OAI22_X1 U3959 ( .A1(n3172), .A2(n3629), .B1(n3628), .B2(n3167), .ZN(n3162)
         );
  AOI211_X1 U3960 ( .C1(n3631), .C2(n3814), .A(n3163), .B(n3162), .ZN(n3164)
         );
  OAI211_X1 U3961 ( .C1(n3634), .C2(n3175), .A(n3165), .B(n3164), .ZN(U3210)
         );
  INV_X1 U3962 ( .A(n3166), .ZN(n3168) );
  OAI211_X1 U3963 ( .C1(n3168), .C2(n3167), .A(n4285), .B(n3286), .ZN(n4548)
         );
  XNOR2_X1 U3964 ( .A(n3169), .B(n3731), .ZN(n3174) );
  AOI22_X1 U3965 ( .A1(n3814), .A2(n4291), .B1(n4290), .B2(n3170), .ZN(n3171)
         );
  OAI21_X1 U3966 ( .B1(n3172), .B2(n4329), .A(n3171), .ZN(n3173) );
  AOI21_X1 U3967 ( .B1(n3174), .B2(n4098), .A(n3173), .ZN(n4549) );
  OAI21_X1 U3968 ( .B1(n4412), .B2(n4548), .A(n4549), .ZN(n3179) );
  OAI22_X1 U3969 ( .A1(n4516), .A2(n2361), .B1(n3175), .B2(n4513), .ZN(n3178)
         );
  AND2_X1 U3970 ( .A1(n3176), .A2(n3731), .ZN(n4545) );
  NOR3_X1 U3971 ( .A1(n4547), .A2(n4545), .A3(n4105), .ZN(n3177) );
  AOI211_X1 U3972 ( .C1(n4516), .C2(n3179), .A(n3178), .B(n3177), .ZN(n3180)
         );
  INV_X1 U3973 ( .A(n3180), .ZN(U3283) );
  NAND2_X1 U3974 ( .A1(n3813), .A2(n3462), .ZN(n3184) );
  NAND2_X1 U3975 ( .A1(n3251), .A2(n3461), .ZN(n3183) );
  NAND2_X1 U3976 ( .A1(n3184), .A2(n3183), .ZN(n3185) );
  XNOR2_X1 U3977 ( .A(n3185), .B(n3508), .ZN(n3237) );
  NOR2_X1 U3978 ( .A1(n3195), .A2(n3505), .ZN(n3186) );
  AOI21_X1 U3979 ( .B1(n3813), .B2(n3464), .A(n3186), .ZN(n3238) );
  XNOR2_X1 U3980 ( .A(n3237), .B(n3238), .ZN(n3235) );
  XNOR2_X1 U3981 ( .A(n3236), .B(n3235), .ZN(n3187) );
  NAND2_X1 U3982 ( .A1(n3187), .A2(n3625), .ZN(n3190) );
  AND2_X1 U3983 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4440) );
  OAI22_X1 U3984 ( .A1(n3254), .A2(n3629), .B1(n3628), .B2(n3195), .ZN(n3188)
         );
  AOI211_X1 U3985 ( .C1(n3631), .C2(n4172), .A(n4440), .B(n3188), .ZN(n3189)
         );
  OAI211_X1 U3986 ( .C1(n3634), .C2(n3197), .A(n3190), .B(n3189), .ZN(U3228)
         );
  INV_X1 U3987 ( .A(n3192), .ZN(n3676) );
  AND2_X1 U3988 ( .A1(n3676), .A2(n3671), .ZN(n3744) );
  XNOR2_X1 U3989 ( .A(n3191), .B(n3744), .ZN(n3256) );
  XOR2_X1 U3990 ( .A(n3744), .B(n3193), .Z(n3194) );
  NAND2_X1 U3991 ( .A1(n3194), .A2(n4098), .ZN(n3253) );
  NOR2_X1 U3992 ( .A1(n3253), .A2(n4525), .ZN(n3202) );
  NOR2_X1 U3993 ( .A1(n3285), .A2(n3195), .ZN(n3196) );
  OR2_X1 U3994 ( .A1(n3264), .A2(n3196), .ZN(n3257) );
  OAI22_X1 U3995 ( .A1(n3197), .A2(n4513), .B1(n3204), .B2(n4516), .ZN(n3198)
         );
  AOI21_X1 U3996 ( .B1(n4182), .B2(n3251), .A(n3198), .ZN(n3200) );
  AOI22_X1 U3997 ( .A1(n4191), .A2(n4172), .B1(n4190), .B2(n3814), .ZN(n3199)
         );
  OAI211_X1 U3998 ( .C1(n3257), .C2(n4196), .A(n3200), .B(n3199), .ZN(n3201)
         );
  AOI211_X1 U3999 ( .C1(n3256), .C2(n4153), .A(n3202), .B(n3201), .ZN(n3203)
         );
  INV_X1 U4000 ( .A(n3203), .ZN(U3281) );
  NOR2_X1 U4001 ( .A1(n3232), .A2(n4150), .ZN(n3857) );
  AOI21_X1 U4002 ( .B1(n4150), .B2(n3232), .A(n3857), .ZN(n3213) );
  NAND2_X1 U4003 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3214), .ZN(n3209) );
  INV_X1 U4004 ( .A(n3214), .ZN(n4533) );
  AOI22_X1 U4005 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3214), .B1(n4533), .B2(
        n4166), .ZN(n4456) );
  NAND2_X1 U4006 ( .A1(n3215), .A2(REG2_REG_9__SCAN_IN), .ZN(n3206) );
  MUX2_X1 U4007 ( .A(REG2_REG_9__SCAN_IN), .B(n3204), .S(n3215), .Z(n4431) );
  NAND2_X1 U4008 ( .A1(n4431), .A2(n4432), .ZN(n4430) );
  NAND2_X1 U4009 ( .A1(n3222), .A2(n3207), .ZN(n3208) );
  NAND2_X1 U4010 ( .A1(n4462), .A2(n3210), .ZN(n3211) );
  OAI21_X1 U4011 ( .B1(n3213), .B2(n3858), .A(n4464), .ZN(n3212) );
  AOI21_X1 U4012 ( .B1(n3213), .B2(n3858), .A(n3212), .ZN(n3234) );
  NAND2_X1 U4013 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3214), .ZN(n3225) );
  AOI22_X1 U4014 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3214), .B1(n4533), .B2(
        n4334), .ZN(n4453) );
  NAND2_X1 U4015 ( .A1(n3215), .A2(REG1_REG_9__SCAN_IN), .ZN(n3221) );
  MUX2_X1 U4016 ( .A(n2386), .B(REG1_REG_9__SCAN_IN), .S(n3215), .Z(n3216) );
  INV_X1 U4017 ( .A(n3216), .ZN(n4434) );
  OAI22_X1 U4018 ( .A1(n3220), .A2(n3219), .B1(n3218), .B2(n3217), .ZN(n4435)
         );
  NAND2_X1 U4019 ( .A1(n4434), .A2(n4435), .ZN(n4433) );
  NAND2_X1 U4020 ( .A1(n3221), .A2(n4433), .ZN(n3223) );
  NAND2_X1 U4021 ( .A1(n3222), .A2(n3223), .ZN(n3224) );
  XOR2_X1 U4022 ( .A(n3223), .B(n3222), .Z(n4448) );
  NAND2_X1 U4023 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4448), .ZN(n4447) );
  NAND2_X1 U4024 ( .A1(n4462), .A2(n3226), .ZN(n3227) );
  NAND2_X1 U4025 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4470), .ZN(n4469) );
  NOR2_X1 U4026 ( .A1(n3232), .A2(n4314), .ZN(n3842) );
  AOI21_X1 U4027 ( .B1(n4314), .B2(n3232), .A(n3842), .ZN(n3228) );
  OAI211_X1 U4028 ( .C1(n3229), .C2(n3228), .A(n4507), .B(n3843), .ZN(n3231)
         );
  NOR2_X1 U4029 ( .A1(STATE_REG_SCAN_IN), .A2(n2435), .ZN(n3590) );
  AOI21_X1 U4030 ( .B1(n4505), .B2(ADDR_REG_13__SCAN_IN), .A(n3590), .ZN(n3230) );
  OAI211_X1 U4031 ( .C1(n4512), .C2(n3232), .A(n3231), .B(n3230), .ZN(n3233)
         );
  OR2_X1 U4032 ( .A1(n3234), .A2(n3233), .ZN(U3253) );
  INV_X1 U4033 ( .A(n3237), .ZN(n3239) );
  OAI22_X1 U4034 ( .A1(n4330), .A2(n3505), .B1(n3503), .B2(n3294), .ZN(n3240)
         );
  XNOR2_X1 U4035 ( .A(n3240), .B(n3508), .ZN(n3305) );
  OR2_X1 U4036 ( .A1(n4330), .A2(n3506), .ZN(n3242) );
  NAND2_X1 U4037 ( .A1(n3267), .A2(n3462), .ZN(n3241) );
  NAND2_X1 U4038 ( .A1(n3242), .A2(n3241), .ZN(n3304) );
  XNOR2_X1 U4039 ( .A(n3305), .B(n3304), .ZN(n3244) );
  AOI21_X1 U4040 ( .B1(n3243), .B2(n3244), .A(n3582), .ZN(n3246) );
  NAND2_X1 U4041 ( .A1(n3246), .A2(n3307), .ZN(n3250) );
  NAND2_X1 U4042 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4444) );
  INV_X1 U40430 ( .A(n4444), .ZN(n3248) );
  OAI22_X1 U4044 ( .A1(n3272), .A2(n3629), .B1(n3628), .B2(n3294), .ZN(n3247)
         );
  AOI211_X1 U4045 ( .C1(n3631), .C2(n3812), .A(n3248), .B(n3247), .ZN(n3249)
         );
  OAI211_X1 U4046 ( .C1(n3634), .C2(n3268), .A(n3250), .B(n3249), .ZN(U3214)
         );
  AOI22_X1 U4047 ( .A1(n4172), .A2(n4291), .B1(n4290), .B2(n3251), .ZN(n3252)
         );
  OAI211_X1 U4048 ( .C1(n3254), .C2(n4329), .A(n3253), .B(n3252), .ZN(n3255)
         );
  AOI21_X1 U4049 ( .B1(n3256), .B2(n4325), .A(n3255), .ZN(n3261) );
  INV_X1 U4050 ( .A(n3257), .ZN(n3259) );
  AOI22_X1 U4051 ( .A1(n3259), .A2(n4346), .B1(REG0_REG_9__SCAN_IN), .B2(n4551), .ZN(n3258) );
  OAI21_X1 U4052 ( .B1(n3261), .B2(n4551), .A(n3258), .ZN(U3485) );
  AOI22_X1 U4053 ( .A1(n3259), .A2(n4221), .B1(REG1_REG_9__SCAN_IN), .B2(n4557), .ZN(n3260) );
  OAI21_X1 U4054 ( .B1(n3261), .B2(n4557), .A(n3260), .ZN(U3527) );
  AND2_X1 U4055 ( .A1(n3645), .A2(n3678), .ZN(n3742) );
  XOR2_X1 U4056 ( .A(n3742), .B(n3262), .Z(n3297) );
  XNOR2_X1 U4057 ( .A(n3263), .B(n3742), .ZN(n3299) );
  NAND2_X1 U4058 ( .A1(n3299), .A2(n4153), .ZN(n3275) );
  INV_X1 U4059 ( .A(n3264), .ZN(n3266) );
  INV_X1 U4060 ( .A(n3265), .ZN(n4169) );
  AOI21_X1 U4061 ( .B1(n3267), .B2(n3266), .A(n4169), .ZN(n3301) );
  AOI22_X1 U4062 ( .A1(n4182), .A2(n3267), .B1(n4191), .B2(n3812), .ZN(n3271)
         );
  INV_X1 U4063 ( .A(n3268), .ZN(n3269) );
  AOI22_X1 U4064 ( .A1(n4525), .A2(REG2_REG_10__SCAN_IN), .B1(n3269), .B2(
        n4180), .ZN(n3270) );
  OAI211_X1 U4065 ( .C1(n3272), .C2(n4131), .A(n3271), .B(n3270), .ZN(n3273)
         );
  AOI21_X1 U4066 ( .B1(n3301), .B2(n4519), .A(n3273), .ZN(n3274) );
  OAI211_X1 U4067 ( .C1(n3297), .C2(n4136), .A(n3275), .B(n3274), .ZN(U3280)
         );
  INV_X1 U4068 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3290) );
  AND2_X1 U4069 ( .A1(n3670), .A2(n3667), .ZN(n3734) );
  XOR2_X1 U4070 ( .A(n3276), .B(n3734), .Z(n4521) );
  INV_X1 U4071 ( .A(n4521), .ZN(n3284) );
  XNOR2_X1 U4072 ( .A(n3277), .B(n3734), .ZN(n3282) );
  OAI22_X1 U4073 ( .A1(n3279), .A2(n4329), .B1(n3278), .B2(n4323), .ZN(n3280)
         );
  AOI21_X1 U4074 ( .B1(n4291), .B2(n3813), .A(n3280), .ZN(n3281) );
  OAI21_X1 U4075 ( .B1(n3282), .B2(n4306), .A(n3281), .ZN(n3283) );
  AOI21_X1 U4076 ( .B1(n4521), .B2(n4162), .A(n3283), .ZN(n4524) );
  OAI21_X1 U4077 ( .B1(n4537), .B2(n3284), .A(n4524), .ZN(n3291) );
  NAND2_X1 U4078 ( .A1(n3291), .A2(n4553), .ZN(n3289) );
  AOI21_X1 U4079 ( .B1(n3287), .B2(n3286), .A(n3285), .ZN(n4518) );
  NAND2_X1 U4080 ( .A1(n4518), .A2(n4346), .ZN(n3288) );
  OAI211_X1 U4081 ( .C1(n4553), .C2(n3290), .A(n3289), .B(n3288), .ZN(U3483)
         );
  NAND2_X1 U4082 ( .A1(n3291), .A2(n4559), .ZN(n3293) );
  NAND2_X1 U4083 ( .A1(n4518), .A2(n4221), .ZN(n3292) );
  OAI211_X1 U4084 ( .C1(n4559), .C2(n3217), .A(n3293), .B(n3292), .ZN(U3526)
         );
  OAI22_X1 U4085 ( .A1(n4318), .A2(n4316), .B1(n4323), .B2(n3294), .ZN(n3295)
         );
  AOI21_X1 U4086 ( .B1(n4304), .B2(n3813), .A(n3295), .ZN(n3296) );
  OAI21_X1 U4087 ( .B1(n3297), .B2(n4306), .A(n3296), .ZN(n3298) );
  AOI21_X1 U4088 ( .B1(n3299), .B2(n4325), .A(n3298), .ZN(n3303) );
  AOI22_X1 U4089 ( .A1(n3301), .A2(n4346), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4551), .ZN(n3300) );
  OAI21_X1 U4090 ( .B1(n3303), .B2(n4551), .A(n3300), .ZN(U3487) );
  AOI22_X1 U4091 ( .A1(n3301), .A2(n4221), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4557), .ZN(n3302) );
  OAI21_X1 U4092 ( .B1(n3303), .B2(n4557), .A(n3302), .ZN(U3528) );
  NAND2_X1 U4093 ( .A1(n3305), .A2(n3304), .ZN(n3306) );
  NAND2_X1 U4094 ( .A1(n3307), .A2(n3306), .ZN(n3319) );
  OAI22_X1 U4095 ( .A1(n4318), .A2(n3505), .B1(n3503), .B2(n4168), .ZN(n3308)
         );
  XNOR2_X1 U4096 ( .A(n3308), .B(n3508), .ZN(n3317) );
  OR2_X1 U4097 ( .A1(n4318), .A2(n3506), .ZN(n3311) );
  NAND2_X1 U4098 ( .A1(n3309), .A2(n3462), .ZN(n3310) );
  NAND2_X1 U4099 ( .A1(n3311), .A2(n3310), .ZN(n3318) );
  XNOR2_X1 U4100 ( .A(n3317), .B(n3318), .ZN(n3312) );
  XNOR2_X1 U4101 ( .A(n3319), .B(n3312), .ZN(n3313) );
  NAND2_X1 U4102 ( .A1(n3313), .A2(n3625), .ZN(n3316) );
  AND2_X1 U4103 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4460) );
  OAI22_X1 U4104 ( .A1(n4330), .A2(n3629), .B1(n3628), .B2(n4168), .ZN(n3314)
         );
  AOI211_X1 U4105 ( .C1(n3631), .C2(n4141), .A(n4460), .B(n3314), .ZN(n3315)
         );
  OAI211_X1 U4106 ( .C1(n3634), .C2(n4165), .A(n3316), .B(n3315), .ZN(U3233)
         );
  OAI21_X1 U4107 ( .B1(n3319), .B2(n3318), .A(n3317), .ZN(n3321) );
  NAND2_X1 U4108 ( .A1(n3319), .A2(n3318), .ZN(n3320) );
  NAND2_X1 U4109 ( .A1(n4141), .A2(n3462), .ZN(n3323) );
  NAND2_X1 U4110 ( .A1(n3346), .A2(n3461), .ZN(n3322) );
  NAND2_X1 U4111 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  XNOR2_X1 U4112 ( .A(n3324), .B(n3508), .ZN(n3330) );
  INV_X1 U4113 ( .A(n3330), .ZN(n3328) );
  NAND2_X1 U4114 ( .A1(n4141), .A2(n3464), .ZN(n3326) );
  NAND2_X1 U4115 ( .A1(n3346), .A2(n3462), .ZN(n3325) );
  NAND2_X1 U4116 ( .A1(n3326), .A2(n3325), .ZN(n3329) );
  INV_X1 U4117 ( .A(n3329), .ZN(n3327) );
  NAND2_X1 U4118 ( .A1(n3328), .A2(n3327), .ZN(n3375) );
  NOR2_X1 U4119 ( .A1(n2174), .A2(n3376), .ZN(n3331) );
  XNOR2_X1 U4120 ( .A(n3377), .B(n3331), .ZN(n3336) );
  INV_X1 U4121 ( .A(n3343), .ZN(n3334) );
  AOI22_X1 U4122 ( .A1(n3595), .A2(n3346), .B1(n3617), .B2(n3812), .ZN(n3332)
         );
  NAND2_X1 U4123 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4466) );
  OAI211_X1 U4124 ( .C1(n4317), .C2(n3578), .A(n3332), .B(n4466), .ZN(n3333)
         );
  AOI21_X1 U4125 ( .B1(n3334), .B2(n3618), .A(n3333), .ZN(n3335) );
  OAI21_X1 U4126 ( .B1(n3336), .B2(n3582), .A(n3335), .ZN(U3221) );
  INV_X1 U4127 ( .A(n4137), .ZN(n3337) );
  OR2_X1 U4128 ( .A1(n3337), .A2(n4138), .ZN(n3340) );
  XNOR2_X1 U4129 ( .A(n3338), .B(n3340), .ZN(n4326) );
  INV_X1 U4130 ( .A(n3340), .ZN(n3732) );
  XNOR2_X1 U4131 ( .A(n3339), .B(n3732), .ZN(n3341) );
  NAND2_X1 U4132 ( .A1(n3341), .A2(n4098), .ZN(n4321) );
  NOR2_X1 U4133 ( .A1(n4321), .A2(n4525), .ZN(n3350) );
  AND2_X1 U4134 ( .A1(n4167), .A2(n3346), .ZN(n3342) );
  OR2_X1 U4135 ( .A1(n3342), .A2(n4146), .ZN(n4402) );
  OAI22_X1 U4136 ( .A1(n4516), .A2(n3344), .B1(n3343), .B2(n4513), .ZN(n3345)
         );
  AOI21_X1 U4137 ( .B1(n3346), .B2(n4182), .A(n3345), .ZN(n3348) );
  AOI22_X1 U4138 ( .A1(n4191), .A2(n4303), .B1(n4190), .B2(n3812), .ZN(n3347)
         );
  OAI211_X1 U4139 ( .C1(n4402), .C2(n4196), .A(n3348), .B(n3347), .ZN(n3349)
         );
  AOI211_X1 U4140 ( .C1(n4326), .C2(n4153), .A(n3350), .B(n3349), .ZN(n3351)
         );
  INV_X1 U4141 ( .A(n3351), .ZN(U3278) );
  INV_X1 U4142 ( .A(n3353), .ZN(n3362) );
  INV_X1 U4143 ( .A(n3807), .ZN(n3644) );
  INV_X1 U4144 ( .A(n3516), .ZN(n3356) );
  INV_X1 U4145 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3354) );
  OAI22_X1 U4146 ( .A1(n4197), .A2(n3515), .B1(n3354), .B2(n4516), .ZN(n3355)
         );
  AOI21_X1 U4147 ( .B1(n3356), .B2(n4180), .A(n3355), .ZN(n3358) );
  NAND2_X1 U4148 ( .A1(n3919), .A2(n4190), .ZN(n3357) );
  OAI211_X1 U4149 ( .C1(n3644), .C2(n4083), .A(n3358), .B(n3357), .ZN(n3361)
         );
  NOR2_X1 U4150 ( .A1(n3359), .A2(n4525), .ZN(n3360) );
  AOI211_X1 U4151 ( .C1(n4519), .C2(n3362), .A(n3361), .B(n3360), .ZN(n3363)
         );
  OAI21_X1 U4152 ( .B1(n3352), .B2(n4105), .A(n3363), .ZN(U3262) );
  XNOR2_X1 U4153 ( .A(n3364), .B(n3787), .ZN(n4219) );
  AOI21_X1 U4154 ( .B1(n4213), .B2(n3922), .A(n3365), .ZN(n4347) );
  AOI22_X1 U4155 ( .A1(n4182), .A2(n4213), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4525), .ZN(n3366) );
  OAI21_X1 U4156 ( .B1(n3467), .B2(n4513), .A(n3366), .ZN(n3367) );
  AOI21_X1 U4157 ( .B1(n4190), .B2(n3808), .A(n3367), .ZN(n3368) );
  OAI21_X1 U4158 ( .B1(n3507), .B2(n4083), .A(n3368), .ZN(n3373) );
  OAI21_X1 U4159 ( .B1(n3787), .B2(n3370), .A(n3369), .ZN(n3371) );
  NAND2_X1 U4160 ( .A1(n3371), .A2(n4098), .ZN(n4217) );
  NOR2_X1 U4161 ( .A1(n4217), .A2(n4525), .ZN(n3372) );
  AOI211_X1 U4162 ( .C1(n4519), .C2(n4347), .A(n3373), .B(n3372), .ZN(n3374)
         );
  OAI21_X1 U4163 ( .B1(n4219), .B2(n4105), .A(n3374), .ZN(U3263) );
  OAI22_X1 U4164 ( .A1(n4317), .A2(n3505), .B1(n3503), .B2(n4145), .ZN(n3378)
         );
  XNOR2_X1 U4165 ( .A(n3378), .B(n3451), .ZN(n3585) );
  OR2_X1 U4166 ( .A1(n4317), .A2(n3506), .ZN(n3381) );
  NAND2_X1 U4167 ( .A1(n3379), .A2(n3462), .ZN(n3380) );
  NAND2_X1 U4168 ( .A1(n3381), .A2(n3380), .ZN(n3584) );
  OAI22_X1 U4169 ( .A1(n4295), .A2(n3505), .B1(n3503), .B2(n4300), .ZN(n3382)
         );
  XNOR2_X1 U4170 ( .A(n3382), .B(n3508), .ZN(n3385) );
  OR2_X1 U4171 ( .A1(n4295), .A2(n3506), .ZN(n3384) );
  NAND2_X1 U4172 ( .A1(n4127), .A2(n3462), .ZN(n3383) );
  NAND2_X1 U4173 ( .A1(n3384), .A2(n3383), .ZN(n3386) );
  AND2_X1 U4174 ( .A1(n3385), .A2(n3386), .ZN(n3473) );
  INV_X1 U4175 ( .A(n3385), .ZN(n3388) );
  INV_X1 U4176 ( .A(n3386), .ZN(n3387) );
  NAND2_X1 U4177 ( .A1(n3388), .A2(n3387), .ZN(n3472) );
  OAI22_X1 U4178 ( .A1(n4301), .A2(n3505), .B1(n3503), .B2(n4118), .ZN(n3389)
         );
  XNOR2_X1 U4179 ( .A(n3389), .B(n3451), .ZN(n3393) );
  OR2_X1 U4180 ( .A1(n4301), .A2(n3506), .ZN(n3391) );
  NAND2_X1 U4181 ( .A1(n2467), .A2(n3462), .ZN(n3390) );
  NAND2_X1 U4182 ( .A1(n3391), .A2(n3390), .ZN(n3623) );
  OAI22_X1 U4183 ( .A1(n4084), .A2(n3504), .B1(n3503), .B2(n4097), .ZN(n3394)
         );
  XNOR2_X1 U4184 ( .A(n3394), .B(n3508), .ZN(n3397) );
  OAI22_X1 U4185 ( .A1(n4084), .A2(n3506), .B1(n3505), .B2(n4097), .ZN(n3396)
         );
  XNOR2_X1 U4186 ( .A(n3397), .B(n3396), .ZN(n3543) );
  INV_X1 U4187 ( .A(n3396), .ZN(n3399) );
  INV_X1 U4188 ( .A(n3397), .ZN(n3398) );
  OAI22_X1 U4189 ( .A1(n2498), .A2(n3505), .B1(n3503), .B2(n2497), .ZN(n3401)
         );
  XOR2_X1 U4190 ( .A(n3508), .B(n3401), .Z(n3553) );
  NOR2_X1 U4191 ( .A1(n2497), .A2(n3505), .ZN(n3402) );
  AOI21_X1 U4192 ( .B1(n4282), .B2(n3464), .A(n3402), .ZN(n3403) );
  INV_X1 U4193 ( .A(n3553), .ZN(n3404) );
  INV_X1 U4194 ( .A(n3403), .ZN(n3552) );
  OAI21_X1 U4195 ( .B1(n3550), .B2(n2063), .A(n3405), .ZN(n3406) );
  OAI22_X1 U4196 ( .A1(n4277), .A2(n3505), .B1(n3503), .B2(n4058), .ZN(n3407)
         );
  XNOR2_X1 U4197 ( .A(n3407), .B(n3451), .ZN(n3412) );
  INV_X1 U4198 ( .A(n3412), .ZN(n3410) );
  NOR2_X1 U4199 ( .A1(n4058), .A2(n3505), .ZN(n3408) );
  AOI21_X1 U4200 ( .B1(n3811), .B2(n3464), .A(n3408), .ZN(n3411) );
  INV_X1 U4201 ( .A(n3411), .ZN(n3409) );
  AND2_X1 U4202 ( .A1(n3412), .A2(n3411), .ZN(n3602) );
  NAND2_X1 U4203 ( .A1(n4022), .A2(n3462), .ZN(n3414) );
  NAND2_X1 U4204 ( .A1(n3494), .A2(n3461), .ZN(n3413) );
  NAND2_X1 U4205 ( .A1(n3414), .A2(n3413), .ZN(n3415) );
  XNOR2_X1 U4206 ( .A(n3415), .B(n3508), .ZN(n3416) );
  OAI22_X1 U4207 ( .A1(n4062), .A2(n3506), .B1(n3505), .B2(n4050), .ZN(n3417)
         );
  XNOR2_X1 U4208 ( .A(n3416), .B(n3417), .ZN(n3493) );
  NAND2_X1 U4209 ( .A1(n4255), .A2(n3462), .ZN(n3422) );
  NAND2_X1 U4210 ( .A1(n3461), .A2(n4030), .ZN(n3421) );
  NAND2_X1 U4211 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  XNOR2_X1 U4212 ( .A(n3423), .B(n3451), .ZN(n3426) );
  NOR2_X1 U4213 ( .A1(n3505), .A2(n3577), .ZN(n3424) );
  AOI21_X1 U4214 ( .B1(n4255), .B2(n3464), .A(n3424), .ZN(n3425) );
  OR2_X1 U4215 ( .A1(n3426), .A2(n3425), .ZN(n3572) );
  NAND2_X1 U4216 ( .A1(n3426), .A2(n3425), .ZN(n3574) );
  NAND2_X1 U4217 ( .A1(n3570), .A2(n3574), .ZN(n3521) );
  NAND2_X1 U4218 ( .A1(n3984), .A2(n3462), .ZN(n3428) );
  INV_X1 U4219 ( .A(n4009), .ZN(n4254) );
  NAND2_X1 U4220 ( .A1(n3461), .A2(n4254), .ZN(n3427) );
  NAND2_X1 U4221 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U4222 ( .A(n3429), .B(n3451), .ZN(n3523) );
  NOR2_X1 U4223 ( .A1(n3505), .A2(n4009), .ZN(n3430) );
  AOI21_X1 U4224 ( .B1(n3984), .B2(n3464), .A(n3430), .ZN(n3522) );
  INV_X1 U4225 ( .A(n3523), .ZN(n3432) );
  INV_X1 U4226 ( .A(n3522), .ZN(n3431) );
  OAI22_X1 U4227 ( .A1(n4258), .A2(n3506), .B1(n3505), .B2(n3994), .ZN(n3437)
         );
  OAI22_X1 U4228 ( .A1(n4258), .A2(n3505), .B1(n3503), .B2(n3994), .ZN(n3434)
         );
  XNOR2_X1 U4229 ( .A(n3434), .B(n3508), .ZN(n3436) );
  XOR2_X1 U4230 ( .A(n3437), .B(n3436), .Z(n3594) );
  OAI22_X1 U4231 ( .A1(n3987), .A2(n3505), .B1(n3503), .B2(n3975), .ZN(n3435)
         );
  XNOR2_X1 U4232 ( .A(n3435), .B(n3451), .ZN(n3443) );
  OAI22_X1 U4233 ( .A1(n3987), .A2(n3506), .B1(n3505), .B2(n3975), .ZN(n3444)
         );
  XNOR2_X1 U4234 ( .A(n3443), .B(n3444), .ZN(n3483) );
  INV_X1 U4235 ( .A(n3436), .ZN(n3439) );
  INV_X1 U4236 ( .A(n3437), .ZN(n3438) );
  NAND2_X1 U4237 ( .A1(n3439), .A2(n3438), .ZN(n3484) );
  OR2_X1 U4238 ( .A1(n3486), .A2(n3506), .ZN(n3442) );
  NAND2_X1 U4239 ( .A1(n3462), .A2(n4236), .ZN(n3441) );
  AND2_X1 U4240 ( .A1(n3442), .A2(n3441), .ZN(n3447) );
  INV_X1 U4241 ( .A(n3443), .ZN(n3445) );
  NAND2_X1 U4242 ( .A1(n3445), .A2(n3444), .ZN(n3448) );
  NAND3_X1 U4243 ( .A1(n3481), .A2(n3447), .A3(n3448), .ZN(n3560) );
  OAI22_X1 U4244 ( .A1(n3486), .A2(n3505), .B1(n3503), .B2(n3954), .ZN(n3446)
         );
  XNOR2_X1 U4245 ( .A(n3446), .B(n3508), .ZN(n3563) );
  NAND2_X1 U4246 ( .A1(n3809), .A2(n3462), .ZN(n3450) );
  NAND2_X1 U4247 ( .A1(n3461), .A2(n4227), .ZN(n3449) );
  NAND2_X1 U4248 ( .A1(n3450), .A2(n3449), .ZN(n3452) );
  XNOR2_X1 U4249 ( .A(n3452), .B(n3451), .ZN(n3455) );
  NOR2_X1 U4250 ( .A1(n3505), .A2(n3937), .ZN(n3453) );
  AOI21_X1 U4251 ( .B1(n3809), .B2(n3464), .A(n3453), .ZN(n3454) );
  AND2_X1 U4252 ( .A1(n3455), .A2(n3454), .ZN(n3531) );
  OR2_X1 U4253 ( .A1(n3455), .A2(n3454), .ZN(n3532) );
  OAI22_X1 U4254 ( .A1(n4231), .A2(n3504), .B1(n3503), .B2(n3923), .ZN(n3456)
         );
  XNOR2_X1 U4255 ( .A(n3456), .B(n3508), .ZN(n3457) );
  OAI22_X1 U4256 ( .A1(n4231), .A2(n3506), .B1(n3505), .B2(n3923), .ZN(n3458)
         );
  AND2_X1 U4257 ( .A1(n3457), .A2(n3458), .ZN(n3609) );
  INV_X1 U4258 ( .A(n3457), .ZN(n3460) );
  INV_X1 U4259 ( .A(n3458), .ZN(n3459) );
  NAND2_X1 U4260 ( .A1(n3460), .A2(n3459), .ZN(n3610) );
  AOI22_X1 U4261 ( .A1(n3919), .A2(n3462), .B1(n4213), .B2(n3461), .ZN(n3463)
         );
  XNOR2_X1 U4262 ( .A(n3463), .B(n3508), .ZN(n3499) );
  AOI22_X1 U4263 ( .A1(n3919), .A2(n3464), .B1(n4213), .B2(n3462), .ZN(n3500)
         );
  XNOR2_X1 U4264 ( .A(n3499), .B(n3500), .ZN(n3501) );
  XNOR2_X1 U4265 ( .A(n3502), .B(n3501), .ZN(n3470) );
  NAND2_X1 U4266 ( .A1(n3808), .A2(n3617), .ZN(n3466) );
  AOI22_X1 U4267 ( .A1(n3595), .A2(n4213), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3465) );
  OAI211_X1 U4268 ( .C1(n3634), .C2(n3467), .A(n3466), .B(n3465), .ZN(n3468)
         );
  AOI21_X1 U4269 ( .B1(n4216), .B2(n3631), .A(n3468), .ZN(n3469) );
  OAI21_X1 U4270 ( .B1(n3470), .B2(n3582), .A(n3469), .ZN(U3211) );
  INV_X1 U4271 ( .A(n3472), .ZN(n3474) );
  NOR2_X1 U4272 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  XNOR2_X1 U4273 ( .A(n3471), .B(n3475), .ZN(n3480) );
  INV_X1 U4274 ( .A(n3476), .ZN(n4128) );
  AOI22_X1 U4275 ( .A1(n3595), .A2(n4127), .B1(n3617), .B2(n4303), .ZN(n3477)
         );
  NAND2_X1 U4276 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4473) );
  OAI211_X1 U4277 ( .C1(n4301), .C2(n3578), .A(n3477), .B(n4473), .ZN(n3478)
         );
  AOI21_X1 U4278 ( .B1(n4128), .B2(n3618), .A(n3478), .ZN(n3479) );
  OAI21_X1 U4279 ( .B1(n3480), .B2(n3582), .A(n3479), .ZN(U3212) );
  NAND2_X1 U4280 ( .A1(n3481), .A2(n3625), .ZN(n3491) );
  AOI21_X1 U4281 ( .B1(n3482), .B2(n3484), .A(n3483), .ZN(n3490) );
  INV_X1 U4282 ( .A(n3485), .ZN(n3977) );
  OAI22_X1 U4283 ( .A1(n4258), .A2(n3629), .B1(STATE_REG_SCAN_IN), .B2(n4565), 
        .ZN(n3488) );
  OAI22_X1 U4284 ( .A1(n3486), .A2(n3578), .B1(n3628), .B2(n3975), .ZN(n3487)
         );
  AOI211_X1 U4285 ( .C1(n3977), .C2(n3618), .A(n3488), .B(n3487), .ZN(n3489)
         );
  OAI21_X1 U4286 ( .B1(n3491), .B2(n3490), .A(n3489), .ZN(U3213) );
  XOR2_X1 U4287 ( .A(n3493), .B(n3492), .Z(n3498) );
  INV_X1 U4288 ( .A(n4255), .ZN(n4010) );
  AOI22_X1 U4289 ( .A1(n3595), .A2(n3494), .B1(n3811), .B2(n3617), .ZN(n3495)
         );
  NAND2_X1 U4290 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3886) );
  OAI211_X1 U4291 ( .C1(n4010), .C2(n3578), .A(n3495), .B(n3886), .ZN(n3496)
         );
  AOI21_X1 U4292 ( .B1(n4052), .B2(n3618), .A(n3496), .ZN(n3497) );
  OAI21_X1 U4293 ( .B1(n3498), .B2(n3582), .A(n3497), .ZN(U3216) );
  OAI22_X1 U4294 ( .A1(n3507), .A2(n3504), .B1(n3503), .B2(n3515), .ZN(n3511)
         );
  OAI22_X1 U4295 ( .A1(n3507), .A2(n3506), .B1(n3505), .B2(n3515), .ZN(n3509)
         );
  XNOR2_X1 U4296 ( .A(n3509), .B(n3508), .ZN(n3510) );
  XOR2_X1 U4297 ( .A(n3511), .B(n3510), .Z(n3512) );
  XNOR2_X1 U4298 ( .A(n3513), .B(n3512), .ZN(n3520) );
  OAI22_X1 U4299 ( .A1(n3628), .A2(n3515), .B1(STATE_REG_SCAN_IN), .B2(n3514), 
        .ZN(n3518) );
  OAI22_X1 U4300 ( .A1(n3644), .A2(n3578), .B1(n3634), .B2(n3516), .ZN(n3517)
         );
  AOI211_X1 U4301 ( .C1(n3617), .C2(n3919), .A(n3518), .B(n3517), .ZN(n3519)
         );
  OAI21_X1 U4302 ( .B1(n3520), .B2(n3582), .A(n3519), .ZN(U3217) );
  XNOR2_X1 U4303 ( .A(n3523), .B(n3522), .ZN(n3524) );
  XNOR2_X1 U4304 ( .A(n3521), .B(n3524), .ZN(n3529) );
  OAI22_X1 U4305 ( .A1(n4010), .A2(n3629), .B1(n3628), .B2(n4009), .ZN(n3527)
         );
  OAI22_X1 U4306 ( .A1(n4258), .A2(n3578), .B1(STATE_REG_SCAN_IN), .B2(n3525), 
        .ZN(n3526) );
  AOI211_X1 U4307 ( .C1(n4007), .C2(n3618), .A(n3527), .B(n3526), .ZN(n3528)
         );
  OAI21_X1 U4308 ( .B1(n3529), .B2(n3582), .A(n3528), .ZN(U3220) );
  INV_X1 U4309 ( .A(n3531), .ZN(n3533) );
  NAND2_X1 U4310 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  XNOR2_X1 U4311 ( .A(n3530), .B(n3534), .ZN(n3539) );
  NOR2_X1 U4312 ( .A1(n3939), .A2(n3634), .ZN(n3537) );
  AOI22_X1 U4313 ( .A1(n4228), .A2(n3617), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3535) );
  OAI21_X1 U4314 ( .B1(n3628), .B2(n3937), .A(n3535), .ZN(n3536) );
  AOI211_X1 U4315 ( .C1(n3631), .C2(n3808), .A(n3537), .B(n3536), .ZN(n3538)
         );
  OAI21_X1 U4316 ( .B1(n3539), .B2(n3582), .A(n3538), .ZN(U3222) );
  INV_X1 U4317 ( .A(n3540), .ZN(n3542) );
  OAI21_X1 U4318 ( .B1(n3542), .B2(n3623), .A(n3541), .ZN(n3544) );
  XNOR2_X1 U4319 ( .A(n3544), .B(n3543), .ZN(n3549) );
  INV_X1 U4320 ( .A(n3545), .ZN(n4094) );
  AOI22_X1 U4321 ( .A1(n3595), .A2(n4281), .B1(n3617), .B2(n2468), .ZN(n3546)
         );
  NAND2_X1 U4322 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4492) );
  OAI211_X1 U4323 ( .C1(n2498), .C2(n3578), .A(n3546), .B(n4492), .ZN(n3547)
         );
  AOI21_X1 U4324 ( .B1(n4094), .B2(n3618), .A(n3547), .ZN(n3548) );
  OAI21_X1 U4325 ( .B1(n3549), .B2(n3582), .A(n3548), .ZN(U3223) );
  XNOR2_X1 U4326 ( .A(n3553), .B(n3552), .ZN(n3554) );
  XNOR2_X1 U4327 ( .A(n3551), .B(n3554), .ZN(n3559) );
  INV_X1 U4328 ( .A(n3555), .ZN(n4081) );
  AOI22_X1 U4329 ( .A1(n3595), .A2(n4274), .B1(n3617), .B2(n4292), .ZN(n3556)
         );
  NAND2_X1 U4330 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3868) );
  OAI211_X1 U4331 ( .C1(n4277), .C2(n3578), .A(n3556), .B(n3868), .ZN(n3557)
         );
  AOI21_X1 U4332 ( .B1(n4081), .B2(n3618), .A(n3557), .ZN(n3558) );
  OAI21_X1 U4333 ( .B1(n3559), .B2(n3582), .A(n3558), .ZN(U3225) );
  INV_X1 U4334 ( .A(n3560), .ZN(n3561) );
  NOR2_X1 U4335 ( .A1(n3562), .A2(n3561), .ZN(n3564) );
  XNOR2_X1 U4336 ( .A(n3564), .B(n3563), .ZN(n3569) );
  NOR2_X1 U4337 ( .A1(n3957), .A2(n3634), .ZN(n3567) );
  AOI22_X1 U4338 ( .A1(n4237), .A2(n3617), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3565) );
  OAI21_X1 U4339 ( .B1(n3628), .B2(n3954), .A(n3565), .ZN(n3566) );
  AOI211_X1 U4340 ( .C1(n3631), .C2(n3809), .A(n3567), .B(n3566), .ZN(n3568)
         );
  OAI21_X1 U4341 ( .B1(n3569), .B2(n3582), .A(n3568), .ZN(U3226) );
  INV_X1 U4342 ( .A(n3570), .ZN(n3575) );
  AOI21_X1 U4343 ( .B1(n3574), .B2(n3572), .A(n3571), .ZN(n3573) );
  AOI21_X1 U4344 ( .B1(n3575), .B2(n3574), .A(n3573), .ZN(n3583) );
  INV_X1 U4345 ( .A(n3576), .ZN(n4033) );
  OAI22_X1 U4346 ( .A1(n4062), .A2(n3629), .B1(STATE_REG_SCAN_IN), .B2(n4564), 
        .ZN(n3580) );
  OAI22_X1 U4347 ( .A1(n4024), .A2(n3578), .B1(n3628), .B2(n3577), .ZN(n3579)
         );
  AOI211_X1 U4348 ( .C1(n4033), .C2(n3618), .A(n3580), .B(n3579), .ZN(n3581)
         );
  OAI21_X1 U4349 ( .B1(n3583), .B2(n3582), .A(n3581), .ZN(U3230) );
  XNOR2_X1 U4350 ( .A(n3585), .B(n3584), .ZN(n3586) );
  XNOR2_X1 U4351 ( .A(n3587), .B(n3586), .ZN(n3588) );
  NAND2_X1 U4352 ( .A1(n3588), .A2(n3625), .ZN(n3592) );
  INV_X1 U4353 ( .A(n4141), .ZN(n4160) );
  OAI22_X1 U4354 ( .A1(n4160), .A2(n3629), .B1(n3628), .B2(n4145), .ZN(n3589)
         );
  AOI211_X1 U4355 ( .C1(n3631), .C2(n4113), .A(n3590), .B(n3589), .ZN(n3591)
         );
  OAI211_X1 U4356 ( .C1(n3634), .C2(n4149), .A(n3592), .B(n3591), .ZN(U3231)
         );
  OAI21_X1 U4357 ( .B1(n3594), .B2(n3593), .A(n3482), .ZN(n3599) );
  AOI22_X1 U4358 ( .A1(n4237), .A2(n3631), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3597) );
  AOI22_X1 U4359 ( .A1(n3984), .A2(n3617), .B1(n3983), .B2(n3595), .ZN(n3596)
         );
  OAI211_X1 U4360 ( .C1(n3634), .C2(n3996), .A(n3597), .B(n3596), .ZN(n3598)
         );
  AOI21_X1 U4361 ( .B1(n3599), .B2(n3625), .A(n3598), .ZN(n3600) );
  INV_X1 U4362 ( .A(n3600), .ZN(U3232) );
  NOR2_X1 U4363 ( .A1(n2066), .A2(n3602), .ZN(n3603) );
  XNOR2_X1 U4364 ( .A(n3601), .B(n3603), .ZN(n3604) );
  NAND2_X1 U4365 ( .A1(n3604), .A2(n3625), .ZN(n3608) );
  NOR2_X1 U4366 ( .A1(n3605), .A2(STATE_REG_SCAN_IN), .ZN(n4504) );
  OAI22_X1 U4367 ( .A1(n2498), .A2(n3629), .B1(n3628), .B2(n4058), .ZN(n3606)
         );
  AOI211_X1 U4368 ( .C1(n3631), .C2(n4022), .A(n4504), .B(n3606), .ZN(n3607)
         );
  OAI211_X1 U4369 ( .C1(n3634), .C2(n4065), .A(n3608), .B(n3607), .ZN(U3235)
         );
  INV_X1 U4370 ( .A(n3609), .ZN(n3611) );
  NAND2_X1 U4371 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  XNOR2_X1 U4372 ( .A(n3613), .B(n3612), .ZN(n3614) );
  NAND2_X1 U4373 ( .A1(n3614), .A2(n3625), .ZN(n3622) );
  OAI22_X1 U4374 ( .A1(n3628), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n3615), 
        .ZN(n3616) );
  AOI21_X1 U4375 ( .B1(n3809), .B2(n3617), .A(n3616), .ZN(n3621) );
  NAND2_X1 U4376 ( .A1(n3924), .A2(n3618), .ZN(n3620) );
  NAND2_X1 U4377 ( .A1(n3919), .A2(n3631), .ZN(n3619) );
  NAND4_X1 U4378 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(U3237)
         );
  NAND2_X1 U4379 ( .A1(n3540), .A2(n3541), .ZN(n3624) );
  XNOR2_X1 U4380 ( .A(n3624), .B(n3623), .ZN(n3626) );
  NAND2_X1 U4381 ( .A1(n3626), .A2(n3625), .ZN(n3633) );
  NOR2_X1 U4382 ( .A1(n3627), .A2(STATE_REG_SCAN_IN), .ZN(n4486) );
  OAI22_X1 U4383 ( .A1(n4295), .A2(n3629), .B1(n3628), .B2(n4118), .ZN(n3630)
         );
  AOI211_X1 U4384 ( .C1(n3631), .C2(n4292), .A(n4486), .B(n3630), .ZN(n3632)
         );
  OAI211_X1 U4385 ( .C1(n3634), .C2(n4114), .A(n3633), .B(n3632), .ZN(U3238)
         );
  INV_X1 U4386 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U4387 ( .A1(n3635), .A2(REG2_REG_31__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4388 ( .A1(n3636), .A2(REG0_REG_31__SCAN_IN), .ZN(n3637) );
  OAI211_X1 U4389 ( .C1(n3639), .C2(n4204), .A(n3638), .B(n3637), .ZN(n3895)
         );
  NAND2_X1 U4390 ( .A1(n2539), .A2(DATAI_31_), .ZN(n3892) );
  NAND2_X1 U4391 ( .A1(n3895), .A2(n3892), .ZN(n3708) );
  INV_X1 U4392 ( .A(n3708), .ZN(n3716) );
  INV_X1 U4393 ( .A(DATAI_30_), .ZN(n4709) );
  NOR2_X1 U4394 ( .A1(n2560), .A2(n4709), .ZN(n4209) );
  NOR2_X1 U4395 ( .A1(n3707), .A2(n4209), .ZN(n3792) );
  INV_X1 U4396 ( .A(n3792), .ZN(n3641) );
  OR2_X1 U4397 ( .A1(n3895), .A2(n3892), .ZN(n3640) );
  NAND2_X1 U4398 ( .A1(n3641), .A2(n3640), .ZN(n3740) );
  INV_X1 U4399 ( .A(n3740), .ZN(n3715) );
  INV_X1 U4400 ( .A(n3902), .ZN(n3643) );
  OAI21_X1 U4401 ( .B1(n3644), .B2(n3643), .A(n3642), .ZN(n3784) );
  INV_X1 U4402 ( .A(n3645), .ZN(n3677) );
  NAND2_X1 U4403 ( .A1(n3647), .A2(n3646), .ZN(n3672) );
  NAND2_X1 U4404 ( .A1(n3672), .A2(n3682), .ZN(n3765) );
  INV_X1 U4405 ( .A(n3765), .ZN(n3688) );
  INV_X1 U4406 ( .A(n3648), .ZN(n3649) );
  NAND4_X1 U4407 ( .A1(n3649), .A2(n3668), .A3(n3667), .A4(n3661), .ZN(n3674)
         );
  OAI211_X1 U4408 ( .C1(n3795), .C2(n2110), .A(n3652), .B(n3651), .ZN(n3653)
         );
  NAND3_X1 U4409 ( .A1(n3654), .A2(n2637), .A3(n3653), .ZN(n3655) );
  NAND3_X1 U4410 ( .A1(n3650), .A2(n3656), .A3(n3655), .ZN(n3657) );
  NAND3_X1 U4411 ( .A1(n3659), .A2(n3658), .A3(n3657), .ZN(n3660) );
  NAND4_X1 U4412 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3664)
         );
  NAND3_X1 U4413 ( .A1(n3731), .A2(n3665), .A3(n3664), .ZN(n3666) );
  NAND3_X1 U4414 ( .A1(n3668), .A2(n3667), .A3(n3666), .ZN(n3669) );
  AND3_X1 U4415 ( .A1(n3671), .A2(n3670), .A3(n3669), .ZN(n3673) );
  OAI22_X1 U4416 ( .A1(n3688), .A2(n3674), .B1(n3673), .B2(n3672), .ZN(n3675)
         );
  AOI22_X1 U4417 ( .A1(n3677), .A2(n3765), .B1(n3676), .B2(n3675), .ZN(n3690)
         );
  NAND3_X1 U4418 ( .A1(n3685), .A2(n3679), .A3(n3678), .ZN(n3689) );
  INV_X1 U4419 ( .A(n3680), .ZN(n3686) );
  INV_X1 U4420 ( .A(n3681), .ZN(n3684) );
  NAND2_X1 U4421 ( .A1(n3683), .A2(n3682), .ZN(n3766) );
  AOI211_X1 U4422 ( .C1(n3686), .C2(n3685), .A(n3684), .B(n3766), .ZN(n3687)
         );
  OAI22_X1 U4423 ( .A1(n3690), .A2(n3689), .B1(n3688), .B2(n3687), .ZN(n3692)
         );
  INV_X1 U4424 ( .A(n3770), .ZN(n3691) );
  AOI21_X1 U4425 ( .B1(n3767), .B2(n3692), .A(n3691), .ZN(n3695) );
  OR3_X1 U4426 ( .A1(n3694), .A2(n3726), .A3(n3693), .ZN(n3768) );
  OAI21_X1 U4427 ( .B1(n3695), .B2(n3768), .A(n3772), .ZN(n3696) );
  INV_X1 U4428 ( .A(n3696), .ZN(n3697) );
  OAI21_X1 U4429 ( .B1(n3965), .B2(n3697), .A(n3773), .ZN(n3698) );
  INV_X1 U4430 ( .A(n3698), .ZN(n3701) );
  INV_X1 U4431 ( .A(n3723), .ZN(n3699) );
  NOR2_X1 U4432 ( .A1(n3699), .A2(n3720), .ZN(n3777) );
  OAI211_X1 U4433 ( .C1(n3701), .C2(n3700), .A(n2660), .B(n3777), .ZN(n3702)
         );
  OAI211_X1 U4434 ( .C1(n3704), .C2(n4213), .A(n3703), .B(n3702), .ZN(n3713)
         );
  NAND2_X1 U4435 ( .A1(n3706), .A2(n3705), .ZN(n3781) );
  INV_X1 U4436 ( .A(n3781), .ZN(n3711) );
  NAND2_X1 U4437 ( .A1(n3707), .A2(n4209), .ZN(n3709) );
  AND2_X1 U4438 ( .A1(n3709), .A2(n3708), .ZN(n3738) );
  OAI21_X1 U4439 ( .B1(n3807), .B2(n3902), .A(n3738), .ZN(n3779) );
  INV_X1 U4440 ( .A(n3779), .ZN(n3710) );
  OAI21_X1 U4441 ( .B1(n3711), .B2(n3784), .A(n3710), .ZN(n3785) );
  INV_X1 U4442 ( .A(n3785), .ZN(n3712) );
  OAI21_X1 U4443 ( .B1(n3784), .B2(n3713), .A(n3712), .ZN(n3714) );
  OAI21_X1 U4444 ( .B1(n3716), .B2(n3715), .A(n3714), .ZN(n3799) );
  INV_X1 U4445 ( .A(n3787), .ZN(n3718) );
  NOR2_X1 U4446 ( .A1(n3718), .A2(n3717), .ZN(n3763) );
  XNOR2_X1 U4447 ( .A(n4231), .B(n3923), .ZN(n3915) );
  INV_X1 U4448 ( .A(n3929), .ZN(n3719) );
  OR2_X1 U4449 ( .A1(n3720), .A2(n3719), .ZN(n3948) );
  INV_X1 U4450 ( .A(n3948), .ZN(n3949) );
  INV_X1 U4451 ( .A(n3721), .ZN(n3966) );
  NOR2_X1 U4452 ( .A1(n3966), .A2(n3965), .ZN(n4004) );
  XNOR2_X1 U4453 ( .A(n4255), .B(n4030), .ZN(n4020) );
  AND2_X1 U4454 ( .A1(n3992), .A2(n4020), .ZN(n3758) );
  NAND2_X1 U4455 ( .A1(n3723), .A2(n3722), .ZN(n3969) );
  NAND2_X1 U4456 ( .A1(n3725), .A2(n3724), .ZN(n4045) );
  NAND2_X1 U4457 ( .A1(n2147), .A2(n4039), .ZN(n4077) );
  INV_X1 U4458 ( .A(n3727), .ZN(n3729) );
  OR2_X1 U4459 ( .A1(n3729), .A2(n3728), .ZN(n4144) );
  OR2_X1 U4460 ( .A1(n4077), .A2(n4144), .ZN(n3730) );
  NOR2_X1 U4461 ( .A1(n4045), .A2(n3730), .ZN(n3755) );
  NAND4_X1 U4462 ( .A1(n3732), .A2(n4100), .A3(n3731), .A4(n4538), .ZN(n3737)
         );
  NAND4_X1 U4463 ( .A1(n2648), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3736)
         );
  NOR2_X1 U4464 ( .A1(n3737), .A2(n3736), .ZN(n3754) );
  INV_X1 U4465 ( .A(n3738), .ZN(n3739) );
  NOR2_X1 U4466 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  AND2_X1 U4467 ( .A1(n4069), .A2(n3741), .ZN(n3753) );
  NAND4_X1 U4468 ( .A1(n2219), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3751)
         );
  INV_X1 U4469 ( .A(n4159), .ZN(n3749) );
  INV_X1 U4470 ( .A(n3745), .ZN(n3748) );
  NAND4_X1 U4471 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3750)
         );
  NOR2_X1 U4472 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  NAND4_X1 U4473 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3756)
         );
  NOR2_X1 U4474 ( .A1(n3969), .A2(n3756), .ZN(n3757) );
  NAND4_X1 U4475 ( .A1(n3949), .A2(n4004), .A3(n3758), .A4(n3757), .ZN(n3760)
         );
  NAND2_X1 U4476 ( .A1(n3912), .A2(n3759), .ZN(n3933) );
  NOR2_X1 U4477 ( .A1(n3760), .A2(n3933), .ZN(n3761) );
  NAND4_X1 U4478 ( .A1(n3763), .A2(n3762), .A3(n3915), .A4(n3761), .ZN(n3797)
         );
  OAI21_X1 U4479 ( .B1(n3764), .B2(n3766), .A(n3765), .ZN(n3771) );
  INV_X1 U4480 ( .A(n3767), .ZN(n3769) );
  AOI211_X1 U4481 ( .C1(n3771), .C2(n3770), .A(n3769), .B(n3768), .ZN(n3776)
         );
  NAND2_X1 U4482 ( .A1(n3773), .A2(n3772), .ZN(n3775) );
  OAI21_X1 U4483 ( .B1(n3776), .B2(n3775), .A(n3774), .ZN(n3778) );
  AOI21_X1 U4484 ( .B1(n3778), .B2(n3777), .A(n3913), .ZN(n3782) );
  NOR4_X1 U4485 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3790)
         );
  NOR2_X1 U4486 ( .A1(n3784), .A2(n3783), .ZN(n3786) );
  AOI21_X1 U4487 ( .B1(n3787), .B2(n3786), .A(n3785), .ZN(n3789) );
  INV_X1 U4488 ( .A(n4209), .ZN(n3788) );
  OAI22_X1 U4489 ( .A1(n3790), .A2(n3789), .B1(n3788), .B2(n3895), .ZN(n3794)
         );
  INV_X1 U4490 ( .A(n3895), .ZN(n3791) );
  INV_X1 U4491 ( .A(n3892), .ZN(n3896) );
  OAI21_X1 U4492 ( .B1(n3792), .B2(n3791), .A(n3896), .ZN(n3793) );
  NAND2_X1 U4493 ( .A1(n3794), .A2(n3793), .ZN(n3796) );
  MUX2_X1 U4494 ( .A(n3797), .B(n3796), .S(n3795), .Z(n3798) );
  MUX2_X1 U4495 ( .A(n3799), .B(n3798), .S(n4411), .Z(n3800) );
  XNOR2_X1 U4496 ( .A(n3800), .B(n3887), .ZN(n3806) );
  NAND2_X1 U4497 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  OAI211_X1 U4498 ( .C1(n4410), .C2(n3805), .A(n3803), .B(B_REG_SCAN_IN), .ZN(
        n3804) );
  OAI21_X1 U4499 ( .B1(n3806), .B2(n3805), .A(n3804), .ZN(U3239) );
  MUX2_X1 U4500 ( .A(DATAO_REG_31__SCAN_IN), .B(n3895), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4501 ( .A(DATAO_REG_29__SCAN_IN), .B(n3807), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4502 ( .A(DATAO_REG_28__SCAN_IN), .B(n4216), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4503 ( .A(DATAO_REG_27__SCAN_IN), .B(n3919), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4504 ( .A(DATAO_REG_26__SCAN_IN), .B(n3808), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4505 ( .A(DATAO_REG_25__SCAN_IN), .B(n3809), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4506 ( .A(DATAO_REG_24__SCAN_IN), .B(n4228), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4507 ( .A(DATAO_REG_23__SCAN_IN), .B(n4237), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4508 ( .A(DATAO_REG_22__SCAN_IN), .B(n3810), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4509 ( .A(DATAO_REG_21__SCAN_IN), .B(n3984), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4510 ( .A(n4255), .B(DATAO_REG_20__SCAN_IN), .S(n3819), .Z(U3570)
         );
  MUX2_X1 U4511 ( .A(n4022), .B(DATAO_REG_19__SCAN_IN), .S(n3819), .Z(U3569)
         );
  MUX2_X1 U4512 ( .A(DATAO_REG_18__SCAN_IN), .B(n3811), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4513 ( .A(n4282), .B(DATAO_REG_17__SCAN_IN), .S(n3819), .Z(U3567)
         );
  MUX2_X1 U4514 ( .A(DATAO_REG_16__SCAN_IN), .B(n4292), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4515 ( .A(DATAO_REG_15__SCAN_IN), .B(n2468), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4516 ( .A(DATAO_REG_14__SCAN_IN), .B(n4113), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4517 ( .A(DATAO_REG_13__SCAN_IN), .B(n4303), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4518 ( .A(n4141), .B(DATAO_REG_12__SCAN_IN), .S(n3819), .Z(U3562)
         );
  MUX2_X1 U4519 ( .A(DATAO_REG_11__SCAN_IN), .B(n3812), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4520 ( .A(DATAO_REG_10__SCAN_IN), .B(n4172), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4521 ( .A(n3813), .B(DATAO_REG_9__SCAN_IN), .S(n3819), .Z(U3559) );
  MUX2_X1 U4522 ( .A(n3814), .B(DATAO_REG_8__SCAN_IN), .S(n3819), .Z(U3558) );
  MUX2_X1 U4523 ( .A(DATAO_REG_7__SCAN_IN), .B(n3815), .S(U4043), .Z(U3557) );
  MUX2_X1 U4524 ( .A(DATAO_REG_6__SCAN_IN), .B(n3816), .S(U4043), .Z(U3556) );
  MUX2_X1 U4525 ( .A(DATAO_REG_5__SCAN_IN), .B(n3817), .S(U4043), .Z(U3555) );
  MUX2_X1 U4526 ( .A(DATAO_REG_4__SCAN_IN), .B(n3818), .S(U4043), .Z(U3554) );
  MUX2_X1 U4527 ( .A(n4183), .B(DATAO_REG_3__SCAN_IN), .S(n3819), .Z(U3553) );
  MUX2_X1 U4528 ( .A(DATAO_REG_2__SCAN_IN), .B(n2977), .S(U4043), .Z(U3552) );
  MUX2_X1 U4529 ( .A(DATAO_REG_1__SCAN_IN), .B(n2300), .S(U4043), .Z(U3551) );
  MUX2_X1 U4530 ( .A(n2834), .B(DATAO_REG_0__SCAN_IN), .S(n3819), .Z(U3550) );
  INV_X1 U4531 ( .A(n4512), .ZN(n3833) );
  OAI211_X1 U4532 ( .C1(n3822), .C2(n3821), .A(n4507), .B(n3820), .ZN(n3830)
         );
  INV_X1 U4533 ( .A(n3823), .ZN(n3827) );
  INV_X1 U4534 ( .A(n3824), .ZN(n3825) );
  OAI211_X1 U4535 ( .C1(n3827), .C2(n3826), .A(n4464), .B(n3825), .ZN(n3829)
         );
  AOI22_X1 U4536 ( .A1(n4505), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3828) );
  NAND4_X1 U4537 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(U3241)
         );
  NAND2_X1 U4538 ( .A1(n3833), .A2(n3832), .ZN(n3841) );
  OAI211_X1 U4539 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3835), .A(n4507), .B(n3834), 
        .ZN(n3840) );
  AOI22_X1 U4540 ( .A1(n4505), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3839) );
  XNOR2_X1 U4541 ( .A(n3836), .B(REG2_REG_3__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4542 ( .A1(n4464), .A2(n3837), .ZN(n3838) );
  NAND4_X1 U4543 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(U3243)
         );
  INV_X1 U4544 ( .A(n3876), .ZN(n3872) );
  NAND2_X1 U4545 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3862), .ZN(n3847) );
  AOI22_X1 U4546 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3862), .B1(n4530), .B2(
        n4298), .ZN(n4489) );
  INV_X1 U4547 ( .A(n3842), .ZN(n3844) );
  NAND2_X1 U4548 ( .A1(n3855), .A2(n3845), .ZN(n3846) );
  NAND2_X1 U4549 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U4550 ( .A1(n3846), .A2(n4478), .ZN(n4488) );
  NAND2_X1 U4551 ( .A1(n4489), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U4552 ( .A1(n3847), .A2(n4487), .ZN(n3848) );
  NOR2_X1 U4553 ( .A1(n3863), .A2(n3848), .ZN(n3849) );
  XNOR2_X1 U4554 ( .A(n3848), .B(n3863), .ZN(n4497) );
  NOR2_X1 U4555 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4497), .ZN(n4498) );
  NOR2_X1 U4556 ( .A1(n3849), .A2(n4498), .ZN(n3853) );
  INV_X1 U4557 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3851) );
  NOR2_X1 U4558 ( .A1(n3876), .A2(REG1_REG_17__SCAN_IN), .ZN(n3881) );
  INV_X1 U4559 ( .A(n3881), .ZN(n3850) );
  OAI21_X1 U4560 ( .B1(n3851), .B2(n3872), .A(n3850), .ZN(n3852) );
  AND2_X1 U4561 ( .A1(n3853), .A2(n3852), .ZN(n3854) );
  OAI21_X1 U4562 ( .B1(n3854), .B2(n3880), .A(n4507), .ZN(n3871) );
  XNOR2_X1 U4563 ( .A(n3872), .B(REG2_REG_17__SCAN_IN), .ZN(n3866) );
  INV_X1 U4564 ( .A(n3855), .ZN(n4531) );
  NOR2_X1 U4565 ( .A1(n4531), .A2(n3859), .ZN(n3860) );
  NOR2_X1 U4566 ( .A1(n3860), .A2(n4474), .ZN(n4484) );
  NAND2_X1 U4567 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3862), .ZN(n3861) );
  OAI21_X1 U4568 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3862), .A(n3861), .ZN(n4483) );
  NOR2_X1 U4569 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  INV_X1 U4570 ( .A(n3863), .ZN(n4529) );
  NAND2_X1 U4571 ( .A1(n3864), .A2(n4529), .ZN(n3865) );
  NAND2_X1 U4572 ( .A1(n3868), .A2(n3867), .ZN(n3869) );
  AOI21_X1 U4573 ( .B1(n4505), .B2(ADDR_REG_17__SCAN_IN), .A(n3869), .ZN(n3870) );
  OAI211_X1 U4574 ( .C1(n4512), .C2(n3872), .A(n3871), .B(n3870), .ZN(U3257)
         );
  INV_X1 U4575 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3873) );
  MUX2_X1 U4576 ( .A(REG2_REG_19__SCAN_IN), .B(n3873), .S(n4412), .Z(n3878) );
  INV_X1 U4577 ( .A(n3879), .ZN(n4528) );
  INV_X1 U4578 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4579 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4528), .B1(n3879), .B2(
        n3874), .ZN(n4503) );
  AOI21_X1 U4580 ( .B1(n3879), .B2(REG2_REG_18__SCAN_IN), .A(n4502), .ZN(n3877) );
  XOR2_X1 U4581 ( .A(n3878), .B(n3877), .Z(n3891) );
  INV_X1 U4582 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4583 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3879), .B1(n4528), .B2(
        n3882), .ZN(n4509) );
  MUX2_X1 U4584 ( .A(n4269), .B(REG1_REG_19__SCAN_IN), .S(n4412), .Z(n3883) );
  XNOR2_X1 U4585 ( .A(n3884), .B(n3883), .ZN(n3889) );
  NAND2_X1 U4586 ( .A1(n4505), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3885) );
  OAI211_X1 U4587 ( .C1(n4512), .C2(n3887), .A(n3886), .B(n3885), .ZN(n3888)
         );
  AOI21_X1 U4588 ( .B1(n3889), .B2(n4507), .A(n3888), .ZN(n3890) );
  OAI21_X1 U4589 ( .B1(n3891), .B2(n4501), .A(n3890), .ZN(U3259) );
  NOR2_X2 U4590 ( .A1(n4208), .A2(n4209), .ZN(n4207) );
  XNOR2_X1 U4591 ( .A(n4207), .B(n3892), .ZN(n4340) );
  INV_X1 U4592 ( .A(n3893), .ZN(n3894) );
  NAND2_X1 U4593 ( .A1(n3895), .A2(n3894), .ZN(n4211) );
  NAND2_X1 U4594 ( .A1(n4290), .A2(n3896), .ZN(n3897) );
  NAND2_X1 U4595 ( .A1(n4211), .A2(n3897), .ZN(n4337) );
  NAND2_X1 U4596 ( .A1(n4516), .A2(n4337), .ZN(n3899) );
  NAND2_X1 U4597 ( .A1(n4525), .A2(REG2_REG_31__SCAN_IN), .ZN(n3898) );
  OAI211_X1 U4598 ( .C1(n4340), .C2(n4196), .A(n3899), .B(n3898), .ZN(U3260)
         );
  INV_X1 U4599 ( .A(n3900), .ZN(n3910) );
  INV_X1 U4600 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3901) );
  OAI22_X1 U4601 ( .A1(n4197), .A2(n3902), .B1(n3901), .B2(n4516), .ZN(n3903)
         );
  AOI21_X1 U4602 ( .B1(n4216), .B2(n4190), .A(n3903), .ZN(n3909) );
  OAI22_X1 U4603 ( .A1(n3905), .A2(n4196), .B1(n3904), .B2(n4513), .ZN(n3906)
         );
  OAI21_X1 U4604 ( .B1(n3907), .B2(n3906), .A(n4516), .ZN(n3908) );
  OAI211_X1 U4605 ( .C1(n3910), .C2(n4105), .A(n3909), .B(n3908), .ZN(U3354)
         );
  XNOR2_X1 U4606 ( .A(n3911), .B(n3915), .ZN(n4224) );
  INV_X1 U4607 ( .A(n4224), .ZN(n3928) );
  OAI21_X1 U4608 ( .B1(n3914), .B2(n3913), .A(n3912), .ZN(n3917) );
  INV_X1 U4609 ( .A(n3915), .ZN(n3916) );
  XNOR2_X1 U4610 ( .A(n3917), .B(n3916), .ZN(n3921) );
  OAI22_X1 U4611 ( .A1(n4240), .A2(n4329), .B1(n3923), .B2(n4323), .ZN(n3918)
         );
  AOI21_X1 U4612 ( .B1(n3919), .B2(n4291), .A(n3918), .ZN(n3920) );
  OAI21_X1 U4613 ( .B1(n3921), .B2(n4306), .A(n3920), .ZN(n4223) );
  OAI21_X1 U4614 ( .B1(n3936), .B2(n3923), .A(n3922), .ZN(n4352) );
  AOI22_X1 U4615 ( .A1(n3924), .A2(n4180), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4525), .ZN(n3925) );
  OAI21_X1 U4616 ( .B1(n4352), .B2(n4196), .A(n3925), .ZN(n3926) );
  AOI21_X1 U4617 ( .B1(n4223), .B2(n4516), .A(n3926), .ZN(n3927) );
  OAI21_X1 U4618 ( .B1(n3928), .B2(n4105), .A(n3927), .ZN(U3264) );
  NAND2_X1 U4619 ( .A1(n3930), .A2(n3929), .ZN(n3931) );
  XNOR2_X1 U4620 ( .A(n3931), .B(n3933), .ZN(n3932) );
  NAND2_X1 U4621 ( .A1(n3932), .A2(n4098), .ZN(n4230) );
  XNOR2_X1 U4622 ( .A(n3934), .B(n3933), .ZN(n4233) );
  NAND2_X1 U4623 ( .A1(n4233), .A2(n4153), .ZN(n3946) );
  NOR2_X1 U4624 ( .A1(n3952), .A2(n3937), .ZN(n3935) );
  OR2_X1 U4625 ( .A1(n3936), .A2(n3935), .ZN(n4356) );
  INV_X1 U4626 ( .A(n4356), .ZN(n3944) );
  NOR2_X1 U4627 ( .A1(n4197), .A2(n3937), .ZN(n3941) );
  INV_X1 U4628 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3938) );
  OAI22_X1 U4629 ( .A1(n3939), .A2(n4513), .B1(n3938), .B2(n4516), .ZN(n3940)
         );
  AOI211_X1 U4630 ( .C1(n4190), .C2(n4228), .A(n3941), .B(n3940), .ZN(n3942)
         );
  OAI21_X1 U4631 ( .B1(n4231), .B2(n4083), .A(n3942), .ZN(n3943) );
  AOI21_X1 U4632 ( .B1(n3944), .B2(n4519), .A(n3943), .ZN(n3945) );
  OAI211_X1 U4633 ( .C1(n4525), .C2(n4230), .A(n3946), .B(n3945), .ZN(U3265)
         );
  XOR2_X1 U4634 ( .A(n3948), .B(n3947), .Z(n4242) );
  XNOR2_X1 U4635 ( .A(n3950), .B(n3949), .ZN(n3951) );
  NAND2_X1 U4636 ( .A1(n3951), .A2(n4098), .ZN(n4239) );
  NOR2_X1 U4637 ( .A1(n4239), .A2(n4525), .ZN(n3962) );
  INV_X1 U4638 ( .A(n3974), .ZN(n3955) );
  INV_X1 U4639 ( .A(n3952), .ZN(n3953) );
  OAI21_X1 U4640 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n4360) );
  INV_X1 U4641 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3956) );
  OAI22_X1 U4642 ( .A1(n3957), .A2(n4513), .B1(n3956), .B2(n4516), .ZN(n3959)
         );
  OAI22_X1 U4643 ( .A1(n4240), .A2(n4083), .B1(n3987), .B2(n4131), .ZN(n3958)
         );
  AOI211_X1 U4644 ( .C1(n4236), .C2(n4182), .A(n3959), .B(n3958), .ZN(n3960)
         );
  OAI21_X1 U4645 ( .B1(n4360), .B2(n4196), .A(n3960), .ZN(n3961) );
  AOI211_X1 U4646 ( .C1(n4242), .C2(n4153), .A(n3962), .B(n3961), .ZN(n3963)
         );
  INV_X1 U4647 ( .A(n3963), .ZN(U3266) );
  XOR2_X1 U4648 ( .A(n3969), .B(n3964), .Z(n4246) );
  INV_X1 U4649 ( .A(n4246), .ZN(n3981) );
  INV_X1 U4650 ( .A(n3965), .ZN(n3967) );
  AOI21_X1 U4651 ( .B1(n4001), .B2(n3967), .A(n3966), .ZN(n3982) );
  OAI21_X1 U4652 ( .B1(n3982), .B2(n2550), .A(n3968), .ZN(n3970) );
  XNOR2_X1 U4653 ( .A(n3970), .B(n3969), .ZN(n3973) );
  OAI22_X1 U4654 ( .A1(n4258), .A2(n4329), .B1(n4323), .B2(n3975), .ZN(n3971)
         );
  AOI21_X1 U4655 ( .B1(n4228), .B2(n4291), .A(n3971), .ZN(n3972) );
  OAI21_X1 U4656 ( .B1(n3973), .B2(n4306), .A(n3972), .ZN(n4245) );
  INV_X1 U4657 ( .A(n3993), .ZN(n3976) );
  OAI21_X1 U4658 ( .B1(n3976), .B2(n3975), .A(n3974), .ZN(n4364) );
  AOI22_X1 U4659 ( .A1(n3977), .A2(n4180), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4525), .ZN(n3978) );
  OAI21_X1 U4660 ( .B1(n4364), .B2(n4196), .A(n3978), .ZN(n3979) );
  AOI21_X1 U4661 ( .B1(n4245), .B2(n4516), .A(n3979), .ZN(n3980) );
  OAI21_X1 U4662 ( .B1(n3981), .B2(n4105), .A(n3980), .ZN(U3267) );
  XNOR2_X1 U4663 ( .A(n3982), .B(n2550), .ZN(n3989) );
  NAND2_X1 U4664 ( .A1(n4290), .A2(n3983), .ZN(n3986) );
  NAND2_X1 U4665 ( .A1(n3984), .A2(n4304), .ZN(n3985) );
  OAI211_X1 U4666 ( .C1(n3987), .C2(n4316), .A(n3986), .B(n3985), .ZN(n3988)
         );
  AOI21_X1 U4667 ( .B1(n3989), .B2(n4098), .A(n3988), .ZN(n4250) );
  NAND2_X1 U4668 ( .A1(n3991), .A2(n3992), .ZN(n4249) );
  NAND3_X1 U4669 ( .A1(n3990), .A2(n4249), .A3(n4153), .ZN(n4000) );
  OAI21_X1 U4670 ( .B1(n4005), .B2(n3994), .A(n3993), .ZN(n4368) );
  INV_X1 U4671 ( .A(n4368), .ZN(n3998) );
  INV_X1 U4672 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3995) );
  OAI22_X1 U4673 ( .A1(n3996), .A2(n4513), .B1(n3995), .B2(n4516), .ZN(n3997)
         );
  AOI21_X1 U4674 ( .B1(n3998), .B2(n4519), .A(n3997), .ZN(n3999) );
  OAI211_X1 U4675 ( .C1(n4525), .C2(n4250), .A(n4000), .B(n3999), .ZN(U3268)
         );
  XNOR2_X1 U4676 ( .A(n4001), .B(n4004), .ZN(n4002) );
  NAND2_X1 U4677 ( .A1(n4002), .A2(n4098), .ZN(n4257) );
  XNOR2_X1 U4678 ( .A(n4003), .B(n4004), .ZN(n4260) );
  NAND2_X1 U4679 ( .A1(n4260), .A2(n4153), .ZN(n4015) );
  INV_X1 U4680 ( .A(n4005), .ZN(n4006) );
  OAI21_X1 U4681 ( .B1(n4031), .B2(n4009), .A(n4006), .ZN(n4372) );
  INV_X1 U4682 ( .A(n4372), .ZN(n4013) );
  AOI22_X1 U4683 ( .A1(n4007), .A2(n4180), .B1(n4525), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4008) );
  OAI21_X1 U4684 ( .B1(n4009), .B2(n4197), .A(n4008), .ZN(n4012) );
  OAI22_X1 U4685 ( .A1(n4258), .A2(n4083), .B1(n4010), .B2(n4131), .ZN(n4011)
         );
  AOI211_X1 U4686 ( .C1(n4013), .C2(n4519), .A(n4012), .B(n4011), .ZN(n4014)
         );
  OAI211_X1 U4687 ( .C1(n4525), .C2(n4257), .A(n4015), .B(n4014), .ZN(U3269)
         );
  XNOR2_X1 U4688 ( .A(n4016), .B(n4020), .ZN(n4029) );
  INV_X1 U4689 ( .A(n4017), .ZN(n4018) );
  NAND2_X1 U4690 ( .A1(n4019), .A2(n4018), .ZN(n4021) );
  XNOR2_X1 U4691 ( .A(n4021), .B(n4020), .ZN(n4026) );
  AOI22_X1 U4692 ( .A1(n4022), .A2(n4304), .B1(n4030), .B2(n4290), .ZN(n4023)
         );
  OAI21_X1 U4693 ( .B1(n4024), .B2(n4316), .A(n4023), .ZN(n4025) );
  AOI21_X1 U4694 ( .B1(n4026), .B2(n4098), .A(n4025), .ZN(n4027) );
  OAI21_X1 U4695 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4263) );
  INV_X1 U4696 ( .A(n4263), .ZN(n4037) );
  INV_X1 U4697 ( .A(n4029), .ZN(n4264) );
  AND2_X1 U4698 ( .A1(n4049), .A2(n4030), .ZN(n4032) );
  OR2_X1 U4699 ( .A1(n4032), .A2(n4031), .ZN(n4376) );
  AOI22_X1 U4700 ( .A1(n4033), .A2(n4180), .B1(n4525), .B2(
        REG2_REG_20__SCAN_IN), .ZN(n4034) );
  OAI21_X1 U4701 ( .B1(n4376), .B2(n4196), .A(n4034), .ZN(n4035) );
  AOI21_X1 U4702 ( .B1(n4264), .B2(n4520), .A(n4035), .ZN(n4036) );
  OAI21_X1 U4703 ( .B1(n4037), .B2(n4525), .A(n4036), .ZN(U3270) );
  XNOR2_X1 U4704 ( .A(n4038), .B(n4045), .ZN(n4268) );
  INV_X1 U4705 ( .A(n4268), .ZN(n4056) );
  NAND2_X1 U4706 ( .A1(n4040), .A2(n4039), .ZN(n4059) );
  INV_X1 U4707 ( .A(n4041), .ZN(n4043) );
  OAI21_X1 U4708 ( .B1(n4059), .B2(n4043), .A(n4042), .ZN(n4044) );
  XOR2_X1 U4709 ( .A(n4045), .B(n4044), .Z(n4048) );
  OAI22_X1 U4710 ( .A1(n4277), .A2(n4329), .B1(n4323), .B2(n4050), .ZN(n4046)
         );
  AOI21_X1 U4711 ( .B1(n4291), .B2(n4255), .A(n4046), .ZN(n4047) );
  OAI21_X1 U4712 ( .B1(n4048), .B2(n4306), .A(n4047), .ZN(n4267) );
  INV_X1 U4713 ( .A(n4057), .ZN(n4051) );
  OAI21_X1 U4714 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4380) );
  AOI22_X1 U4715 ( .A1(n4525), .A2(REG2_REG_19__SCAN_IN), .B1(n4052), .B2(
        n4180), .ZN(n4053) );
  OAI21_X1 U4716 ( .B1(n4380), .B2(n4196), .A(n4053), .ZN(n4054) );
  AOI21_X1 U4717 ( .B1(n4267), .B2(n4516), .A(n4054), .ZN(n4055) );
  OAI21_X1 U4718 ( .B1(n4056), .B2(n4105), .A(n4055), .ZN(U3271) );
  OAI211_X1 U4719 ( .C1(n4079), .C2(n4058), .A(n4057), .B(n4285), .ZN(n4271)
         );
  XNOR2_X1 U4720 ( .A(n4059), .B(n4069), .ZN(n4064) );
  AOI22_X1 U4721 ( .A1(n4282), .A2(n4304), .B1(n4060), .B2(n4290), .ZN(n4061)
         );
  OAI21_X1 U4722 ( .B1(n4062), .B2(n4316), .A(n4061), .ZN(n4063) );
  AOI21_X1 U4723 ( .B1(n4064), .B2(n4098), .A(n4063), .ZN(n4272) );
  OAI21_X1 U4724 ( .B1(n4412), .B2(n4271), .A(n4272), .ZN(n4072) );
  OAI22_X1 U4725 ( .A1(n4516), .A2(n3874), .B1(n4065), .B2(n4513), .ZN(n4071)
         );
  INV_X1 U4726 ( .A(n4067), .ZN(n4068) );
  AOI21_X1 U4727 ( .B1(n4069), .B2(n4066), .A(n4068), .ZN(n4273) );
  NOR2_X1 U4728 ( .A1(n4273), .A2(n4105), .ZN(n4070) );
  AOI211_X1 U4729 ( .C1(n4516), .C2(n4072), .A(n4071), .B(n4070), .ZN(n4073)
         );
  INV_X1 U4730 ( .A(n4073), .ZN(U3272) );
  XNOR2_X1 U4731 ( .A(n4074), .B(n4077), .ZN(n4075) );
  NAND2_X1 U4732 ( .A1(n4075), .A2(n4098), .ZN(n4276) );
  XOR2_X1 U4733 ( .A(n4077), .B(n4076), .Z(n4279) );
  NAND2_X1 U4734 ( .A1(n4279), .A2(n4153), .ZN(n4089) );
  INV_X1 U4735 ( .A(n4078), .ZN(n4093) );
  INV_X1 U4736 ( .A(n4079), .ZN(n4080) );
  OAI21_X1 U4737 ( .B1(n4093), .B2(n2497), .A(n4080), .ZN(n4385) );
  INV_X1 U4738 ( .A(n4385), .ZN(n4087) );
  AOI22_X1 U4739 ( .A1(n4525), .A2(REG2_REG_17__SCAN_IN), .B1(n4081), .B2(
        n4180), .ZN(n4082) );
  OAI21_X1 U4740 ( .B1(n2497), .B2(n4197), .A(n4082), .ZN(n4086) );
  OAI22_X1 U4741 ( .A1(n4131), .A2(n4084), .B1(n4277), .B2(n4083), .ZN(n4085)
         );
  AOI211_X1 U4742 ( .C1(n4087), .C2(n4519), .A(n4086), .B(n4085), .ZN(n4088)
         );
  OAI211_X1 U4743 ( .C1(n4525), .C2(n4276), .A(n4089), .B(n4088), .ZN(U3273)
         );
  INV_X1 U4744 ( .A(n4100), .ZN(n4091) );
  OAI21_X1 U4745 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4289) );
  AOI21_X1 U4746 ( .B1(n4281), .B2(n4111), .A(n4093), .ZN(n4286) );
  AOI22_X1 U4747 ( .A1(n4191), .A2(n4282), .B1(n4190), .B2(n2468), .ZN(n4096)
         );
  AOI22_X1 U4748 ( .A1(n4525), .A2(REG2_REG_16__SCAN_IN), .B1(n4094), .B2(
        n4180), .ZN(n4095) );
  OAI211_X1 U4749 ( .C1(n4097), .C2(n4197), .A(n4096), .B(n4095), .ZN(n4103)
         );
  OAI211_X1 U4750 ( .C1(n4101), .C2(n4100), .A(n4099), .B(n4098), .ZN(n4287)
         );
  NOR2_X1 U4751 ( .A1(n4287), .A2(n4525), .ZN(n4102) );
  AOI211_X1 U4752 ( .C1(n4286), .C2(n4519), .A(n4103), .B(n4102), .ZN(n4104)
         );
  OAI21_X1 U4753 ( .B1(n4289), .B2(n4105), .A(n4104), .ZN(U3274) );
  AOI21_X1 U4754 ( .B1(n4106), .B2(n4109), .A(n4306), .ZN(n4108) );
  NAND2_X1 U4755 ( .A1(n4108), .A2(n4107), .ZN(n4294) );
  XNOR2_X1 U4756 ( .A(n4110), .B(n4109), .ZN(n4297) );
  NAND2_X1 U4757 ( .A1(n4297), .A2(n4153), .ZN(n4122) );
  INV_X1 U4758 ( .A(n4126), .ZN(n4112) );
  OAI21_X1 U4759 ( .B1(n4112), .B2(n4118), .A(n4111), .ZN(n4390) );
  INV_X1 U4760 ( .A(n4390), .ZN(n4120) );
  AOI22_X1 U4761 ( .A1(n4191), .A2(n4292), .B1(n4190), .B2(n4113), .ZN(n4117)
         );
  INV_X1 U4762 ( .A(n4114), .ZN(n4115) );
  AOI22_X1 U4763 ( .A1(n4525), .A2(REG2_REG_15__SCAN_IN), .B1(n4115), .B2(
        n4180), .ZN(n4116) );
  OAI211_X1 U4764 ( .C1(n4118), .C2(n4197), .A(n4117), .B(n4116), .ZN(n4119)
         );
  AOI21_X1 U4765 ( .B1(n4120), .B2(n4519), .A(n4119), .ZN(n4121) );
  OAI211_X1 U4766 ( .C1(n4525), .C2(n4294), .A(n4122), .B(n4121), .ZN(U3275)
         );
  XNOR2_X1 U4767 ( .A(n3764), .B(n4124), .ZN(n4307) );
  OAI21_X1 U4768 ( .B1(n4125), .B2(n4124), .A(n4123), .ZN(n4309) );
  NAND2_X1 U4769 ( .A1(n4309), .A2(n4153), .ZN(n4135) );
  OAI21_X1 U4770 ( .B1(n4148), .B2(n4300), .A(n4126), .ZN(n4394) );
  INV_X1 U4771 ( .A(n4394), .ZN(n4133) );
  AOI22_X1 U4772 ( .A1(n4182), .A2(n4127), .B1(n4191), .B2(n2468), .ZN(n4130)
         );
  AOI22_X1 U4773 ( .A1(n4525), .A2(REG2_REG_14__SCAN_IN), .B1(n4128), .B2(
        n4180), .ZN(n4129) );
  OAI211_X1 U4774 ( .C1(n4317), .C2(n4131), .A(n4130), .B(n4129), .ZN(n4132)
         );
  AOI21_X1 U4775 ( .B1(n4133), .B2(n4519), .A(n4132), .ZN(n4134) );
  OAI211_X1 U4776 ( .C1(n4307), .C2(n4136), .A(n4135), .B(n4134), .ZN(U3276)
         );
  OAI21_X1 U4777 ( .B1(n3339), .B2(n4138), .A(n4137), .ZN(n4139) );
  XOR2_X1 U4778 ( .A(n4144), .B(n4139), .Z(n4143) );
  OAI22_X1 U4779 ( .A1(n4295), .A2(n4316), .B1(n4323), .B2(n4145), .ZN(n4140)
         );
  AOI21_X1 U4780 ( .B1(n4304), .B2(n4141), .A(n4140), .ZN(n4142) );
  OAI21_X1 U4781 ( .B1(n4143), .B2(n4306), .A(n4142), .ZN(n4312) );
  INV_X1 U4782 ( .A(n4312), .ZN(n4155) );
  XOR2_X1 U4783 ( .A(n4144), .B(n2064), .Z(n4313) );
  NOR2_X1 U4784 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  OR2_X1 U4785 ( .A1(n4148), .A2(n4147), .ZN(n4398) );
  NOR2_X1 U4786 ( .A1(n4398), .A2(n4196), .ZN(n4152) );
  OAI22_X1 U4787 ( .A1(n4516), .A2(n4150), .B1(n4149), .B2(n4513), .ZN(n4151)
         );
  AOI211_X1 U4788 ( .C1(n4313), .C2(n4153), .A(n4152), .B(n4151), .ZN(n4154)
         );
  OAI21_X1 U4789 ( .B1(n4525), .B2(n4155), .A(n4154), .ZN(U3277) );
  OAI21_X1 U4790 ( .B1(n4157), .B2(n4159), .A(n4156), .ZN(n4333) );
  INV_X1 U4791 ( .A(n4333), .ZN(n4176) );
  XNOR2_X1 U4792 ( .A(n4158), .B(n4159), .ZN(n4164) );
  OAI22_X1 U4793 ( .A1(n4160), .A2(n4316), .B1(n4323), .B2(n4168), .ZN(n4161)
         );
  AOI21_X1 U4794 ( .B1(n4333), .B2(n4162), .A(n4161), .ZN(n4163) );
  OAI21_X1 U4795 ( .B1(n4306), .B2(n4164), .A(n4163), .ZN(n4331) );
  NAND2_X1 U4796 ( .A1(n4331), .A2(n4516), .ZN(n4174) );
  OAI22_X1 U4797 ( .A1(n4516), .A2(n4166), .B1(n4165), .B2(n4513), .ZN(n4171)
         );
  OAI21_X1 U4798 ( .B1(n4169), .B2(n4168), .A(n4167), .ZN(n4407) );
  NOR2_X1 U4799 ( .A1(n4407), .A2(n4196), .ZN(n4170) );
  AOI211_X1 U4800 ( .C1(n4190), .C2(n4172), .A(n4171), .B(n4170), .ZN(n4173)
         );
  OAI211_X1 U4801 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4173), .ZN(U3279)
         );
  MUX2_X1 U4802 ( .A(n4178), .B(n4177), .S(n4525), .Z(n4188) );
  AOI22_X1 U4803 ( .A1(n4179), .A2(n4520), .B1(n4190), .B2(n2300), .ZN(n4187)
         );
  AOI22_X1 U4804 ( .A1(n4182), .A2(n4181), .B1(REG3_REG_2__SCAN_IN), .B2(n4180), .ZN(n4186) );
  AOI22_X1 U4805 ( .A1(n4519), .A2(n4184), .B1(n4191), .B2(n4183), .ZN(n4185)
         );
  NAND4_X1 U4806 ( .A1(n4188), .A2(n4187), .A3(n4186), .A4(n4185), .ZN(U3288)
         );
  MUX2_X1 U4807 ( .A(n4189), .B(n2763), .S(n4525), .Z(n4203) );
  AOI22_X1 U4808 ( .A1(n4191), .A2(n2977), .B1(n4190), .B2(n2834), .ZN(n4202)
         );
  NAND2_X1 U4809 ( .A1(n4192), .A2(n4520), .ZN(n4193) );
  OAI21_X1 U4810 ( .B1(n4513), .B2(n4194), .A(n4193), .ZN(n4200) );
  OAI22_X1 U4811 ( .A1(n4198), .A2(n4197), .B1(n4196), .B2(n4195), .ZN(n4199)
         );
  NOR2_X1 U4812 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  NAND3_X1 U4813 ( .A1(n4203), .A2(n4202), .A3(n4201), .ZN(U3289) );
  NOR2_X1 U4814 ( .A1(n4559), .A2(n4204), .ZN(n4205) );
  AOI21_X1 U4815 ( .B1(n4559), .B2(n4337), .A(n4205), .ZN(n4206) );
  OAI21_X1 U4816 ( .B1(n4340), .B2(n4336), .A(n4206), .ZN(U3549) );
  AOI21_X1 U4817 ( .B1(n4209), .B2(n4208), .A(n4207), .ZN(n4420) );
  INV_X1 U4818 ( .A(n4420), .ZN(n4343) );
  NAND2_X1 U4819 ( .A1(n4290), .A2(n4209), .ZN(n4210) );
  AND2_X1 U4820 ( .A1(n4211), .A2(n4210), .ZN(n4422) );
  MUX2_X1 U4821 ( .A(n2721), .B(n4422), .S(n4559), .Z(n4212) );
  OAI21_X1 U4822 ( .B1(n4343), .B2(n4336), .A(n4212), .ZN(U3548) );
  INV_X1 U4823 ( .A(n4213), .ZN(n4214) );
  OAI22_X1 U4824 ( .A1(n4231), .A2(n4329), .B1(n4214), .B2(n4323), .ZN(n4215)
         );
  AOI21_X1 U4825 ( .B1(n4216), .B2(n4291), .A(n4215), .ZN(n4218) );
  OAI211_X1 U4826 ( .C1(n4219), .C2(n4546), .A(n4218), .B(n4217), .ZN(n4344)
         );
  MUX2_X1 U4827 ( .A(REG1_REG_27__SCAN_IN), .B(n4344), .S(n4559), .Z(n4220) );
  INV_X1 U4828 ( .A(n4222), .ZN(U3545) );
  AOI21_X1 U4829 ( .B1(n4224), .B2(n4325), .A(n4223), .ZN(n4349) );
  MUX2_X1 U4830 ( .A(n4225), .B(n4349), .S(n4559), .Z(n4226) );
  OAI21_X1 U4831 ( .B1(n4336), .B2(n4352), .A(n4226), .ZN(U3544) );
  AOI22_X1 U4832 ( .A1(n4228), .A2(n4304), .B1(n4227), .B2(n4290), .ZN(n4229)
         );
  OAI211_X1 U4833 ( .C1(n4231), .C2(n4316), .A(n4230), .B(n4229), .ZN(n4232)
         );
  AOI21_X1 U4834 ( .B1(n4233), .B2(n4325), .A(n4232), .ZN(n4353) );
  MUX2_X1 U4835 ( .A(n4234), .B(n4353), .S(n4559), .Z(n4235) );
  OAI21_X1 U4836 ( .B1(n4336), .B2(n4356), .A(n4235), .ZN(U3543) );
  AOI22_X1 U4837 ( .A1(n4237), .A2(n4304), .B1(n4290), .B2(n4236), .ZN(n4238)
         );
  OAI211_X1 U4838 ( .C1(n4240), .C2(n4316), .A(n4239), .B(n4238), .ZN(n4241)
         );
  AOI21_X1 U4839 ( .B1(n4242), .B2(n4325), .A(n4241), .ZN(n4357) );
  MUX2_X1 U4840 ( .A(n4243), .B(n4357), .S(n4559), .Z(n4244) );
  OAI21_X1 U4841 ( .B1(n4336), .B2(n4360), .A(n4244), .ZN(U3542) );
  AOI21_X1 U4842 ( .B1(n4246), .B2(n4325), .A(n4245), .ZN(n4361) );
  MUX2_X1 U4843 ( .A(n4247), .B(n4361), .S(n4559), .Z(n4248) );
  OAI21_X1 U4844 ( .B1(n4336), .B2(n4364), .A(n4248), .ZN(U3541) );
  NAND3_X1 U4845 ( .A1(n3990), .A2(n4249), .A3(n4325), .ZN(n4251) );
  AND2_X1 U4846 ( .A1(n4251), .A2(n4250), .ZN(n4365) );
  MUX2_X1 U4847 ( .A(n4252), .B(n4365), .S(n4559), .Z(n4253) );
  OAI21_X1 U4848 ( .B1(n4336), .B2(n4368), .A(n4253), .ZN(U3540) );
  AOI22_X1 U4849 ( .A1(n4255), .A2(n4304), .B1(n4254), .B2(n4290), .ZN(n4256)
         );
  OAI211_X1 U4850 ( .C1(n4258), .C2(n4316), .A(n4257), .B(n4256), .ZN(n4259)
         );
  AOI21_X1 U4851 ( .B1(n4260), .B2(n4325), .A(n4259), .ZN(n4369) );
  MUX2_X1 U4852 ( .A(n4261), .B(n4369), .S(n4559), .Z(n4262) );
  OAI21_X1 U4853 ( .B1(n4336), .B2(n4372), .A(n4262), .ZN(U3539) );
  AOI21_X1 U4854 ( .B1(n4543), .B2(n4264), .A(n4263), .ZN(n4373) );
  MUX2_X1 U4855 ( .A(n4265), .B(n4373), .S(n4559), .Z(n4266) );
  OAI21_X1 U4856 ( .B1(n4336), .B2(n4376), .A(n4266), .ZN(U3538) );
  AOI21_X1 U4857 ( .B1(n4268), .B2(n4325), .A(n4267), .ZN(n4377) );
  MUX2_X1 U4858 ( .A(n4269), .B(n4377), .S(n4559), .Z(n4270) );
  OAI21_X1 U4859 ( .B1(n4336), .B2(n4380), .A(n4270), .ZN(U3537) );
  OAI211_X1 U4860 ( .C1(n4273), .C2(n4546), .A(n4272), .B(n4271), .ZN(n4381)
         );
  MUX2_X1 U4861 ( .A(REG1_REG_18__SCAN_IN), .B(n4381), .S(n4559), .Z(U3536) );
  AOI22_X1 U4862 ( .A1(n4292), .A2(n4304), .B1(n4274), .B2(n4290), .ZN(n4275)
         );
  OAI211_X1 U4863 ( .C1(n4277), .C2(n4316), .A(n4276), .B(n4275), .ZN(n4278)
         );
  AOI21_X1 U4864 ( .B1(n4279), .B2(n4325), .A(n4278), .ZN(n4382) );
  MUX2_X1 U4865 ( .A(n3851), .B(n4382), .S(n4559), .Z(n4280) );
  OAI21_X1 U4866 ( .B1(n4336), .B2(n4385), .A(n4280), .ZN(U3535) );
  AOI22_X1 U4867 ( .A1(n4282), .A2(n4291), .B1(n4290), .B2(n4281), .ZN(n4283)
         );
  OAI21_X1 U4868 ( .B1(n4301), .B2(n4329), .A(n4283), .ZN(n4284) );
  AOI21_X1 U4869 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4288) );
  OAI211_X1 U4870 ( .C1(n4289), .C2(n4546), .A(n4288), .B(n4287), .ZN(n4386)
         );
  MUX2_X1 U4871 ( .A(REG1_REG_16__SCAN_IN), .B(n4386), .S(n4559), .Z(U3534) );
  AOI22_X1 U4872 ( .A1(n4292), .A2(n4291), .B1(n2467), .B2(n4290), .ZN(n4293)
         );
  OAI211_X1 U4873 ( .C1(n4295), .C2(n4329), .A(n4294), .B(n4293), .ZN(n4296)
         );
  AOI21_X1 U4874 ( .B1(n4297), .B2(n4325), .A(n4296), .ZN(n4387) );
  MUX2_X1 U4875 ( .A(n4298), .B(n4387), .S(n4559), .Z(n4299) );
  OAI21_X1 U4876 ( .B1(n4336), .B2(n4390), .A(n4299), .ZN(U3533) );
  OAI22_X1 U4877 ( .A1(n4301), .A2(n4316), .B1(n4323), .B2(n4300), .ZN(n4302)
         );
  AOI21_X1 U4878 ( .B1(n4304), .B2(n4303), .A(n4302), .ZN(n4305) );
  OAI21_X1 U4879 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(n4308) );
  AOI21_X1 U4880 ( .B1(n4309), .B2(n4325), .A(n4308), .ZN(n4391) );
  MUX2_X1 U4881 ( .A(n4310), .B(n4391), .S(n4559), .Z(n4311) );
  OAI21_X1 U4882 ( .B1(n4336), .B2(n4394), .A(n4311), .ZN(U3532) );
  AOI21_X1 U4883 ( .B1(n4313), .B2(n4325), .A(n4312), .ZN(n4395) );
  MUX2_X1 U4884 ( .A(n4314), .B(n4395), .S(n4559), .Z(n4315) );
  OAI21_X1 U4885 ( .B1(n4336), .B2(n4398), .A(n4315), .ZN(U3531) );
  OAI22_X1 U4886 ( .A1(n4318), .A2(n4329), .B1(n4317), .B2(n4316), .ZN(n4319)
         );
  INV_X1 U4887 ( .A(n4319), .ZN(n4320) );
  OAI211_X1 U4888 ( .C1(n4323), .C2(n4322), .A(n4321), .B(n4320), .ZN(n4324)
         );
  AOI21_X1 U4889 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(n4399) );
  MUX2_X1 U4890 ( .A(n4327), .B(n4399), .S(n4559), .Z(n4328) );
  OAI21_X1 U4891 ( .B1(n4336), .B2(n4402), .A(n4328), .ZN(U3530) );
  NOR2_X1 U4892 ( .A1(n4330), .A2(n4329), .ZN(n4332) );
  AOI211_X1 U4893 ( .C1(n4543), .C2(n4333), .A(n4332), .B(n4331), .ZN(n4403)
         );
  MUX2_X1 U4894 ( .A(n4334), .B(n4403), .S(n4559), .Z(n4335) );
  OAI21_X1 U4895 ( .B1(n4336), .B2(n4407), .A(n4335), .ZN(U3529) );
  NAND2_X1 U4896 ( .A1(n4553), .A2(n4337), .ZN(n4339) );
  NAND2_X1 U4897 ( .A1(n4551), .A2(REG0_REG_31__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U4898 ( .C1(n4340), .C2(n4406), .A(n4339), .B(n4338), .ZN(U3517)
         );
  INV_X1 U4899 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4341) );
  MUX2_X1 U4900 ( .A(n4341), .B(n4422), .S(n4553), .Z(n4342) );
  OAI21_X1 U4901 ( .B1(n4343), .B2(n4406), .A(n4342), .ZN(U3516) );
  MUX2_X1 U4902 ( .A(REG0_REG_27__SCAN_IN), .B(n4344), .S(n4553), .Z(n4345) );
  INV_X1 U4903 ( .A(n4348), .ZN(U3513) );
  INV_X1 U4904 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4350) );
  MUX2_X1 U4905 ( .A(n4350), .B(n4349), .S(n4553), .Z(n4351) );
  OAI21_X1 U4906 ( .B1(n4352), .B2(n4406), .A(n4351), .ZN(U3512) );
  INV_X1 U4907 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4354) );
  MUX2_X1 U4908 ( .A(n4354), .B(n4353), .S(n4553), .Z(n4355) );
  OAI21_X1 U4909 ( .B1(n4356), .B2(n4406), .A(n4355), .ZN(U3511) );
  INV_X1 U4910 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4358) );
  MUX2_X1 U4911 ( .A(n4358), .B(n4357), .S(n4553), .Z(n4359) );
  OAI21_X1 U4912 ( .B1(n4360), .B2(n4406), .A(n4359), .ZN(U3510) );
  INV_X1 U4913 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4362) );
  MUX2_X1 U4914 ( .A(n4362), .B(n4361), .S(n4553), .Z(n4363) );
  OAI21_X1 U4915 ( .B1(n4364), .B2(n4406), .A(n4363), .ZN(U3509) );
  INV_X1 U4916 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4366) );
  MUX2_X1 U4917 ( .A(n4366), .B(n4365), .S(n4553), .Z(n4367) );
  OAI21_X1 U4918 ( .B1(n4368), .B2(n4406), .A(n4367), .ZN(U3508) );
  INV_X1 U4919 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4370) );
  MUX2_X1 U4920 ( .A(n4370), .B(n4369), .S(n4553), .Z(n4371) );
  OAI21_X1 U4921 ( .B1(n4372), .B2(n4406), .A(n4371), .ZN(U3507) );
  INV_X1 U4922 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4374) );
  MUX2_X1 U4923 ( .A(n4374), .B(n4373), .S(n4553), .Z(n4375) );
  OAI21_X1 U4924 ( .B1(n4376), .B2(n4406), .A(n4375), .ZN(U3506) );
  INV_X1 U4925 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4378) );
  MUX2_X1 U4926 ( .A(n4378), .B(n4377), .S(n4553), .Z(n4379) );
  OAI21_X1 U4927 ( .B1(n4380), .B2(n4406), .A(n4379), .ZN(U3505) );
  MUX2_X1 U4928 ( .A(REG0_REG_18__SCAN_IN), .B(n4381), .S(n4553), .Z(U3503) );
  INV_X1 U4929 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4383) );
  MUX2_X1 U4930 ( .A(n4383), .B(n4382), .S(n4553), .Z(n4384) );
  OAI21_X1 U4931 ( .B1(n4385), .B2(n4406), .A(n4384), .ZN(U3501) );
  MUX2_X1 U4932 ( .A(REG0_REG_16__SCAN_IN), .B(n4386), .S(n4553), .Z(U3499) );
  INV_X1 U4933 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4388) );
  MUX2_X1 U4934 ( .A(n4388), .B(n4387), .S(n4553), .Z(n4389) );
  OAI21_X1 U4935 ( .B1(n4390), .B2(n4406), .A(n4389), .ZN(U3497) );
  INV_X1 U4936 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4392) );
  MUX2_X1 U4937 ( .A(n4392), .B(n4391), .S(n4553), .Z(n4393) );
  OAI21_X1 U4938 ( .B1(n4394), .B2(n4406), .A(n4393), .ZN(U3495) );
  INV_X1 U4939 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U4940 ( .A(n4396), .B(n4395), .S(n4553), .Z(n4397) );
  OAI21_X1 U4941 ( .B1(n4398), .B2(n4406), .A(n4397), .ZN(U3493) );
  INV_X1 U4942 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4400) );
  MUX2_X1 U4943 ( .A(n4400), .B(n4399), .S(n4553), .Z(n4401) );
  OAI21_X1 U4944 ( .B1(n4402), .B2(n4406), .A(n4401), .ZN(U3491) );
  INV_X1 U4945 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U4946 ( .A(n4404), .B(n4403), .S(n4553), .Z(n4405) );
  OAI21_X1 U4947 ( .B1(n4407), .B2(n4406), .A(n4405), .ZN(U3489) );
  MUX2_X1 U4948 ( .A(DATAI_30_), .B(n4408), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4949 ( .A(n4409), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4950 ( .A(n2690), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4951 ( .A(DATAI_22_), .B(n4410), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4952 ( .A(DATAI_20_), .B(n4411), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4953 ( .A(n4412), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4954 ( .A(DATAI_8_), .B(n4413), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4955 ( .A(DATAI_7_), .B(n4414), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4956 ( .A(n4415), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4957 ( .A(n4416), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4958 ( .A(DATAI_4_), .B(n4417), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4959 ( .A(DATAI_2_), .B(n4418), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  AOI22_X1 U4960 ( .A1(STATE_REG_SCAN_IN), .A2(n4419), .B1(n4687), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4961 ( .A1(n4420), .A2(n4519), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4525), .ZN(n4421) );
  OAI21_X1 U4962 ( .B1(n4525), .B2(n4422), .A(n4421), .ZN(U3261) );
  INV_X1 U4963 ( .A(n4425), .ZN(n4423) );
  OAI211_X1 U4964 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4424), .A(n4426), .B(n4423), 
        .ZN(n4429) );
  INV_X1 U4965 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U4966 ( .A1(n4426), .A2(n4425), .B1(n4507), .B2(n4554), .ZN(n4428)
         );
  AOI22_X1 U4967 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4505), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4427) );
  OAI221_X1 U4968 ( .B1(IR_REG_0__SCAN_IN), .B2(n4429), .C1(n2764), .C2(n4428), 
        .A(n4427), .ZN(U3240) );
  OAI211_X1 U4969 ( .C1(n4432), .C2(n4431), .A(n4464), .B(n4430), .ZN(n4437)
         );
  OAI211_X1 U4970 ( .C1(n4435), .C2(n4434), .A(n4507), .B(n4433), .ZN(n4436)
         );
  OAI211_X1 U4971 ( .C1(n4512), .C2(n4438), .A(n4437), .B(n4436), .ZN(n4439)
         );
  AOI211_X1 U4972 ( .C1(n4505), .C2(ADDR_REG_9__SCAN_IN), .A(n4440), .B(n4439), 
        .ZN(n4441) );
  INV_X1 U4973 ( .A(n4441), .ZN(U3249) );
  OAI211_X1 U4974 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4443), .A(n4464), .B(n4442), .ZN(n4445) );
  NAND2_X1 U4975 ( .A1(n4445), .A2(n4444), .ZN(n4446) );
  AOI21_X1 U4976 ( .B1(n4505), .B2(ADDR_REG_10__SCAN_IN), .A(n4446), .ZN(n4450) );
  OAI211_X1 U4977 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4448), .A(n4507), .B(n4447), .ZN(n4449) );
  OAI211_X1 U4978 ( .C1(n4512), .C2(n4534), .A(n4450), .B(n4449), .ZN(U3250)
         );
  OAI211_X1 U4979 ( .C1(n4453), .C2(n4452), .A(n4507), .B(n4451), .ZN(n4458)
         );
  OAI211_X1 U4980 ( .C1(n4456), .C2(n4455), .A(n4464), .B(n4454), .ZN(n4457)
         );
  OAI211_X1 U4981 ( .C1(n4512), .C2(n4533), .A(n4458), .B(n4457), .ZN(n4459)
         );
  AOI211_X1 U4982 ( .C1(n4505), .C2(ADDR_REG_11__SCAN_IN), .A(n4460), .B(n4459), .ZN(n4461) );
  INV_X1 U4983 ( .A(n4461), .ZN(U3251) );
  OAI211_X1 U4984 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4465), .A(n4464), .B(n4463), .ZN(n4467) );
  NAND2_X1 U4985 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AOI21_X1 U4986 ( .B1(n4505), .B2(ADDR_REG_12__SCAN_IN), .A(n4468), .ZN(n4472) );
  OAI211_X1 U4987 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4470), .A(n4507), .B(n4469), .ZN(n4471) );
  OAI211_X1 U4988 ( .C1(n4512), .C2(n2167), .A(n4472), .B(n4471), .ZN(U3252)
         );
  INV_X1 U4989 ( .A(n4473), .ZN(n4477) );
  AOI211_X1 U4990 ( .C1(n2451), .C2(n4475), .A(n4474), .B(n4501), .ZN(n4476)
         );
  AOI211_X1 U4991 ( .C1(n4505), .C2(ADDR_REG_14__SCAN_IN), .A(n4477), .B(n4476), .ZN(n4481) );
  OAI211_X1 U4992 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4479), .A(n4507), .B(n4478), .ZN(n4480) );
  OAI211_X1 U4993 ( .C1(n4512), .C2(n4531), .A(n4481), .B(n4480), .ZN(U3254)
         );
  AOI211_X1 U4994 ( .C1(n4484), .C2(n4483), .A(n4482), .B(n4501), .ZN(n4485)
         );
  AOI211_X1 U4995 ( .C1(n4505), .C2(ADDR_REG_15__SCAN_IN), .A(n4486), .B(n4485), .ZN(n4491) );
  OAI211_X1 U4996 ( .C1(n4489), .C2(n4488), .A(n4507), .B(n4487), .ZN(n4490)
         );
  OAI211_X1 U4997 ( .C1(n4512), .C2(n4530), .A(n4491), .B(n4490), .ZN(U3255)
         );
  INV_X1 U4998 ( .A(n4492), .ZN(n4496) );
  AOI221_X1 U4999 ( .B1(n4494), .B2(n4493), .C1(n2470), .C2(n4493), .A(n4501), 
        .ZN(n4495) );
  AOI211_X1 U5000 ( .C1(n4505), .C2(ADDR_REG_16__SCAN_IN), .A(n4496), .B(n4495), .ZN(n4500) );
  OAI221_X1 U5001 ( .B1(n4498), .B2(REG1_REG_16__SCAN_IN), .C1(n4498), .C2(
        n4497), .A(n4507), .ZN(n4499) );
  OAI211_X1 U5002 ( .C1(n4512), .C2(n4529), .A(n4500), .B(n4499), .ZN(U3256)
         );
  OAI211_X1 U5003 ( .C1(n4509), .C2(n4508), .A(n4507), .B(n4506), .ZN(n4510)
         );
  OAI211_X1 U5004 ( .C1(n4512), .C2(n4528), .A(n4511), .B(n4510), .ZN(U3258)
         );
  OAI22_X1 U5005 ( .A1(n4516), .A2(n4515), .B1(n4514), .B2(n4513), .ZN(n4517)
         );
  INV_X1 U5006 ( .A(n4517), .ZN(n4523) );
  AOI22_X1 U5007 ( .A1(n4521), .A2(n4520), .B1(n4519), .B2(n4518), .ZN(n4522)
         );
  OAI211_X1 U5008 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(U3282)
         );
  AND2_X1 U5009 ( .A1(D_REG_31__SCAN_IN), .A2(n4526), .ZN(U3291) );
  AND2_X1 U5010 ( .A1(D_REG_30__SCAN_IN), .A2(n4526), .ZN(U3292) );
  AND2_X1 U5011 ( .A1(D_REG_29__SCAN_IN), .A2(n4526), .ZN(U3293) );
  AND2_X1 U5012 ( .A1(D_REG_28__SCAN_IN), .A2(n4526), .ZN(U3294) );
  AND2_X1 U5013 ( .A1(D_REG_27__SCAN_IN), .A2(n4526), .ZN(U3295) );
  AND2_X1 U5014 ( .A1(D_REG_26__SCAN_IN), .A2(n4526), .ZN(U3296) );
  AND2_X1 U5015 ( .A1(D_REG_25__SCAN_IN), .A2(n4526), .ZN(U3297) );
  AND2_X1 U5016 ( .A1(D_REG_24__SCAN_IN), .A2(n4526), .ZN(U3298) );
  AND2_X1 U5017 ( .A1(D_REG_23__SCAN_IN), .A2(n4526), .ZN(U3299) );
  AND2_X1 U5018 ( .A1(D_REG_22__SCAN_IN), .A2(n4526), .ZN(U3300) );
  AND2_X1 U5019 ( .A1(D_REG_21__SCAN_IN), .A2(n4526), .ZN(U3301) );
  AND2_X1 U5020 ( .A1(D_REG_20__SCAN_IN), .A2(n4526), .ZN(U3302) );
  AND2_X1 U5021 ( .A1(D_REG_19__SCAN_IN), .A2(n4526), .ZN(U3303) );
  AND2_X1 U5022 ( .A1(D_REG_18__SCAN_IN), .A2(n4526), .ZN(U3304) );
  AND2_X1 U5023 ( .A1(D_REG_17__SCAN_IN), .A2(n4526), .ZN(U3305) );
  AND2_X1 U5024 ( .A1(D_REG_16__SCAN_IN), .A2(n4526), .ZN(U3306) );
  AND2_X1 U5025 ( .A1(D_REG_15__SCAN_IN), .A2(n4526), .ZN(U3307) );
  AND2_X1 U5026 ( .A1(D_REG_14__SCAN_IN), .A2(n4526), .ZN(U3308) );
  AND2_X1 U5027 ( .A1(D_REG_13__SCAN_IN), .A2(n4526), .ZN(U3309) );
  AND2_X1 U5028 ( .A1(D_REG_12__SCAN_IN), .A2(n4526), .ZN(U3310) );
  AND2_X1 U5029 ( .A1(D_REG_11__SCAN_IN), .A2(n4526), .ZN(U3311) );
  AND2_X1 U5030 ( .A1(D_REG_10__SCAN_IN), .A2(n4526), .ZN(U3312) );
  AND2_X1 U5031 ( .A1(D_REG_9__SCAN_IN), .A2(n4526), .ZN(U3313) );
  AND2_X1 U5032 ( .A1(D_REG_8__SCAN_IN), .A2(n4526), .ZN(U3314) );
  AND2_X1 U5033 ( .A1(D_REG_7__SCAN_IN), .A2(n4526), .ZN(U3315) );
  AND2_X1 U5034 ( .A1(D_REG_6__SCAN_IN), .A2(n4526), .ZN(U3316) );
  AND2_X1 U5035 ( .A1(D_REG_5__SCAN_IN), .A2(n4526), .ZN(U3317) );
  AND2_X1 U5036 ( .A1(D_REG_4__SCAN_IN), .A2(n4526), .ZN(U3318) );
  AND2_X1 U5037 ( .A1(D_REG_3__SCAN_IN), .A2(n4526), .ZN(U3319) );
  AND2_X1 U5038 ( .A1(D_REG_2__SCAN_IN), .A2(n4526), .ZN(U3320) );
  INV_X1 U5039 ( .A(DATAI_23_), .ZN(n4683) );
  AOI21_X1 U5040 ( .B1(U3149), .B2(n4683), .A(n4527), .ZN(U3329) );
  INV_X1 U5041 ( .A(DATAI_18_), .ZN(n4584) );
  AOI22_X1 U5042 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .B1(n4584), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5043 ( .A(DATAI_16_), .ZN(n4601) );
  AOI22_X1 U5044 ( .A1(STATE_REG_SCAN_IN), .A2(n4529), .B1(n4601), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n4530), .B1(n2466), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5046 ( .A(DATAI_14_), .ZN(n4589) );
  AOI22_X1 U5047 ( .A1(STATE_REG_SCAN_IN), .A2(n4531), .B1(n4589), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5048 ( .A(DATAI_12_), .ZN(n4574) );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n2167), .B1(n4574), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5050 ( .A(DATAI_11_), .ZN(n4532) );
  AOI22_X1 U5051 ( .A1(STATE_REG_SCAN_IN), .A2(n4533), .B1(n4532), .B2(U3149), 
        .ZN(U3341) );
  AOI22_X1 U5052 ( .A1(STATE_REG_SCAN_IN), .A2(n4534), .B1(n4721), .B2(U3149), 
        .ZN(U3342) );
  OAI211_X1 U5053 ( .C1(n4538), .C2(n4537), .A(n4536), .B(n4535), .ZN(n4539)
         );
  INV_X1 U5054 ( .A(n4539), .ZN(n4555) );
  AOI22_X1 U5055 ( .A1(n4553), .A2(n4555), .B1(n2295), .B2(n4551), .ZN(U3467)
         );
  INV_X1 U5056 ( .A(n4540), .ZN(n4542) );
  AOI211_X1 U5057 ( .C1(n4544), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4556)
         );
  AOI22_X1 U5058 ( .A1(n4553), .A2(n4556), .B1(n2328), .B2(n4551), .ZN(U3475)
         );
  OR3_X1 U5059 ( .A1(n4547), .A2(n4546), .A3(n4545), .ZN(n4550) );
  AND3_X1 U5060 ( .A1(n4550), .A2(n4549), .A3(n4548), .ZN(n4558) );
  INV_X1 U5061 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4552) );
  AOI22_X1 U5062 ( .A1(n4553), .A2(n4558), .B1(n4552), .B2(n4551), .ZN(U3481)
         );
  AOI22_X1 U5063 ( .A1(n4559), .A2(n4555), .B1(n4554), .B2(n4557), .ZN(U3518)
         );
  AOI22_X1 U5064 ( .A1(n4559), .A2(n4556), .B1(n2325), .B2(n4557), .ZN(U3522)
         );
  AOI22_X1 U5065 ( .A1(n4559), .A2(n4558), .B1(n2365), .B2(n4557), .ZN(U3525)
         );
  AOI22_X1 U5066 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4744) );
  INV_X1 U5067 ( .A(DATAI_19_), .ZN(n4561) );
  AOI22_X1 U5068 ( .A1(n4561), .A2(keyinput_g12), .B1(n2764), .B2(keyinput_g55), .ZN(n4560) );
  OAI221_X1 U5069 ( .B1(n4561), .B2(keyinput_g12), .C1(n2764), .C2(
        keyinput_g55), .A(n4560), .ZN(n4571) );
  AOI22_X1 U5070 ( .A1(n2446), .A2(keyinput_g18), .B1(n4684), .B2(keyinput_g45), .ZN(n4562) );
  OAI221_X1 U5071 ( .B1(n2446), .B2(keyinput_g18), .C1(n4684), .C2(
        keyinput_g45), .A(n4562), .ZN(n4570) );
  AOI22_X1 U5072 ( .A1(n4565), .A2(keyinput_g36), .B1(keyinput_g53), .B2(n4564), .ZN(n4563) );
  OAI221_X1 U5073 ( .B1(n4565), .B2(keyinput_g36), .C1(n4564), .C2(
        keyinput_g53), .A(n4563), .ZN(n4569) );
  XNOR2_X1 U5074 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_g42), .ZN(n4567) );
  XNOR2_X1 U5075 ( .A(DATAI_31_), .B(keyinput_g0), .ZN(n4566) );
  NAND2_X1 U5076 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  NOR4_X1 U5077 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4609)
         );
  AOI22_X1 U5078 ( .A1(DATAI_30_), .A2(keyinput_g1), .B1(DATAI_6_), .B2(
        keyinput_g25), .ZN(n4572) );
  OAI221_X1 U5079 ( .B1(DATAI_30_), .B2(keyinput_g1), .C1(DATAI_6_), .C2(
        keyinput_g25), .A(n4572), .ZN(n4582) );
  INV_X1 U5080 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5081 ( .A1(n4575), .A2(keyinput_g41), .B1(keyinput_g19), .B2(n4574), .ZN(n4573) );
  OAI221_X1 U5082 ( .B1(n4575), .B2(keyinput_g41), .C1(n4574), .C2(
        keyinput_g19), .A(n4573), .ZN(n4581) );
  AOI22_X1 U5083 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_g38), .ZN(n4576) );
  OAI221_X1 U5084 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(REG3_REG_3__SCAN_IN), 
        .C2(keyinput_g38), .A(n4576), .ZN(n4580) );
  XNOR2_X1 U5085 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4578) );
  XNOR2_X1 U5086 ( .A(DATAI_4_), .B(keyinput_g27), .ZN(n4577) );
  NAND2_X1 U5087 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  NOR4_X1 U5088 ( .A1(n4582), .A2(n4581), .A3(n4580), .A4(n4579), .ZN(n4608)
         );
  AOI22_X1 U5089 ( .A1(n3525), .A2(keyinput_g43), .B1(keyinput_g13), .B2(n4584), .ZN(n4583) );
  OAI221_X1 U5090 ( .B1(n3525), .B2(keyinput_g43), .C1(n4584), .C2(
        keyinput_g13), .A(n4583), .ZN(n4593) );
  AOI22_X1 U5091 ( .A1(n2604), .A2(keyinput_g4), .B1(keyinput_g11), .B2(n4586), 
        .ZN(n4585) );
  OAI221_X1 U5092 ( .B1(n2604), .B2(keyinput_g4), .C1(n4586), .C2(keyinput_g11), .A(n4585), .ZN(n4592) );
  INV_X1 U5093 ( .A(DATAI_0_), .ZN(n4722) );
  AOI22_X1 U5094 ( .A1(n4718), .A2(keyinput_g46), .B1(keyinput_g31), .B2(n4722), .ZN(n4587) );
  OAI221_X1 U5095 ( .B1(n4718), .B2(keyinput_g46), .C1(n4722), .C2(
        keyinput_g31), .A(n4587), .ZN(n4591) );
  AOI22_X1 U5096 ( .A1(n4589), .A2(keyinput_g17), .B1(U3149), .B2(keyinput_g32), .ZN(n4588) );
  OAI221_X1 U5097 ( .B1(n4589), .B2(keyinput_g17), .C1(U3149), .C2(
        keyinput_g32), .A(n4588), .ZN(n4590) );
  NOR4_X1 U5098 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4607)
         );
  AOI22_X1 U5099 ( .A1(n4596), .A2(keyinput_g2), .B1(keyinput_g9), .B2(n4595), 
        .ZN(n4594) );
  OAI221_X1 U5100 ( .B1(n4596), .B2(keyinput_g2), .C1(n4595), .C2(keyinput_g9), 
        .A(n4594), .ZN(n4605) );
  AOI22_X1 U5101 ( .A1(n4683), .A2(keyinput_g8), .B1(keyinput_g14), .B2(n4598), 
        .ZN(n4597) );
  OAI221_X1 U5102 ( .B1(n4683), .B2(keyinput_g8), .C1(n4598), .C2(keyinput_g14), .A(n4597), .ZN(n4604) );
  AOI22_X1 U5103 ( .A1(n2362), .A2(keyinput_g33), .B1(n3514), .B2(keyinput_g40), .ZN(n4599) );
  OAI221_X1 U5104 ( .B1(n2362), .B2(keyinput_g33), .C1(n3514), .C2(
        keyinput_g40), .A(n4599), .ZN(n4603) );
  AOI22_X1 U5105 ( .A1(n4601), .A2(keyinput_g15), .B1(keyinput_g16), .B2(n2466), .ZN(n4600) );
  OAI221_X1 U5106 ( .B1(n4601), .B2(keyinput_g15), .C1(n2466), .C2(
        keyinput_g16), .A(n4600), .ZN(n4602) );
  NOR4_X1 U5107 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4606)
         );
  NAND4_X1 U5108 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4742)
         );
  AOI22_X1 U5109 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_g47), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .ZN(n4610) );
  OAI221_X1 U5110 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_g47), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_g51), .A(n4610), .ZN(n4617) );
  AOI22_X1 U5111 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .ZN(n4611) );
  OAI221_X1 U5112 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_g44), .A(n4611), .ZN(n4616) );
  AOI22_X1 U5113 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n4612) );
  OAI221_X1 U5114 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n4612), .ZN(n4615) );
  AOI22_X1 U5115 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput_g35), .ZN(n4613) );
  OAI221_X1 U5116 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_g35), .A(n4613), .ZN(n4614) );
  NOR4_X1 U5117 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4644)
         );
  XOR2_X1 U5118 ( .A(DATAI_5_), .B(keyinput_g26), .Z(n4624) );
  AOI22_X1 U5119 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n4618) );
  OAI221_X1 U5120 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4618), .ZN(n4623) );
  AOI22_X1 U5121 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(DATAI_25_), .B2(
        keyinput_g6), .ZN(n4619) );
  OAI221_X1 U5122 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(DATAI_25_), .C2(
        keyinput_g6), .A(n4619), .ZN(n4622) );
  AOI22_X1 U5123 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n4620) );
  OAI221_X1 U5124 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n4620), .ZN(n4621) );
  NOR4_X1 U5125 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4643)
         );
  AOI22_X1 U5126 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(REG3_REG_17__SCAN_IN), 
        .B2(keyinput_g48), .ZN(n4625) );
  OAI221_X1 U5127 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(REG3_REG_17__SCAN_IN), .C2(keyinput_g48), .A(n4625), .ZN(n4632) );
  AOI22_X1 U5128 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n4626) );
  OAI221_X1 U5129 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_g63), .A(n4626), .ZN(n4631) );
  AOI22_X1 U5130 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n4627) );
  OAI221_X1 U5131 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n4627), .ZN(n4630) );
  AOI22_X1 U5132 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .ZN(n4628) );
  OAI221_X1 U5133 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_g34), .A(n4628), .ZN(n4629) );
  NOR4_X1 U5134 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(n4642)
         );
  AOI22_X1 U5135 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_g56), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4633) );
  OAI221_X1 U5136 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_g56), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4633), .ZN(n4640) );
  AOI22_X1 U5137 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n4634) );
  OAI221_X1 U5138 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_g62), .A(n4634), .ZN(n4639) );
  AOI22_X1 U5139 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_g50), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4635) );
  OAI221_X1 U5140 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4635), .ZN(n4638) );
  AOI22_X1 U5141 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_g58), .ZN(n4636) );
  OAI221_X1 U5142 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_g58), .A(n4636), .ZN(n4637) );
  NOR4_X1 U5143 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641)
         );
  NAND4_X1 U5144 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4741)
         );
  AOI22_X1 U5145 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4645) );
  OAI221_X1 U5146 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4645), .ZN(n4652) );
  AOI22_X1 U5147 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(DATAI_17_), .B2(
        keyinput_f14), .ZN(n4646) );
  OAI221_X1 U5148 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(DATAI_17_), .C2(
        keyinput_f14), .A(n4646), .ZN(n4651) );
  AOI22_X1 U5149 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(DATAI_15_), .B2(
        keyinput_f16), .ZN(n4647) );
  OAI221_X1 U5150 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(DATAI_15_), .C2(
        keyinput_f16), .A(n4647), .ZN(n4650) );
  AOI22_X1 U5151 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_f47), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4648) );
  OAI221_X1 U5152 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_f47), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4648), .ZN(n4649) );
  NOR4_X1 U5153 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4679)
         );
  XOR2_X1 U5154 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .Z(n4659) );
  AOI22_X1 U5155 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n4653) );
  OAI221_X1 U5156 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_f49), .A(n4653), .ZN(n4658) );
  AOI22_X1 U5157 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n4654) );
  OAI221_X1 U5158 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n4654), .ZN(n4657) );
  AOI22_X1 U5159 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4655) );
  OAI221_X1 U5160 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4655), .ZN(n4656) );
  NOR4_X1 U5161 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4678)
         );
  AOI22_X1 U5162 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .ZN(n4660) );
  OAI221_X1 U5163 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_f43), .A(n4660), .ZN(n4667) );
  AOI22_X1 U5164 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_f39), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4661) );
  OAI221_X1 U5165 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4661), .ZN(n4666) );
  AOI22_X1 U5166 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_f41), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .ZN(n4662) );
  OAI221_X1 U5167 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_f41), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4662), .ZN(n4665) );
  AOI22_X1 U5168 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4663) );
  OAI221_X1 U5169 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4663), .ZN(n4664) );
  NOR4_X1 U5170 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4677)
         );
  AOI22_X1 U5171 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_f33), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_f57), .ZN(n4668) );
  OAI221_X1 U5172 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_f33), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_f57), .A(n4668), .ZN(n4675) );
  AOI22_X1 U5173 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4669) );
  OAI221_X1 U5174 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4669), .ZN(n4674) );
  AOI22_X1 U5175 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(IR_REG_5__SCAN_IN), 
        .B2(keyinput_f60), .ZN(n4670) );
  OAI221_X1 U5176 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(IR_REG_5__SCAN_IN), 
        .C2(keyinput_f60), .A(n4670), .ZN(n4673) );
  AOI22_X1 U5177 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(IR_REG_3__SCAN_IN), 
        .B2(keyinput_f58), .ZN(n4671) );
  OAI221_X1 U5178 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(IR_REG_3__SCAN_IN), 
        .C2(keyinput_f58), .A(n4671), .ZN(n4672) );
  NOR4_X1 U5179 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4676)
         );
  NAND4_X1 U5180 ( .A1(n4679), .A2(n4678), .A3(n4677), .A4(n4676), .ZN(n4735)
         );
  AOI22_X1 U5181 ( .A1(n4681), .A2(keyinput_f48), .B1(keyinput_f18), .B2(n2446), .ZN(n4680) );
  OAI221_X1 U5182 ( .B1(n4681), .B2(keyinput_f48), .C1(n2446), .C2(
        keyinput_f18), .A(n4680), .ZN(n4693) );
  AOI22_X1 U5183 ( .A1(n4684), .A2(keyinput_f45), .B1(keyinput_f8), .B2(n4683), 
        .ZN(n4682) );
  OAI221_X1 U5184 ( .B1(n4684), .B2(keyinput_f45), .C1(n4683), .C2(keyinput_f8), .A(n4682), .ZN(n4692) );
  INV_X1 U5185 ( .A(DATAI_24_), .ZN(n4686) );
  AOI22_X1 U5186 ( .A1(n4687), .A2(keyinput_f3), .B1(keyinput_f7), .B2(n4686), 
        .ZN(n4685) );
  OAI221_X1 U5187 ( .B1(n4687), .B2(keyinput_f3), .C1(n4686), .C2(keyinput_f7), 
        .A(n4685), .ZN(n4691) );
  XNOR2_X1 U5188 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4689) );
  XNOR2_X1 U5189 ( .A(keyinput_f24), .B(DATAI_7_), .ZN(n4688) );
  NAND2_X1 U5190 ( .A1(n4689), .A2(n4688), .ZN(n4690) );
  NOR4_X1 U5191 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4733)
         );
  AOI22_X1 U5192 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(n3514), .B2(
        keyinput_f40), .ZN(n4694) );
  OAI221_X1 U5193 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(n3514), .C2(
        keyinput_f40), .A(n4694), .ZN(n4702) );
  AOI22_X1 U5194 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput_f32), .ZN(n4695) );
  OAI221_X1 U5195 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput_f32), .A(n4695), .ZN(n4701) );
  AOI22_X1 U5196 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n4696) );
  OAI221_X1 U5197 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_f62), .A(n4696), .ZN(n4700) );
  XNOR2_X1 U5198 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_f52), .ZN(n4698) );
  XNOR2_X1 U5199 ( .A(DATAI_26_), .B(keyinput_f5), .ZN(n4697) );
  NAND2_X1 U5200 ( .A1(n4698), .A2(n4697), .ZN(n4699) );
  NOR4_X1 U5201 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4732)
         );
  AOI22_X1 U5202 ( .A1(n4704), .A2(keyinput_f37), .B1(keyinput_f26), .B2(n2349), .ZN(n4703) );
  OAI221_X1 U5203 ( .B1(n4704), .B2(keyinput_f37), .C1(n2349), .C2(
        keyinput_f26), .A(n4703), .ZN(n4716) );
  INV_X1 U5204 ( .A(IR_REG_8__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5205 ( .A1(n4707), .A2(keyinput_f63), .B1(keyinput_f0), .B2(n4706), 
        .ZN(n4705) );
  OAI221_X1 U5206 ( .B1(n4707), .B2(keyinput_f63), .C1(n4706), .C2(keyinput_f0), .A(n4705), .ZN(n4715) );
  INV_X1 U5207 ( .A(DATAI_8_), .ZN(n4710) );
  AOI22_X1 U5208 ( .A1(n4710), .A2(keyinput_f23), .B1(keyinput_f1), .B2(n4709), 
        .ZN(n4708) );
  OAI221_X1 U5209 ( .B1(n4710), .B2(keyinput_f23), .C1(n4709), .C2(keyinput_f1), .A(n4708), .ZN(n4714) );
  XOR2_X1 U5210 ( .A(n2582), .B(keyinput_f6), .Z(n4712) );
  XNOR2_X1 U5211 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4711) );
  NAND2_X1 U5212 ( .A1(n4712), .A2(n4711), .ZN(n4713) );
  NOR4_X1 U5213 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4731)
         );
  AOI22_X1 U5214 ( .A1(n4718), .A2(keyinput_f46), .B1(keyinput_f54), .B2(n2435), .ZN(n4717) );
  OAI221_X1 U5215 ( .B1(n4718), .B2(keyinput_f46), .C1(n2435), .C2(
        keyinput_f54), .A(n4717), .ZN(n4729) );
  AOI22_X1 U5216 ( .A1(n4721), .A2(keyinput_f21), .B1(n4720), .B2(keyinput_f10), .ZN(n4719) );
  OAI221_X1 U5217 ( .B1(n4721), .B2(keyinput_f21), .C1(n4720), .C2(
        keyinput_f10), .A(n4719), .ZN(n4728) );
  XOR2_X1 U5218 ( .A(n4722), .B(keyinput_f31), .Z(n4726) );
  XNOR2_X1 U5219 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4725) );
  XNOR2_X1 U5220 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_f35), .ZN(n4724) );
  XNOR2_X1 U5221 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4723) );
  NAND4_X1 U5222 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4727)
         );
  NOR3_X1 U5223 ( .A1(n4729), .A2(n4728), .A3(n4727), .ZN(n4730) );
  NAND4_X1 U5224 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4734)
         );
  OAI22_X1 U5225 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(n4735), .B2(n4734), 
        .ZN(n4737) );
  NAND2_X1 U5226 ( .A1(n4737), .A2(keyinput_g30), .ZN(n4739) );
  INV_X1 U5227 ( .A(keyinput_g30), .ZN(n4736) );
  OAI211_X1 U5228 ( .C1(n4737), .C2(keyinput_f30), .A(DATAI_1_), .B(n4736), 
        .ZN(n4738) );
  OAI21_X1 U5229 ( .B1(DATAI_1_), .B2(n4739), .A(n4738), .ZN(n4740) );
  OAI21_X1 U5230 ( .B1(n4742), .B2(n4741), .A(n4740), .ZN(n4743) );
  XOR2_X1 U5231 ( .A(n4744), .B(n4743), .Z(U3352) );
  CLKBUF_X3 U2293 ( .A(n2887), .Z(n3462) );
  NAND2_X2 U2299 ( .A1(n2836), .A2(n2835), .ZN(n3503) );
  CLKBUF_X1 U2300 ( .A(n2314), .Z(n2488) );
  AND2_X1 U2310 ( .A1(n3003), .A2(n2335), .ZN(n3066) );
  CLKBUF_X2 U2317 ( .A(n2450), .Z(n2610) );
endmodule

