

module b17_C_SARLock_k_128_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9760, n9761, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9794, n9795, n9796, n9798, n9799, n9800,
         n9801, n9802, n9805, n9808, n9809, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461;

  AOI211_X1 U11192 ( .C1(n16265), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14607) );
  INV_X1 U11194 ( .A(n20210), .ZN(n20218) );
  NOR2_X1 U11195 ( .A1(n9876), .A2(n14974), .ZN(n14975) );
  XNOR2_X1 U11196 ( .A(n12843), .B(n12839), .ZN(n14981) );
  INV_X2 U11197 ( .A(n10005), .ZN(n18405) );
  NAND2_X1 U11198 ( .A1(n10180), .A2(n10178), .ZN(n19141) );
  OR2_X1 U11199 ( .A1(n14152), .A2(n20408), .ZN(n14120) );
  XNOR2_X1 U11200 ( .A(n12320), .B(n12319), .ZN(n15126) );
  OR2_X1 U11201 ( .A1(n11731), .A2(n11714), .ZN(n19507) );
  NAND2_X1 U11204 ( .A1(n12330), .A2(n10294), .ZN(n12325) );
  XNOR2_X1 U11205 ( .A(n13261), .B(n12670), .ZN(n13283) );
  BUF_X1 U11206 ( .A(n10416), .Z(n17381) );
  INV_X2 U11207 ( .A(n11638), .ZN(n11860) );
  BUF_X2 U11208 ( .A(n11817), .Z(n12731) );
  INV_X2 U11209 ( .A(n17427), .ZN(n15843) );
  BUF_X2 U11210 ( .A(n15914), .Z(n17433) );
  AND2_X1 U11211 ( .A1(n12766), .A2(n11754), .ZN(n11768) );
  AND2_X1 U11212 ( .A1(n15661), .A2(n12766), .ZN(n12500) );
  AND2_X1 U11213 ( .A1(n9968), .A2(n9972), .ZN(n10641) );
  INV_X4 U11214 ( .A(n9873), .ZN(n9763) );
  CLKBUF_X2 U11215 ( .A(n10505), .Z(n11399) );
  CLKBUF_X2 U11216 ( .A(n10525), .Z(n11402) );
  CLKBUF_X1 U11217 ( .A(n11023), .Z(n11478) );
  INV_X2 U11219 ( .A(n17473), .ZN(n15874) );
  INV_X2 U11220 ( .A(n17450), .ZN(n15877) );
  INV_X1 U11221 ( .A(n10496), .ZN(n9760) );
  AND4_X1 U11222 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10550) );
  NAND4_X2 U11223 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10552) );
  AND4_X1 U11224 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10482) );
  NAND2_X1 U11226 ( .A1(n13563), .A2(n21260), .ZN(n10544) );
  AND2_X2 U11228 ( .A1(n11753), .A2(n16597), .ZN(n11551) );
  AND2_X1 U11230 ( .A1(n9971), .A2(n20412), .ZN(n9969) );
  CLKBUF_X3 U11231 ( .A(n11327), .Z(n11300) );
  AOI22_X1 U11232 ( .A1(n21336), .A2(keyinput68), .B1(n21335), .B2(keyinput78), 
        .ZN(n21334) );
  AOI21_X1 U11233 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21335), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11189) );
  NOR2_X1 U11234 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  NAND2_X1 U11235 ( .A1(n10893), .A2(n10755), .ZN(n10881) );
  NOR2_X1 U11236 ( .A1(n12027), .A2(n10246), .ZN(n12040) );
  AND2_X1 U11237 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11753) );
  OAI221_X1 U11238 ( .B1(n21336), .B2(keyinput68), .C1(n21335), .C2(keyinput78), .A(n21334), .ZN(n21340) );
  AND2_X1 U11239 ( .A1(n13563), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10525) );
  AND2_X1 U11240 ( .A1(n11883), .A2(n11884), .ZN(n11874) );
  NAND2_X2 U11241 ( .A1(n11626), .A2(n13285), .ZN(n12175) );
  CLKBUF_X3 U11242 ( .A(n11602), .Z(n12926) );
  AND2_X1 U11243 ( .A1(n11755), .A2(n12766), .ZN(n11769) );
  AND2_X1 U11244 ( .A1(n11506), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15661) );
  AND2_X2 U11245 ( .A1(n11744), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12141) );
  AOI22_X1 U11246 ( .A1(n21139), .A2(keyinput49), .B1(keyinput124), .B2(n21138), .ZN(n21137) );
  AND4_X1 U11247 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10520) );
  INV_X1 U11248 ( .A(n14120), .ZN(n14139) );
  INV_X2 U11249 ( .A(n12175), .ZN(n14870) );
  OR2_X1 U11250 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  XNOR2_X1 U11251 ( .A(n12797), .B(n12821), .ZN(n15061) );
  OR2_X1 U11252 ( .A1(n11708), .A2(n10117), .ZN(n19876) );
  INV_X1 U11254 ( .A(n17130), .ZN(n17156) );
  NOR3_X1 U11255 ( .A1(n19121), .A2(n19108), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13964) );
  OAI221_X1 U11256 ( .B1(n21139), .B2(keyinput49), .C1(n21138), .C2(
        keyinput124), .A(n21137), .ZN(n21140) );
  NAND2_X1 U11257 ( .A1(n18091), .A2(n18092), .ZN(n18090) );
  AND2_X2 U11258 ( .A1(n20398), .A2(n20408), .ZN(n14149) );
  NAND2_X1 U11259 ( .A1(n14412), .A2(n10359), .ZN(n14395) );
  INV_X1 U11260 ( .A(n14582), .ZN(n16212) );
  AND2_X1 U11261 ( .A1(n10917), .A2(n9935), .ZN(n14560) );
  NAND2_X1 U11262 ( .A1(n11615), .A2(n11611), .ZN(n20143) );
  CLKBUF_X3 U11263 ( .A(n11862), .Z(n9789) );
  NAND2_X1 U11264 ( .A1(n10111), .A2(n10402), .ZN(n12843) );
  NAND2_X1 U11265 ( .A1(n12667), .A2(n12666), .ZN(n13261) );
  AND2_X1 U11266 ( .A1(n14363), .A2(n14215), .ZN(n20257) );
  OR2_X1 U11267 ( .A1(n9781), .A2(n9782), .ZN(n14246) );
  BUF_X1 U11268 ( .A(n10215), .Z(n9755) );
  AND2_X1 U11270 ( .A1(n10391), .A2(n14956), .ZN(n14966) );
  NAND2_X1 U11271 ( .A1(n14991), .A2(n14994), .ZN(n14993) );
  NOR2_X1 U11272 ( .A1(n10037), .A2(n9951), .ZN(n15163) );
  AND2_X1 U11273 ( .A1(n10049), .A2(n10048), .ZN(n15223) );
  NAND2_X1 U11274 ( .A1(n15642), .A2(n12303), .ZN(n15320) );
  NOR2_X1 U11275 ( .A1(n19949), .A2(n19662), .ZN(n19711) );
  INV_X2 U11276 ( .A(n17449), .ZN(n17365) );
  INV_X2 U11277 ( .A(n9947), .ZN(n17436) );
  INV_X1 U11278 ( .A(n20257), .ZN(n20285) );
  OAI21_X1 U11279 ( .B1(n14257), .B2(n14258), .A(n14246), .ZN(n14603) );
  INV_X1 U11280 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21027) );
  OR2_X1 U11282 ( .A1(n18047), .A2(n15909), .ZN(n9747) );
  AND2_X1 U11283 ( .A1(n10729), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9748) );
  AND2_X2 U11284 ( .A1(n11954), .A2(n11953), .ZN(n11969) );
  AND2_X2 U11285 ( .A1(n11610), .A2(n12955), .ZN(n11615) );
  AND2_X1 U11286 ( .A1(n9976), .A2(n10441), .ZN(n9749) );
  AND2_X1 U11287 ( .A1(n9976), .A2(n10441), .ZN(n10505) );
  AND3_X1 U11290 ( .A1(n11859), .A2(n11858), .A3(n11857), .ZN(n9750) );
  INV_X4 U11291 ( .A(n10416), .ZN(n17468) );
  NAND2_X2 U11292 ( .A1(n11619), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11649) );
  NAND3_X1 U11293 ( .A1(n13565), .A2(n10928), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11371) );
  AND2_X2 U11294 ( .A1(n10928), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U11295 ( .A1(n9982), .A2(n9981), .ZN(n11992) );
  NAND2_X4 U11296 ( .A1(n10550), .A2(n10549), .ZN(n20408) );
  INV_X2 U11297 ( .A(n13961), .ZN(n17449) );
  OAI21_X1 U11299 ( .B1(n15126), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10307), 
        .ZN(n13788) );
  OR2_X4 U11300 ( .A1(n18939), .A2(n13955), .ZN(n15718) );
  BUF_X1 U11301 ( .A(n11023), .Z(n9752) );
  CLKBUF_X1 U11302 ( .A(n11023), .Z(n9796) );
  OAI21_X2 U11303 ( .B1(n13603), .B2(n10374), .A(n10769), .ZN(n13531) );
  XNOR2_X2 U11304 ( .A(n10685), .B(n10642), .ZN(n20496) );
  AOI221_X2 U11305 ( .B1(n14810), .B2(n14847), .C1(n14701), .C2(n14847), .A(
        n14700), .ZN(n14801) );
  NOR2_X2 U11306 ( .A1(n14395), .A2(n14396), .ZN(n14293) );
  OAI21_X1 U11307 ( .B1(n15320), .B2(n10263), .A(n10260), .ZN(n16539) );
  CLKBUF_X1 U11308 ( .A(n12304), .Z(n9772) );
  NAND2_X1 U11309 ( .A1(n15014), .A2(n12541), .ZN(n14886) );
  NOR2_X1 U11310 ( .A1(n19912), .A2(n20103), .ZN(n19832) );
  INV_X4 U11312 ( .A(n10070), .ZN(n9753) );
  AOI211_X1 U11313 ( .C1(n13887), .C2(n20110), .A(n19491), .B(n20102), .ZN(
        n13879) );
  OR2_X1 U11314 ( .A1(n11725), .A2(n10117), .ZN(n19847) );
  NAND2_X2 U11315 ( .A1(n13200), .A2(n9908), .ZN(n10289) );
  XNOR2_X1 U11316 ( .A(n12164), .B(n12165), .ZN(n12654) );
  NAND2_X2 U11317 ( .A1(n18952), .A2(n18929), .ZN(n10005) );
  NAND2_X1 U11318 ( .A1(n12047), .A2(n12049), .ZN(n12053) );
  INV_X2 U11319 ( .A(n9747), .ZN(n9788) );
  NAND2_X1 U11320 ( .A1(n10641), .A2(n10630), .ZN(n13129) );
  AND4_X1 U11321 ( .A1(n9841), .A2(n11549), .A3(n11550), .A4(n10266), .ZN(
        n11625) );
  NAND2_X1 U11322 ( .A1(n20152), .A2(n20155), .ZN(n11624) );
  INV_X1 U11323 ( .A(n17666), .ZN(n18479) );
  CLKBUF_X1 U11324 ( .A(n11641), .Z(n9785) );
  INV_X1 U11325 ( .A(n9805), .ZN(n9761) );
  INV_X1 U11326 ( .A(n11402), .ZN(n9756) );
  INV_X2 U11327 ( .A(n11373), .ZN(n11453) );
  INV_X4 U11328 ( .A(n9878), .ZN(n17349) );
  INV_X1 U11329 ( .A(n10661), .ZN(n9805) );
  INV_X4 U11330 ( .A(n17483), .ZN(n17417) );
  INV_X1 U11332 ( .A(n11473), .ZN(n9757) );
  CLKBUF_X1 U11333 ( .A(n11551), .Z(n12901) );
  AND2_X2 U11334 ( .A1(n11752), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U11335 ( .A1(n10439), .A2(n10438), .ZN(n11446) );
  NAND2_X2 U11336 ( .A1(n13565), .A2(n10424), .ZN(n11369) );
  NAND3_X1 U11337 ( .A1(n16597), .A2(n11506), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11601) );
  NOR2_X1 U11339 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17190) );
  AND2_X1 U11340 ( .A1(n10033), .A2(n15489), .ZN(n16515) );
  AND2_X1 U11341 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  OR2_X1 U11342 ( .A1(n12649), .A2(n16558), .ZN(n12314) );
  OAI21_X1 U11343 ( .B1(n10034), .B2(n21229), .A(n12097), .ZN(n10033) );
  AOI21_X1 U11344 ( .B1(n14196), .B2(n20378), .A(n11503), .ZN(n11504) );
  AOI211_X1 U11345 ( .C1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n20271), .A(
        n16093), .B(n16092), .ZN(n16094) );
  NAND2_X1 U11346 ( .A1(n14981), .A2(n14980), .ZN(n14979) );
  NAND3_X1 U11347 ( .A1(n10347), .A2(n10346), .A3(n10348), .ZN(n14196) );
  NOR2_X1 U11348 ( .A1(n15257), .A2(n15246), .ZN(n15245) );
  OR2_X1 U11349 ( .A1(n15489), .A2(n15525), .ZN(n15260) );
  NOR2_X1 U11350 ( .A1(n10037), .A2(n10038), .ZN(n15174) );
  AND2_X1 U11351 ( .A1(n10018), .A2(n10070), .ZN(n14559) );
  INV_X1 U11352 ( .A(n14631), .ZN(n16091) );
  NAND2_X1 U11353 ( .A1(n15622), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15621) );
  NAND2_X1 U11354 ( .A1(n15622), .A2(n12623), .ZN(n15424) );
  OAI22_X1 U11355 ( .A1(n15312), .A2(n10058), .B1(n10124), .B2(n10059), .ZN(
        n15538) );
  AND2_X1 U11356 ( .A1(n14395), .A2(n16103), .ZN(n16204) );
  NAND2_X1 U11357 ( .A1(n10068), .A2(n10072), .ZN(n10020) );
  NAND2_X1 U11358 ( .A1(n10341), .A2(n9928), .ZN(n9988) );
  NAND2_X1 U11359 ( .A1(n10913), .A2(n10070), .ZN(n14627) );
  AND2_X1 U11360 ( .A1(n15072), .A2(n12821), .ZN(n12798) );
  OR2_X1 U11361 ( .A1(n14307), .A2(n11171), .ZN(n14419) );
  AND2_X1 U11362 ( .A1(n10201), .A2(n9901), .ZN(n10060) );
  AOI21_X1 U11363 ( .B1(n10264), .B2(n10262), .A(n10261), .ZN(n10260) );
  NOR2_X1 U11364 ( .A1(n14950), .A2(n12563), .ZN(n14875) );
  OR2_X1 U11365 ( .A1(n15318), .A2(n16569), .ZN(n10264) );
  INV_X1 U11366 ( .A(n15361), .ZN(n16433) );
  NAND2_X1 U11367 ( .A1(n12297), .A2(n13826), .ZN(n10270) );
  XNOR2_X1 U11368 ( .A(n12306), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16540) );
  NAND2_X1 U11369 ( .A1(n10045), .A2(n11905), .ZN(n13836) );
  NAND2_X1 U11370 ( .A1(n11020), .A2(n11019), .ZN(n13935) );
  NAND2_X1 U11371 ( .A1(n14886), .A2(n12542), .ZN(n15343) );
  NAND2_X1 U11372 ( .A1(n10093), .A2(n10311), .ZN(n10310) );
  NAND2_X1 U11373 ( .A1(n10312), .A2(n10313), .ZN(n16709) );
  NOR2_X1 U11374 ( .A1(n9872), .A2(n12633), .ZN(n15012) );
  NAND2_X1 U11375 ( .A1(n12985), .A2(n12227), .ZN(n13018) );
  AND2_X1 U11376 ( .A1(n12296), .A2(n12295), .ZN(n13826) );
  NOR2_X1 U11377 ( .A1(n16006), .A2(n21361), .ZN(n10311) );
  NOR2_X1 U11378 ( .A1(n15171), .A2(n10131), .ZN(n10130) );
  NOR2_X1 U11379 ( .A1(n10345), .A2(n10344), .ZN(n10343) );
  AND2_X1 U11380 ( .A1(n12277), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13828) );
  NAND2_X1 U11381 ( .A1(n12014), .A2(n12298), .ZN(n12304) );
  NOR3_X1 U11382 ( .A1(n14645), .A2(n16230), .A3(n14647), .ZN(n10904) );
  NAND2_X1 U11383 ( .A1(n15264), .A2(n15263), .ZN(n15266) );
  AND2_X1 U11384 ( .A1(n12120), .A2(n10255), .ZN(n14915) );
  NOR2_X1 U11385 ( .A1(n10385), .A2(n10384), .ZN(n10383) );
  NOR2_X1 U11386 ( .A1(n13751), .A2(n13750), .ZN(n13730) );
  NAND2_X1 U11387 ( .A1(n10828), .A2(n10827), .ZN(n16262) );
  NOR3_X1 U11388 ( .A1(n17827), .A2(n16004), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U11389 ( .A1(n9877), .A2(n13665), .ZN(n15300) );
  XNOR2_X1 U11390 ( .A(n14150), .B(n10200), .ZN(n14689) );
  AND2_X1 U11391 ( .A1(n12013), .A2(n12012), .ZN(n12298) );
  AND2_X1 U11392 ( .A1(n10151), .A2(n10150), .ZN(n16859) );
  NAND2_X1 U11393 ( .A1(n10982), .A2(n10981), .ZN(n13802) );
  NAND2_X1 U11394 ( .A1(n13731), .A2(n11001), .ZN(n10344) );
  OAI211_X1 U11395 ( .C1(n11112), .C2(n20322), .A(n10973), .B(n10972), .ZN(
        n13731) );
  NAND2_X1 U11396 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18068), .ZN(n17985) );
  OR2_X1 U11397 ( .A1(n10906), .A2(n16330), .ZN(n14654) );
  NAND2_X1 U11398 ( .A1(n10883), .A2(n10895), .ZN(n10906) );
  INV_X2 U11399 ( .A(n18136), .ZN(n18122) );
  OR2_X1 U11400 ( .A1(n11799), .A2(n11798), .ZN(n11802) );
  OAI22_X1 U11401 ( .A1(n11733), .A2(n11992), .B1(n11980), .B2(n11732), .ZN(
        n11739) );
  OR2_X1 U11402 ( .A1(n11706), .A2(n11705), .ZN(n11713) );
  NAND2_X1 U11403 ( .A1(n10821), .A2(n9855), .ZN(n10871) );
  NOR2_X1 U11404 ( .A1(n13444), .A2(n13445), .ZN(n13775) );
  AND2_X1 U11405 ( .A1(n13535), .A2(n13534), .ZN(n14842) );
  AND2_X1 U11406 ( .A1(n12664), .A2(n12684), .ZN(n13350) );
  NAND2_X1 U11407 ( .A1(n10821), .A2(n9860), .ZN(n10883) );
  NAND2_X1 U11408 ( .A1(n15590), .A2(n13424), .ZN(n15569) );
  INV_X1 U11409 ( .A(n13818), .ZN(n14844) );
  NAND2_X1 U11410 ( .A1(n11717), .A2(n11716), .ZN(n19916) );
  NOR2_X1 U11411 ( .A1(n13702), .A2(n13343), .ZN(n13395) );
  NAND2_X1 U11412 ( .A1(n10354), .A2(n14258), .ZN(n10353) );
  OR2_X1 U11413 ( .A1(n12681), .A2(n12680), .ZN(n13311) );
  NAND2_X1 U11414 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NAND2_X1 U11415 ( .A1(n13373), .A2(n13403), .ZN(n13390) );
  BUF_X2 U11416 ( .A(n12654), .Z(n9839) );
  NOR2_X1 U11417 ( .A1(n14440), .A2(n14434), .ZN(n14436) );
  NOR2_X1 U11418 ( .A1(n18949), .A2(n17521), .ZN(n17653) );
  AND2_X1 U11419 ( .A1(n13830), .A2(n12415), .ZN(n13200) );
  NAND3_X1 U11420 ( .A1(n9985), .A2(n9983), .A3(n10330), .ZN(n12164) );
  NAND2_X1 U11421 ( .A1(n10239), .A2(n10238), .ZN(n12081) );
  NAND2_X1 U11422 ( .A1(n10921), .A2(n10922), .ZN(n10725) );
  AOI21_X1 U11423 ( .B1(n20680), .B2(n21027), .A(n10076), .ZN(n13653) );
  INV_X1 U11424 ( .A(n12053), .ZN(n10239) );
  XNOR2_X1 U11425 ( .A(n10717), .B(n10722), .ZN(n10921) );
  NOR2_X2 U11426 ( .A1(n19468), .A2(n19917), .ZN(n19469) );
  OR2_X1 U11427 ( .A1(n16353), .A2(n16352), .ZN(n16355) );
  XNOR2_X1 U11428 ( .A(n10142), .B(n20535), .ZN(n20680) );
  INV_X1 U11429 ( .A(n16056), .ZN(n13368) );
  NAND2_X1 U11430 ( .A1(n10732), .A2(n10731), .ZN(n10142) );
  AND2_X1 U11431 ( .A1(n10274), .A2(n10276), .ZN(n13606) );
  AOI21_X1 U11432 ( .B1(n10718), .B2(n10721), .A(n10720), .ZN(n10922) );
  OR2_X1 U11433 ( .A1(n12399), .A2(n13296), .ZN(n10274) );
  NAND2_X1 U11434 ( .A1(n10278), .A2(n10277), .ZN(n10276) );
  NAND4_X1 U11435 ( .A1(n10105), .A2(n11657), .A3(n11658), .A4(n11649), .ZN(
        n11689) );
  AND2_X1 U11436 ( .A1(n16392), .A2(n13909), .ZN(n16378) );
  AND2_X1 U11437 ( .A1(n13669), .A2(n12040), .ZN(n12048) );
  AOI21_X1 U11438 ( .B1(n9801), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11670), .ZN(n11675) );
  INV_X1 U11439 ( .A(n15938), .ZN(n10308) );
  OR2_X1 U11440 ( .A1(n13277), .A2(n13276), .ZN(n13279) );
  OR2_X1 U11441 ( .A1(n13624), .A2(n13625), .ZN(n13739) );
  NAND2_X2 U11442 ( .A1(n17725), .A2(n17724), .ZN(n17752) );
  AOI21_X1 U11443 ( .B1(n10053), .B2(n10052), .A(n9885), .ZN(n11688) );
  OR2_X1 U11444 ( .A1(n13545), .A2(n13544), .ZN(n13624) );
  AND2_X1 U11445 ( .A1(n15948), .A2(n10170), .ZN(n18928) );
  AOI21_X1 U11446 ( .B1(n15673), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10107), 
        .ZN(n10106) );
  AND2_X1 U11447 ( .A1(n13208), .A2(n13207), .ZN(n13210) );
  NOR2_X2 U11448 ( .A1(n19157), .A2(n15946), .ZN(n18947) );
  NAND2_X1 U11449 ( .A1(n18106), .A2(n18105), .ZN(n18104) );
  AND2_X1 U11450 ( .A1(n11656), .A2(n11655), .ZN(n11657) );
  NOR2_X1 U11451 ( .A1(n11906), .A2(n10235), .ZN(n10234) );
  XNOR2_X1 U11452 ( .A(n15931), .B(n18422), .ZN(n18106) );
  INV_X1 U11453 ( .A(n12052), .ZN(n10238) );
  NOR2_X2 U11454 ( .A1(n11861), .A2(n11879), .ZN(n11884) );
  INV_X1 U11455 ( .A(n12175), .ZN(n9758) );
  NAND2_X1 U11456 ( .A1(n10236), .A2(n10237), .ZN(n11873) );
  INV_X1 U11457 ( .A(n14103), .ZN(n14146) );
  AND2_X1 U11458 ( .A1(n10638), .A2(n13233), .ZN(n10630) );
  CLKBUF_X2 U11459 ( .A(n11625), .Z(n13285) );
  AND2_X1 U11460 ( .A1(n14143), .A2(n14149), .ZN(n14103) );
  NAND2_X1 U11461 ( .A1(n13224), .A2(n14197), .ZN(n13378) );
  AND2_X2 U11462 ( .A1(n12587), .A2(n11651), .ZN(n14869) );
  INV_X1 U11463 ( .A(n19141), .ZN(n18484) );
  NOR2_X2 U11464 ( .A1(n11624), .A2(n12578), .ZN(n11626) );
  NOR2_X2 U11465 ( .A1(n12352), .A2(n19191), .ZN(n12334) );
  NAND3_X2 U11466 ( .A1(n12390), .A2(n16624), .A3(n11860), .ZN(n14883) );
  AND3_X1 U11467 ( .A1(n13382), .A2(n21102), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10637) );
  AND4_X2 U11468 ( .A1(n9890), .A2(n10554), .A3(n10625), .A4(n10633), .ZN(
        n13246) );
  AND2_X1 U11469 ( .A1(n10880), .A2(n13128), .ZN(n10606) );
  INV_X1 U11470 ( .A(n11624), .ZN(n11651) );
  NAND2_X1 U11471 ( .A1(n11548), .A2(n11638), .ZN(n12389) );
  NAND2_X1 U11472 ( .A1(n12353), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12352) );
  AND2_X1 U11473 ( .A1(n10627), .A2(n9890), .ZN(n13132) );
  AND2_X1 U11474 ( .A1(n10553), .A2(n20424), .ZN(n10633) );
  NOR2_X1 U11475 ( .A1(n12629), .A2(n11623), .ZN(n11611) );
  INV_X2 U11476 ( .A(n20155), .ZN(n16624) );
  AND2_X1 U11477 ( .A1(n15888), .A2(n10408), .ZN(n17660) );
  AND2_X1 U11478 ( .A1(n10628), .A2(n13361), .ZN(n13564) );
  NAND2_X1 U11479 ( .A1(n13338), .A2(n14152), .ZN(n13229) );
  OAI211_X1 U11480 ( .C1(n17483), .C2(n17490), .A(n13973), .B(n13972), .ZN(
        n17625) );
  AND2_X1 U11481 ( .A1(n10623), .A2(n20424), .ZN(n14197) );
  INV_X1 U11482 ( .A(n19476), .ZN(n12580) );
  OR2_X1 U11483 ( .A1(n11917), .A2(n11916), .ZN(n12411) );
  INV_X1 U11484 ( .A(n9765), .ZN(n10623) );
  OR2_X1 U11485 ( .A1(n11786), .A2(n11785), .ZN(n12394) );
  INV_X1 U11486 ( .A(n10552), .ZN(n13324) );
  AND2_X1 U11487 ( .A1(n15926), .A2(n15927), .ZN(n18134) );
  AND2_X2 U11488 ( .A1(n10620), .A2(n10552), .ZN(n13216) );
  OAI211_X1 U11489 ( .C1(n15718), .C2(n17509), .A(n15873), .B(n15872), .ZN(
        n17652) );
  OR2_X1 U11490 ( .A1(n11827), .A2(n11826), .ZN(n12402) );
  MUX2_X1 U11491 ( .A(n11573), .B(n11572), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12362) );
  INV_X2 U11492 ( .A(U212), .ZN(n16773) );
  NAND2_X1 U11493 ( .A1(n11595), .A2(n11594), .ZN(n12629) );
  AND2_X1 U11494 ( .A1(n10448), .A2(n10447), .ZN(n10620) );
  NAND4_X2 U11495 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n20424) );
  AND4_X1 U11496 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  AND4_X1 U11497 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10569) );
  AND4_X1 U11498 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11511) );
  AND4_X1 U11499 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10566) );
  AND4_X1 U11500 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10481) );
  AND4_X1 U11501 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10535) );
  AND4_X1 U11502 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10502) );
  AND4_X1 U11503 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10503) );
  AND4_X1 U11504 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10504) );
  AND4_X1 U11505 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10547) );
  AND4_X1 U11506 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10480) );
  AND4_X1 U11508 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  AND2_X1 U11509 ( .A1(n11600), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U11510 ( .A1(n12347), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12346) );
  CLKBUF_X3 U11511 ( .A(n11327), .Z(n11404) );
  INV_X4 U11512 ( .A(n17230), .ZN(n15875) );
  AND2_X2 U11513 ( .A1(n11744), .A2(n15689), .ZN(n12783) );
  INV_X2 U11514 ( .A(n20304), .ZN(n20332) );
  NAND2_X2 U11515 ( .A1(n20092), .A2(n20045), .ZN(n20094) );
  NAND2_X2 U11516 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20092), .ZN(n20091) );
  OR2_X1 U11517 ( .A1(n19096), .A2(n13965), .ZN(n10416) );
  INV_X2 U11518 ( .A(n16808), .ZN(U215) );
  BUF_X4 U11519 ( .A(n10491), .Z(n11406) );
  NOR2_X1 U11520 ( .A1(n12343), .A2(n16564), .ZN(n12347) );
  NAND2_X2 U11521 ( .A1(n19083), .A2(n19016), .ZN(n19073) );
  NAND2_X1 U11522 ( .A1(n10014), .A2(n10013), .ZN(n17450) );
  CLKBUF_X1 U11523 ( .A(n11744), .Z(n9774) );
  NAND2_X1 U11526 ( .A1(n9976), .A2(n10436), .ZN(n11470) );
  INV_X2 U11528 ( .A(n11446), .ZN(n9818) );
  NAND2_X2 U11529 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13954), .ZN(
        n17427) );
  INV_X2 U11530 ( .A(n16812), .ZN(n16814) );
  INV_X1 U11531 ( .A(n11444), .ZN(n9820) );
  NAND2_X1 U11532 ( .A1(n19096), .A2(n13964), .ZN(n17230) );
  INV_X1 U11533 ( .A(n11371), .ZN(n9799) );
  INV_X1 U11534 ( .A(n11369), .ZN(n9808) );
  OR2_X1 U11535 ( .A1(n13955), .A2(n13959), .ZN(n9878) );
  AND2_X1 U11536 ( .A1(n13563), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9794) );
  INV_X1 U11537 ( .A(n11444), .ZN(n9819) );
  INV_X1 U11538 ( .A(n11601), .ZN(n11745) );
  INV_X1 U11539 ( .A(n11200), .ZN(n9764) );
  NAND4_X2 U11540 ( .A1(n19096), .A2(n19114), .A3(n19108), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17473) );
  NAND2_X1 U11541 ( .A1(n19121), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13958) );
  AND2_X2 U11542 ( .A1(n12766), .A2(n11753), .ZN(n11767) );
  NAND2_X1 U11543 ( .A1(n9976), .A2(n10442), .ZN(n11444) );
  AND2_X1 U11544 ( .A1(n10015), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U11545 ( .A1(n11754), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12799) );
  AND2_X1 U11546 ( .A1(n10438), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13563) );
  AND2_X1 U11547 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10442) );
  NOR2_X1 U11548 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10424) );
  NOR2_X2 U11549 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10439) );
  INV_X1 U11550 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19114) );
  AND2_X1 U11551 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18942) );
  AND2_X2 U11552 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10438) );
  OR2_X2 U11553 ( .A1(n10456), .A2(n10455), .ZN(n9766) );
  NAND2_X1 U11554 ( .A1(n10122), .A2(n9979), .ZN(n13699) );
  NOR2_X4 U11555 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  NAND4_X1 U11556 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n9767) );
  OR2_X2 U11557 ( .A1(n15037), .A2(n15028), .ZN(n9872) );
  NOR2_X2 U11558 ( .A1(n13671), .A2(n13672), .ZN(n13670) );
  CLKBUF_X1 U11559 ( .A(n13638), .Z(n9768) );
  NAND2_X1 U11560 ( .A1(n10729), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9769) );
  CLKBUF_X1 U11561 ( .A(n10144), .Z(n9770) );
  NAND2_X2 U11562 ( .A1(n10683), .A2(n10631), .ZN(n10729) );
  AND2_X2 U11563 ( .A1(n12142), .A2(n13861), .ZN(n11523) );
  NAND2_X1 U11564 ( .A1(n16255), .A2(n10145), .ZN(n10144) );
  BUF_X1 U11565 ( .A(n11970), .Z(n9771) );
  MUX2_X2 U11566 ( .A(n11573), .B(n11572), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n9773) );
  XNOR2_X1 U11567 ( .A(n11638), .B(n13263), .ZN(n12583) );
  CLKBUF_X1 U11568 ( .A(n16255), .Z(n9775) );
  INV_X1 U11569 ( .A(n10724), .ZN(n9776) );
  NAND2_X1 U11570 ( .A1(n9777), .A2(n10725), .ZN(n10797) );
  NOR2_X1 U11571 ( .A1(n10759), .A2(n9776), .ZN(n9777) );
  CLKBUF_X1 U11572 ( .A(n13376), .Z(n9778) );
  INV_X1 U11573 ( .A(n10625), .ZN(n9779) );
  NAND2_X1 U11574 ( .A1(n16257), .A2(n16256), .ZN(n16255) );
  NAND2_X1 U11575 ( .A1(n13620), .A2(n9780), .ZN(n13751) );
  AND2_X1 U11576 ( .A1(n13619), .A2(n10961), .ZN(n9780) );
  NAND2_X1 U11577 ( .A1(n14412), .A2(n10359), .ZN(n9781) );
  OR2_X1 U11578 ( .A1(n10353), .A2(n14396), .ZN(n9782) );
  XNOR2_X1 U11579 ( .A(n10921), .B(n10922), .ZN(n13604) );
  NAND2_X1 U11582 ( .A1(n10110), .A2(n11689), .ZN(n11694) );
  NAND2_X2 U11583 ( .A1(n15671), .A2(n13861), .ZN(n12774) );
  INV_X2 U11584 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13861) );
  AND2_X1 U11585 ( .A1(n12576), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20152) );
  BUF_X2 U11586 ( .A(n11746), .Z(n9823) );
  INV_X1 U11588 ( .A(n9798), .ZN(n9787) );
  INV_X4 U11589 ( .A(n13788), .ZN(n19312) );
  NAND2_X1 U11590 ( .A1(n9988), .A2(n12038), .ZN(n15312) );
  OR2_X1 U11591 ( .A1(n9772), .A2(n15119), .ZN(n12306) );
  NOR2_X1 U11592 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  NAND2_X2 U11593 ( .A1(n13676), .A2(n9861), .ZN(n13521) );
  NAND2_X2 U11594 ( .A1(n13349), .A2(n12685), .ZN(n13676) );
  AND2_X4 U11595 ( .A1(n10440), .A2(n10442), .ZN(n10491) );
  NAND2_X2 U11596 ( .A1(n12765), .A2(n12764), .ZN(n12797) );
  NAND4_X2 U11597 ( .A1(n10552), .A2(n20412), .A3(n20424), .A4(n9765), .ZN(
        n10622) );
  NAND2_X1 U11598 ( .A1(n9748), .A2(n10728), .ZN(n9963) );
  INV_X2 U11599 ( .A(n9822), .ZN(n9833) );
  NAND2_X2 U11600 ( .A1(n10144), .A2(n10143), .ZN(n14674) );
  NAND2_X1 U11601 ( .A1(n11612), .A2(n12576), .ZN(n11862) );
  XNOR2_X2 U11602 ( .A(n10770), .B(n13541), .ZN(n13532) );
  XNOR2_X2 U11603 ( .A(n9960), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14711) );
  NAND2_X2 U11604 ( .A1(n12304), .A2(n12017), .ZN(n12276) );
  NAND2_X2 U11605 ( .A1(n20495), .A2(n10686), .ZN(n20861) );
  AND2_X1 U11606 ( .A1(n10441), .A2(n10438), .ZN(n9790) );
  AND2_X1 U11607 ( .A1(n10441), .A2(n10438), .ZN(n9791) );
  NAND2_X1 U11608 ( .A1(n11676), .A2(n11675), .ZN(n10330) );
  NAND2_X1 U11609 ( .A1(n10108), .A2(n10106), .ZN(n11664) );
  INV_X2 U11610 ( .A(n10695), .ZN(n9792) );
  INV_X1 U11612 ( .A(n10695), .ZN(n11448) );
  INV_X1 U11613 ( .A(n10695), .ZN(n10461) );
  AND2_X2 U11614 ( .A1(n10441), .A2(n10440), .ZN(n10466) );
  NAND2_X1 U11615 ( .A1(n11688), .A2(n11690), .ZN(n11695) );
  CLKBUF_X1 U11616 ( .A(n11023), .Z(n9795) );
  INV_X1 U11618 ( .A(n11369), .ZN(n9798) );
  INV_X1 U11619 ( .A(n9818), .ZN(n9800) );
  INV_X1 U11620 ( .A(n11446), .ZN(n11266) );
  INV_X1 U11621 ( .A(n11446), .ZN(n9817) );
  INV_X1 U11622 ( .A(n12244), .ZN(n9801) );
  INV_X2 U11623 ( .A(n12244), .ZN(n11671) );
  INV_X2 U11624 ( .A(n13263), .ZN(n11548) );
  AND2_X1 U11625 ( .A1(n13263), .A2(n13287), .ZN(n12955) );
  INV_X1 U11626 ( .A(n11297), .ZN(n9802) );
  INV_X1 U11628 ( .A(n11297), .ZN(n11454) );
  AND2_X1 U11631 ( .A1(n10441), .A2(n10438), .ZN(n10661) );
  OAI21_X1 U11632 ( .B1(n13603), .B2(n11095), .A(n10938), .ZN(n10939) );
  INV_X1 U11633 ( .A(n11470), .ZN(n11405) );
  NAND2_X2 U11634 ( .A1(n11637), .A2(n11862), .ZN(n12602) );
  AOI21_X1 U11635 ( .B1(n10729), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10730), .ZN(n10735) );
  AND2_X2 U11637 ( .A1(n9989), .A2(n10124), .ZN(n9846) );
  NAND2_X1 U11638 ( .A1(n15183), .A2(n10336), .ZN(n10132) );
  INV_X1 U11639 ( .A(n13887), .ZN(n11979) );
  INV_X2 U11640 ( .A(n16213), .ZN(n9973) );
  NAND2_X2 U11641 ( .A1(n10380), .A2(n10381), .ZN(n16213) );
  INV_X1 U11642 ( .A(n10656), .ZN(n9814) );
  INV_X1 U11643 ( .A(n19570), .ZN(n11980) );
  OAI21_X2 U11644 ( .B1(n12276), .B2(n15120), .A(n19307), .ZN(n12020) );
  AND2_X1 U11645 ( .A1(n10439), .A2(n9976), .ZN(n9815) );
  AND2_X1 U11646 ( .A1(n10439), .A2(n9976), .ZN(n10425) );
  AOI22_X2 U11647 ( .A1(n15194), .A2(n15195), .B1(n12997), .B2(n12118), .ZN(
        n15183) );
  NOR2_X4 U11648 ( .A1(n13219), .A2(n10624), .ZN(n13051) );
  NAND3_X2 U11649 ( .A1(n10066), .A2(n9897), .A3(n10065), .ZN(n13219) );
  OR2_X1 U11650 ( .A1(n10717), .A2(n10723), .ZN(n10724) );
  NOR2_X2 U11651 ( .A1(n13935), .A2(n10362), .ZN(n14431) );
  XNOR2_X2 U11652 ( .A(n10801), .B(n13725), .ZN(n13632) );
  AOI21_X2 U11653 ( .B1(n14221), .B2(n14220), .A(n14205), .ZN(n14574) );
  AND2_X2 U11654 ( .A1(n14231), .A2(n10351), .ZN(n14205) );
  XNOR2_X2 U11655 ( .A(n13356), .B(n10709), .ZN(n13509) );
  AND3_X1 U11656 ( .A1(n20412), .A2(n9755), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10880) );
  INV_X2 U11657 ( .A(n11444), .ZN(n11200) );
  AND2_X4 U11658 ( .A1(n10437), .A2(n10439), .ZN(n11327) );
  NAND2_X2 U11659 ( .A1(n12600), .A2(n12611), .ZN(n15669) );
  NOR2_X4 U11660 ( .A1(n11633), .A2(n11632), .ZN(n12600) );
  INV_X1 U11661 ( .A(n11601), .ZN(n9821) );
  INV_X1 U11662 ( .A(n11746), .ZN(n9822) );
  INV_X1 U11663 ( .A(n9823), .ZN(n9824) );
  INV_X1 U11664 ( .A(n9823), .ZN(n9825) );
  INV_X1 U11665 ( .A(n9823), .ZN(n9826) );
  INV_X2 U11666 ( .A(n11523), .ZN(n9827) );
  INV_X1 U11667 ( .A(n9827), .ZN(n9828) );
  INV_X1 U11668 ( .A(n9827), .ZN(n9829) );
  INV_X1 U11669 ( .A(n9827), .ZN(n9830) );
  INV_X1 U11670 ( .A(n9833), .ZN(n9831) );
  INV_X1 U11671 ( .A(n9827), .ZN(n9832) );
  INV_X1 U11672 ( .A(n9833), .ZN(n9834) );
  INV_X1 U11673 ( .A(n9833), .ZN(n9835) );
  INV_X1 U11674 ( .A(n9833), .ZN(n9836) );
  BUF_X2 U11675 ( .A(n12654), .Z(n9837) );
  INV_X1 U11676 ( .A(n10544), .ZN(n10496) );
  NAND2_X1 U11677 ( .A1(n10796), .A2(n10022), .ZN(n10845) );
  AND2_X1 U11678 ( .A1(n10795), .A2(n10820), .ZN(n10022) );
  NAND2_X1 U11679 ( .A1(n10257), .A2(n10256), .ZN(n11673) );
  INV_X1 U11680 ( .A(n11672), .ZN(n10256) );
  AOI211_X1 U11681 ( .C1(n12883), .C2(n12881), .A(n12880), .B(n14957), .ZN(
        n12882) );
  NAND2_X1 U11682 ( .A1(n17782), .A2(n18920), .ZN(n16719) );
  INV_X1 U11683 ( .A(n10762), .ZN(n10713) );
  OAI21_X2 U11684 ( .B1(n14186), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10703), 
        .ZN(n10717) );
  OR2_X1 U11685 ( .A1(n10893), .A2(n10713), .ZN(n10703) );
  NAND2_X1 U11686 ( .A1(n11636), .A2(n11651), .ZN(n10051) );
  NAND2_X1 U11687 ( .A1(n12627), .A2(n9931), .ZN(n10109) );
  OR2_X1 U11688 ( .A1(n10622), .A2(n21027), .ZN(n11488) );
  OR2_X1 U11689 ( .A1(n13935), .A2(n10368), .ZN(n14322) );
  AOI21_X1 U11690 ( .B1(n9753), .B2(n10073), .A(n21316), .ZN(n10072) );
  INV_X1 U11691 ( .A(n14697), .ZN(n10073) );
  NAND2_X1 U11692 ( .A1(n13129), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10631) );
  INV_X1 U11693 ( .A(n10794), .ZN(n10076) );
  INV_X1 U11694 ( .A(n15052), .ZN(n10281) );
  NAND2_X1 U11695 ( .A1(n12861), .A2(n10394), .ZN(n10393) );
  INV_X1 U11696 ( .A(n12863), .ZN(n10394) );
  AND3_X1 U11697 ( .A1(n12432), .A2(n12431), .A3(n12430), .ZN(n13779) );
  AOI21_X1 U11698 ( .B1(n13199), .B2(n9908), .A(n10292), .ZN(n10291) );
  INV_X1 U11699 ( .A(n13197), .ZN(n10292) );
  NAND2_X1 U11700 ( .A1(n20155), .A2(n12660), .ZN(n12880) );
  AND3_X1 U11701 ( .A1(n11623), .A2(n9773), .A3(n19467), .ZN(n10216) );
  NAND2_X1 U11702 ( .A1(n11533), .A2(n15689), .ZN(n10025) );
  NAND2_X1 U11703 ( .A1(n11538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10024) );
  INV_X1 U11704 ( .A(n13684), .ZN(n10227) );
  INV_X1 U11705 ( .A(n15622), .ZN(n10037) );
  INV_X1 U11706 ( .A(n10125), .ZN(n10124) );
  OAI21_X1 U11707 ( .B1(n9883), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12057), .ZN(n10125) );
  INV_X1 U11708 ( .A(n11673), .ZN(n11676) );
  INV_X1 U11709 ( .A(n14883), .ZN(n12534) );
  NAND2_X1 U11710 ( .A1(n12655), .A2(n20110), .ZN(n12676) );
  NOR2_X1 U11711 ( .A1(n11723), .A2(n10117), .ZN(n11716) );
  AOI211_X1 U11712 ( .C1(n17468), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n14012), .B(n14011), .ZN(n14013) );
  INV_X1 U11713 ( .A(n17190), .ZN(n13959) );
  NOR2_X1 U11714 ( .A1(n15819), .A2(n14058), .ZN(n16077) );
  NOR3_X1 U11715 ( .A1(n15794), .A2(n17625), .A3(n15812), .ZN(n14058) );
  NAND2_X1 U11716 ( .A1(n19096), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13962) );
  INV_X1 U11717 ( .A(n17467), .ZN(n15914) );
  NAND2_X1 U11718 ( .A1(n16007), .A2(n9956), .ZN(n10312) );
  NOR2_X1 U11719 ( .A1(n16821), .A2(n15944), .ZN(n15795) );
  NOR2_X1 U11720 ( .A1(n15817), .A2(n10171), .ZN(n15948) );
  NAND2_X1 U11721 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  NAND2_X1 U11722 ( .A1(n15804), .A2(n15803), .ZN(n10172) );
  INV_X1 U11723 ( .A(n15816), .ZN(n10173) );
  NAND2_X1 U11724 ( .A1(n17625), .A2(n15803), .ZN(n15947) );
  NAND2_X1 U11725 ( .A1(n18112), .A2(n15930), .ZN(n15931) );
  AND2_X1 U11726 ( .A1(n16053), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U11727 ( .A1(n14245), .A2(n14233), .ZN(n14235) );
  NAND2_X1 U11728 ( .A1(n10147), .A2(n9896), .ZN(n10913) );
  AND2_X1 U11729 ( .A1(n14114), .A2(n14795), .ZN(n10148) );
  NAND2_X1 U11730 ( .A1(n10382), .A2(n14640), .ZN(n10381) );
  INV_X1 U11731 ( .A(n10383), .ZN(n10382) );
  AND4_X1 U11732 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  NAND2_X1 U11733 ( .A1(n11688), .A2(n11634), .ZN(n10110) );
  NAND2_X1 U11734 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10336) );
  INV_X1 U11735 ( .A(n15181), .ZN(n10337) );
  INV_X1 U11736 ( .A(n12362), .ZN(n11612) );
  NAND2_X1 U11737 ( .A1(n12596), .A2(n20165), .ZN(n12648) );
  AND2_X1 U11738 ( .A1(n19504), .A2(n20133), .ZN(n19661) );
  AOI21_X1 U11739 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(n15982) );
  OR2_X1 U11740 ( .A1(n16920), .A2(n9898), .ZN(n10156) );
  NOR2_X1 U11741 ( .A1(n13985), .A2(n10179), .ZN(n10178) );
  INV_X1 U11742 ( .A(n13984), .ZN(n10180) );
  AND2_X1 U11743 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10179) );
  NOR2_X1 U11744 ( .A1(n15795), .A2(n10003), .ZN(n15949) );
  OR2_X1 U11745 ( .A1(n15796), .A2(n15950), .ZN(n10003) );
  AOI21_X1 U11746 ( .B1(n10092), .B2(n10089), .A(n10083), .ZN(n10082) );
  NAND2_X1 U11747 ( .A1(n10085), .A2(n18090), .ZN(n10084) );
  NOR2_X1 U11748 ( .A1(n15943), .A2(n15942), .ZN(n18920) );
  NAND2_X1 U11749 ( .A1(n13061), .A2(n13337), .ZN(n21117) );
  INV_X1 U11750 ( .A(n10822), .ZN(n10820) );
  INV_X1 U11751 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U11752 ( .A1(n11872), .A2(n11871), .ZN(n11899) );
  OAI21_X1 U11753 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19108), .A(
        n14047), .ZN(n14048) );
  AND2_X1 U11754 ( .A1(n10818), .A2(n10817), .ZN(n10848) );
  OR2_X1 U11755 ( .A1(n10655), .A2(n10654), .ZN(n10896) );
  INV_X1 U11756 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10433) );
  INV_X1 U11757 ( .A(n10880), .ZN(n10754) );
  INV_X1 U11758 ( .A(n12798), .ZN(n10113) );
  INV_X1 U11759 ( .A(n10398), .ZN(n10397) );
  AND2_X1 U11760 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11543) );
  INV_X1 U11761 ( .A(n11626), .ZN(n10050) );
  NAND2_X1 U11762 ( .A1(n9977), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10108) );
  NAND2_X1 U11763 ( .A1(n12389), .A2(n12609), .ZN(n11630) );
  AOI21_X1 U11764 ( .B1(n9828), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10419), .ZN(n11584) );
  NAND2_X1 U11765 ( .A1(n10004), .A2(n15813), .ZN(n15790) );
  NOR2_X1 U11766 ( .A1(n18934), .A2(n14045), .ZN(n10004) );
  NOR2_X1 U11767 ( .A1(n15932), .A2(n17648), .ZN(n15911) );
  NOR2_X1 U11768 ( .A1(n18134), .A2(n17660), .ZN(n15961) );
  NAND2_X1 U11769 ( .A1(n10622), .A2(n20408), .ZN(n10066) );
  NOR2_X1 U11770 ( .A1(n14221), .A2(n10352), .ZN(n10351) );
  INV_X1 U11771 ( .A(n14232), .ZN(n10352) );
  NOR2_X1 U11772 ( .A1(n14284), .A2(n10357), .ZN(n10356) );
  INV_X1 U11773 ( .A(n14294), .ZN(n10357) );
  OR2_X1 U11774 ( .A1(n11096), .A2(n10365), .ZN(n10364) );
  AND2_X1 U11775 ( .A1(n10368), .A2(n10366), .ZN(n10365) );
  OR2_X1 U11776 ( .A1(n14337), .A2(n10367), .ZN(n10366) );
  AND2_X1 U11777 ( .A1(n21030), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11494) );
  NOR2_X1 U11778 ( .A1(n10021), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10019) );
  OR2_X1 U11779 ( .A1(n10072), .A2(n10070), .ZN(n10069) );
  OR2_X1 U11780 ( .A1(n16213), .A2(n10070), .ZN(n10067) );
  NAND2_X1 U11782 ( .A1(n14097), .A2(n10205), .ZN(n10204) );
  NOR2_X1 U11783 ( .A1(n9950), .A2(n14339), .ZN(n10205) );
  NAND2_X1 U11784 ( .A1(n10704), .A2(n20398), .ZN(n10708) );
  NOR2_X1 U11785 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NAND2_X1 U11786 ( .A1(n10576), .A2(n10575), .ZN(n10608) );
  OR2_X1 U11787 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20376), .ZN(
        n10607) );
  NOR2_X1 U11788 ( .A1(n15278), .A2(n10300), .ZN(n10299) );
  INV_X1 U11789 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U11790 ( .A1(n11873), .A2(n11874), .ZN(n11907) );
  NAND2_X1 U11791 ( .A1(n10404), .A2(n9918), .ZN(n10400) );
  NOR2_X1 U11792 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12766) );
  INV_X1 U11793 ( .A(n14906), .ZN(n10280) );
  AND2_X1 U11794 ( .A1(n10116), .A2(n15004), .ZN(n10115) );
  NOR2_X1 U11795 ( .A1(n15175), .A2(n10296), .ZN(n10295) );
  INV_X1 U11796 ( .A(n15011), .ZN(n10279) );
  NAND2_X1 U11797 ( .A1(n12999), .A2(n14988), .ZN(n10223) );
  NOR2_X1 U11798 ( .A1(n15266), .A2(n10217), .ZN(n12985) );
  OR3_X1 U11799 ( .A1(n14933), .A2(n10218), .A3(n14917), .ZN(n10217) );
  NAND2_X1 U11800 ( .A1(n10219), .A2(n14997), .ZN(n10218) );
  INV_X1 U11801 ( .A(n15006), .ZN(n10219) );
  INV_X1 U11802 ( .A(n14869), .ZN(n12559) );
  NAND2_X1 U11803 ( .A1(n15206), .A2(n15535), .ZN(n10056) );
  NOR2_X1 U11804 ( .A1(n15568), .A2(n10286), .ZN(n10285) );
  INV_X1 U11805 ( .A(n13588), .ZN(n10286) );
  INV_X1 U11806 ( .A(n15569), .ZN(n10284) );
  NAND2_X1 U11807 ( .A1(n15312), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12044) );
  INV_X1 U11808 ( .A(n13779), .ZN(n10288) );
  XNOR2_X1 U11809 ( .A(n11964), .B(n9771), .ZN(n12277) );
  INV_X1 U11810 ( .A(n12277), .ZN(n12296) );
  INV_X1 U11811 ( .A(n9771), .ZN(n11965) );
  NAND2_X1 U11812 ( .A1(n10044), .A2(n10043), .ZN(n11831) );
  INV_X1 U11813 ( .A(n9754), .ZN(n12482) );
  AND2_X1 U11814 ( .A1(n21322), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12673) );
  AND2_X1 U11815 ( .A1(n11623), .A2(n19467), .ZN(n12611) );
  INV_X1 U11816 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21259) );
  NAND2_X1 U11817 ( .A1(n19141), .A2(n17666), .ZN(n15792) );
  NAND2_X1 U11818 ( .A1(n17775), .A2(n9864), .ZN(n16681) );
  NAND2_X1 U11819 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13955) );
  NOR2_X1 U11820 ( .A1(n18247), .A2(n16000), .ZN(n17867) );
  OAI21_X1 U11821 ( .B1(n18055), .B2(n18054), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15977) );
  OR2_X1 U11822 ( .A1(n18079), .A2(n10090), .ZN(n10087) );
  NAND2_X1 U11823 ( .A1(n15911), .A2(n15951), .ZN(n15910) );
  XNOR2_X1 U11824 ( .A(n15961), .B(n10011), .ZN(n15962) );
  INV_X1 U11825 ( .A(n17652), .ZN(n10011) );
  XNOR2_X1 U11826 ( .A(n17652), .B(n15965), .ZN(n15929) );
  NAND2_X1 U11827 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15922) );
  INV_X1 U11828 ( .A(n15920), .ZN(n15924) );
  INV_X1 U11829 ( .A(n15805), .ZN(n10170) );
  NOR2_X1 U11830 ( .A1(n10190), .A2(n10185), .ZN(n10184) );
  INV_X1 U11831 ( .A(n14040), .ZN(n10190) );
  INV_X1 U11832 ( .A(n14043), .ZN(n10191) );
  AND2_X1 U11833 ( .A1(n13245), .A2(n13244), .ZN(n13402) );
  INV_X1 U11834 ( .A(n13229), .ZN(n10371) );
  INV_X1 U11835 ( .A(n20398), .ZN(n13338) );
  AND2_X1 U11836 ( .A1(n10350), .A2(n11495), .ZN(n10349) );
  AND2_X1 U11837 ( .A1(n10351), .A2(n14206), .ZN(n10350) );
  AND2_X1 U11838 ( .A1(n11439), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11440) );
  NAND2_X1 U11839 ( .A1(n11440), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11499) );
  AND2_X1 U11840 ( .A1(n14293), .A2(n10354), .ZN(n14257) );
  NAND2_X1 U11841 ( .A1(n11314), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11339) );
  NAND2_X1 U11842 ( .A1(n14293), .A2(n14294), .ZN(n14283) );
  AND2_X1 U11843 ( .A1(n11232), .A2(n11231), .ZN(n14401) );
  AND2_X1 U11844 ( .A1(n14445), .A2(n14446), .ZN(n14447) );
  INV_X1 U11845 ( .A(n13936), .ZN(n11019) );
  INV_X1 U11846 ( .A(n10952), .ZN(n10960) );
  NAND2_X1 U11847 ( .A1(n13591), .A2(n10942), .ZN(n13620) );
  INV_X2 U11848 ( .A(n14149), .ZN(n14208) );
  AND2_X1 U11849 ( .A1(n14261), .A2(n14243), .ZN(n14245) );
  NOR2_X2 U11850 ( .A1(n14399), .A2(n10210), .ZN(n14261) );
  NAND2_X1 U11851 ( .A1(n10212), .A2(n10211), .ZN(n10210) );
  INV_X1 U11852 ( .A(n10213), .ZN(n10212) );
  NOR2_X1 U11853 ( .A1(n10214), .A2(n14259), .ZN(n10211) );
  INV_X1 U11854 ( .A(n14820), .ZN(n10385) );
  NOR2_X1 U11855 ( .A1(n9753), .A2(n10905), .ZN(n10384) );
  AND2_X1 U11856 ( .A1(n10904), .A2(n10387), .ZN(n10386) );
  NAND2_X1 U11857 ( .A1(n16212), .A2(n14092), .ZN(n14666) );
  NOR2_X1 U11858 ( .A1(n10389), .A2(n10146), .ZN(n10145) );
  INV_X1 U11859 ( .A(n10892), .ZN(n10146) );
  INV_X1 U11860 ( .A(n9927), .ZN(n10389) );
  OR2_X1 U11861 ( .A1(n13363), .A2(n13362), .ZN(n13372) );
  NAND2_X1 U11862 ( .A1(n10778), .A2(n10777), .ZN(n20535) );
  NAND2_X1 U11863 ( .A1(n21027), .A2(n20383), .ZN(n20544) );
  AND2_X1 U11864 ( .A1(n20889), .A2(n20427), .ZN(n20755) );
  NOR2_X1 U11865 ( .A1(n20748), .A2(n20544), .ZN(n20900) );
  INV_X1 U11866 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20957) );
  INV_X1 U11867 ( .A(n20544), .ZN(n20427) );
  AND2_X1 U11868 ( .A1(n21324), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16053) );
  NOR2_X1 U11869 ( .A1(n19374), .A2(n19373), .ZN(n12687) );
  AND2_X1 U11870 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10114) );
  NAND2_X1 U11871 ( .A1(n10390), .A2(n12882), .ZN(n14956) );
  NAND2_X1 U11872 ( .A1(n10289), .A2(n10291), .ZN(n13778) );
  NAND2_X1 U11873 ( .A1(n9997), .A2(n15689), .ZN(n9996) );
  NAND2_X1 U11874 ( .A1(n9995), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9994) );
  NAND2_X1 U11875 ( .A1(n9991), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9990) );
  NAND2_X1 U11876 ( .A1(n9993), .A2(n15689), .ZN(n9992) );
  NOR2_X2 U11877 ( .A1(n12325), .A2(n12163), .ZN(n12322) );
  AND2_X1 U11878 ( .A1(n15300), .A2(n9936), .ZN(n15264) );
  NAND2_X1 U11879 ( .A1(n12351), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12350) );
  NAND2_X1 U11880 ( .A1(n13395), .A2(n13396), .ZN(n13444) );
  CLKBUF_X1 U11881 ( .A(n12244), .Z(n14873) );
  NAND2_X1 U11882 ( .A1(n14975), .A2(n9942), .ZN(n14950) );
  INV_X1 U11883 ( .A(n14947), .ZN(n10228) );
  NAND2_X1 U11884 ( .A1(n14975), .A2(n10229), .ZN(n14948) );
  NAND2_X1 U11885 ( .A1(n14975), .A2(n14968), .ZN(n14967) );
  INV_X1 U11886 ( .A(n10335), .ZN(n10131) );
  NAND2_X1 U11887 ( .A1(n15181), .A2(n21149), .ZN(n10335) );
  AND2_X1 U11888 ( .A1(n14915), .A2(n10254), .ZN(n15170) );
  NOR2_X1 U11889 ( .A1(n15119), .A2(n15397), .ZN(n10254) );
  NOR2_X1 U11890 ( .A1(n15212), .A2(n15233), .ZN(n10049) );
  NAND2_X1 U11891 ( .A1(n15244), .A2(n15213), .ZN(n10048) );
  NOR3_X1 U11892 ( .A1(n15266), .A2(n14933), .A3(n15006), .ZN(n14998) );
  OR2_X1 U11893 ( .A1(n9888), .A2(n10059), .ZN(n10058) );
  INV_X1 U11894 ( .A(n15283), .ZN(n10059) );
  AND3_X1 U11895 ( .A1(n12377), .A2(n12376), .A3(n12375), .ZN(n13841) );
  NAND2_X1 U11896 ( .A1(n10284), .A2(n10285), .ZN(n13842) );
  INV_X1 U11897 ( .A(n15617), .ZN(n10340) );
  INV_X1 U11898 ( .A(n10264), .ZN(n10263) );
  INV_X1 U11899 ( .A(n10265), .ZN(n10262) );
  NAND2_X1 U11900 ( .A1(n15318), .A2(n16569), .ZN(n10265) );
  NAND2_X1 U11901 ( .A1(n15643), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15642) );
  AND2_X1 U11902 ( .A1(n12417), .A2(n12416), .ZN(n13199) );
  NAND2_X1 U11903 ( .A1(n13699), .A2(n13698), .ZN(n10045) );
  AND2_X1 U11904 ( .A1(n10231), .A2(n12166), .ZN(n13701) );
  NAND2_X1 U11905 ( .A1(n12164), .A2(n12165), .ZN(n10231) );
  AND2_X1 U11906 ( .A1(n11677), .A2(n10330), .ZN(n11692) );
  NAND2_X1 U11907 ( .A1(n11615), .A2(n11614), .ZN(n11661) );
  NAND2_X1 U11908 ( .A1(n20106), .A2(n19501), .ZN(n19883) );
  INV_X1 U11909 ( .A(n19952), .ZN(n19917) );
  OAI21_X1 U11910 ( .B1(n15810), .B2(n15809), .A(n15808), .ZN(n18921) );
  AND2_X1 U11911 ( .A1(n10153), .A2(n17130), .ZN(n10150) );
  NAND2_X1 U11912 ( .A1(n10182), .A2(n10181), .ZN(n14072) );
  NOR2_X1 U11913 ( .A1(n15792), .A2(n18985), .ZN(n10181) );
  INV_X1 U11914 ( .A(n16077), .ZN(n10182) );
  INV_X1 U11915 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17477) );
  OAI22_X1 U11916 ( .A1(n16079), .A2(n16078), .B1(n16077), .B2(n16076), .ZN(
        n16080) );
  INV_X1 U11917 ( .A(n17634), .ZN(n10176) );
  INV_X1 U11918 ( .A(n17633), .ZN(n10175) );
  NAND3_X2 U11919 ( .A1(n17190), .A2(n19096), .A3(n19108), .ZN(n17483) );
  NOR3_X1 U11920 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n19121), .ZN(n13954) );
  NAND2_X1 U11921 ( .A1(n10096), .A2(n9894), .ZN(n10095) );
  NAND2_X1 U11922 ( .A1(n15914), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10096) );
  NOR2_X1 U11923 ( .A1(n9875), .A2(n10098), .ZN(n10097) );
  INV_X1 U11924 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10098) );
  AOI21_X1 U11925 ( .B1(n17436), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n15883), .ZN(n15886) );
  INV_X1 U11926 ( .A(n16681), .ZN(n16671) );
  AND2_X1 U11927 ( .A1(n17887), .A2(n9938), .ZN(n17811) );
  INV_X1 U11928 ( .A(n16658), .ZN(n17856) );
  INV_X1 U11929 ( .A(n10326), .ZN(n10321) );
  INV_X1 U11930 ( .A(n17779), .ZN(n18150) );
  NAND2_X1 U11931 ( .A1(n10325), .A2(n10322), .ZN(n17817) );
  NOR2_X1 U11932 ( .A1(n10324), .A2(n10323), .ZN(n10322) );
  NAND2_X1 U11933 ( .A1(n10002), .A2(n15948), .ZN(n18932) );
  NAND2_X1 U11934 ( .A1(n15949), .A2(n9919), .ZN(n10002) );
  OR2_X1 U11935 ( .A1(n9788), .A2(n10317), .ZN(n10316) );
  INV_X1 U11936 ( .A(n18014), .ZN(n10317) );
  NOR2_X1 U11937 ( .A1(n16004), .A2(n18330), .ZN(n18023) );
  NAND2_X1 U11938 ( .A1(n18104), .A2(n15933), .ZN(n18091) );
  XNOR2_X1 U11939 ( .A(n15929), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18114) );
  XNOR2_X1 U11940 ( .A(n17660), .B(n10078), .ZN(n18125) );
  NAND2_X1 U11941 ( .A1(n18133), .A2(n18125), .ZN(n18124) );
  INV_X1 U11942 ( .A(n18942), .ZN(n18939) );
  AND2_X1 U11943 ( .A1(n14214), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14215) );
  INV_X1 U11944 ( .A(n20276), .ZN(n20261) );
  INV_X1 U11945 ( .A(n14151), .ZN(n10200) );
  NAND2_X1 U11946 ( .A1(n10142), .A2(n10737), .ZN(n20831) );
  INV_X1 U11947 ( .A(n21101), .ZN(n14862) );
  OR2_X1 U11948 ( .A1(n12027), .A2(n10249), .ZN(n12039) );
  NOR2_X1 U11949 ( .A1(n12468), .A2(n12467), .ZN(n13662) );
  NAND2_X1 U11950 ( .A1(n12942), .A2(n20165), .ZN(n19419) );
  INV_X1 U11951 ( .A(n15141), .ZN(n10221) );
  NAND2_X1 U11952 ( .A1(n16517), .A2(n16549), .ZN(n10032) );
  NAND2_X1 U11953 ( .A1(n16516), .A2(n16561), .ZN(n10031) );
  INV_X1 U11954 ( .A(n16555), .ZN(n16554) );
  NAND2_X1 U11955 ( .A1(n13038), .A2(n12160), .ZN(n16565) );
  AND2_X1 U11956 ( .A1(n16565), .A2(n14079), .ZN(n16555) );
  INV_X1 U11957 ( .A(n16565), .ZN(n16546) );
  INV_X1 U11958 ( .A(n16558), .ZN(n16550) );
  INV_X1 U11959 ( .A(n15342), .ZN(n15350) );
  XNOR2_X1 U11960 ( .A(n15137), .B(n15136), .ZN(n15354) );
  OR2_X1 U11961 ( .A1(n12648), .A2(n12632), .ZN(n16581) );
  OR2_X1 U11962 ( .A1(n12648), .A2(n12628), .ZN(n15600) );
  AND2_X1 U11963 ( .A1(n12598), .A2(n12597), .ZN(n16592) );
  INV_X1 U11964 ( .A(n19501), .ZN(n20133) );
  XNOR2_X1 U11965 ( .A(n13283), .B(n13284), .ZN(n20127) );
  NAND2_X1 U11966 ( .A1(n13349), .A2(n13352), .ZN(n19504) );
  AND2_X1 U11967 ( .A1(n10159), .A2(n17130), .ZN(n16907) );
  INV_X1 U11968 ( .A(n17187), .ZN(n17171) );
  INV_X2 U11969 ( .A(n17625), .ZN(n18511) );
  INV_X1 U11970 ( .A(n17332), .ZN(n17317) );
  AND2_X1 U11971 ( .A1(n15695), .A2(n17411), .ZN(n17363) );
  NOR2_X1 U11972 ( .A1(n17432), .A2(n17464), .ZN(n17431) );
  NAND2_X1 U11973 ( .A1(n17486), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17464) );
  INV_X1 U11974 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17490) );
  NOR2_X2 U11975 ( .A1(n14072), .A2(n18511), .ZN(n17517) );
  NOR2_X1 U11976 ( .A1(n17625), .A2(n17559), .ZN(n17555) );
  NAND2_X1 U11977 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17606), .ZN(n17601) );
  NAND2_X1 U11978 ( .A1(n16692), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10138) );
  OR2_X1 U11979 ( .A1(n16690), .A2(n16689), .ZN(n10139) );
  NOR2_X1 U11980 ( .A1(n17846), .A2(n18195), .ZN(n10001) );
  AND2_X1 U11981 ( .A1(n17933), .A2(n9999), .ZN(n17844) );
  NOR2_X1 U11982 ( .A1(n17851), .A2(n18211), .ZN(n9999) );
  NAND2_X1 U11983 ( .A1(n17887), .A2(n9842), .ZN(n17835) );
  AND2_X1 U11984 ( .A1(n18045), .A2(n18047), .ZN(n17998) );
  NOR2_X1 U11985 ( .A1(n16822), .A2(n18484), .ZN(n18045) );
  INV_X1 U11986 ( .A(n18127), .ZN(n18140) );
  XNOR2_X1 U11987 ( .A(n16009), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16688) );
  OAI21_X1 U11988 ( .B1(n16719), .B2(n16004), .A(n9851), .ZN(n10080) );
  NOR2_X1 U11989 ( .A1(n18457), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10079) );
  OAI21_X1 U11990 ( .B1(n16719), .B2(n10320), .A(n10318), .ZN(n16717) );
  AND2_X1 U11991 ( .A1(n16715), .A2(n10319), .ZN(n10318) );
  OR2_X1 U11992 ( .A1(n16711), .A2(n18047), .ZN(n10320) );
  NAND2_X1 U11993 ( .A1(n18152), .A2(n21361), .ZN(n10006) );
  NAND2_X1 U11994 ( .A1(n10008), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10007) );
  OR2_X1 U11995 ( .A1(n18159), .A2(n10009), .ZN(n10008) );
  AND2_X1 U11996 ( .A1(n18458), .A2(n18151), .ZN(n10009) );
  NOR2_X1 U11997 ( .A1(n16708), .A2(n16709), .ZN(n17789) );
  OR3_X1 U11998 ( .A1(n17905), .A2(n16001), .A3(n18211), .ZN(n17841) );
  NOR2_X1 U11999 ( .A1(n18457), .A2(n15992), .ZN(n18454) );
  INV_X1 U12000 ( .A(n10823), .ZN(n10821) );
  INV_X1 U12001 ( .A(n10844), .ZN(n10843) );
  NOR2_X1 U12002 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10430), .ZN(
        n10436) );
  NAND2_X1 U12003 ( .A1(n10440), .A2(n10439), .ZN(n10695) );
  OR2_X1 U12004 ( .A1(n14337), .A2(n10369), .ZN(n10368) );
  INV_X1 U12005 ( .A(n14321), .ZN(n10369) );
  OR2_X1 U12006 ( .A1(n10842), .A2(n10841), .ZN(n10872) );
  INV_X1 U12007 ( .A(n10896), .ZN(n10719) );
  INV_X1 U12008 ( .A(n13653), .ZN(n10795) );
  AND3_X1 U12009 ( .A1(n10716), .A2(n10715), .A3(n10714), .ZN(n10722) );
  NAND2_X1 U12010 ( .A1(n10673), .A2(n10764), .ZN(n10017) );
  OAI211_X1 U12011 ( .C1(n10544), .C2(n10516), .A(n10515), .B(n10514), .ZN(
        n10517) );
  AND2_X1 U12012 ( .A1(n21258), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12135) );
  AOI21_X1 U12013 ( .B1(n9836), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A(n11518), .ZN(n11522) );
  AND2_X1 U12014 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11518) );
  OR2_X1 U12015 ( .A1(n12175), .A2(n11650), .ZN(n11656) );
  INV_X1 U12016 ( .A(n15310), .ZN(n10331) );
  AND2_X1 U12017 ( .A1(n9859), .A2(n12407), .ZN(n10338) );
  NAND2_X1 U12018 ( .A1(n11649), .A2(n10051), .ZN(n9977) );
  NOR2_X1 U12019 ( .A1(n11901), .A2(n11900), .ZN(n11902) );
  INV_X1 U12020 ( .A(n11899), .ZN(n11901) );
  INV_X1 U12021 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11715) );
  INV_X1 U12022 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11733) );
  INV_X1 U12023 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11724) );
  INV_X1 U12024 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11726) );
  NOR2_X1 U12025 ( .A1(n11638), .A2(n13263), .ZN(n11628) );
  NOR2_X1 U12026 ( .A1(n21214), .A2(n18128), .ZN(n10163) );
  AND2_X1 U12027 ( .A1(n15790), .A2(n15986), .ZN(n15804) );
  AND2_X1 U12028 ( .A1(n15944), .A2(n18488), .ZN(n15815) );
  INV_X1 U12029 ( .A(n15813), .ZN(n14044) );
  NOR2_X1 U12030 ( .A1(n9891), .A2(n14041), .ZN(n10189) );
  INV_X1 U12031 ( .A(n10187), .ZN(n10186) );
  OAI21_X1 U12032 ( .B1(n17381), .B2(n18814), .A(n10188), .ZN(n10187) );
  NAND2_X1 U12033 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10188) );
  NOR2_X1 U12034 ( .A1(n15804), .A2(n15947), .ZN(n15788) );
  NOR2_X1 U12035 ( .A1(n14270), .A2(n10355), .ZN(n10354) );
  INV_X1 U12036 ( .A(n10356), .ZN(n10355) );
  OR2_X1 U12037 ( .A1(n14295), .A2(n14271), .ZN(n10213) );
  INV_X1 U12038 ( .A(n14281), .ZN(n10214) );
  INV_X1 U12039 ( .A(n14414), .ZN(n10208) );
  NAND2_X1 U12040 ( .A1(n9753), .A2(n10911), .ZN(n10387) );
  OAI22_X1 U12041 ( .A1(n10952), .A2(n10374), .B1(n10825), .B2(n16044), .ZN(
        n10826) );
  NAND2_X1 U12042 ( .A1(n14143), .A2(n14208), .ZN(n14134) );
  NAND2_X1 U12043 ( .A1(n13532), .A2(n13531), .ZN(n10772) );
  NAND2_X1 U12044 ( .A1(n10671), .A2(n10670), .ZN(n10763) );
  AND4_X1 U12045 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10671) );
  AND4_X1 U12046 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10670) );
  NOR2_X1 U12047 ( .A1(n10375), .A2(n10374), .ZN(n10373) );
  INV_X1 U12048 ( .A(n10377), .ZN(n10375) );
  NOR2_X1 U12049 ( .A1(n10370), .A2(n13229), .ZN(n13224) );
  NOR2_X1 U12050 ( .A1(n10435), .A2(n10434), .ZN(n10448) );
  OAI21_X1 U12051 ( .B1(n21123), .B2(n16411), .A(n14862), .ZN(n20383) );
  NAND2_X1 U12052 ( .A1(n14152), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10755) );
  OR3_X1 U12053 ( .A1(n10602), .A2(n10601), .A3(n13053), .ZN(n10603) );
  OR2_X1 U12054 ( .A1(n16439), .A2(n12126), .ZN(n15115) );
  OR2_X1 U12055 ( .A1(n12065), .A2(n10242), .ZN(n10241) );
  NAND2_X1 U12056 ( .A1(n12061), .A2(n10243), .ZN(n10242) );
  NAND2_X1 U12057 ( .A1(n12106), .A2(n12107), .ZN(n12115) );
  NAND2_X1 U12058 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  INV_X1 U12059 ( .A(n10249), .ZN(n10248) );
  NAND2_X1 U12060 ( .A1(n10253), .A2(n12023), .ZN(n10252) );
  OR2_X1 U12061 ( .A1(n12027), .A2(n10252), .ZN(n12032) );
  INV_X1 U12062 ( .A(n11906), .ZN(n10233) );
  NAND2_X1 U12063 ( .A1(n11860), .A2(n13798), .ZN(n10237) );
  NAND2_X1 U12064 ( .A1(n12150), .A2(n13885), .ZN(n10236) );
  NAND2_X1 U12065 ( .A1(n9863), .A2(n14985), .ZN(n10402) );
  NAND2_X1 U12066 ( .A1(n15061), .A2(n15062), .ZN(n10112) );
  NAND2_X1 U12067 ( .A1(n12720), .A2(n9955), .ZN(n10398) );
  NOR2_X1 U12068 ( .A1(n9933), .A2(n19368), .ZN(n10116) );
  INV_X1 U12069 ( .A(n19353), .ZN(n10399) );
  AOI21_X1 U12070 ( .B1(n9831), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11543), .ZN(n11544) );
  AND2_X1 U12071 ( .A1(n9916), .A2(n10226), .ZN(n10225) );
  INV_X1 U12072 ( .A(n13844), .ZN(n10226) );
  NOR2_X1 U12073 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  OR2_X1 U12074 ( .A1(n10306), .A2(n16532), .ZN(n10305) );
  NAND2_X1 U12075 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12076 ( .A1(n12175), .A2(n13861), .ZN(n10052) );
  NOR2_X1 U12077 ( .A1(n12251), .A2(n10230), .ZN(n10229) );
  INV_X1 U12078 ( .A(n14968), .ZN(n10230) );
  NAND2_X1 U12079 ( .A1(n10132), .A2(n10127), .ZN(n15113) );
  INV_X1 U12080 ( .A(n10130), .ZN(n10129) );
  INV_X1 U12081 ( .A(n15162), .ZN(n10128) );
  NAND2_X1 U12082 ( .A1(n15113), .A2(n15111), .ZN(n12124) );
  NAND2_X1 U12083 ( .A1(n9867), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10038) );
  NAND2_X1 U12084 ( .A1(n9988), .A2(n9986), .ZN(n9989) );
  NOR2_X1 U12085 ( .A1(n9888), .A2(n9987), .ZN(n9986) );
  INV_X1 U12086 ( .A(n12038), .ZN(n9987) );
  INV_X1 U12087 ( .A(n13841), .ZN(n10283) );
  INV_X1 U12088 ( .A(n16540), .ZN(n10261) );
  AND2_X1 U12089 ( .A1(n12183), .A2(n12182), .ZN(n13445) );
  INV_X1 U12090 ( .A(n12297), .ZN(n10027) );
  NAND2_X1 U12091 ( .A1(n10272), .A2(n12301), .ZN(n10271) );
  INV_X1 U12092 ( .A(n13826), .ZN(n10272) );
  INV_X1 U12093 ( .A(n13828), .ZN(n12300) );
  OR2_X1 U12094 ( .A1(n12010), .A2(n12009), .ZN(n12414) );
  OAI21_X1 U12095 ( .B1(n10126), .B2(n9940), .A(n12287), .ZN(n12292) );
  AOI21_X1 U12096 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10406), .ZN(n11684) );
  OR2_X1 U12097 ( .A1(n12880), .A2(n13899), .ZN(n12670) );
  INV_X1 U12098 ( .A(n11729), .ZN(n9981) );
  NAND2_X1 U12099 ( .A1(n11588), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11595) );
  AOI22_X1 U12100 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11507) );
  AOI21_X1 U12101 ( .B1(n9829), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A(n11505), .ZN(n11510) );
  AND2_X1 U12102 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11505) );
  AOI21_X1 U12103 ( .B1(n20159), .B2(n12273), .A(n15655), .ZN(n13884) );
  AOI21_X1 U12104 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18958), .A(
        n14046), .ZN(n14055) );
  AND2_X1 U12105 ( .A1(n15807), .A2(n15806), .ZN(n14046) );
  NOR2_X1 U12106 ( .A1(n19121), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n15806) );
  NAND2_X1 U12107 ( .A1(n19108), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13960) );
  INV_X1 U12108 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21139) );
  AND3_X1 U12109 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17925), .ZN(n16991) );
  NOR2_X1 U12110 ( .A1(n18135), .A2(n18122), .ZN(n16658) );
  NOR2_X1 U12111 ( .A1(n16001), .A2(n10327), .ZN(n10326) );
  NAND2_X1 U12112 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U12113 ( .A1(n16004), .A2(n10326), .ZN(n10323) );
  NAND2_X1 U12114 ( .A1(n10329), .A2(n9915), .ZN(n10328) );
  NAND2_X1 U12115 ( .A1(n15999), .A2(n17828), .ZN(n10329) );
  NOR2_X1 U12116 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10315) );
  NAND2_X1 U12117 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  INV_X1 U12118 ( .A(n10089), .ZN(n10086) );
  INV_X1 U12119 ( .A(n15982), .ZN(n15809) );
  AOI21_X1 U12120 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18967), .A(
        n14049), .ZN(n15808) );
  NAND2_X1 U12121 ( .A1(n18934), .A2(n15788), .ZN(n15946) );
  OAI211_X1 U12122 ( .C1(n9873), .C2(n21364), .A(n14026), .B(n14025), .ZN(
        n14045) );
  AOI211_X1 U12123 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n14024), .B(n14023), .ZN(n14025) );
  OAI211_X1 U12124 ( .C1(n17381), .C2(n21166), .A(n14036), .B(n14035), .ZN(
        n15803) );
  AOI211_X1 U12125 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n14034), .B(n14033), .ZN(n14035) );
  NOR2_X1 U12126 ( .A1(n15946), .A2(n16645), .ZN(n15819) );
  NAND2_X1 U12127 ( .A1(n17723), .A2(n15823), .ZN(n16075) );
  NAND2_X1 U12128 ( .A1(n15791), .A2(n18978), .ZN(n17663) );
  NAND2_X1 U12129 ( .A1(n18499), .A2(n15788), .ZN(n15793) );
  NAND2_X1 U12130 ( .A1(n11002), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11022) );
  INV_X1 U12131 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11021) );
  NOR2_X1 U12132 ( .A1(n10964), .A2(n16269), .ZN(n10971) );
  OR2_X1 U12133 ( .A1(n21117), .A2(n14158), .ZN(n14363) );
  NOR2_X1 U12134 ( .A1(n16190), .A2(n13410), .ZN(n14193) );
  NOR2_X1 U12135 ( .A1(n11389), .A2(n14602), .ZN(n11390) );
  NAND2_X1 U12136 ( .A1(n11390), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11438) );
  AND2_X1 U12137 ( .A1(n11316), .A2(n11315), .ZN(n14294) );
  NOR2_X1 U12138 ( .A1(n16101), .A2(n10361), .ZN(n10359) );
  NAND2_X1 U12139 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11254), .ZN(
        n11276) );
  NAND2_X1 U12140 ( .A1(n14412), .A2(n10360), .ZN(n16102) );
  AND2_X1 U12141 ( .A1(n14412), .A2(n14404), .ZN(n14406) );
  NAND2_X1 U12142 ( .A1(n11211), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U12143 ( .A1(n11172), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11173) );
  NOR2_X1 U12144 ( .A1(n21335), .A2(n11173), .ZN(n11211) );
  INV_X1 U12145 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21335) );
  AND2_X1 U12146 ( .A1(n11152), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11172) );
  AND2_X1 U12147 ( .A1(n11132), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11152) );
  AND2_X1 U12148 ( .A1(n11116), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11132) );
  NOR2_X1 U12149 ( .A1(n11097), .A2(n14332), .ZN(n11116) );
  OR2_X1 U12150 ( .A1(n10364), .A2(n10363), .ZN(n10362) );
  INV_X1 U12151 ( .A(n14438), .ZN(n10363) );
  INV_X1 U12152 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14332) );
  NAND2_X1 U12153 ( .A1(n11041), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11042) );
  NOR2_X1 U12154 ( .A1(n11042), .A2(n16179), .ZN(n11090) );
  NOR2_X1 U12155 ( .A1(n11022), .A2(n11021), .ZN(n11041) );
  AND3_X1 U12156 ( .A1(n11000), .A2(n10999), .A3(n10998), .ZN(n13902) );
  NOR2_X1 U12157 ( .A1(n10345), .A2(n10342), .ZN(n13803) );
  INV_X1 U12158 ( .A(n13731), .ZN(n10342) );
  INV_X1 U12159 ( .A(n13689), .ZN(n10961) );
  NAND2_X1 U12160 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10944) );
  NOR2_X1 U12161 ( .A1(n10944), .A2(n10943), .ZN(n10955) );
  INV_X1 U12162 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10943) );
  INV_X1 U12163 ( .A(n13593), .ZN(n10941) );
  INV_X1 U12164 ( .A(n14135), .ZN(n14145) );
  AND2_X1 U12165 ( .A1(n14133), .A2(n14132), .ZN(n14259) );
  NAND2_X1 U12166 ( .A1(n9973), .A2(n9753), .ZN(n10068) );
  NOR2_X1 U12167 ( .A1(n14399), .A2(n14295), .ZN(n14297) );
  AND2_X1 U12168 ( .A1(n10147), .A2(n9850), .ZN(n14633) );
  NOR2_X1 U12169 ( .A1(n14426), .A2(n14414), .ZN(n14415) );
  NOR3_X1 U12170 ( .A1(n14426), .A2(n10209), .A3(n14414), .ZN(n14409) );
  OR2_X1 U12171 ( .A1(n14424), .A2(n14423), .ZN(n14426) );
  NAND2_X1 U12172 ( .A1(n14664), .A2(n10904), .ZN(n14821) );
  NAND2_X1 U12173 ( .A1(n14436), .A2(n14310), .ZN(n14424) );
  AND2_X1 U12174 ( .A1(n16212), .A2(n21199), .ZN(n16230) );
  AND3_X1 U12175 ( .A1(n14095), .A2(n14094), .A3(n14093), .ZN(n14450) );
  INV_X1 U12176 ( .A(n14769), .ZN(n14847) );
  NOR2_X1 U12177 ( .A1(n16355), .A2(n10203), .ZN(n14456) );
  INV_X1 U12178 ( .A(n10205), .ZN(n10203) );
  AND2_X1 U12179 ( .A1(n13928), .A2(n10412), .ZN(n10143) );
  AND2_X1 U12180 ( .A1(n14090), .A2(n14089), .ZN(n14339) );
  NOR2_X1 U12181 ( .A1(n16355), .A2(n14339), .ZN(n14455) );
  NOR2_X1 U12182 ( .A1(n14844), .A2(n13538), .ZN(n14695) );
  NAND2_X1 U12183 ( .A1(n21102), .A2(n21027), .ZN(n11501) );
  AND2_X1 U12184 ( .A1(n14208), .A2(n14120), .ZN(n14135) );
  AND2_X1 U12185 ( .A1(n13229), .A2(n10588), .ZN(n13130) );
  NAND2_X1 U12186 ( .A1(n10721), .A2(n10379), .ZN(n10377) );
  NAND2_X1 U12187 ( .A1(n10675), .A2(n9893), .ZN(n10378) );
  NAND2_X1 U12188 ( .A1(n10736), .A2(n10734), .ZN(n10732) );
  NAND2_X1 U12189 ( .A1(n10823), .A2(n13656), .ZN(n20380) );
  NAND2_X1 U12190 ( .A1(n9975), .A2(n16039), .ZN(n13584) );
  INV_X1 U12191 ( .A(n9976), .ZN(n14858) );
  INV_X1 U12192 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21260) );
  AND2_X1 U12193 ( .A1(n13328), .A2(n13255), .ZN(n16026) );
  AND2_X1 U12194 ( .A1(n20380), .A2(n13603), .ZN(n20494) );
  OR2_X1 U12195 ( .A1(n13604), .A2(n20381), .ZN(n20724) );
  INV_X1 U12196 ( .A(n20724), .ZN(n20860) );
  NAND2_X1 U12197 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  INV_X1 U12198 ( .A(n20745), .ZN(n20887) );
  AND3_X1 U12199 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21027), .A3(n20383), 
        .ZN(n20425) );
  AND2_X1 U12200 ( .A1(n10578), .A2(n10607), .ZN(n13057) );
  OR2_X1 U12201 ( .A1(n10608), .A2(n10577), .ZN(n10578) );
  NAND2_X1 U12202 ( .A1(n16454), .A2(n16441), .ZN(n16439) );
  NOR2_X1 U12203 ( .A1(n14911), .A2(n19312), .ZN(n16449) );
  NAND2_X1 U12204 ( .A1(n13002), .A2(n9939), .ZN(n15055) );
  NOR2_X1 U12205 ( .A1(n19242), .A2(n9874), .ZN(n13855) );
  NAND2_X1 U12206 ( .A1(n19253), .A2(n19254), .ZN(n19242) );
  NOR2_X1 U12207 ( .A1(n19265), .A2(n19266), .ZN(n19253) );
  NAND2_X1 U12208 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  INV_X1 U12209 ( .A(n10252), .ZN(n10251) );
  NAND2_X1 U12210 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10307) );
  NOR2_X1 U12211 ( .A1(n19328), .A2(n19330), .ZN(n19311) );
  NAND2_X1 U12212 ( .A1(n13757), .A2(n13756), .ZN(n19328) );
  NOR2_X1 U12213 ( .A1(n13789), .A2(n13791), .ZN(n13757) );
  AND2_X1 U12214 ( .A1(n12226), .A2(n12225), .ZN(n12986) );
  OR2_X1 U12215 ( .A1(n12442), .A2(n12441), .ZN(n12686) );
  AND2_X1 U12216 ( .A1(n13675), .A2(n9941), .ZN(n10401) );
  NAND2_X1 U12217 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10245) );
  INV_X1 U12218 ( .A(n12882), .ZN(n10392) );
  NAND2_X1 U12219 ( .A1(n13002), .A2(n9944), .ZN(n15037) );
  XNOR2_X1 U12220 ( .A(n12861), .B(n12863), .ZN(n14973) );
  INV_X1 U12221 ( .A(n10112), .ZN(n15063) );
  INV_X1 U12222 ( .A(n13002), .ZN(n13021) );
  CLKBUF_X1 U12223 ( .A(n14991), .Z(n14992) );
  AND2_X1 U12224 ( .A1(n12516), .A2(n12515), .ZN(n15085) );
  AND2_X1 U12225 ( .A1(n12514), .A2(n12513), .ZN(n14935) );
  OR2_X1 U12226 ( .A1(n15099), .A2(n14935), .ZN(n15086) );
  AND2_X1 U12227 ( .A1(n15509), .A2(n15510), .ZN(n15512) );
  NAND2_X1 U12228 ( .A1(n15512), .A2(n15097), .ZN(n15099) );
  OR2_X1 U12229 ( .A1(n12709), .A2(n12708), .ZN(n15004) );
  AND3_X1 U12230 ( .A1(n12458), .A2(n12457), .A3(n12456), .ZN(n15588) );
  AND2_X1 U12231 ( .A1(n13147), .A2(n20151), .ZN(n19429) );
  AND2_X1 U12232 ( .A1(n9858), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10294) );
  NOR3_X1 U12233 ( .A1(n13018), .A2(n13017), .A3(n10224), .ZN(n14989) );
  CLKBUF_X1 U12234 ( .A(n12352), .Z(n12355) );
  AND2_X1 U12235 ( .A1(n9848), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10298) );
  AND2_X1 U12236 ( .A1(n15300), .A2(n10225), .ZN(n13846) );
  AND2_X1 U12237 ( .A1(n12201), .A2(n12200), .ZN(n13684) );
  NAND2_X1 U12238 ( .A1(n15300), .A2(n9916), .ZN(n13845) );
  NAND2_X1 U12239 ( .A1(n15300), .A2(n15299), .ZN(n15302) );
  AND2_X1 U12240 ( .A1(n12194), .A2(n12193), .ZN(n13665) );
  CLKBUF_X1 U12241 ( .A(n12339), .Z(n12348) );
  AND2_X1 U12242 ( .A1(n12174), .A2(n12173), .ZN(n13343) );
  NAND2_X1 U12243 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12344) );
  INV_X1 U12244 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13793) );
  OR2_X1 U12245 ( .A1(n11761), .A2(n11760), .ZN(n13203) );
  NOR2_X1 U12246 ( .A1(n15013), .A2(n15014), .ZN(n15361) );
  NAND2_X1 U12247 ( .A1(n15163), .A2(n9959), .ZN(n15147) );
  NOR2_X1 U12248 ( .A1(n14899), .A2(n15119), .ZN(n15109) );
  XNOR2_X1 U12249 ( .A(n12124), .B(n15106), .ZN(n15154) );
  AND2_X1 U12250 ( .A1(n15163), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15152) );
  OR2_X1 U12251 ( .A1(n10223), .A2(n14904), .ZN(n10222) );
  NAND2_X1 U12252 ( .A1(n15622), .A2(n9867), .ZN(n15185) );
  NAND2_X1 U12253 ( .A1(n13002), .A2(n10409), .ZN(n15053) );
  NOR2_X1 U12254 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  AND2_X1 U12255 ( .A1(n12213), .A2(n12212), .ZN(n15006) );
  NAND2_X1 U12256 ( .A1(n10057), .A2(n10054), .ZN(n15262) );
  AND2_X1 U12257 ( .A1(n10055), .A2(n15274), .ZN(n10054) );
  OR2_X1 U12258 ( .A1(n15207), .A2(n10056), .ZN(n10055) );
  NOR2_X2 U12259 ( .A1(n15569), .A2(n10282), .ZN(n15509) );
  NAND2_X1 U12260 ( .A1(n9856), .A2(n13627), .ZN(n10282) );
  NAND2_X1 U12261 ( .A1(n12046), .A2(n12045), .ZN(n10333) );
  NAND2_X1 U12262 ( .A1(n12044), .A2(n15310), .ZN(n10334) );
  AND2_X1 U12263 ( .A1(n9921), .A2(n13319), .ZN(n10287) );
  AND2_X1 U12264 ( .A1(n10289), .A2(n9921), .ZN(n13777) );
  NAND2_X1 U12265 ( .A1(n13836), .A2(n13835), .ZN(n11968) );
  OR2_X1 U12266 ( .A1(n13825), .A2(n13826), .ZN(n13829) );
  NOR3_X1 U12267 ( .A1(n16583), .A2(n16594), .A3(n16582), .ZN(n15645) );
  AND3_X1 U12268 ( .A1(n12410), .A2(n12409), .A3(n12408), .ZN(n13672) );
  NAND2_X1 U12269 ( .A1(n9978), .A2(n13636), .ZN(n9979) );
  NAND2_X1 U12270 ( .A1(n10042), .A2(n9920), .ZN(n9978) );
  NAND2_X1 U12271 ( .A1(n11831), .A2(n12289), .ZN(n10126) );
  NAND2_X1 U12272 ( .A1(n11677), .A2(n9984), .ZN(n9983) );
  INV_X1 U12273 ( .A(n11667), .ZN(n9984) );
  NAND2_X1 U12274 ( .A1(n10042), .A2(n13794), .ZN(n13638) );
  INV_X1 U12275 ( .A(n12397), .ZN(n10277) );
  NAND2_X1 U12276 ( .A1(n13279), .A2(n10423), .ZN(n10278) );
  INV_X1 U12277 ( .A(n10276), .ZN(n10273) );
  OR2_X1 U12278 ( .A1(n15494), .A2(n15500), .ZN(n15498) );
  INV_X1 U12279 ( .A(n12544), .ZN(n20140) );
  XNOR2_X1 U12280 ( .A(n13210), .B(n12393), .ZN(n13277) );
  INV_X1 U12281 ( .A(n19504), .ZN(n20106) );
  NAND2_X1 U12282 ( .A1(n12682), .A2(n13310), .ZN(n13351) );
  INV_X1 U12283 ( .A(n12659), .ZN(n10395) );
  AND2_X1 U12284 ( .A1(n20117), .A2(n20124), .ZN(n19500) );
  INV_X1 U12285 ( .A(n11992), .ZN(n19603) );
  INV_X1 U12286 ( .A(n11943), .ZN(n19634) );
  INV_X1 U12287 ( .A(n11735), .ZN(n9980) );
  NOR2_X2 U12288 ( .A1(n13881), .A2(n13882), .ZN(n19493) );
  NAND2_X1 U12289 ( .A1(n20106), .A2(n20133), .ZN(n19912) );
  OR2_X1 U12290 ( .A1(n20117), .A2(n20127), .ZN(n19882) );
  INV_X2 U12291 ( .A(n12629), .ZN(n19467) );
  NAND2_X1 U12292 ( .A1(n9882), .A2(n15689), .ZN(n11608) );
  INV_X1 U12293 ( .A(n19494), .ZN(n19488) );
  INV_X1 U12294 ( .A(n19493), .ZN(n19487) );
  OR2_X1 U12295 ( .A1(n19912), .A2(n19949), .ZN(n19919) );
  OR2_X1 U12296 ( .A1(n20117), .A2(n20124), .ZN(n19949) );
  AND2_X1 U12297 ( .A1(n13873), .A2(n13872), .ZN(n16611) );
  OR2_X1 U12298 ( .A1(n12550), .A2(n20132), .ZN(n13874) );
  INV_X1 U12299 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15656) );
  NOR2_X1 U12300 ( .A1(n15793), .A2(n15799), .ZN(n15796) );
  NOR2_X1 U12301 ( .A1(n18488), .A2(n15805), .ZN(n15811) );
  NAND2_X1 U12302 ( .A1(n18479), .A2(n19141), .ZN(n15944) );
  NAND2_X1 U12303 ( .A1(n17156), .A2(n16682), .ZN(n10153) );
  NAND2_X1 U12304 ( .A1(n10152), .A2(n9865), .ZN(n10151) );
  OR2_X1 U12305 ( .A1(n16920), .A2(n17831), .ZN(n10159) );
  NOR2_X1 U12306 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17016), .ZN(n17004) );
  AND2_X1 U12307 ( .A1(n17431), .A2(n10193), .ZN(n17319) );
  AND2_X1 U12308 ( .A1(n10195), .A2(n10194), .ZN(n10193) );
  NOR2_X1 U12309 ( .A1(n17344), .A2(n17345), .ZN(n10194) );
  NOR2_X1 U12310 ( .A1(n21223), .A2(n17065), .ZN(n10197) );
  NOR2_X1 U12311 ( .A1(n17676), .A2(n10168), .ZN(n10167) );
  OAI211_X1 U12312 ( .C1(n17473), .C2(n21259), .A(n14006), .B(n14005), .ZN(
        n17523) );
  AOI211_X1 U12313 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14004), .B(n14003), .ZN(n14005) );
  NAND4_X1 U12314 ( .A1(n14016), .A2(n14015), .A3(n14014), .A4(n14013), .ZN(
        n17527) );
  INV_X1 U12315 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15773) );
  INV_X1 U12316 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21244) );
  NOR2_X1 U12317 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10013) );
  INV_X1 U12318 ( .A(n13958), .ZN(n10014) );
  NAND2_X1 U12319 ( .A1(n18942), .A2(n13963), .ZN(n17467) );
  NAND2_X1 U12320 ( .A1(n16080), .A2(n19149), .ZN(n17521) );
  OAI211_X1 U12321 ( .C1(n17483), .C2(n17477), .A(n13996), .B(n13995), .ZN(
        n17666) );
  AOI22_X1 U12322 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15875), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13996) );
  AOI211_X1 U12323 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13994), .B(n13993), .ZN(n13995) );
  NOR2_X1 U12324 ( .A1(n17665), .A2(n17664), .ZN(n17693) );
  NAND2_X1 U12325 ( .A1(n19140), .A2(n17663), .ZN(n17664) );
  OR2_X1 U12326 ( .A1(n15793), .A2(n15792), .ZN(n17723) );
  AND2_X1 U12327 ( .A1(n17771), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17775) );
  NAND2_X1 U12328 ( .A1(n10310), .A2(n10309), .ZN(n16710) );
  AND3_X1 U12329 ( .A1(n10312), .A2(n10313), .A3(n9788), .ZN(n10309) );
  NAND2_X1 U12330 ( .A1(n17783), .A2(n17784), .ZN(n17782) );
  NAND2_X1 U12331 ( .A1(n17775), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16851) );
  NOR2_X1 U12332 ( .A1(n17800), .A2(n17801), .ZN(n17771) );
  NOR2_X1 U12333 ( .A1(n10161), .A2(n10162), .ZN(n10160) );
  INV_X1 U12334 ( .A(n16848), .ZN(n17854) );
  NOR2_X1 U12335 ( .A1(n17899), .A2(n17888), .ZN(n16980) );
  NAND2_X1 U12336 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16991), .ZN(
        n17888) );
  NOR2_X1 U12337 ( .A1(n17910), .A2(n17909), .ZN(n17887) );
  NOR3_X1 U12338 ( .A1(n17970), .A2(n17972), .A3(n17957), .ZN(n17924) );
  OR2_X1 U12339 ( .A1(n17972), .A2(n17055), .ZN(n17035) );
  NOR2_X1 U12340 ( .A1(n17057), .A2(n17070), .ZN(n17969) );
  INV_X1 U12341 ( .A(n17969), .ZN(n17055) );
  NOR2_X1 U12342 ( .A1(n17069), .A2(n18013), .ZN(n17955) );
  NOR2_X1 U12343 ( .A1(n17954), .A2(n18066), .ZN(n18038) );
  NAND2_X1 U12344 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18088) );
  AND2_X1 U12345 ( .A1(n9788), .A2(n16708), .ZN(n16711) );
  AOI21_X1 U12346 ( .B1(n16712), .B2(n18331), .A(n16713), .ZN(n10319) );
  INV_X1 U12347 ( .A(n18275), .ZN(n18207) );
  NOR2_X1 U12348 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15993), .ZN(
        n17868) );
  INV_X1 U12349 ( .A(n17867), .ZN(n10094) );
  AOI21_X1 U12350 ( .B1(n17920), .B2(n16004), .A(n15998), .ZN(n17916) );
  OAI22_X1 U12351 ( .A1(n15999), .A2(n15997), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16004), .ZN(n15998) );
  NAND2_X1 U12352 ( .A1(n17916), .A2(n18250), .ZN(n17915) );
  NAND2_X1 U12353 ( .A1(n15995), .A2(n10141), .ZN(n17940) );
  NOR2_X1 U12354 ( .A1(n10314), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10141) );
  INV_X1 U12355 ( .A(n10315), .ZN(n10314) );
  NAND2_X1 U12356 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17960), .ZN(
        n18278) );
  NAND2_X1 U12357 ( .A1(n18036), .A2(n15979), .ZN(n17962) );
  INV_X1 U12358 ( .A(n15977), .ZN(n15975) );
  NOR2_X1 U12359 ( .A1(n18291), .A2(n17961), .ZN(n17960) );
  NOR2_X1 U12360 ( .A1(n17940), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17952) );
  INV_X1 U12361 ( .A(n17962), .ZN(n18332) );
  NOR2_X1 U12362 ( .A1(n18009), .A2(n9788), .ZN(n18022) );
  NAND2_X1 U12363 ( .A1(n18069), .A2(n15974), .ZN(n18055) );
  NAND2_X1 U12364 ( .A1(n18094), .A2(n15970), .ZN(n18076) );
  NAND2_X1 U12365 ( .A1(n18076), .A2(n18077), .ZN(n18075) );
  XNOR2_X1 U12366 ( .A(n15968), .B(n10012), .ZN(n18095) );
  INV_X1 U12367 ( .A(n15969), .ZN(n10012) );
  NAND2_X1 U12368 ( .A1(n18095), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18094) );
  XNOR2_X1 U12369 ( .A(n15962), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18117) );
  NOR3_X1 U12370 ( .A1(n15925), .A2(n15924), .A3(n15923), .ZN(n15926) );
  INV_X1 U12371 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18958) );
  INV_X1 U12372 ( .A(n15949), .ZN(n18927) );
  NAND2_X1 U12373 ( .A1(n18928), .A2(n15949), .ZN(n15823) );
  INV_X1 U12374 ( .A(n14045), .ZN(n18488) );
  NOR2_X1 U12375 ( .A1(n10192), .A2(n10183), .ZN(n18495) );
  INV_X1 U12376 ( .A(n14039), .ZN(n10192) );
  INV_X1 U12377 ( .A(n17527), .ZN(n18499) );
  OR2_X1 U12378 ( .A1(n15945), .A2(n15793), .ZN(n18978) );
  OAI22_X1 U12379 ( .A1(n13368), .A2(n10371), .B1(n13139), .B2(n13138), .ZN(
        n20172) );
  AND2_X1 U12380 ( .A1(n14173), .A2(n14153), .ZN(n20260) );
  INV_X1 U12381 ( .A(n20260), .ZN(n20279) );
  NAND2_X1 U12382 ( .A1(n14173), .A2(n14171), .ZN(n20273) );
  NAND2_X1 U12383 ( .A1(n21117), .A2(n10371), .ZN(n14357) );
  NAND2_X1 U12384 ( .A1(n14173), .A2(n14172), .ZN(n20276) );
  INV_X1 U12385 ( .A(n20288), .ZN(n20298) );
  INV_X1 U12386 ( .A(n20302), .ZN(n14458) );
  AND2_X2 U12387 ( .A1(n13329), .A2(n13403), .ZN(n20302) );
  INV_X1 U12388 ( .A(n16196), .ZN(n14537) );
  INV_X1 U12389 ( .A(n14465), .ZN(n16191) );
  NAND2_X1 U12390 ( .A1(n14193), .A2(n20379), .ZN(n14540) );
  INV_X1 U12391 ( .A(n14553), .ZN(n16193) );
  OR2_X1 U12392 ( .A1(n16191), .A2(n14193), .ZN(n14555) );
  AND2_X1 U12393 ( .A1(n13404), .A2(n13403), .ZN(n14546) );
  NAND2_X1 U12394 ( .A1(n13402), .A2(n13401), .ZN(n13404) );
  NAND2_X1 U12395 ( .A1(n13400), .A2(n10371), .ZN(n13401) );
  INV_X1 U12396 ( .A(n14555), .ZN(n14548) );
  INV_X2 U12397 ( .A(n13452), .ZN(n20363) );
  XNOR2_X1 U12398 ( .A(n11500), .B(n14174), .ZN(n14214) );
  OR2_X1 U12399 ( .A1(n10350), .A2(n11495), .ZN(n10348) );
  OR2_X1 U12400 ( .A1(n14231), .A2(n11495), .ZN(n10347) );
  NAND2_X1 U12401 ( .A1(n10071), .A2(n9753), .ZN(n14626) );
  INV_X1 U12402 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16117) );
  AOI21_X1 U12403 ( .B1(n14449), .B2(n14448), .A(n14447), .ZN(n16240) );
  INV_X1 U12404 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16261) );
  INV_X1 U12405 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16269) );
  INV_X1 U12406 ( .A(n20369), .ZN(n16244) );
  INV_X1 U12407 ( .A(n16268), .ZN(n20367) );
  NAND2_X1 U12408 ( .A1(n14600), .A2(n9962), .ZN(n9961) );
  AND2_X1 U12409 ( .A1(n14235), .A2(n14234), .ZN(n14737) );
  NAND2_X1 U12410 ( .A1(n10147), .A2(n10383), .ZN(n14641) );
  NAND2_X1 U12411 ( .A1(n14654), .A2(n10901), .ZN(n14668) );
  NAND2_X1 U12412 ( .A1(n9770), .A2(n13928), .ZN(n14684) );
  NAND2_X1 U12413 ( .A1(n9775), .A2(n10892), .ZN(n13930) );
  INV_X1 U12414 ( .A(n16319), .ZN(n16400) );
  INV_X1 U12415 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21321) );
  INV_X1 U12416 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20679) );
  NOR2_X1 U12417 ( .A1(n13656), .A2(n13655), .ZN(n20637) );
  INV_X1 U12418 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20376) );
  NOR2_X1 U12419 ( .A1(n14862), .A2(n9974), .ZN(n14863) );
  NOR2_X1 U12420 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21102) );
  OAI211_X1 U12421 ( .C1(n20536), .C2(n21030), .A(n20755), .B(n20389), .ZN(
        n20430) );
  OAI221_X1 U12422 ( .B1(n20546), .B2(n20840), .C1(n20546), .C2(n20545), .A(
        n20900), .ZN(n20571) );
  NAND2_X1 U12423 ( .A1(n20637), .A2(n20860), .ZN(n20630) );
  OAI211_X1 U12424 ( .C1(n20689), .C2(n20840), .A(n20755), .B(n20688), .ZN(
        n20714) );
  OR2_X1 U12425 ( .A1(n20797), .A2(n20724), .ZN(n20773) );
  OAI211_X1 U12426 ( .C1(n10410), .C2(n20840), .A(n20900), .B(n20839), .ZN(
        n20856) );
  OAI211_X1 U12427 ( .C1(n20945), .C2(n20901), .A(n20900), .B(n20899), .ZN(
        n20949) );
  INV_X1 U12428 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21324) );
  OAI21_X1 U12429 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n15656), .A(n12253), 
        .ZN(n20159) );
  NOR2_X1 U12430 ( .A1(n16421), .A2(n16420), .ZN(n16418) );
  NOR2_X1 U12431 ( .A1(n14894), .A2(n19312), .ZN(n16421) );
  NOR2_X1 U12432 ( .A1(n14896), .A2(n14895), .ZN(n14894) );
  CLKBUF_X1 U12433 ( .A(n16449), .Z(n16450) );
  NOR2_X1 U12434 ( .A1(n16466), .A2(n19312), .ZN(n14912) );
  NOR2_X1 U12435 ( .A1(n14912), .A2(n15177), .ZN(n14911) );
  NOR2_X1 U12436 ( .A1(n16464), .A2(n16467), .ZN(n16466) );
  CLKBUF_X1 U12437 ( .A(n16464), .Z(n16465) );
  CLKBUF_X1 U12438 ( .A(n12994), .Z(n12995) );
  CLKBUF_X1 U12439 ( .A(n13010), .Z(n13011) );
  AOI21_X1 U12440 ( .B1(n10307), .B2(n10103), .A(n10100), .ZN(n19197) );
  NOR2_X1 U12441 ( .A1(n10102), .A2(n10101), .ZN(n10100) );
  NAND2_X1 U12442 ( .A1(n10104), .A2(n21322), .ZN(n10103) );
  INV_X1 U12443 ( .A(n15126), .ZN(n10104) );
  NAND2_X1 U12444 ( .A1(n13855), .A2(n16520), .ZN(n19227) );
  NAND2_X1 U12445 ( .A1(n19311), .A2(n19313), .ZN(n19294) );
  AND2_X1 U12446 ( .A1(n19166), .A2(n12361), .ZN(n19339) );
  OAI21_X1 U12447 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A(n10099), .ZN(n19352) );
  NAND2_X1 U12448 ( .A1(n13273), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10099) );
  INV_X1 U12449 ( .A(n19282), .ZN(n19349) );
  OR2_X1 U12450 ( .A1(n12374), .A2(n12373), .ZN(n19360) );
  OR2_X1 U12451 ( .A1(n12429), .A2(n12428), .ZN(n19379) );
  NAND2_X1 U12452 ( .A1(n13676), .A2(n10401), .ZN(n13443) );
  NAND2_X1 U12453 ( .A1(n13676), .A2(n13675), .ZN(n13342) );
  INV_X1 U12454 ( .A(n19380), .ZN(n19386) );
  INV_X1 U12455 ( .A(n15096), .ZN(n19396) );
  NAND2_X1 U12456 ( .A1(n10290), .A2(n9908), .ZN(n13198) );
  OR2_X1 U12457 ( .A1(n13200), .A2(n13199), .ZN(n10290) );
  AND2_X1 U12458 ( .A1(n19400), .A2(n19422), .ZN(n19428) );
  NOR2_X1 U12459 ( .A1(n13261), .A2(n13266), .ZN(n19501) );
  INV_X1 U12460 ( .A(n19422), .ZN(n16501) );
  NAND2_X1 U12461 ( .A1(n15094), .A2(n13196), .ZN(n13679) );
  INV_X1 U12462 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15215) );
  INV_X1 U12463 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19191) );
  INV_X1 U12464 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16564) );
  OR2_X1 U12465 ( .A1(n12313), .A2(n12544), .ZN(n16558) );
  AND2_X1 U12466 ( .A1(n12159), .A2(n20141), .ZN(n16549) );
  NOR2_X1 U12467 ( .A1(n10269), .A2(n15333), .ZN(n10267) );
  AND2_X1 U12468 ( .A1(n9784), .A2(n10130), .ZN(n15160) );
  NAND2_X1 U12469 ( .A1(n9784), .A2(n10335), .ZN(n15172) );
  XNOR2_X1 U12470 ( .A(n10046), .B(n15214), .ZN(n15440) );
  NAND2_X1 U12471 ( .A1(n10047), .A2(n15221), .ZN(n10046) );
  NAND2_X1 U12472 ( .A1(n15223), .A2(n15222), .ZN(n10047) );
  OAI21_X1 U12473 ( .B1(n15538), .B2(n15206), .A(n15535), .ZN(n15275) );
  NOR2_X1 U12474 ( .A1(n15569), .A2(n15568), .ZN(n13589) );
  AND2_X1 U12475 ( .A1(n10339), .A2(n9917), .ZN(n15605) );
  NAND2_X1 U12476 ( .A1(n10339), .A2(n12030), .ZN(n15620) );
  NAND2_X1 U12477 ( .A1(n10259), .A2(n10264), .ZN(n16541) );
  NAND2_X1 U12478 ( .A1(n15320), .A2(n10265), .ZN(n10259) );
  INV_X1 U12479 ( .A(n16581), .ZN(n15602) );
  INV_X1 U12480 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21258) );
  INV_X1 U12481 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20121) );
  NOR2_X2 U12482 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20102) );
  INV_X1 U12483 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16074) );
  INV_X1 U12484 ( .A(n20127), .ZN(n20124) );
  INV_X1 U12485 ( .A(n10118), .ZN(n16598) );
  INV_X1 U12486 ( .A(n15677), .ZN(n10119) );
  INV_X1 U12487 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15830) );
  NOR2_X1 U12488 ( .A1(n19750), .A2(n19698), .ZN(n19554) );
  AND2_X1 U12489 ( .A1(n19661), .A2(n19537), .ZN(n19589) );
  INV_X1 U12490 ( .A(n19773), .ZN(n19774) );
  NOR2_X1 U12491 ( .A1(n19883), .A2(n19750), .ZN(n19800) );
  INV_X1 U12492 ( .A(n20012), .ZN(n19842) );
  NOR2_X1 U12493 ( .A1(n19883), .A2(n20103), .ZN(n19870) );
  OR2_X1 U12494 ( .A1(n19883), .A2(n19882), .ZN(n19913) );
  OAI21_X1 U12495 ( .B1(n19924), .B2(n19923), .A(n19922), .ZN(n19943) );
  INV_X1 U12496 ( .A(n19913), .ZN(n19942) );
  INV_X1 U12497 ( .A(n19823), .ZN(n19970) );
  INV_X1 U12498 ( .A(n19512), .ZN(n19967) );
  OAI22_X1 U12499 ( .A1(n16744), .A2(n19488), .B1(n21230), .B2(n19487), .ZN(
        n19996) );
  INV_X1 U12500 ( .A(n19901), .ZN(n19997) );
  INV_X1 U12501 ( .A(n19521), .ZN(n19994) );
  INV_X1 U12502 ( .A(n19905), .ZN(n20004) );
  NOR2_X2 U12503 ( .A1(n19883), .A2(n19949), .ZN(n20015) );
  OAI22_X1 U12504 ( .A1(n19489), .A2(n19488), .B1(n21238), .B2(n19487), .ZN(
        n20012) );
  INV_X1 U12505 ( .A(n19911), .ZN(n20014) );
  INV_X1 U12506 ( .A(n19919), .ZN(n20013) );
  INV_X1 U12507 ( .A(n13874), .ZN(n20165) );
  INV_X1 U12508 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20110) );
  NAND2_X1 U12509 ( .A1(n18922), .A2(n17724), .ZN(n19158) );
  NOR2_X1 U12510 ( .A1(n15796), .A2(n15811), .ZN(n16821) );
  INV_X1 U12511 ( .A(n19158), .ZN(n19162) );
  OR2_X1 U12512 ( .A1(n18985), .A2(n16646), .ZN(n16822) );
  AND2_X1 U12513 ( .A1(n10156), .A2(n10155), .ZN(n16901) );
  NOR2_X1 U12514 ( .A1(n17156), .A2(n10164), .ZN(n16960) );
  NOR2_X1 U12515 ( .A1(n17890), .A2(n10165), .ZN(n10164) );
  INV_X1 U12516 ( .A(n16849), .ZN(n10165) );
  NOR2_X1 U12517 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16994), .ZN(n16985) );
  NOR2_X1 U12518 ( .A1(n17156), .A2(n16849), .ZN(n16967) );
  NOR2_X1 U12519 ( .A1(n16967), .A2(n17890), .ZN(n16966) );
  NOR2_X1 U12520 ( .A1(n19160), .A2(n18977), .ZN(n17160) );
  INV_X1 U12521 ( .A(n17160), .ZN(n17195) );
  INV_X1 U12522 ( .A(n17186), .ZN(n17205) );
  NOR2_X1 U12523 ( .A1(n17220), .A2(n17219), .ZN(n17247) );
  NOR2_X1 U12524 ( .A1(n17212), .A2(n17256), .ZN(n17261) );
  NOR2_X1 U12525 ( .A1(n17210), .A2(n17265), .ZN(n17270) );
  NOR3_X1 U12526 ( .A1(n10198), .A2(n10199), .A3(n10196), .ZN(n10195) );
  INV_X1 U12527 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n10199) );
  INV_X1 U12528 ( .A(n10197), .ZN(n10196) );
  INV_X1 U12529 ( .A(n15695), .ZN(n10198) );
  NAND2_X1 U12530 ( .A1(n17431), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17428) );
  AND2_X1 U12531 ( .A1(n17487), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17486) );
  NOR3_X1 U12532 ( .A1(n9909), .A2(n17112), .A3(n17493), .ZN(n17487) );
  NOR2_X1 U12533 ( .A1(n14072), .A2(n17502), .ZN(n17499) );
  NAND2_X1 U12534 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17499), .ZN(n17498) );
  INV_X1 U12535 ( .A(n14072), .ZN(n17520) );
  INV_X1 U12536 ( .A(n17537), .ZN(n17533) );
  AND2_X1 U12537 ( .A1(n17555), .A2(n10166), .ZN(n17541) );
  AND2_X1 U12538 ( .A1(n9870), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U12539 ( .A1(n17555), .A2(n9870), .ZN(n17546) );
  NAND2_X1 U12540 ( .A1(n17555), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17554) );
  NOR2_X1 U12541 ( .A1(n17681), .A2(n17564), .ZN(n17560) );
  AOI22_X1 U12542 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15874), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13973) );
  AOI211_X1 U12543 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n13971), .B(n13970), .ZN(n13972) );
  NOR2_X1 U12544 ( .A1(n17692), .A2(n17601), .ZN(n17596) );
  INV_X1 U12545 ( .A(n17593), .ZN(n17594) );
  AND2_X1 U12546 ( .A1(n16080), .A2(n9953), .ZN(n17606) );
  NOR2_X1 U12547 ( .A1(n17522), .A2(n10177), .ZN(n10174) );
  NAND3_X1 U12548 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U12549 ( .A1(n17521), .A2(n18511), .ZN(n17607) );
  OR2_X1 U12550 ( .A1(n15863), .A2(n10135), .ZN(n10134) );
  AND2_X1 U12551 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10135) );
  AND2_X1 U12552 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17647), .ZN(n17650) );
  INV_X1 U12553 ( .A(n17607), .ZN(n17651) );
  AOI211_X1 U12554 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n15871), .B(n15870), .ZN(n15872) );
  OR2_X1 U12555 ( .A1(n17633), .A2(n17632), .ZN(n17656) );
  NOR2_X1 U12556 ( .A1(n10097), .A2(n10095), .ZN(n15885) );
  INV_X1 U12557 ( .A(n17653), .ZN(n17661) );
  INV_X1 U12558 ( .A(n17662), .ZN(n17654) );
  CLKBUF_X1 U12559 ( .A(n17744), .Z(n21457) );
  INV_X1 U12560 ( .A(n17762), .ZN(n21455) );
  NOR2_X1 U12561 ( .A1(n17752), .A2(n18484), .ZN(n17767) );
  NAND2_X1 U12562 ( .A1(n16671), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16656) );
  INV_X1 U12563 ( .A(n17998), .ZN(n17977) );
  INV_X1 U12564 ( .A(n17933), .ZN(n17850) );
  NAND2_X1 U12565 ( .A1(n17887), .A2(n10417), .ZN(n17877) );
  INV_X1 U12566 ( .A(n17985), .ZN(n17927) );
  INV_X1 U12567 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17909) );
  INV_X1 U12568 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17957) );
  NOR2_X1 U12569 ( .A1(n18122), .A2(n18089), .ZN(n18068) );
  INV_X1 U12570 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18013) );
  AOI22_X1 U12571 ( .A1(n18127), .A2(n17962), .B1(n17998), .B2(n16668), .ZN(
        n18035) );
  INV_X1 U12572 ( .A(n18330), .ZN(n16668) );
  AND2_X1 U12573 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18041) );
  INV_X1 U12574 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21294) );
  NOR2_X1 U12575 ( .A1(n18088), .A2(n18100), .ZN(n18085) );
  INV_X1 U12576 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18100) );
  NOR2_X2 U12577 ( .A1(n18516), .A2(n18828), .ZN(n18866) );
  NOR2_X2 U12578 ( .A1(n19141), .A2(n16822), .ZN(n18127) );
  OAI21_X2 U12579 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19148), .A(n16822), 
        .ZN(n18136) );
  OR2_X1 U12580 ( .A1(n18150), .A2(n18306), .ZN(n10010) );
  NAND2_X1 U12581 ( .A1(n18405), .A2(n18923), .ZN(n18367) );
  NAND2_X1 U12582 ( .A1(n17962), .A2(n16718), .ZN(n18275) );
  INV_X1 U12583 ( .A(n18929), .ZN(n18950) );
  NAND2_X1 U12584 ( .A1(n15995), .A2(n10133), .ZN(n17995) );
  INV_X1 U12585 ( .A(n10316), .ZN(n10133) );
  INV_X1 U12586 ( .A(n15995), .ZN(n10077) );
  INV_X1 U12587 ( .A(n18302), .ZN(n18373) );
  AND2_X1 U12588 ( .A1(n10091), .A2(n10088), .ZN(n18065) );
  NAND2_X1 U12589 ( .A1(n18080), .A2(n18079), .ZN(n18078) );
  NAND2_X1 U12590 ( .A1(n18090), .A2(n15934), .ZN(n18080) );
  INV_X1 U12591 ( .A(n18952), .ZN(n18458) );
  INV_X1 U12592 ( .A(n18431), .ZN(n18456) );
  INV_X1 U12593 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18967) );
  INV_X1 U12594 ( .A(n19122), .ZN(n19119) );
  INV_X1 U12595 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18710) );
  INV_X1 U12596 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n21166) );
  INV_X1 U12597 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18814) );
  NAND2_X1 U12598 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18990), .ZN(n18985) );
  NOR2_X1 U12599 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19146), .ZN(n18990) );
  INV_X1 U12600 ( .A(n20379), .ZN(n20377) );
  OAI21_X1 U12602 ( .B1(n14710), .B2(n16319), .A(n10060), .ZN(P1_U3000) );
  NOR2_X1 U12603 ( .A1(n14708), .A2(n14709), .ZN(n10201) );
  NOR2_X1 U12604 ( .A1(n9889), .A2(n10221), .ZN(n10040) );
  NAND2_X1 U12605 ( .A1(n15352), .A2(n16550), .ZN(n10041) );
  AOI21_X1 U12606 ( .B1(n16515), .B2(n16550), .A(n10030), .ZN(n16518) );
  NAND2_X1 U12607 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  OAI211_X1 U12608 ( .C1(n15350), .C2(n15600), .A(n9847), .B(n15349), .ZN(
        n15351) );
  AND2_X1 U12609 ( .A1(n15348), .A2(n15347), .ZN(n15349) );
  OR2_X1 U12610 ( .A1(n16874), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10149) );
  AOI211_X1 U12611 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n17171), .A(
        n16863), .B(n16862), .ZN(n16866) );
  NAND2_X1 U12612 ( .A1(n17317), .A2(n9869), .ZN(n17287) );
  AND2_X1 U12613 ( .A1(n17317), .A2(n9954), .ZN(n17302) );
  NAND2_X1 U12614 ( .A1(n17431), .A2(n10195), .ZN(n17360) );
  AOI21_X1 U12615 ( .B1(n16688), .B2(n18032), .A(n10136), .ZN(n16693) );
  OR2_X1 U12616 ( .A1(n16691), .A2(n10137), .ZN(n10136) );
  NAND2_X1 U12617 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  NAND2_X1 U12618 ( .A1(n17844), .A2(n18195), .ZN(n9998) );
  AOI21_X1 U12619 ( .B1(n18199), .B2(n18032), .A(n10001), .ZN(n10000) );
  INV_X1 U12620 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18062) );
  NAND2_X1 U12621 ( .A1(n16717), .A2(n16716), .ZN(n16724) );
  NAND2_X1 U12622 ( .A1(n10080), .A2(n10079), .ZN(n16723) );
  NAND2_X1 U12623 ( .A1(n10007), .A2(n10006), .ZN(n18153) );
  INV_X1 U12624 ( .A(n11470), .ZN(n10696) );
  INV_X1 U12625 ( .A(n11601), .ZN(n11579) );
  NOR2_X1 U12626 ( .A1(n15003), .A2(n16490), .ZN(n9840) );
  OR2_X1 U12627 ( .A1(n19476), .A2(n13287), .ZN(n9841) );
  AND2_X1 U12628 ( .A1(n9857), .A2(n10160), .ZN(n9842) );
  INV_X1 U12629 ( .A(n9880), .ZN(n12788) );
  INV_X1 U12630 ( .A(n9880), .ZN(n12736) );
  INV_X1 U12631 ( .A(n10388), .ZN(n14644) );
  INV_X1 U12632 ( .A(n11523), .ZN(n11746) );
  INV_X1 U12633 ( .A(n10425), .ZN(n11373) );
  NAND2_X1 U12634 ( .A1(n10215), .A2(n20398), .ZN(n14082) );
  INV_X1 U12635 ( .A(n10906), .ZN(n14582) );
  INV_X1 U12636 ( .A(n9837), .ZN(n10035) );
  INV_X4 U12637 ( .A(n11860), .ZN(n13885) );
  OR2_X1 U12638 ( .A1(n12346), .A2(n10306), .ZN(n9843) );
  NOR2_X1 U12639 ( .A1(n13935), .A2(n14337), .ZN(n14320) );
  AND2_X1 U12640 ( .A1(n12351), .A2(n10299), .ZN(n9844) );
  AND2_X1 U12641 ( .A1(n19366), .A2(n10404), .ZN(n9845) );
  INV_X2 U12642 ( .A(n10656), .ZN(n10746) );
  INV_X2 U12643 ( .A(n12576), .ZN(n11627) );
  NAND2_X1 U12644 ( .A1(n10625), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10893) );
  OR2_X1 U12645 ( .A1(n16581), .A2(n15343), .ZN(n9847) );
  AND2_X1 U12646 ( .A1(n10299), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9848) );
  INV_X1 U12647 ( .A(n14152), .ZN(n10215) );
  NOR2_X1 U12648 ( .A1(n14984), .A2(n14985), .ZN(n9849) );
  INV_X1 U12649 ( .A(n15934), .ZN(n10090) );
  AND2_X1 U12650 ( .A1(n10383), .A2(n9957), .ZN(n9850) );
  OR2_X1 U12651 ( .A1(n18196), .A2(n16720), .ZN(n9851) );
  OR2_X1 U12652 ( .A1(n10332), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9852) );
  AND2_X1 U12653 ( .A1(n12021), .A2(n9913), .ZN(n9853) );
  NAND2_X1 U12654 ( .A1(n16080), .A2(n9949), .ZN(n9854) );
  NAND2_X1 U12655 ( .A1(n13663), .A2(n10115), .ZN(n15003) );
  AND2_X1 U12656 ( .A1(n10843), .A2(n10820), .ZN(n9855) );
  AND2_X1 U12657 ( .A1(n10285), .A2(n10283), .ZN(n9856) );
  AND2_X1 U12658 ( .A1(n10417), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9857) );
  NAND2_X1 U12659 ( .A1(n12330), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12328) );
  INV_X1 U12660 ( .A(n11918), .ZN(n10235) );
  AND2_X1 U12661 ( .A1(n10295), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9858) );
  AND2_X1 U12662 ( .A1(n11829), .A2(n11787), .ZN(n9859) );
  OR2_X1 U12663 ( .A1(n12480), .A2(n12479), .ZN(n12689) );
  AND2_X1 U12664 ( .A1(n9855), .A2(n10869), .ZN(n9860) );
  AND2_X1 U12665 ( .A1(n10114), .A2(n19379), .ZN(n9861) );
  INV_X1 U12666 ( .A(n11752), .ZN(n15681) );
  AND2_X1 U12667 ( .A1(n17775), .A2(n10163), .ZN(n9862) );
  NAND2_X1 U12668 ( .A1(n12821), .A2(n12820), .ZN(n9863) );
  AOI21_X2 U12669 ( .B1(n15990), .B2(n15989), .A(n18985), .ZN(n18439) );
  AND2_X1 U12670 ( .A1(n10163), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9864) );
  AND2_X1 U12671 ( .A1(n16682), .A2(n10154), .ZN(n9865) );
  AND2_X1 U12672 ( .A1(n9939), .A2(n10280), .ZN(n9866) );
  AND2_X1 U12673 ( .A1(n12623), .A2(n10039), .ZN(n9867) );
  NOR2_X1 U12674 ( .A1(n19208), .A2(n19209), .ZN(n14941) );
  INV_X1 U12675 ( .A(n14941), .ZN(n10102) );
  AND3_X1 U12676 ( .A1(n9952), .A2(n10176), .A3(n10175), .ZN(n9868) );
  AND2_X1 U12677 ( .A1(n9954), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n9869) );
  AND2_X1 U12678 ( .A1(n10167), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n9870) );
  AND2_X1 U12679 ( .A1(n9869), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9871) );
  INV_X2 U12680 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15689) );
  AND2_X2 U12681 ( .A1(n11551), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11762) );
  OR2_X1 U12682 ( .A1(n13959), .A2(n13962), .ZN(n9873) );
  NOR2_X1 U12683 ( .A1(n12351), .A2(n12338), .ZN(n9874) );
  OR2_X1 U12684 ( .A1(n13960), .A2(n13958), .ZN(n9875) );
  OR3_X1 U12685 ( .A1(n13018), .A2(n13017), .A3(n10222), .ZN(n9876) );
  OR2_X1 U12686 ( .A1(n15593), .A2(n15592), .ZN(n9877) );
  NOR2_X1 U12687 ( .A1(n13960), .A2(n13959), .ZN(n13961) );
  OR3_X1 U12688 ( .A1(n14426), .A2(n10207), .A3(n14790), .ZN(n9879) );
  NAND2_X1 U12689 ( .A1(n12922), .A2(n15689), .ZN(n9880) );
  AND2_X1 U12690 ( .A1(n10077), .A2(n18330), .ZN(n9881) );
  NOR2_X1 U12691 ( .A1(n13935), .A2(n10364), .ZN(n14323) );
  NOR2_X1 U12692 ( .A1(n12339), .A2(n19263), .ZN(n12340) );
  NOR2_X1 U12693 ( .A1(n12346), .A2(n10305), .ZN(n12341) );
  NOR2_X1 U12694 ( .A1(n12346), .A2(n21274), .ZN(n12342) );
  AND3_X1 U12695 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12345) );
  INV_X1 U12696 ( .A(n10310), .ZN(n16708) );
  INV_X1 U12697 ( .A(n10034), .ZN(n15533) );
  OR2_X1 U12698 ( .A1(n15309), .A2(n15298), .ZN(n10034) );
  AND2_X1 U12699 ( .A1(n12340), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12337) );
  AND2_X1 U12700 ( .A1(n14674), .A2(n10900), .ZN(n10388) );
  AND4_X1 U12701 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n9882) );
  OR2_X1 U12702 ( .A1(n10332), .A2(n10331), .ZN(n9883) );
  NAND4_X1 U12703 ( .A1(n15204), .A2(n15213), .A3(n12105), .A4(n15221), .ZN(
        n9884) );
  NOR2_X1 U12704 ( .A1(n15669), .A2(n21322), .ZN(n9885) );
  AND2_X1 U12705 ( .A1(n13002), .A2(n9866), .ZN(n9886) );
  OR3_X1 U12706 ( .A1(n13018), .A2(n13017), .A3(n10223), .ZN(n9887) );
  AND2_X1 U12707 ( .A1(n9883), .A2(n9852), .ZN(n9888) );
  NAND2_X1 U12708 ( .A1(n11694), .A2(n11696), .ZN(n11687) );
  INV_X1 U12709 ( .A(n18032), .ZN(n17967) );
  NOR2_X2 U12710 ( .A1(n18139), .A2(n18047), .ZN(n18032) );
  AND2_X1 U12711 ( .A1(n15342), .A2(n16561), .ZN(n9889) );
  AND3_X1 U12712 ( .A1(n13361), .A2(n9765), .A3(n20408), .ZN(n9890) );
  AND2_X1 U12713 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n9891) );
  AND2_X1 U12714 ( .A1(n13861), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11755) );
  INV_X1 U12715 ( .A(n13287), .ZN(n10266) );
  AND3_X1 U12716 ( .A1(n14640), .A2(n10900), .A3(n10387), .ZN(n9892) );
  NAND2_X2 U12717 ( .A1(n9996), .A2(n9994), .ZN(n13263) );
  NOR2_X1 U12718 ( .A1(n10721), .A2(n10379), .ZN(n9893) );
  OR2_X1 U12719 ( .A1(n9873), .A2(n15884), .ZN(n9894) );
  NAND2_X1 U12720 ( .A1(n14293), .A2(n10356), .ZN(n10358) );
  NOR2_X1 U12721 ( .A1(n10914), .A2(n9961), .ZN(n9895) );
  NAND2_X1 U12722 ( .A1(n11687), .A2(n11699), .ZN(n15665) );
  AND2_X1 U12723 ( .A1(n9850), .A2(n10148), .ZN(n9896) );
  AND2_X1 U12724 ( .A1(n10621), .A2(n20424), .ZN(n9897) );
  NAND2_X1 U12725 ( .A1(n11694), .A2(n11695), .ZN(n12665) );
  OR2_X1 U12726 ( .A1(n16908), .A2(n17831), .ZN(n9898) );
  INV_X1 U12727 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21274) );
  NAND2_X1 U12728 ( .A1(n14979), .A2(n12844), .ZN(n12861) );
  INV_X1 U12729 ( .A(n13361), .ZN(n10063) );
  OR2_X1 U12730 ( .A1(n12125), .A2(n15106), .ZN(n9899) );
  INV_X1 U12731 ( .A(n20412), .ZN(n10625) );
  AND2_X2 U12732 ( .A1(n12922), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11832) );
  AND3_X1 U12733 ( .A1(n10020), .A2(n14627), .A3(n16284), .ZN(n9900) );
  OAI211_X1 U12734 ( .C1(n10754), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10721) );
  OR2_X1 U12735 ( .A1(n14689), .A2(n16383), .ZN(n9901) );
  NOR2_X1 U12736 ( .A1(n16877), .A2(n17156), .ZN(n9902) );
  NOR2_X1 U12737 ( .A1(n17905), .A2(n16001), .ZN(n9903) );
  AND2_X1 U12738 ( .A1(n9966), .A2(n10684), .ZN(n9904) );
  AND2_X1 U12739 ( .A1(n10328), .A2(n10140), .ZN(n9905) );
  INV_X1 U12740 ( .A(n10158), .ZN(n10157) );
  NOR2_X1 U12741 ( .A1(n16908), .A2(n17130), .ZN(n10158) );
  AND2_X1 U12742 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9906) );
  INV_X2 U12743 ( .A(n9773), .ZN(n20155) );
  AND2_X1 U12744 ( .A1(n17431), .A2(n10197), .ZN(n9907) );
  OR2_X1 U12745 ( .A1(n12482), .A2(n15119), .ZN(n9908) );
  INV_X1 U12746 ( .A(n16383), .ZN(n16395) );
  OR2_X1 U12747 ( .A1(n13390), .A2(n13381), .ZN(n16383) );
  NOR2_X1 U12748 ( .A1(n13683), .A2(n10400), .ZN(n13742) );
  OR2_X1 U12749 ( .A1(n17498), .A2(n17494), .ZN(n9909) );
  AND2_X1 U12750 ( .A1(n10554), .A2(n10633), .ZN(n9910) );
  AND2_X1 U12751 ( .A1(n17555), .A2(n10167), .ZN(n9911) );
  AND2_X1 U12752 ( .A1(n15995), .A2(n10315), .ZN(n9912) );
  AND2_X1 U12753 ( .A1(n16535), .A2(n16533), .ZN(n9913) );
  AND2_X1 U12754 ( .A1(n12217), .A2(n12216), .ZN(n14933) );
  AND2_X1 U12755 ( .A1(n13663), .A2(n10116), .ZN(n15002) );
  NAND2_X1 U12756 ( .A1(n12351), .A2(n9848), .ZN(n12335) );
  AND2_X1 U12757 ( .A1(n10284), .A2(n9856), .ZN(n9914) );
  OR3_X1 U12758 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17847), .ZN(n9915) );
  INV_X1 U12759 ( .A(n12026), .ZN(n10253) );
  AND2_X1 U12760 ( .A1(n10227), .A2(n15299), .ZN(n9916) );
  AND2_X1 U12761 ( .A1(n12030), .A2(n10340), .ZN(n9917) );
  OR2_X1 U12762 ( .A1(n12506), .A2(n12505), .ZN(n9918) );
  AND2_X1 U12763 ( .A1(n19141), .A2(n15947), .ZN(n9919) );
  AND2_X1 U12764 ( .A1(n13794), .A2(n16594), .ZN(n9920) );
  NAND2_X1 U12765 ( .A1(n12334), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12332) );
  AND2_X1 U12766 ( .A1(n10291), .A2(n10288), .ZN(n9921) );
  OR3_X1 U12767 ( .A1(n14399), .A2(n10214), .A3(n14295), .ZN(n9922) );
  OR3_X1 U12768 ( .A1(n15266), .A2(n14933), .A3(n10218), .ZN(n9923) );
  OR2_X1 U12769 ( .A1(n15003), .A2(n10398), .ZN(n9924) );
  NOR2_X1 U12770 ( .A1(n15063), .A2(n12798), .ZN(n14984) );
  NAND2_X1 U12771 ( .A1(n13663), .A2(n12689), .ZN(n13683) );
  OR3_X1 U12772 ( .A1(n14399), .A2(n10213), .A3(n10214), .ZN(n9925) );
  OR2_X1 U12773 ( .A1(n14426), .A2(n10207), .ZN(n9926) );
  OR2_X1 U12774 ( .A1(n10899), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9927) );
  OAI21_X1 U12775 ( .B1(n14154), .B2(n14613), .A(n11365), .ZN(n14270) );
  AND2_X1 U12776 ( .A1(n20398), .A2(n10552), .ZN(n13128) );
  INV_X1 U12777 ( .A(n13128), .ZN(n10374) );
  AND2_X1 U12778 ( .A1(n9917), .A2(n15607), .ZN(n9928) );
  OR2_X1 U12779 ( .A1(n10752), .A2(n10751), .ZN(n10764) );
  AND2_X1 U12780 ( .A1(n17317), .A2(n9871), .ZN(n9929) );
  INV_X1 U12781 ( .A(n13900), .ZN(n11020) );
  AND2_X1 U12782 ( .A1(n10397), .A2(n12743), .ZN(n9930) );
  AND2_X1 U12783 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n9931) );
  AND4_X1 U12784 ( .A1(n14654), .A2(n14666), .A3(n10901), .A4(n14663), .ZN(
        n9932) );
  NOR2_X1 U12785 ( .A1(n15266), .A2(n15006), .ZN(n10220) );
  OR2_X1 U12786 ( .A1(n10400), .A2(n10399), .ZN(n9933) );
  AND2_X1 U12787 ( .A1(n14101), .A2(n14100), .ZN(n14442) );
  INV_X1 U12788 ( .A(n10361), .ZN(n10360) );
  NAND2_X1 U12789 ( .A1(n14401), .A2(n14404), .ZN(n10361) );
  NAND2_X1 U12790 ( .A1(n12033), .A2(n13885), .ZN(n12122) );
  INV_X1 U12791 ( .A(n12122), .ZN(n10240) );
  NOR2_X1 U12792 ( .A1(n12662), .A2(n10395), .ZN(n9934) );
  AND2_X1 U12793 ( .A1(n9753), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9935) );
  AND2_X1 U12794 ( .A1(n10225), .A2(n13744), .ZN(n9936) );
  AND2_X1 U12795 ( .A1(n10115), .A2(n9930), .ZN(n9937) );
  AND2_X1 U12796 ( .A1(n9842), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9938) );
  INV_X1 U12797 ( .A(n12407), .ZN(n12288) );
  OR2_X1 U12798 ( .A1(n11898), .A2(n11897), .ZN(n12407) );
  AND3_X1 U12799 ( .A1(n12615), .A2(n12614), .A3(n12613), .ZN(n15660) );
  INV_X1 U12800 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19203) );
  INV_X4 U12801 ( .A(n12799), .ZN(n12922) );
  INV_X2 U12802 ( .A(n19356), .ZN(n19385) );
  INV_X2 U12803 ( .A(n17517), .ZN(n17511) );
  NAND2_X1 U12804 ( .A1(n12330), .A2(n9858), .ZN(n12324) );
  INV_X1 U12805 ( .A(n10121), .ZN(n19721) );
  AND2_X1 U12806 ( .A1(n10281), .A2(n10409), .ZN(n9939) );
  XOR2_X1 U12807 ( .A(n12286), .B(n16594), .Z(n9940) );
  INV_X1 U12808 ( .A(n16718), .ZN(n18255) );
  INV_X1 U12809 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10928) );
  AND2_X1 U12810 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9941) );
  AND2_X1 U12811 ( .A1(n10229), .A2(n10228), .ZN(n9942) );
  NOR3_X1 U12812 ( .A1(n16355), .A2(n10204), .A3(n14442), .ZN(n10202) );
  NAND2_X1 U12813 ( .A1(n13676), .A2(n10114), .ZN(n9943) );
  AND2_X1 U12814 ( .A1(n9866), .A2(n15038), .ZN(n9944) );
  INV_X1 U12815 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21322) );
  INV_X1 U12816 ( .A(n10206), .ZN(n14441) );
  NOR2_X1 U12817 ( .A1(n16355), .A2(n10204), .ZN(n10206) );
  INV_X1 U12818 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20114) );
  AND2_X1 U12819 ( .A1(n12330), .A2(n10295), .ZN(n9945) );
  OR2_X1 U12820 ( .A1(n10274), .A2(n10273), .ZN(n9946) );
  INV_X1 U12821 ( .A(n14407), .ZN(n10209) );
  INV_X1 U12822 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10015) );
  OR2_X2 U12823 ( .A1(n18939), .A2(n13960), .ZN(n9947) );
  INV_X1 U12824 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10078) );
  INV_X1 U12825 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10161) );
  INV_X1 U12826 ( .A(n17774), .ZN(n10154) );
  INV_X1 U12827 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10162) );
  AND2_X1 U12828 ( .A1(n17887), .A2(n9857), .ZN(n9948) );
  INV_X1 U12829 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10301) );
  INV_X1 U12830 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10247) );
  INV_X1 U12831 ( .A(n14453), .ZN(n10367) );
  AND2_X1 U12832 ( .A1(n19149), .A2(n9868), .ZN(n9949) );
  INV_X1 U12833 ( .A(n15119), .ZN(n15120) );
  NAND2_X1 U12834 ( .A1(n10420), .A2(n14091), .ZN(n9950) );
  OR2_X1 U12835 ( .A1(n10038), .A2(n10036), .ZN(n9951) );
  AND4_X1 U12836 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n9952) );
  AND2_X1 U12837 ( .A1(n9949), .A2(n10174), .ZN(n9953) );
  AND2_X1 U12838 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .ZN(n9954) );
  OR2_X1 U12839 ( .A1(n12730), .A2(n12729), .ZN(n9955) );
  INV_X1 U12840 ( .A(n15247), .ZN(n10101) );
  AND2_X1 U12841 ( .A1(n10440), .A2(n10436), .ZN(n10787) );
  INV_X1 U12842 ( .A(n10787), .ZN(n10656) );
  AND2_X1 U12843 ( .A1(n21361), .A2(n18151), .ZN(n9956) );
  AND2_X1 U12844 ( .A1(n14818), .A2(n10912), .ZN(n9957) );
  INV_X1 U12845 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10296) );
  INV_X1 U12846 ( .A(n10269), .ZN(n10268) );
  NAND2_X1 U12847 ( .A1(n9959), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10269) );
  AND2_X1 U12848 ( .A1(n9871), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n9958) );
  INV_X1 U12849 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10036) );
  INV_X1 U12850 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10140) );
  AND2_X1 U12851 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9959) );
  INV_X1 U12852 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10169) );
  INV_X1 U12853 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n10168) );
  INV_X1 U12854 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10243) );
  INV_X1 U12855 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10297) );
  INV_X1 U12856 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10304) );
  INV_X1 U12857 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10250) );
  NOR2_X2 U12858 ( .A1(n19490), .A2(n19476), .ZN(n19987) );
  NOR2_X2 U12859 ( .A1(n19490), .A2(n19467), .ZN(n19974) );
  NOR2_X2 U12860 ( .A1(n14560), .A2(n9895), .ZN(n9960) );
  NOR3_X1 U12861 ( .A1(n9753), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14738), .ZN(n9962) );
  NOR2_X2 U12862 ( .A1(n14590), .A2(n14739), .ZN(n10917) );
  NAND3_X1 U12863 ( .A1(n9964), .A2(n9963), .A3(n9966), .ZN(n20495) );
  NAND4_X1 U12864 ( .A1(n9963), .A2(n9904), .A3(n10685), .A4(n9964), .ZN(
        n10736) );
  NAND2_X1 U12865 ( .A1(n9769), .A2(n9965), .ZN(n9964) );
  NOR2_X1 U12866 ( .A1(n10728), .A2(n10682), .ZN(n9965) );
  NAND2_X1 U12867 ( .A1(n10728), .A2(n10682), .ZN(n9966) );
  NAND2_X2 U12868 ( .A1(n9967), .A2(n10632), .ZN(n10685) );
  NAND2_X1 U12869 ( .A1(n10729), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9967) );
  INV_X1 U12870 ( .A(n10683), .ZN(n10728) );
  NAND3_X1 U12871 ( .A1(n13383), .A2(n13215), .A3(n14358), .ZN(n9970) );
  INV_X2 U12872 ( .A(n16044), .ZN(n9971) );
  NAND2_X1 U12873 ( .A1(n13219), .A2(n14152), .ZN(n9972) );
  NAND2_X1 U12874 ( .A1(n16213), .A2(n14697), .ZN(n10071) );
  INV_X2 U12875 ( .A(n10906), .ZN(n10070) );
  NOR2_X4 U12876 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12877 ( .A1(n14857), .A2(n14858), .ZN(n9974) );
  OR2_X1 U12878 ( .A1(n16040), .A2(n9976), .ZN(n9975) );
  NAND2_X1 U12879 ( .A1(n9977), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10257) );
  AOI21_X1 U12880 ( .B1(n9977), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11681), .ZN(n11685) );
  NAND2_X2 U12881 ( .A1(n9982), .A2(n9980), .ZN(n11936) );
  NAND2_X2 U12882 ( .A1(n9982), .A2(n11730), .ZN(n11941) );
  NAND2_X2 U12883 ( .A1(n9982), .A2(n11707), .ZN(n11943) );
  AND2_X2 U12884 ( .A1(n10258), .A2(n10035), .ZN(n9982) );
  NAND4_X1 U12885 ( .A1(n11677), .A2(n10330), .A3(n11696), .A4(n11694), .ZN(
        n9985) );
  XNOR2_X2 U12886 ( .A(n11664), .B(n11665), .ZN(n11696) );
  NAND2_X1 U12887 ( .A1(n11674), .A2(n11673), .ZN(n11677) );
  NAND2_X2 U12888 ( .A1(n9992), .A2(n9990), .ZN(n13287) );
  NAND4_X1 U12889 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11527), .ZN(
        n9991) );
  NAND4_X1 U12890 ( .A1(n11522), .A2(n11521), .A3(n11519), .A4(n11520), .ZN(
        n9993) );
  NAND4_X1 U12891 ( .A1(n11544), .A2(n11547), .A3(n11545), .A4(n11546), .ZN(
        n9995) );
  NAND4_X1 U12892 ( .A1(n11540), .A2(n11539), .A3(n11542), .A4(n11541), .ZN(
        n9997) );
  NAND3_X1 U12893 ( .A1(n17845), .A2(n10000), .A3(n9998), .ZN(P3_U2807) );
  INV_X2 U12894 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19096) );
  NOR2_X2 U12895 ( .A1(n18367), .A2(n19141), .ZN(n18974) );
  NAND3_X1 U12896 ( .A1(n18149), .A2(n18169), .A3(n10010), .ZN(n18159) );
  NAND2_X1 U12897 ( .A1(n10016), .A2(n10017), .ZN(n10757) );
  NAND3_X1 U12898 ( .A1(n10142), .A2(n21027), .A3(n10737), .ZN(n10016) );
  NAND3_X1 U12899 ( .A1(n10020), .A2(n14627), .A3(n10019), .ZN(n10018) );
  NAND2_X2 U12900 ( .A1(n10020), .A2(n14627), .ZN(n16199) );
  INV_X1 U12901 ( .A(n14581), .ZN(n10021) );
  NAND2_X1 U12902 ( .A1(n10796), .A2(n10795), .ZN(n10823) );
  NAND2_X1 U12903 ( .A1(n10824), .A2(n10845), .ZN(n10952) );
  NAND3_X1 U12904 ( .A1(n10554), .A2(n10625), .A3(n10633), .ZN(n13214) );
  NAND2_X1 U12905 ( .A1(n10023), .A2(n19476), .ZN(n11620) );
  INV_X1 U12906 ( .A(n12583), .ZN(n10023) );
  NAND2_X2 U12907 ( .A1(n10025), .A2(n10024), .ZN(n11638) );
  INV_X1 U12908 ( .A(n13825), .ZN(n10029) );
  NAND3_X1 U12909 ( .A1(n10028), .A2(n12299), .A3(n10026), .ZN(n15643) );
  NAND3_X1 U12910 ( .A1(n10270), .A2(n13825), .A3(n10027), .ZN(n10026) );
  NAND3_X1 U12911 ( .A1(n10029), .A2(n10270), .A3(n10271), .ZN(n10028) );
  NOR2_X2 U12912 ( .A1(n15621), .A2(n15610), .ZN(n15587) );
  NAND2_X2 U12913 ( .A1(n16539), .A2(n12308), .ZN(n15622) );
  NAND2_X2 U12914 ( .A1(n10117), .A2(n10035), .ZN(n11731) );
  INV_X1 U12915 ( .A(n15381), .ZN(n10039) );
  AND3_X2 U12916 ( .A1(n11830), .A2(n11788), .A3(n10338), .ZN(n11970) );
  NAND3_X1 U12917 ( .A1(n10041), .A2(n10123), .A3(n10040), .ZN(P2_U2984) );
  NAND3_X1 U12918 ( .A1(n11831), .A2(n12289), .A3(n15119), .ZN(n10042) );
  NAND3_X1 U12919 ( .A1(n11830), .A2(n11788), .A3(n9859), .ZN(n12289) );
  NAND2_X1 U12920 ( .A1(n11788), .A2(n11787), .ZN(n10043) );
  NAND2_X1 U12921 ( .A1(n11830), .A2(n11829), .ZN(n10044) );
  OAI21_X2 U12922 ( .B1(n15252), .B2(n15253), .A(n15211), .ZN(n15244) );
  NAND3_X1 U12923 ( .A1(n11649), .A2(n10050), .A3(n10051), .ZN(n10053) );
  NAND3_X1 U12924 ( .A1(n15538), .A2(n15535), .A3(n15273), .ZN(n10057) );
  NAND2_X1 U12925 ( .A1(n9839), .A2(n9816), .ZN(n11722) );
  NAND3_X1 U12926 ( .A1(n11723), .A2(n9816), .A3(n9839), .ZN(n11725) );
  AND2_X2 U12927 ( .A1(n10430), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10441) );
  NAND3_X1 U12928 ( .A1(n10064), .A2(n10062), .A3(n10061), .ZN(n10065) );
  NAND2_X1 U12929 ( .A1(n9765), .A2(n13361), .ZN(n10061) );
  NAND2_X1 U12930 ( .A1(n13216), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U12931 ( .A1(n13324), .A2(n13361), .ZN(n10064) );
  NAND2_X1 U12932 ( .A1(n10067), .A2(n10069), .ZN(n14608) );
  NAND3_X1 U12933 ( .A1(n10075), .A2(n14654), .A3(n10074), .ZN(n14645) );
  AND2_X1 U12934 ( .A1(n14663), .A2(n10903), .ZN(n10074) );
  AND2_X1 U12935 ( .A1(n14666), .A2(n10901), .ZN(n10075) );
  NAND2_X2 U12936 ( .A1(n18044), .A2(n18009), .ZN(n17979) );
  NAND2_X2 U12937 ( .A1(n9881), .A2(n9788), .ZN(n18044) );
  INV_X2 U12938 ( .A(n17660), .ZN(n15965) );
  AOI21_X1 U12939 ( .B1(n10090), .B2(n18079), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12940 ( .A1(n10081), .A2(n18090), .ZN(n10091) );
  INV_X1 U12941 ( .A(n10087), .ZN(n10081) );
  NAND2_X1 U12942 ( .A1(n10084), .A2(n10082), .ZN(n18063) );
  INV_X1 U12943 ( .A(n18064), .ZN(n10083) );
  OAI21_X1 U12944 ( .B1(n18090), .B2(n10092), .A(n10089), .ZN(n10088) );
  INV_X1 U12945 ( .A(n18079), .ZN(n10092) );
  INV_X4 U12946 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19108) );
  INV_X1 U12947 ( .A(n17805), .ZN(n16007) );
  OR2_X2 U12948 ( .A1(n17805), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10093) );
  AND2_X2 U12949 ( .A1(n17880), .A2(n10094), .ZN(n17905) );
  NAND2_X2 U12950 ( .A1(n17915), .A2(n16004), .ZN(n17880) );
  NAND2_X1 U12951 ( .A1(n11648), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10105) );
  AND2_X1 U12952 ( .A1(n11680), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10107) );
  AND3_X2 U12953 ( .A1(n11660), .A2(n11659), .A3(n10109), .ZN(n11665) );
  NAND3_X1 U12954 ( .A1(n10113), .A2(n10112), .A3(n9863), .ZN(n10111) );
  INV_X1 U12955 ( .A(n13521), .ZN(n12688) );
  AND2_X2 U12956 ( .A1(n13663), .A2(n9937), .ZN(n14991) );
  INV_X1 U12957 ( .A(n11708), .ZN(n10120) );
  INV_X2 U12958 ( .A(n10258), .ZN(n10117) );
  OR2_X2 U12959 ( .A1(n11702), .A2(n10258), .ZN(n19811) );
  XNOR2_X2 U12960 ( .A(n11693), .B(n11692), .ZN(n10258) );
  NAND2_X1 U12961 ( .A1(n15665), .A2(n10117), .ZN(n11700) );
  OAI21_X1 U12962 ( .B1(n10117), .B2(n15660), .A(n10119), .ZN(n10118) );
  NAND2_X1 U12963 ( .A1(n10120), .A2(n10117), .ZN(n19754) );
  NOR2_X1 U12964 ( .A1(n11725), .A2(n10258), .ZN(n10121) );
  NAND2_X1 U12965 ( .A1(n13638), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10122) );
  OR2_X2 U12966 ( .A1(n15354), .A2(n16557), .ZN(n10123) );
  INV_X1 U12967 ( .A(n15312), .ZN(n12046) );
  XNOR2_X1 U12968 ( .A(n10126), .B(n9940), .ZN(n16589) );
  NOR2_X2 U12969 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15671) );
  NOR2_X2 U12970 ( .A1(n15910), .A2(n15952), .ZN(n15935) );
  NAND2_X1 U12972 ( .A1(n17880), .A2(n10328), .ZN(n17827) );
  AND2_X2 U12973 ( .A1(n17880), .A2(n9905), .ZN(n17826) );
  INV_X2 U12974 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19121) );
  NOR2_X1 U12975 ( .A1(n10142), .A2(n20830), .ZN(n13578) );
  NAND2_X2 U12976 ( .A1(n10797), .A2(n13654), .ZN(n13603) );
  NAND2_X1 U12977 ( .A1(n10388), .A2(n10386), .ZN(n10147) );
  NAND3_X1 U12978 ( .A1(n16866), .A2(n16865), .A3(n10149), .ZN(P3_U2641) );
  NOR2_X1 U12979 ( .A1(n16878), .A2(n17774), .ZN(n16877) );
  NAND2_X1 U12980 ( .A1(n10151), .A2(n10153), .ZN(n16867) );
  INV_X1 U12981 ( .A(n16878), .ZN(n10152) );
  NAND2_X1 U12982 ( .A1(n10156), .A2(n10157), .ZN(n16906) );
  NOR2_X1 U12983 ( .A1(n17156), .A2(n10158), .ZN(n10155) );
  INV_X1 U12984 ( .A(n10159), .ZN(n16919) );
  NOR2_X1 U12985 ( .A1(n16960), .A2(n17879), .ZN(n16959) );
  NAND2_X1 U12986 ( .A1(n17317), .A2(n9958), .ZN(n17265) );
  NAND3_X1 U12987 ( .A1(n10191), .A2(n10184), .A3(n14038), .ZN(n10183) );
  NAND3_X1 U12988 ( .A1(n14042), .A2(n10189), .A3(n10186), .ZN(n10185) );
  INV_X1 U12989 ( .A(n10202), .ZN(n14440) );
  NAND3_X1 U12990 ( .A1(n14407), .A2(n14402), .A3(n10208), .ZN(n10207) );
  NAND2_X1 U12991 ( .A1(n9811), .A2(n9773), .ZN(n11637) );
  AND2_X1 U12992 ( .A1(n9812), .A2(n10216), .ZN(n12604) );
  NAND2_X1 U12993 ( .A1(n12604), .A2(n11639), .ZN(n11663) );
  INV_X1 U12994 ( .A(n10220), .ZN(n15005) );
  INV_X1 U12995 ( .A(n12999), .ZN(n10224) );
  NAND3_X1 U12996 ( .A1(n11873), .A2(n11874), .A3(n10233), .ZN(n10232) );
  AND3_X2 U12997 ( .A1(n11873), .A2(n11874), .A3(n10234), .ZN(n12019) );
  OR2_X2 U12998 ( .A1(n12048), .A2(n10240), .ZN(n12047) );
  NOR2_X2 U12999 ( .A1(n12069), .A2(n10241), .ZN(n10244) );
  OR3_X1 U13000 ( .A1(n12069), .A2(P2_EBX_REG_20__SCAN_IN), .A3(n12065), .ZN(
        n12062) );
  OR2_X2 U13001 ( .A1(n10244), .A2(n10240), .ZN(n12106) );
  NOR2_X1 U13002 ( .A1(n12069), .A2(n12065), .ZN(n12089) );
  INV_X1 U13003 ( .A(n10244), .ZN(n12109) );
  NAND3_X1 U13004 ( .A1(n12924), .A2(n12923), .A3(n10245), .ZN(n12935) );
  NOR2_X2 U13005 ( .A1(n12027), .A2(n12026), .ZN(n12033) );
  AOI21_X1 U13006 ( .B1(n12121), .B2(n14982), .A(n10240), .ZN(n10255) );
  NAND2_X1 U13007 ( .A1(n10258), .A2(n12673), .ZN(n12678) );
  NAND3_X1 U13008 ( .A1(n9841), .A2(n11549), .A3(n11550), .ZN(n11616) );
  AND2_X1 U13009 ( .A1(n15163), .A2(n10268), .ZN(n15146) );
  NAND2_X1 U13010 ( .A1(n15163), .A2(n10267), .ZN(n15125) );
  NAND2_X1 U13011 ( .A1(n10275), .A2(n10276), .ZN(n13297) );
  INV_X1 U13012 ( .A(n12399), .ZN(n10275) );
  NOR3_X4 U13013 ( .A1(n9872), .A2(n12633), .A3(n10279), .ZN(n15014) );
  NAND2_X1 U13014 ( .A1(n10289), .A2(n10287), .ZN(n15589) );
  INV_X1 U13015 ( .A(n12344), .ZN(n10293) );
  NAND2_X1 U13016 ( .A1(n10293), .A2(n9906), .ZN(n12343) );
  INV_X1 U13018 ( .A(n12346), .ZN(n10302) );
  NAND2_X1 U13019 ( .A1(n10302), .A2(n10303), .ZN(n12339) );
  NOR2_X2 U13020 ( .A1(n15994), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15995) );
  NAND2_X2 U13021 ( .A1(n18050), .A2(n15940), .ZN(n15994) );
  NAND2_X2 U13022 ( .A1(n18051), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18050) );
  XNOR2_X2 U13023 ( .A(n15939), .B(n10308), .ZN(n18051) );
  NAND2_X1 U13024 ( .A1(n16006), .A2(n21361), .ZN(n10313) );
  NOR3_X1 U13025 ( .A1(n17826), .A2(n10321), .A3(n17905), .ZN(n16003) );
  NAND2_X1 U13026 ( .A1(n17905), .A2(n9788), .ZN(n10325) );
  NAND2_X1 U13027 ( .A1(n11687), .A2(n11667), .ZN(n11693) );
  NAND2_X1 U13028 ( .A1(n15297), .A2(n15294), .ZN(n15285) );
  NAND2_X1 U13029 ( .A1(n10334), .A2(n10333), .ZN(n15297) );
  INV_X1 U13030 ( .A(n15294), .ZN(n10332) );
  NAND2_X1 U13031 ( .A1(n12022), .A2(n9853), .ZN(n10341) );
  CLKBUF_X1 U13032 ( .A(n10341), .Z(n10339) );
  NAND2_X1 U13033 ( .A1(n12022), .A2(n12021), .ZN(n15321) );
  INV_X1 U13034 ( .A(n13730), .ZN(n10345) );
  NAND2_X1 U13035 ( .A1(n13802), .A2(n10343), .ZN(n13900) );
  NAND2_X1 U13036 ( .A1(n13803), .A2(n13802), .ZN(n13901) );
  NAND2_X1 U13037 ( .A1(n14231), .A2(n10349), .ZN(n10346) );
  NAND2_X1 U13038 ( .A1(n14231), .A2(n14232), .ZN(n14220) );
  INV_X1 U13039 ( .A(n10358), .ZN(n14269) );
  NAND2_X1 U13040 ( .A1(n13564), .A2(n13324), .ZN(n10370) );
  NAND2_X1 U13041 ( .A1(n13219), .A2(n10371), .ZN(n13220) );
  INV_X1 U13042 ( .A(n10675), .ZN(n10372) );
  NAND3_X1 U13043 ( .A1(n10376), .A2(n10377), .A3(n10378), .ZN(n20381) );
  NAND2_X1 U13044 ( .A1(n10372), .A2(n10721), .ZN(n10376) );
  NAND3_X1 U13045 ( .A1(n10376), .A2(n10373), .A3(n10378), .ZN(n10681) );
  NAND2_X1 U13046 ( .A1(n10675), .A2(n10674), .ZN(n10718) );
  INV_X1 U13047 ( .A(n10674), .ZN(n10379) );
  NAND3_X1 U13048 ( .A1(n14674), .A2(n10904), .A3(n9892), .ZN(n10380) );
  OAI21_X2 U13049 ( .B1(n13808), .B2(n13807), .A(n10879), .ZN(n16257) );
  NAND2_X2 U13050 ( .A1(n10853), .A2(n10852), .ZN(n13808) );
  NAND2_X1 U13051 ( .A1(n14971), .A2(n10393), .ZN(n10390) );
  NAND3_X1 U13052 ( .A1(n14971), .A2(n10393), .A3(n10392), .ZN(n10391) );
  NAND2_X1 U13053 ( .A1(n14966), .A2(n14965), .ZN(n14964) );
  NAND2_X1 U13054 ( .A1(n9839), .A2(n12673), .ZN(n10396) );
  NAND2_X1 U13055 ( .A1(n10396), .A2(n12659), .ZN(n12663) );
  NAND2_X1 U13056 ( .A1(n10396), .A2(n9934), .ZN(n12664) );
  CLKBUF_X1 U13057 ( .A(n12331), .Z(n12333) );
  XNOR2_X2 U13058 ( .A(n14886), .B(n14885), .ZN(n19390) );
  NOR2_X1 U13059 ( .A1(n19721), .A2(n11724), .ZN(n11728) );
  XNOR2_X1 U13060 ( .A(n12129), .B(n12128), .ZN(n12599) );
  NAND2_X1 U13061 ( .A1(n15155), .A2(n9899), .ZN(n12129) );
  OR2_X2 U13062 ( .A1(n11722), .A2(n11700), .ZN(n19783) );
  INV_X1 U13063 ( .A(n15130), .ZN(n15131) );
  NOR2_X1 U13064 ( .A1(n19312), .A2(n19195), .ZN(n14927) );
  OAI211_X1 U13065 ( .C1(n16480), .C2(n13882), .A(n15129), .B(n15128), .ZN(
        n15130) );
  INV_X1 U13066 ( .A(n13594), .ZN(n10940) );
  NAND2_X1 U13067 ( .A1(n10871), .A2(n10846), .ZN(n10962) );
  INV_X2 U13068 ( .A(n10620), .ZN(n20412) );
  OAI21_X2 U13069 ( .B1(n15429), .B2(n15425), .A(n15426), .ZN(n15194) );
  AOI21_X2 U13070 ( .B1(n9846), .B2(n10405), .A(n9884), .ZN(n15429) );
  AOI21_X1 U13071 ( .B1(n10969), .B2(n11129), .A(n10968), .ZN(n13750) );
  INV_X1 U13072 ( .A(n10962), .ZN(n10969) );
  NAND2_X1 U13073 ( .A1(n15338), .A2(n16550), .ZN(n15129) );
  OAI21_X1 U13074 ( .B1(n13137), .B2(n13140), .A(n13378), .ZN(n10629) );
  CLKBUF_X1 U13075 ( .A(n14307), .Z(n14432) );
  NAND2_X1 U13076 ( .A1(n13214), .A2(n10622), .ZN(n10638) );
  NAND2_X2 U13077 ( .A1(n10712), .A2(n10711), .ZN(n10770) );
  INV_X1 U13078 ( .A(n14993), .ZN(n12765) );
  AND2_X1 U13079 ( .A1(n13324), .A2(n20424), .ZN(n13409) );
  OR2_X1 U13080 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  OAI211_X1 U13081 ( .C1(n11617), .C2(n11616), .A(n9812), .B(n11661), .ZN(
        n12606) );
  INV_X1 U13082 ( .A(n12797), .ZN(n15072) );
  NOR2_X1 U13083 ( .A1(n13028), .A2(n12546), .ZN(n13040) );
  AND2_X1 U13084 ( .A1(n11638), .A2(n19476), .ZN(n11610) );
  NOR2_X1 U13085 ( .A1(n13028), .A2(n16615), .ZN(n19166) );
  INV_X1 U13086 ( .A(n18407), .ZN(n18451) );
  OR3_X1 U13087 ( .A1(n15345), .A2(n15611), .A3(n15335), .ZN(n10403) );
  NOR2_X1 U13088 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10934) );
  INV_X1 U13089 ( .A(n10934), .ZN(n14154) );
  AND2_X1 U13090 ( .A1(n19361), .A2(n19360), .ZN(n10404) );
  AND4_X1 U13091 ( .A1(n15205), .A2(n12091), .A3(n15261), .A4(n15222), .ZN(
        n10405) );
  NAND2_X1 U13092 ( .A1(n14546), .A2(n13405), .ZN(n14553) );
  NAND2_X1 U13093 ( .A1(n11679), .A2(n11678), .ZN(n10406) );
  AND2_X1 U13094 ( .A1(n11512), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10407) );
  INV_X1 U13095 ( .A(n9788), .ZN(n16004) );
  AND3_X1 U13096 ( .A1(n15887), .A2(n15886), .A3(n15885), .ZN(n10408) );
  AND2_X1 U13097 ( .A1(n13022), .A2(n13001), .ZN(n10409) );
  NOR2_X1 U13098 ( .A1(n20833), .A2(n20956), .ZN(n10410) );
  OR2_X1 U13099 ( .A1(n9873), .A2(n15921), .ZN(n10411) );
  OR2_X1 U13100 ( .A1(n16212), .A2(n16361), .ZN(n10412) );
  NOR2_X1 U13101 ( .A1(n13604), .A2(n20382), .ZN(n10413) );
  OR2_X1 U13102 ( .A1(n15657), .A2(n15656), .ZN(n10414) );
  INV_X1 U13103 ( .A(n11751), .ZN(n12368) );
  INV_X1 U13104 ( .A(n20024), .ZN(n19336) );
  INV_X1 U13105 ( .A(n19346), .ZN(n12566) );
  AND2_X1 U13106 ( .A1(n13287), .A2(n12580), .ZN(n10415) );
  OR3_X1 U13107 ( .A1(n20132), .A2(n15656), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16630) );
  AND2_X1 U13108 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10417) );
  AND2_X1 U13109 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10418) );
  INV_X1 U13110 ( .A(n13881), .ZN(n13103) );
  INV_X1 U13111 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21030) );
  AND2_X1 U13112 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10419) );
  OR2_X1 U13113 ( .A1(n14145), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10420) );
  INV_X1 U13114 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20132) );
  INV_X1 U13115 ( .A(n11623), .ZN(n12609) );
  NAND2_X1 U13116 ( .A1(n20302), .A2(n14194), .ZN(n20288) );
  AND2_X1 U13117 ( .A1(n12389), .A2(n9773), .ZN(n10421) );
  NOR2_X1 U13118 ( .A1(n13210), .A2(n13209), .ZN(n10422) );
  OR2_X1 U13119 ( .A1(n13210), .A2(n12393), .ZN(n10423) );
  INV_X1 U13120 ( .A(n12385), .ZN(n12418) );
  NAND3_X2 U13121 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20102), .A3(n19952), 
        .ZN(n13882) );
  OR2_X1 U13122 ( .A1(n19165), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15303) );
  INV_X1 U13123 ( .A(n15303), .ZN(n19326) );
  NOR2_X1 U13124 ( .A1(n20424), .A2(n21030), .ZN(n10963) );
  NOR2_X1 U13125 ( .A1(n19847), .A2(n11726), .ZN(n11727) );
  NAND2_X1 U13126 ( .A1(n9765), .A2(n10620), .ZN(n10621) );
  OR2_X1 U13127 ( .A1(n10592), .A2(n13338), .ZN(n10610) );
  NOR2_X1 U13128 ( .A1(n11728), .A2(n11727), .ZN(n11741) );
  INV_X1 U13129 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11863) );
  NAND2_X1 U13130 ( .A1(n11574), .A2(n11623), .ZN(n11621) );
  OR2_X1 U13131 ( .A1(n14054), .A2(n14055), .ZN(n14047) );
  INV_X1 U13132 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10574) );
  NAND2_X1 U13133 ( .A1(n9755), .A2(n10063), .ZN(n13215) );
  INV_X1 U13134 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U13135 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  OAI211_X1 U13136 ( .C1(n12943), .C2(n19476), .A(n11620), .B(n13287), .ZN(
        n12607) );
  INV_X1 U13137 ( .A(n10585), .ZN(n10582) );
  INV_X1 U13138 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10516) );
  AND2_X1 U13139 ( .A1(n10867), .A2(n10866), .ZN(n10885) );
  OR2_X1 U13140 ( .A1(n10702), .A2(n10701), .ZN(n10762) );
  INV_X1 U13141 ( .A(n15073), .ZN(n12764) );
  OR2_X1 U13142 ( .A1(n11601), .A2(n11715), .ZN(n11555) );
  INV_X1 U13143 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11506) );
  NOR2_X1 U13144 ( .A1(n10608), .A2(n10607), .ZN(n13055) );
  INV_X1 U13145 ( .A(n13902), .ZN(n11001) );
  INV_X1 U13146 ( .A(n11339), .ZN(n11340) );
  INV_X1 U13147 ( .A(n10764), .ZN(n10760) );
  INV_X1 U13148 ( .A(n13564), .ZN(n13233) );
  AOI21_X1 U13149 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20114), .A(
        n11902), .ZN(n12131) );
  OR2_X1 U13150 ( .A1(n15014), .A2(n12541), .ZN(n12542) );
  INV_X1 U13151 ( .A(n16490), .ZN(n12720) );
  OR2_X1 U13152 ( .A1(n12699), .A2(n12698), .ZN(n19353) );
  AOI22_X1 U13153 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U13154 ( .A1(n11593), .A2(n15689), .ZN(n11594) );
  NAND2_X1 U13155 ( .A1(n12133), .A2(n12132), .ZN(n12268) );
  AOI22_X1 U13156 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18963), .B2(n19108), .ZN(
        n14054) );
  NOR2_X1 U13157 ( .A1(n18495), .A2(n17523), .ZN(n18934) );
  NAND2_X1 U13158 ( .A1(n17652), .A2(n15965), .ZN(n15932) );
  NAND2_X1 U13159 ( .A1(n13132), .A2(n13409), .ZN(n13137) );
  NAND2_X1 U13160 ( .A1(n10971), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10976) );
  OR2_X1 U13161 ( .A1(n11499), .A2(n14562), .ZN(n11500) );
  AND2_X1 U13162 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11340), .ZN(
        n11341) );
  NOR2_X1 U13163 ( .A1(n11253), .A2(n16117), .ZN(n11254) );
  AND2_X1 U13164 ( .A1(n14654), .A2(n10908), .ZN(n16226) );
  NAND2_X1 U13165 ( .A1(n9765), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11095) );
  NOR2_X1 U13166 ( .A1(n10976), .A2(n16261), .ZN(n11002) );
  NAND2_X1 U13167 ( .A1(n10955), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10964) );
  INV_X1 U13168 ( .A(n11095), .ZN(n11129) );
  OR2_X1 U13169 ( .A1(n10793), .A2(n10792), .ZN(n10799) );
  INV_X1 U13170 ( .A(n20381), .ZN(n20382) );
  AOI221_X1 U13171 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12131), 
        .C1(n15830), .C2(n12131), .A(n12130), .ZN(n12271) );
  INV_X1 U13172 ( .A(n12986), .ZN(n12227) );
  INV_X2 U13173 ( .A(n12418), .ZN(n14880) );
  AND4_X1 U13174 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11858) );
  OR2_X1 U13175 ( .A1(n19239), .A2(n12099), .ZN(n15283) );
  NAND2_X1 U13176 ( .A1(n13206), .A2(n12673), .ZN(n12667) );
  OR2_X1 U13177 ( .A1(n15665), .A2(n13206), .ZN(n11729) );
  OAI21_X1 U13178 ( .B1(n15790), .B2(n17666), .A(n15789), .ZN(n15799) );
  AND2_X1 U13179 ( .A1(n16979), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16849) );
  INV_X1 U13180 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21364) );
  NAND2_X1 U13181 ( .A1(n16711), .A2(n16669), .ZN(n16649) );
  NOR2_X1 U13182 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9788), .ZN(
        n17903) );
  NOR3_X1 U13183 ( .A1(n18511), .A2(n15794), .A3(n16076), .ZN(n15950) );
  AND2_X1 U13184 ( .A1(n14111), .A2(n14110), .ZN(n14414) );
  INV_X1 U13185 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16179) );
  NOR2_X1 U13186 ( .A1(n14359), .A2(n14152), .ZN(n14173) );
  AND2_X1 U13187 ( .A1(n11213), .A2(n11212), .ZN(n14404) );
  NAND2_X1 U13188 ( .A1(n13368), .A2(n13058), .ZN(n13337) );
  NAND2_X1 U13189 ( .A1(n11341), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11389) );
  AND2_X1 U13190 ( .A1(n16226), .A2(n10910), .ZN(n14820) );
  NAND2_X1 U13191 ( .A1(n11090), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11097) );
  AND2_X1 U13192 ( .A1(n14802), .A2(n13510), .ZN(n16303) );
  OR2_X1 U13193 ( .A1(n13390), .A2(n13386), .ZN(n14783) );
  OR2_X1 U13194 ( .A1(n13390), .A2(n13387), .ZN(n14769) );
  OR2_X1 U13195 ( .A1(n13390), .A2(n16020), .ZN(n14802) );
  AND2_X1 U13196 ( .A1(n20641), .A2(n20640), .ZN(n20670) );
  AND2_X1 U13197 ( .A1(n20683), .A2(n20682), .ZN(n20710) );
  AND2_X1 U13198 ( .A1(n20791), .A2(n20790), .ZN(n20818) );
  OR2_X1 U13199 ( .A1(n20797), .A2(n20796), .ZN(n20825) );
  INV_X1 U13200 ( .A(n20826), .ZN(n20958) );
  AOI21_X1 U13201 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21321), .A(n20544), 
        .ZN(n20966) );
  AND2_X1 U13202 ( .A1(n10619), .A2(n10618), .ZN(n16056) );
  NAND2_X1 U13203 ( .A1(n11662), .A2(n9813), .ZN(n12574) );
  INV_X1 U13204 ( .A(n19336), .ZN(n16419) );
  INV_X1 U13205 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19263) );
  AOI21_X1 U13206 ( .B1(n15665), .B2(n12673), .A(n12669), .ZN(n13284) );
  INV_X1 U13207 ( .A(n12384), .ZN(n12419) );
  OR2_X1 U13208 ( .A1(n13869), .A2(n12941), .ZN(n12942) );
  INV_X1 U13209 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15278) );
  INV_X1 U13210 ( .A(n12673), .ZN(n12253) );
  OR3_X1 U13211 ( .A1(n12100), .A2(n15119), .A3(n15525), .ZN(n15273) );
  OR3_X1 U13212 ( .A1(n19251), .A2(n15119), .A3(n15298), .ZN(n15294) );
  OR2_X1 U13213 ( .A1(n12300), .A2(n12298), .ZN(n12299) );
  INV_X1 U13214 ( .A(n19326), .ZN(n19305) );
  AND2_X1 U13215 ( .A1(n12571), .A2(n12272), .ZN(n16614) );
  INV_X1 U13216 ( .A(n19661), .ZN(n19662) );
  NAND2_X1 U13217 ( .A1(n19504), .A2(n19501), .ZN(n19698) );
  NAND2_X1 U13218 ( .A1(n20117), .A2(n20127), .ZN(n20103) );
  OR2_X1 U13219 ( .A1(n16642), .A2(n13884), .ZN(n19490) );
  NOR2_X1 U13220 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16952), .ZN(n16940) );
  NOR2_X1 U13221 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17042), .ZN(n17029) );
  NOR2_X1 U13222 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17137), .ZN(n17117) );
  INV_X1 U13223 ( .A(n17203), .ZN(n17194) );
  INV_X1 U13224 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17305) );
  INV_X1 U13225 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21224) );
  OAI21_X1 U13226 ( .B1(n17723), .B2(n19143), .A(n18978), .ZN(n17725) );
  NAND2_X1 U13227 ( .A1(n17811), .A2(n10418), .ZN(n17801) );
  NOR2_X1 U13228 ( .A1(n17978), .A2(n18330), .ZN(n18307) );
  INV_X1 U13229 ( .A(n17120), .ZN(n17106) );
  INV_X1 U13230 ( .A(n18278), .ZN(n18206) );
  INV_X1 U13231 ( .A(n18346), .ZN(n18340) );
  INV_X1 U13232 ( .A(n18253), .ZN(n18415) );
  INV_X1 U13233 ( .A(n18947), .ZN(n18923) );
  OR2_X1 U13234 ( .A1(n13243), .A2(n20171), .ZN(n13061) );
  AND2_X1 U13235 ( .A1(n14363), .A2(n14159), .ZN(n20210) );
  INV_X1 U13236 ( .A(n20273), .ZN(n20236) );
  INV_X1 U13237 ( .A(n14540), .ZN(n16192) );
  INV_X1 U13238 ( .A(n14546), .ZN(n16190) );
  AND2_X1 U13239 ( .A1(n13163), .A2(n13162), .ZN(n20306) );
  NOR2_X1 U13240 ( .A1(n21139), .A2(n11276), .ZN(n11314) );
  AND2_X1 U13241 ( .A1(n16268), .A2(n20366), .ZN(n16265) );
  AND3_X1 U13242 ( .A1(n16034), .A2(n13403), .A3(n13368), .ZN(n20369) );
  INV_X1 U13243 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10919) );
  AND2_X1 U13244 ( .A1(n14757), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14751) );
  INV_X1 U13245 ( .A(n16303), .ZN(n16364) );
  NOR2_X1 U13246 ( .A1(n13820), .A2(n16340), .ZN(n16366) );
  NOR2_X1 U13247 ( .A1(n20840), .A2(n16056), .ZN(n21101) );
  OAI22_X1 U13248 ( .A1(n20395), .A2(n20394), .B1(n20543), .B2(n20393), .ZN(
        n20429) );
  INV_X1 U13249 ( .A(n20442), .ZN(n20455) );
  OAI22_X1 U13250 ( .A1(n20465), .A2(n20464), .B1(n20543), .B2(n20606), .ZN(
        n20489) );
  INV_X1 U13251 ( .A(n20529), .ZN(n20522) );
  NOR2_X2 U13252 ( .A1(n20504), .A2(n20796), .ZN(n20570) );
  INV_X1 U13253 ( .A(n20630), .ZN(n20595) );
  OAI22_X1 U13254 ( .A1(n20608), .A2(n20607), .B1(n20606), .B2(n20889), .ZN(
        n20632) );
  INV_X1 U13255 ( .A(n20666), .ZN(n20673) );
  INV_X1 U13256 ( .A(n20677), .ZN(n20713) );
  INV_X1 U13257 ( .A(n20773), .ZN(n20780) );
  NAND2_X1 U13258 ( .A1(n13657), .A2(n13603), .ZN(n20797) );
  INV_X1 U13259 ( .A(n20825), .ZN(n20855) );
  AND2_X1 U13260 ( .A1(n20888), .A2(n10413), .ZN(n20883) );
  INV_X1 U13261 ( .A(n20973), .ZN(n20907) );
  INV_X1 U13262 ( .A(n20994), .ZN(n20925) );
  INV_X1 U13263 ( .A(n20902), .ZN(n20948) );
  AND2_X1 U13264 ( .A1(n20888), .A2(n20636), .ZN(n21021) );
  INV_X1 U13265 ( .A(n20403), .ZN(n20423) );
  INV_X1 U13266 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21043) );
  INV_X1 U13267 ( .A(n21076), .ZN(n21089) );
  NOR2_X1 U13268 ( .A1(n20024), .A2(n9751), .ZN(n19241) );
  OR2_X1 U13269 ( .A1(n19166), .A2(n12552), .ZN(n19341) );
  INV_X1 U13270 ( .A(n19341), .ZN(n19327) );
  NAND2_X1 U13271 ( .A1(n12549), .A2(n12548), .ZN(n19344) );
  OR2_X1 U13272 ( .A1(n12493), .A2(n12492), .ZN(n19361) );
  INV_X1 U13273 ( .A(n12686), .ZN(n19374) );
  OR2_X1 U13274 ( .A1(n12753), .A2(n12752), .ZN(n14994) );
  NAND2_X1 U13275 ( .A1(n13670), .A2(n13831), .ZN(n13830) );
  INV_X1 U13276 ( .A(n14888), .ZN(n13098) );
  INV_X1 U13277 ( .A(n13883), .ZN(n13881) );
  OAI211_X1 U13278 ( .C1(n15600), .C2(n16480), .A(n15336), .B(n10403), .ZN(
        n15337) );
  INV_X1 U13279 ( .A(n16588), .ZN(n16574) );
  NOR2_X1 U13280 ( .A1(n12648), .A2(n16620), .ZN(n15494) );
  NOR2_X1 U13281 ( .A1(n16614), .A2(n20110), .ZN(n15655) );
  OAI21_X1 U13282 ( .B1(n13890), .B2(n13889), .A(n13888), .ZN(n19495) );
  INV_X1 U13283 ( .A(n19532), .ZN(n19524) );
  INV_X1 U13284 ( .A(n19582), .ZN(n19594) );
  NOR2_X1 U13285 ( .A1(n19698), .A2(n20103), .ZN(n19621) );
  AND2_X1 U13286 ( .A1(n19661), .A2(n19602), .ZN(n19650) );
  NOR2_X1 U13287 ( .A1(n19698), .A2(n19882), .ZN(n19680) );
  NOR2_X1 U13288 ( .A1(n19698), .A2(n19949), .ZN(n19741) );
  INV_X1 U13289 ( .A(n19500), .ZN(n19750) );
  AND2_X1 U13290 ( .A1(n19815), .A2(n19813), .ZN(n19837) );
  NOR2_X1 U13291 ( .A1(n19912), .A2(n19882), .ZN(n19907) );
  NOR2_X2 U13292 ( .A1(n13883), .A2(n13882), .ZN(n19494) );
  INV_X1 U13293 ( .A(n19820), .ZN(n19963) );
  INV_X1 U13294 ( .A(n19895), .ZN(n19983) );
  OAI22_X1 U13295 ( .A1(n19484), .A2(n19488), .B1(n19483), .B2(n19487), .ZN(
        n20003) );
  NOR2_X2 U13296 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13884), .ZN(n19952) );
  INV_X1 U13297 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20045) );
  NOR2_X1 U13298 ( .A1(n18985), .A2(n18921), .ZN(n17724) );
  NOR2_X1 U13299 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16975), .ZN(n16956) );
  NOR2_X1 U13300 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17064), .ZN(n17047) );
  NOR2_X1 U13301 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17089), .ZN(n17073) );
  NOR2_X1 U13302 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17109), .ZN(n17096) );
  AOI211_X2 U13303 ( .C1(n18990), .C2(n18982), .A(n19162), .B(n17145), .ZN(
        n17186) );
  INV_X1 U13304 ( .A(n17392), .ZN(n17411) );
  INV_X1 U13305 ( .A(n21455), .ZN(n17760) );
  NOR2_X1 U13306 ( .A1(n19141), .A2(n17752), .ZN(n17762) );
  NOR2_X1 U13307 ( .A1(n17853), .A2(n16846), .ZN(n17839) );
  INV_X1 U13308 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18066) );
  INV_X1 U13309 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18128) );
  AND2_X1 U13310 ( .A1(n18207), .A2(n15980), .ZN(n16714) );
  NOR2_X1 U13311 ( .A1(n18451), .A2(n17780), .ZN(n16716) );
  INV_X1 U13312 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21226) );
  NOR2_X1 U13313 ( .A1(n18415), .A2(n18254), .ZN(n18320) );
  INV_X1 U13314 ( .A(n18440), .ZN(n18388) );
  INV_X1 U13315 ( .A(n18407), .ZN(n18446) );
  NAND2_X1 U13316 ( .A1(n19146), .A2(n18477), .ZN(n18516) );
  INV_X1 U13317 ( .A(n19102), .ZN(n19115) );
  INV_X1 U13318 ( .A(n18618), .ZN(n18621) );
  INV_X1 U13319 ( .A(n18695), .ZN(n18720) );
  INV_X1 U13320 ( .A(n18866), .ZN(n18798) );
  NAND2_X2 U13321 ( .A1(n12977), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20379)
         );
  OAI21_X1 U13322 ( .B1(n12952), .B2(n12951), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13883) );
  NOR2_X1 U13323 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12980), .ZN(n16792)
         );
  INV_X1 U13324 ( .A(n21117), .ZN(n14359) );
  INV_X1 U13325 ( .A(n20271), .ZN(n20240) );
  INV_X1 U13326 ( .A(n20306), .ZN(n20334) );
  INV_X1 U13327 ( .A(n20360), .ZN(n13453) );
  OAI21_X1 U13328 ( .B1(n14447), .B2(n14325), .A(n14324), .ZN(n14673) );
  INV_X1 U13329 ( .A(n16265), .ZN(n16254) );
  OR2_X1 U13330 ( .A1(n20369), .A2(n11497), .ZN(n16268) );
  OR2_X1 U13331 ( .A1(n13390), .A2(n13377), .ZN(n16319) );
  NAND2_X1 U13332 ( .A1(n20494), .A2(n10413), .ZN(n20442) );
  NAND2_X1 U13333 ( .A1(n20494), .A2(n20860), .ZN(n20487) );
  NAND2_X1 U13334 ( .A1(n20494), .A2(n20887), .ZN(n20529) );
  AOI22_X1 U13335 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20508), .B1(n20506), 
        .B2(n20503), .ZN(n20534) );
  NAND2_X1 U13336 ( .A1(n20637), .A2(n10413), .ZN(n20599) );
  NAND2_X1 U13337 ( .A1(n20637), .A2(n20887), .ZN(n20666) );
  NAND2_X1 U13338 ( .A1(n20678), .A2(n10413), .ZN(n20744) );
  AOI22_X1 U13339 ( .A1(n20753), .A2(n20751), .B1(n20749), .B2(n20748), .ZN(
        n20784) );
  OR2_X1 U13340 ( .A1(n20797), .A2(n20745), .ZN(n20824) );
  AOI22_X1 U13341 ( .A1(n20838), .A2(n20834), .B1(n20832), .B2(n20835), .ZN(
        n20859) );
  NAND2_X1 U13342 ( .A1(n20888), .A2(n20860), .ZN(n20902) );
  NAND2_X1 U13343 ( .A1(n20888), .A2(n20887), .ZN(n21025) );
  INV_X1 U13344 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20840) );
  INV_X1 U13345 ( .A(n21099), .ZN(n21032) );
  AND2_X1 U13346 ( .A1(n21043), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21116) );
  OR2_X1 U13347 ( .A1(n12313), .A2(n9813), .ZN(n13038) );
  AND2_X1 U13348 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  INV_X1 U13349 ( .A(n19344), .ZN(n19324) );
  INV_X1 U13350 ( .A(n19339), .ZN(n19306) );
  AND2_X1 U13351 ( .A1(n13286), .A2(n20165), .ZN(n19356) );
  XNOR2_X1 U13352 ( .A(n13309), .B(n13312), .ZN(n20117) );
  INV_X1 U13353 ( .A(n19419), .ZN(n15094) );
  INV_X1 U13354 ( .A(n19392), .ZN(n19400) );
  INV_X1 U13355 ( .A(n19429), .ZN(n19460) );
  CLKBUF_X1 U13356 ( .A(n13101), .Z(n13126) );
  NAND2_X1 U13357 ( .A1(n13040), .A2(n16624), .ZN(n14888) );
  INV_X1 U13358 ( .A(n16549), .ZN(n16557) );
  INV_X1 U13359 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16532) );
  AND2_X1 U13360 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  INV_X1 U13361 ( .A(n16592), .ZN(n15632) );
  OR2_X1 U13362 ( .A1(n12648), .A2(n12647), .ZN(n16588) );
  INV_X1 U13363 ( .A(n15498), .ZN(n16583) );
  INV_X1 U13364 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13899) );
  AOI211_X2 U13365 ( .C1(n13880), .C2(n13889), .A(n13879), .B(n19917), .ZN(
        n19499) );
  INV_X1 U13366 ( .A(n19554), .ZN(n19562) );
  AND2_X1 U13367 ( .A1(n19569), .A2(n19568), .ZN(n19582) );
  INV_X1 U13368 ( .A(n19589), .ZN(n19597) );
  INV_X1 U13369 ( .A(n19621), .ZN(n19629) );
  INV_X1 U13370 ( .A(n19650), .ZN(n19658) );
  INV_X1 U13371 ( .A(n19680), .ZN(n19688) );
  INV_X1 U13372 ( .A(n19711), .ZN(n19718) );
  INV_X1 U13373 ( .A(n19741), .ZN(n19749) );
  OR2_X1 U13374 ( .A1(n19912), .A2(n19750), .ZN(n19773) );
  INV_X1 U13375 ( .A(n19800), .ZN(n19808) );
  INV_X1 U13376 ( .A(n20003), .ZN(n19835) );
  INV_X1 U13377 ( .A(n19996), .ZN(n19864) );
  INV_X1 U13378 ( .A(n19907), .ZN(n19904) );
  AOI211_X2 U13379 ( .C1(n19920), .C2(n19923), .A(n19918), .B(n19917), .ZN(
        n19947) );
  INV_X1 U13380 ( .A(n20100), .ZN(n20027) );
  NAND2_X1 U13381 ( .A1(n19162), .A2(n17666), .ZN(n19160) );
  INV_X1 U13382 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19146) );
  NAND2_X1 U13383 ( .A1(n19014), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19155) );
  INV_X1 U13384 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17876) );
  INV_X1 U13385 ( .A(n17204), .ZN(n17161) );
  NAND2_X1 U13386 ( .A1(n17205), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17187) );
  INV_X1 U13387 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21348) );
  AND2_X1 U13388 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17614), .ZN(n17617) );
  NOR4_X1 U13389 ( .A1(n17625), .A2(n9854), .A3(n17704), .A4(n17706), .ZN(
        n17628) );
  NAND2_X1 U13390 ( .A1(n18949), .A2(n17607), .ZN(n17662) );
  NAND2_X1 U13391 ( .A1(n17693), .A2(n17666), .ZN(n17691) );
  INV_X1 U13392 ( .A(n17693), .ZN(n17722) );
  INV_X1 U13393 ( .A(n17767), .ZN(n17744) );
  INV_X1 U13394 ( .A(n18045), .ZN(n18139) );
  OR3_X1 U13395 ( .A1(n16721), .A2(n18302), .A3(n17784), .ZN(n16722) );
  INV_X1 U13396 ( .A(n18439), .ZN(n18457) );
  INV_X1 U13397 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18242) );
  NAND2_X1 U13398 ( .A1(n18046), .A2(n18454), .ZN(n18302) );
  NAND2_X1 U13399 ( .A1(n18407), .A2(n18457), .ZN(n18440) );
  INV_X1 U13400 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18963) );
  NOR2_X1 U13401 ( .A1(n18478), .A2(n15822), .ZN(n19122) );
  INV_X1 U13402 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18705) );
  INV_X1 U13403 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21319) );
  INV_X1 U13404 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n21197) );
  INV_X1 U13405 ( .A(n18862), .ZN(n18834) );
  INV_X1 U13406 ( .A(n18835), .ZN(n18876) );
  INV_X1 U13407 ( .A(n18846), .ZN(n18900) );
  INV_X1 U13408 ( .A(n17157), .ZN(n18993) );
  INV_X1 U13409 ( .A(n19088), .ZN(n18997) );
  INV_X1 U13410 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19014) );
  AND2_X2 U13411 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U13412 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U13413 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10428) );
  NAND2_X1 U13414 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13415 ( .A1(n11448), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10426) );
  NAND4_X1 U13416 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  INV_X1 U13417 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U13418 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13419 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10431) );
  OAI211_X1 U13420 ( .C1(n10544), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        n10434) );
  AOI22_X1 U13421 ( .A1(n10505), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10787), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13422 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10445) );
  AND2_X2 U13423 ( .A1(n10441), .A2(n10437), .ZN(n11023) );
  AOI22_X1 U13424 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13425 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9819), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10443) );
  INV_X2 U13426 ( .A(n11371), .ZN(n11473) );
  AOI22_X1 U13427 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U13428 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13429 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10450) );
  NAND2_X1 U13430 ( .A1(n11448), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10449) );
  NAND4_X1 U13431 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10456) );
  NAND2_X1 U13432 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13433 ( .A1(n9790), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10453) );
  OAI211_X1 U13434 ( .C1(n10544), .C2(n11445), .A(n10454), .B(n10453), .ZN(
        n10455) );
  AOI22_X1 U13435 ( .A1(n10505), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10787), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13436 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13437 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13438 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9820), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13439 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U13440 ( .A1(n9794), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13441 ( .A1(n10425), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U13442 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13443 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13444 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13445 ( .A1(n11266), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13446 ( .A1(n9819), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13447 ( .A1(n10787), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10474) );
  NAND2_X1 U13448 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13449 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13450 ( .A1(n10491), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10471) );
  INV_X1 U13451 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10477) );
  NAND2_X1 U13452 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10476) );
  NAND2_X1 U13453 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10475) );
  OAI211_X1 U13454 ( .C1(n10544), .C2(n10477), .A(n10476), .B(n10475), .ZN(
        n10478) );
  INV_X1 U13455 ( .A(n10478), .ZN(n10479) );
  AOI22_X1 U13456 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13457 ( .A1(n9794), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10485) );
  NAND2_X1 U13458 ( .A1(n10425), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10484) );
  NAND2_X1 U13459 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10483) );
  NAND2_X1 U13460 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13461 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10489) );
  NAND2_X1 U13462 ( .A1(n9817), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13463 ( .A1(n9819), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10487) );
  NAND2_X1 U13464 ( .A1(n10787), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13465 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10494) );
  NAND2_X1 U13466 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10493) );
  NAND2_X1 U13467 ( .A1(n10491), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10492) );
  INV_X1 U13468 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13469 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10498) );
  NAND2_X1 U13470 ( .A1(n10661), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10497) );
  OAI211_X1 U13471 ( .C1(n10544), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n10500) );
  INV_X1 U13472 ( .A(n10500), .ZN(n10501) );
  AOI22_X1 U13473 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10787), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13474 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13475 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13476 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9819), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13477 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13478 ( .A1(n9794), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10512) );
  NAND2_X1 U13479 ( .A1(n10425), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10511) );
  NAND2_X1 U13480 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10510) );
  NAND4_X1 U13481 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10518) );
  NAND2_X1 U13482 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10515) );
  NAND2_X1 U13483 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10514) );
  AND2_X4 U13484 ( .A1(n10520), .A2(n10519), .ZN(n14152) );
  AOI22_X1 U13485 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10787), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13486 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13487 ( .A1(n11023), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13488 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9819), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13489 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U13490 ( .A1(n9794), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10528) );
  NAND2_X1 U13491 ( .A1(n10425), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U13492 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10526) );
  NAND4_X1 U13493 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10533) );
  INV_X1 U13494 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U13495 ( .A1(n10696), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10531) );
  NAND2_X1 U13496 ( .A1(n10661), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10530) );
  OAI211_X1 U13497 ( .C1(n10544), .C2(n11349), .A(n10531), .B(n10530), .ZN(
        n10532) );
  NOR2_X1 U13498 ( .A1(n10533), .A2(n10532), .ZN(n10534) );
  AND2_X2 U13499 ( .A1(n10535), .A2(n10534), .ZN(n13361) );
  AOI22_X1 U13500 ( .A1(n9802), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9790), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13501 ( .A1(n9796), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13502 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11266), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13503 ( .A1(n10505), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10425), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13504 ( .A1(n9814), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U13505 ( .A1(n10461), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13506 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10542) );
  NAND2_X1 U13507 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10541) );
  NAND2_X1 U13508 ( .A1(n9786), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10540) );
  NAND2_X1 U13509 ( .A1(n9794), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10546) );
  INV_X1 U13510 ( .A(n9760), .ZN(n11007) );
  NAND2_X1 U13511 ( .A1(n10496), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10545) );
  NAND2_X1 U13512 ( .A1(n13361), .A2(n20408), .ZN(n10551) );
  AOI21_X1 U13513 ( .B1(n10622), .B2(n14152), .A(n10551), .ZN(n10555) );
  NAND2_X1 U13514 ( .A1(n13216), .A2(n9765), .ZN(n10554) );
  NAND2_X1 U13515 ( .A1(n13324), .A2(n10623), .ZN(n10553) );
  NAND2_X1 U13516 ( .A1(n10555), .A2(n9910), .ZN(n13249) );
  INV_X1 U13517 ( .A(n13216), .ZN(n10588) );
  NOR2_X1 U13518 ( .A1(n13249), .A2(n10588), .ZN(n16034) );
  AOI22_X1 U13519 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10505), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13520 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10661), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13521 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9817), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13522 ( .A1(n10787), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10425), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13523 ( .A1(n10491), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13524 ( .A1(n11448), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13525 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10562) );
  NAND2_X1 U13526 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10561) );
  NAND2_X1 U13527 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U13528 ( .A1(n10525), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13529 ( .A1(n10496), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10564) );
  NAND2_X4 U13530 ( .A1(n10569), .A2(n10568), .ZN(n20398) );
  XNOR2_X1 U13531 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U13532 ( .A1(n21321), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13533 ( .A1(n10581), .A2(n10582), .ZN(n10571) );
  NAND2_X1 U13534 ( .A1(n20957), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U13535 ( .A1(n10571), .A2(n10570), .ZN(n10596) );
  XNOR2_X1 U13536 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13537 ( .A1(n10596), .A2(n10595), .ZN(n10573) );
  NAND2_X1 U13538 ( .A1(n20679), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10572) );
  NAND2_X1 U13539 ( .A1(n10573), .A2(n10572), .ZN(n10580) );
  MUX2_X1 U13540 ( .A(n10574), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10579) );
  NAND2_X1 U13541 ( .A1(n10580), .A2(n10579), .ZN(n10576) );
  NAND2_X1 U13542 ( .A1(n10574), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10575) );
  INV_X1 U13543 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16406) );
  NOR2_X1 U13544 ( .A1(n16406), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13545 ( .A1(n10606), .A2(n13057), .ZN(n10619) );
  NAND2_X1 U13546 ( .A1(n13057), .A2(n10881), .ZN(n10617) );
  XNOR2_X1 U13547 ( .A(n10580), .B(n10579), .ZN(n13054) );
  XNOR2_X1 U13548 ( .A(n10582), .B(n10581), .ZN(n13052) );
  NAND2_X1 U13549 ( .A1(n10881), .A2(n20398), .ZN(n10584) );
  NAND2_X1 U13550 ( .A1(n13324), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13551 ( .A1(n10584), .A2(n10583), .ZN(n10592) );
  NOR2_X1 U13552 ( .A1(n13052), .A2(n10592), .ZN(n10591) );
  INV_X1 U13553 ( .A(n10881), .ZN(n10602) );
  OAI21_X1 U13554 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21321), .A(
        n10585), .ZN(n10586) );
  NOR2_X1 U13555 ( .A1(n10602), .A2(n10586), .ZN(n10590) );
  OAI21_X1 U13556 ( .B1(n14152), .B2(n10552), .A(n13338), .ZN(n10601) );
  INV_X1 U13557 ( .A(n10586), .ZN(n10587) );
  OAI211_X1 U13558 ( .C1(n14152), .C2(n10588), .A(n10601), .B(n10587), .ZN(
        n10589) );
  OAI21_X1 U13559 ( .B1(n10606), .B2(n10590), .A(n10589), .ZN(n10593) );
  NAND2_X1 U13560 ( .A1(n10591), .A2(n10593), .ZN(n10600) );
  INV_X1 U13561 ( .A(n10592), .ZN(n10594) );
  OAI211_X1 U13562 ( .C1(n10594), .C2(n10593), .A(n13052), .B(n10610), .ZN(
        n10599) );
  XNOR2_X1 U13563 ( .A(n10596), .B(n10595), .ZN(n13053) );
  NAND2_X1 U13564 ( .A1(n10880), .A2(n13053), .ZN(n10597) );
  OAI211_X1 U13565 ( .C1(n10602), .C2(n13053), .A(n10597), .B(n10601), .ZN(
        n10598) );
  NAND3_X1 U13566 ( .A1(n10600), .A2(n10599), .A3(n10598), .ZN(n10604) );
  AOI22_X1 U13567 ( .A1(n10754), .A2(n13054), .B1(n10604), .B2(n10603), .ZN(
        n10605) );
  AOI21_X1 U13568 ( .B1(n10606), .B2(n13054), .A(n10605), .ZN(n10614) );
  INV_X1 U13569 ( .A(n13055), .ZN(n10609) );
  NOR2_X1 U13570 ( .A1(n10880), .A2(n10609), .ZN(n10613) );
  INV_X1 U13571 ( .A(n10610), .ZN(n10611) );
  NAND3_X1 U13572 ( .A1(n10880), .A2(n10611), .A3(n13055), .ZN(n10612) );
  OAI21_X1 U13573 ( .B1(n10614), .B2(n10613), .A(n10612), .ZN(n10615) );
  AOI21_X1 U13574 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21027), .A(
        n10615), .ZN(n10616) );
  NAND2_X1 U13575 ( .A1(n10617), .A2(n10616), .ZN(n10618) );
  INV_X1 U13576 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13577 ( .A1(n13216), .A2(n14152), .ZN(n10624) );
  NAND2_X1 U13578 ( .A1(n13051), .A2(n13338), .ZN(n13226) );
  NAND2_X1 U13579 ( .A1(n13246), .A2(n14143), .ZN(n10626) );
  NAND2_X1 U13580 ( .A1(n13226), .A2(n10626), .ZN(n13376) );
  AND2_X1 U13581 ( .A1(n9755), .A2(n10625), .ZN(n10627) );
  XNOR2_X1 U13582 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13140) );
  INV_X1 U13583 ( .A(n20408), .ZN(n10628) );
  OAI21_X1 U13584 ( .B1(n13376), .B2(n10629), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10683) );
  OR2_X2 U13585 ( .A1(n14152), .A2(n20398), .ZN(n16044) );
  NAND2_X1 U13586 ( .A1(n13216), .A2(n14149), .ZN(n13383) );
  NAND2_X1 U13587 ( .A1(n14152), .A2(n20398), .ZN(n14358) );
  MUX2_X1 U13588 ( .A(n11501), .B(n16053), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10632) );
  NAND2_X1 U13589 ( .A1(n13564), .A2(n9765), .ZN(n13382) );
  AND2_X1 U13590 ( .A1(n13229), .A2(n14208), .ZN(n13064) );
  OAI21_X1 U13591 ( .B1(n13324), .B2(n10623), .A(n20408), .ZN(n10635) );
  INV_X1 U13592 ( .A(n10633), .ZN(n10634) );
  AOI22_X1 U13593 ( .A1(n13064), .A2(n10635), .B1(n9971), .B2(n10634), .ZN(
        n10636) );
  OAI211_X1 U13594 ( .C1(n10638), .C2(n13338), .A(n10637), .B(n10636), .ZN(
        n10639) );
  INV_X1 U13595 ( .A(n10639), .ZN(n10640) );
  NAND2_X1 U13596 ( .A1(n10641), .A2(n10640), .ZN(n10684) );
  INV_X1 U13597 ( .A(n10684), .ZN(n10642) );
  NAND2_X1 U13598 ( .A1(n20496), .A2(n21027), .ZN(n10675) );
  INV_X1 U13599 ( .A(n10893), .ZN(n10673) );
  INV_X1 U13600 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U13601 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10644) );
  NAND2_X1 U13602 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10643) );
  OAI211_X1 U13603 ( .C1(n9760), .C2(n11469), .A(n10644), .B(n10643), .ZN(
        n10645) );
  INV_X1 U13604 ( .A(n10645), .ZN(n10649) );
  AOI22_X1 U13605 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13606 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13607 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10646) );
  NAND4_X1 U13608 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10655) );
  AOI22_X1 U13609 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13610 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13611 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13612 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10650) );
  NAND4_X1 U13613 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10654) );
  AOI22_X1 U13614 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13615 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13616 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13617 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13618 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U13619 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10665) );
  NAND2_X1 U13620 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U13621 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10663) );
  NAND2_X1 U13622 ( .A1(n9798), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10662) );
  AND4_X1 U13623 ( .A1(n10665), .A2(n10664), .A3(n10663), .A4(n10662), .ZN(
        n10668) );
  NAND2_X1 U13624 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10667) );
  NAND2_X1 U13625 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10666) );
  XNOR2_X1 U13626 ( .A(n10719), .B(n10763), .ZN(n10672) );
  NAND2_X1 U13627 ( .A1(n10673), .A2(n10672), .ZN(n10674) );
  INV_X1 U13628 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10678) );
  AOI21_X1 U13629 ( .B1(n14152), .B2(n10763), .A(n21027), .ZN(n10677) );
  NAND2_X1 U13630 ( .A1(n10625), .A2(n10896), .ZN(n10676) );
  NAND2_X1 U13631 ( .A1(n14152), .A2(n20408), .ZN(n10766) );
  OAI21_X1 U13632 ( .B1(n16044), .B2(n10763), .A(n10766), .ZN(n10679) );
  INV_X1 U13633 ( .A(n10679), .ZN(n10680) );
  NAND2_X1 U13634 ( .A1(n10681), .A2(n10680), .ZN(n13355) );
  NAND2_X2 U13635 ( .A1(n13355), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13356) );
  NAND2_X1 U13636 ( .A1(n20957), .A2(n21321), .ZN(n20833) );
  NAND2_X1 U13637 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U13638 ( .A1(n20833), .A2(n10773), .ZN(n20747) );
  OR2_X1 U13639 ( .A1(n16053), .A2(n20957), .ZN(n10726) );
  OAI21_X1 U13640 ( .B1(n11501), .B2(n20747), .A(n10726), .ZN(n10682) );
  NAND2_X2 U13641 ( .A1(n10736), .A2(n20861), .ZN(n14186) );
  INV_X1 U13642 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13643 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10688) );
  NAND2_X1 U13644 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10687) );
  OAI211_X1 U13645 ( .C1(n9760), .C2(n10689), .A(n10688), .B(n10687), .ZN(
        n10690) );
  INV_X1 U13646 ( .A(n10690), .ZN(n10694) );
  AOI22_X1 U13647 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13648 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13649 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10691) );
  NAND4_X1 U13650 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10702) );
  AOI22_X1 U13651 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13652 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13653 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13654 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U13655 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  INV_X1 U13656 ( .A(n10717), .ZN(n10704) );
  XNOR2_X1 U13657 ( .A(n10713), .B(n10763), .ZN(n10706) );
  NAND2_X1 U13658 ( .A1(n13361), .A2(n10552), .ZN(n10705) );
  AOI21_X1 U13659 ( .B1(n9971), .B2(n10706), .A(n10705), .ZN(n10707) );
  NAND2_X1 U13660 ( .A1(n10708), .A2(n10707), .ZN(n10709) );
  NAND2_X1 U13661 ( .A1(n13509), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10712) );
  INV_X1 U13662 ( .A(n10709), .ZN(n10710) );
  OR2_X1 U13663 ( .A1(n13356), .A2(n10710), .ZN(n10711) );
  INV_X1 U13664 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U13665 ( .A1(n10880), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10716) );
  OR2_X1 U13666 ( .A1(n10896), .A2(n10893), .ZN(n10715) );
  OR2_X1 U13667 ( .A1(n10755), .A2(n10713), .ZN(n10714) );
  NOR2_X1 U13668 ( .A1(n10893), .A2(n10719), .ZN(n10720) );
  INV_X1 U13669 ( .A(n10722), .ZN(n10723) );
  NAND2_X1 U13670 ( .A1(n10725), .A2(n10724), .ZN(n10758) );
  NAND2_X1 U13671 ( .A1(n10726), .A2(n10015), .ZN(n10727) );
  NAND2_X1 U13672 ( .A1(n10728), .A2(n10727), .ZN(n10734) );
  NOR2_X1 U13673 ( .A1(n16053), .A2(n20679), .ZN(n10730) );
  INV_X1 U13674 ( .A(n11501), .ZN(n10776) );
  XNOR2_X1 U13675 ( .A(n10773), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20392) );
  NAND2_X1 U13676 ( .A1(n10776), .A2(n20392), .ZN(n10733) );
  NAND2_X1 U13677 ( .A1(n10735), .A2(n10733), .ZN(n10731) );
  NAND4_X1 U13678 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n10737) );
  INV_X1 U13679 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13680 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13681 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10738) );
  OAI211_X1 U13682 ( .C1(n9760), .C2(n10740), .A(n10739), .B(n10738), .ZN(
        n10741) );
  INV_X1 U13683 ( .A(n10741), .ZN(n10745) );
  AOI22_X1 U13684 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13685 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13686 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10742) );
  NAND4_X1 U13687 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10752) );
  AOI22_X1 U13688 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13689 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13690 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13691 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10747) );
  NAND4_X1 U13692 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10751) );
  INV_X1 U13693 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10753) );
  OAI22_X1 U13694 ( .A1(n10760), .A2(n10755), .B1(n10754), .B2(n10753), .ZN(
        n10756) );
  XNOR2_X1 U13695 ( .A(n10757), .B(n10756), .ZN(n10759) );
  NAND2_X1 U13696 ( .A1(n10758), .A2(n10759), .ZN(n13654) );
  NAND2_X1 U13697 ( .A1(n10763), .A2(n10762), .ZN(n10761) );
  NAND2_X1 U13698 ( .A1(n10761), .A2(n10760), .ZN(n10798) );
  NAND3_X1 U13699 ( .A1(n10764), .A2(n10763), .A3(n10762), .ZN(n10765) );
  NAND2_X1 U13700 ( .A1(n10798), .A2(n10765), .ZN(n10768) );
  INV_X1 U13701 ( .A(n10766), .ZN(n10767) );
  AOI21_X1 U13702 ( .B1(n9971), .B2(n10768), .A(n10767), .ZN(n10769) );
  NAND2_X1 U13703 ( .A1(n10770), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10771) );
  NAND2_X2 U13704 ( .A1(n10772), .A2(n10771), .ZN(n10801) );
  INV_X1 U13705 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13725) );
  INV_X1 U13706 ( .A(n10797), .ZN(n10796) );
  NAND2_X1 U13707 ( .A1(n10729), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10778) );
  OAI21_X1 U13708 ( .B1(n10773), .B2(n20679), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10775) );
  INV_X1 U13709 ( .A(n10773), .ZN(n20954) );
  NAND2_X1 U13710 ( .A1(n10574), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20600) );
  INV_X1 U13711 ( .A(n20600), .ZN(n10774) );
  NAND2_X1 U13712 ( .A1(n20954), .A2(n10774), .ZN(n20671) );
  NAND2_X1 U13713 ( .A1(n10775), .A2(n20671), .ZN(n20681) );
  INV_X1 U13714 ( .A(n16053), .ZN(n16047) );
  AOI22_X1 U13715 ( .A1(n10776), .A2(n20681), .B1(n16047), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10777) );
  INV_X1 U13716 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13717 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10780) );
  NAND2_X1 U13718 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10779) );
  OAI211_X1 U13719 ( .C1(n9760), .C2(n10781), .A(n10780), .B(n10779), .ZN(
        n10782) );
  INV_X1 U13720 ( .A(n10782), .ZN(n10786) );
  AOI22_X1 U13721 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13722 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13723 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10783) );
  NAND4_X1 U13724 ( .A1(n10786), .A2(n10785), .A3(n10784), .A4(n10783), .ZN(
        n10793) );
  AOI22_X1 U13725 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13726 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13727 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13728 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10788) );
  NAND4_X1 U13729 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10792) );
  AOI22_X1 U13730 ( .A1(n10881), .A2(n10799), .B1(n10880), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U13731 ( .A1(n10797), .A2(n13653), .ZN(n13656) );
  NAND2_X1 U13732 ( .A1(n10798), .A2(n10799), .ZN(n10847) );
  OAI211_X1 U13733 ( .C1(n10799), .C2(n10798), .A(n10847), .B(n9971), .ZN(
        n10800) );
  OAI21_X1 U13734 ( .B1(n20380), .B2(n10374), .A(n10800), .ZN(n13631) );
  NAND2_X1 U13735 ( .A1(n13632), .A2(n13631), .ZN(n10803) );
  NAND2_X1 U13736 ( .A1(n10801), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10802) );
  NAND2_X1 U13737 ( .A1(n10803), .A2(n10802), .ZN(n13715) );
  AOI22_X1 U13738 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13739 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11454), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13740 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13741 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11300), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10804) );
  AND4_X1 U13742 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10818) );
  AOI22_X1 U13743 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U13744 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10810) );
  NAND2_X1 U13745 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10809) );
  NAND2_X1 U13746 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10808) );
  NAND4_X1 U13747 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .ZN(
        n10816) );
  INV_X1 U13748 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13749 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10813) );
  NAND2_X1 U13750 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10812) );
  OAI211_X1 U13751 ( .C1(n9760), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n10815) );
  NOR2_X1 U13752 ( .A1(n10816), .A2(n10815), .ZN(n10817) );
  INV_X1 U13753 ( .A(n10848), .ZN(n10819) );
  AOI22_X1 U13754 ( .A1(n10881), .A2(n10819), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10880), .ZN(n10822) );
  NAND2_X1 U13755 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  XNOR2_X1 U13756 ( .A(n10847), .B(n10848), .ZN(n10825) );
  INV_X1 U13757 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13691) );
  XNOR2_X1 U13758 ( .A(n10826), .B(n13691), .ZN(n13716) );
  NAND2_X1 U13759 ( .A1(n13715), .A2(n13716), .ZN(n10828) );
  NAND2_X1 U13760 ( .A1(n10826), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10827) );
  INV_X1 U13761 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U13762 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10830) );
  NAND2_X1 U13763 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10829) );
  OAI211_X1 U13764 ( .C1(n9760), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        n10832) );
  INV_X1 U13765 ( .A(n10832), .ZN(n10836) );
  AOI22_X1 U13766 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13767 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13768 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10833) );
  NAND4_X1 U13769 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10842) );
  AOI22_X1 U13770 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13771 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13772 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13773 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13774 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  AOI22_X1 U13775 ( .A1(n10881), .A2(n10872), .B1(n10880), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13776 ( .A1(n10845), .A2(n10844), .ZN(n10846) );
  NOR2_X1 U13777 ( .A1(n10848), .A2(n10847), .ZN(n10873) );
  XNOR2_X1 U13778 ( .A(n10872), .B(n10873), .ZN(n10849) );
  OAI22_X1 U13779 ( .A1(n10962), .A2(n10374), .B1(n10849), .B2(n16044), .ZN(
        n10851) );
  INV_X1 U13780 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10850) );
  XNOR2_X1 U13781 ( .A(n10851), .B(n10850), .ZN(n16263) );
  NAND2_X1 U13782 ( .A1(n16262), .A2(n16263), .ZN(n10853) );
  NAND2_X1 U13783 ( .A1(n10851), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10852) );
  AOI22_X1 U13784 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U13785 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10855) );
  AOI22_X1 U13786 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10854) );
  NAND3_X1 U13787 ( .A1(n10856), .A2(n10855), .A3(n10854), .ZN(n10861) );
  NAND2_X1 U13788 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U13789 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10858) );
  NAND2_X1 U13790 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10857) );
  NAND3_X1 U13791 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10860) );
  NOR2_X1 U13792 ( .A1(n10861), .A2(n10860), .ZN(n10867) );
  AOI22_X1 U13793 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13794 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13795 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13796 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10862) );
  AND4_X1 U13797 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n10866) );
  INV_X1 U13798 ( .A(n10885), .ZN(n10868) );
  AOI22_X1 U13799 ( .A1(n10881), .A2(n10868), .B1(n10880), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10870) );
  INV_X1 U13800 ( .A(n10870), .ZN(n10869) );
  NAND2_X1 U13801 ( .A1(n10871), .A2(n10870), .ZN(n10970) );
  NAND3_X1 U13802 ( .A1(n10883), .A2(n13128), .A3(n10970), .ZN(n10877) );
  NAND2_X1 U13803 ( .A1(n10873), .A2(n10872), .ZN(n10884) );
  INV_X1 U13804 ( .A(n10884), .ZN(n10874) );
  XNOR2_X1 U13805 ( .A(n10885), .B(n10874), .ZN(n10875) );
  NAND2_X1 U13806 ( .A1(n9971), .A2(n10875), .ZN(n10876) );
  NAND2_X1 U13807 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  XNOR2_X1 U13808 ( .A(n10878), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13807) );
  OR2_X1 U13809 ( .A1(n10878), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10879) );
  AOI22_X1 U13810 ( .A1(n10881), .A2(n10896), .B1(n10880), .B2(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10882) );
  XNOR2_X1 U13811 ( .A(n10883), .B(n10882), .ZN(n10974) );
  OR2_X1 U13812 ( .A1(n10974), .A2(n10374), .ZN(n10889) );
  NOR2_X1 U13813 ( .A1(n10885), .A2(n10884), .ZN(n10897) );
  INV_X1 U13814 ( .A(n10897), .ZN(n10886) );
  XNOR2_X1 U13815 ( .A(n10896), .B(n10886), .ZN(n10887) );
  NAND2_X1 U13816 ( .A1(n9971), .A2(n10887), .ZN(n10888) );
  NAND2_X1 U13817 ( .A1(n10889), .A2(n10888), .ZN(n10890) );
  INV_X1 U13818 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16387) );
  XNOR2_X1 U13819 ( .A(n10890), .B(n16387), .ZN(n16256) );
  INV_X1 U13820 ( .A(n10890), .ZN(n10891) );
  NAND2_X1 U13821 ( .A1(n10891), .A2(n16387), .ZN(n10892) );
  NAND2_X1 U13822 ( .A1(n13128), .A2(n10896), .ZN(n10894) );
  NOR2_X1 U13823 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  NAND3_X1 U13824 ( .A1(n9971), .A2(n10897), .A3(n10896), .ZN(n10898) );
  NAND2_X1 U13825 ( .A1(n16212), .A2(n10898), .ZN(n10899) );
  NAND2_X1 U13826 ( .A1(n10899), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13928) );
  INV_X1 U13827 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16361) );
  NAND2_X1 U13828 ( .A1(n9753), .A2(n16361), .ZN(n10900) );
  INV_X1 U13829 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16330) );
  NAND2_X1 U13830 ( .A1(n16212), .A2(n16330), .ZN(n10901) );
  INV_X1 U13831 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U13832 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U13833 ( .A1(n16212), .A2(n10902), .ZN(n14663) );
  INV_X1 U13834 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U13835 ( .A1(n16212), .A2(n10907), .ZN(n10903) );
  INV_X1 U13836 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21199) );
  INV_X1 U13837 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16313) );
  XNOR2_X1 U13838 ( .A(n16212), .B(n16313), .ZN(n14647) );
  NOR2_X1 U13839 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10905) );
  OR2_X1 U13840 ( .A1(n10906), .A2(n10907), .ZN(n10908) );
  NOR2_X1 U13841 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14661) );
  AND2_X1 U13842 ( .A1(n14661), .A2(n14092), .ZN(n10909) );
  OR2_X1 U13843 ( .A1(n10906), .A2(n10909), .ZN(n16225) );
  OR2_X1 U13844 ( .A1(n10906), .A2(n21199), .ZN(n16229) );
  AND2_X1 U13845 ( .A1(n16225), .A2(n16229), .ZN(n10910) );
  XNOR2_X1 U13846 ( .A(n9753), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14640) );
  NAND2_X1 U13847 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14789) );
  INV_X1 U13848 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14795) );
  NOR2_X1 U13849 ( .A1(n14789), .A2(n14795), .ZN(n14697) );
  INV_X1 U13850 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14818) );
  INV_X1 U13851 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10912) );
  INV_X1 U13852 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14114) );
  AND2_X1 U13853 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U13854 ( .A1(n14768), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14698) );
  INV_X1 U13855 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14704) );
  AOI211_X2 U13856 ( .C1(n16199), .C2(n14698), .A(n14704), .B(n14608), .ZN(
        n10914) );
  NOR2_X1 U13857 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14581) );
  NOR2_X1 U13858 ( .A1(n10914), .A2(n14559), .ZN(n14590) );
  NAND2_X1 U13859 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14739) );
  INV_X1 U13860 ( .A(n10914), .ZN(n10915) );
  NOR2_X1 U13861 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14558) );
  NAND2_X1 U13862 ( .A1(n10915), .A2(n14558), .ZN(n10916) );
  OAI22_X1 U13863 ( .A1(n10917), .A2(n10070), .B1(n14559), .B2(n10916), .ZN(
        n14569) );
  NOR3_X1 U13864 ( .A1(n16212), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10918) );
  OAI22_X1 U13865 ( .A1(n14569), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n14560), .B2(n10918), .ZN(n10920) );
  XNOR2_X1 U13866 ( .A(n10920), .B(n10919), .ZN(n14710) );
  NAND2_X1 U13867 ( .A1(n13604), .A2(n11129), .ZN(n10926) );
  INV_X2 U13868 ( .A(n11112), .ZN(n11436) );
  AOI22_X1 U13869 ( .A1(n11436), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21030), .ZN(n10924) );
  NAND2_X1 U13870 ( .A1(n14197), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10949) );
  INV_X1 U13871 ( .A(n10949), .ZN(n10953) );
  NAND2_X1 U13872 ( .A1(n10953), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10923) );
  AND2_X1 U13873 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  NAND2_X1 U13874 ( .A1(n10926), .A2(n10925), .ZN(n13450) );
  NAND2_X1 U13875 ( .A1(n20381), .A2(n9765), .ZN(n10927) );
  NAND2_X1 U13876 ( .A1(n10927), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U13877 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21030), .ZN(
        n10930) );
  NAND2_X1 U13878 ( .A1(n10963), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10929) );
  OAI211_X1 U13879 ( .C1(n10949), .C2(n10928), .A(n10930), .B(n10929), .ZN(
        n10931) );
  AOI21_X1 U13880 ( .B1(n20496), .B2(n11129), .A(n10931), .ZN(n10932) );
  OR2_X1 U13881 ( .A1(n13330), .A2(n10932), .ZN(n13331) );
  INV_X1 U13882 ( .A(n10932), .ZN(n13332) );
  OR2_X1 U13883 ( .A1(n13332), .A2(n14154), .ZN(n10933) );
  NAND2_X1 U13884 ( .A1(n13331), .A2(n10933), .ZN(n13449) );
  NAND2_X1 U13885 ( .A1(n13450), .A2(n13449), .ZN(n13593) );
  INV_X1 U13886 ( .A(n14154), .ZN(n11150) );
  XNOR2_X1 U13887 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14361) );
  AOI21_X1 U13888 ( .B1(n11150), .B2(n14361), .A(n11494), .ZN(n10936) );
  NAND2_X1 U13889 ( .A1(n11436), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10935) );
  OAI211_X1 U13890 ( .C1(n10949), .C2(n10430), .A(n10936), .B(n10935), .ZN(
        n10937) );
  INV_X1 U13891 ( .A(n10937), .ZN(n10938) );
  NAND2_X1 U13892 ( .A1(n11494), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10942) );
  NAND2_X1 U13893 ( .A1(n10939), .A2(n10942), .ZN(n13594) );
  NAND2_X1 U13894 ( .A1(n10941), .A2(n10940), .ZN(n13591) );
  INV_X1 U13895 ( .A(n10944), .ZN(n10946) );
  INV_X1 U13896 ( .A(n10955), .ZN(n10945) );
  OAI21_X1 U13897 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10946), .A(
        n10945), .ZN(n20256) );
  AOI22_X1 U13898 ( .A1(n11150), .A2(n20256), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U13899 ( .A1(n11436), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10947) );
  OAI211_X1 U13900 ( .C1(n10949), .C2(n21260), .A(n10948), .B(n10947), .ZN(
        n10950) );
  INV_X1 U13901 ( .A(n10950), .ZN(n10951) );
  OAI21_X1 U13902 ( .B1(n20380), .B2(n11095), .A(n10951), .ZN(n13619) );
  NAND2_X1 U13903 ( .A1(n13620), .A2(n13619), .ZN(n13618) );
  NAND2_X1 U13904 ( .A1(n10953), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10958) );
  INV_X1 U13905 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20239) );
  AOI21_X1 U13906 ( .B1(n20239), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10954) );
  AOI21_X1 U13907 ( .B1(n11436), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10954), .ZN(
        n10957) );
  OAI21_X1 U13908 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10955), .A(
        n10964), .ZN(n20244) );
  NOR2_X1 U13909 ( .A1(n20244), .A2(n14154), .ZN(n10956) );
  AOI21_X1 U13910 ( .B1(n10958), .B2(n10957), .A(n10956), .ZN(n10959) );
  AOI21_X1 U13911 ( .B1(n10960), .B2(n11129), .A(n10959), .ZN(n13689) );
  INV_X1 U13912 ( .A(n10963), .ZN(n11112) );
  INV_X1 U13913 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13753) );
  INV_X1 U13914 ( .A(n10964), .ZN(n10966) );
  INV_X1 U13915 ( .A(n10971), .ZN(n10965) );
  OAI21_X1 U13916 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10966), .A(
        n10965), .ZN(n16264) );
  AOI22_X1 U13917 ( .A1(n11150), .A2(n16264), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10967) );
  OAI21_X1 U13918 ( .B1(n11112), .B2(n13753), .A(n10967), .ZN(n10968) );
  INV_X1 U13919 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20322) );
  NAND2_X1 U13920 ( .A1(n10970), .A2(n11129), .ZN(n10973) );
  OAI21_X1 U13921 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10971), .A(
        n10976), .ZN(n20216) );
  AOI22_X1 U13922 ( .A1(n11150), .A2(n20216), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10972) );
  INV_X1 U13923 ( .A(n10974), .ZN(n10975) );
  NAND2_X1 U13924 ( .A1(n10975), .A2(n11129), .ZN(n10982) );
  INV_X1 U13925 ( .A(n11494), .ZN(n11039) );
  INV_X1 U13926 ( .A(n10976), .ZN(n10978) );
  INV_X1 U13927 ( .A(n11002), .ZN(n10977) );
  OAI21_X1 U13928 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10978), .A(
        n10977), .ZN(n20207) );
  NAND2_X1 U13929 ( .A1(n20207), .A2(n10934), .ZN(n10979) );
  OAI21_X1 U13930 ( .B1(n16261), .B2(n11039), .A(n10979), .ZN(n10980) );
  AOI21_X1 U13931 ( .B1(n11436), .B2(P1_EAX_REG_7__SCAN_IN), .A(n10980), .ZN(
        n10981) );
  NAND2_X1 U13932 ( .A1(n11436), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11000) );
  XNOR2_X1 U13933 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11002), .ZN(
        n14352) );
  AOI22_X1 U13934 ( .A1(n10934), .A2(n14352), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10999) );
  INV_X1 U13935 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U13936 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U13937 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10983) );
  OAI211_X1 U13938 ( .C1(n9760), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n10986) );
  INV_X1 U13939 ( .A(n10986), .ZN(n10990) );
  AOI22_X1 U13940 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U13941 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13942 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10987) );
  NAND4_X1 U13943 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n10996) );
  AOI22_X1 U13944 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13945 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13946 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13947 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10991) );
  NAND4_X1 U13948 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10995) );
  NOR2_X1 U13949 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  OR2_X1 U13950 ( .A1(n11095), .A2(n10997), .ZN(n10998) );
  XOR2_X1 U13951 ( .A(n11021), .B(n11022), .Z(n20194) );
  INV_X1 U13952 ( .A(n20194), .ZN(n14686) );
  INV_X1 U13953 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U13954 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13955 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13956 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13957 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11003) );
  AND4_X1 U13958 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11014) );
  AOI22_X1 U13959 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U13960 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13961 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11009) );
  AOI22_X1 U13962 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11008) );
  AND3_X1 U13963 ( .A1(n11010), .A2(n11009), .A3(n11008), .ZN(n11012) );
  NAND2_X1 U13964 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11011) );
  NAND4_X1 U13965 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11015) );
  NAND2_X1 U13966 ( .A1(n11129), .A2(n11015), .ZN(n11017) );
  NAND2_X1 U13967 ( .A1(n11494), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11016) );
  OAI211_X1 U13968 ( .C1(n13938), .C2(n11112), .A(n11017), .B(n11016), .ZN(
        n11018) );
  AOI21_X1 U13969 ( .B1(n14686), .B2(n10934), .A(n11018), .ZN(n13936) );
  XNOR2_X1 U13970 ( .A(n11041), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14679) );
  INV_X1 U13971 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13972 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9761), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13973 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13974 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13975 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11024) );
  AND4_X1 U13976 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11034) );
  AOI22_X1 U13977 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U13978 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U13979 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U13980 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11028) );
  AND3_X1 U13981 ( .A1(n11030), .A2(n11029), .A3(n11028), .ZN(n11032) );
  NAND2_X1 U13982 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11031) );
  NAND4_X1 U13983 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11035) );
  NAND2_X1 U13984 ( .A1(n11129), .A2(n11035), .ZN(n11037) );
  NAND2_X1 U13985 ( .A1(n11436), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11036) );
  OAI211_X1 U13986 ( .C1(n11039), .C2(n11038), .A(n11037), .B(n11036), .ZN(
        n11040) );
  AOI21_X1 U13987 ( .B1(n14679), .B2(n10934), .A(n11040), .ZN(n14337) );
  NAND2_X1 U13988 ( .A1(n11436), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11046) );
  INV_X1 U13989 ( .A(n11042), .ZN(n11044) );
  INV_X1 U13990 ( .A(n11090), .ZN(n11043) );
  OAI21_X1 U13991 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11044), .A(
        n11043), .ZN(n16253) );
  AOI22_X1 U13992 ( .A1(n10934), .A2(n16253), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U13993 ( .A1(n11046), .A2(n11045), .ZN(n14321) );
  INV_X1 U13994 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U13995 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U13996 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11047) );
  OAI211_X1 U13997 ( .C1(n9760), .C2(n11049), .A(n11048), .B(n11047), .ZN(
        n11050) );
  INV_X1 U13998 ( .A(n11050), .ZN(n11054) );
  AOI22_X1 U13999 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14000 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U14001 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11051) );
  NAND4_X1 U14002 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11060) );
  AOI22_X1 U14003 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14004 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14005 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14006 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11055) );
  NAND4_X1 U14007 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        n11059) );
  NOR2_X1 U14008 ( .A1(n11060), .A2(n11059), .ZN(n11061) );
  NOR2_X1 U14009 ( .A1(n11095), .A2(n11061), .ZN(n14453) );
  XOR2_X1 U14010 ( .A(n14332), .B(n11097), .Z(n14670) );
  AOI22_X1 U14011 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9761), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14012 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14013 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14014 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11062) );
  AND4_X1 U14015 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11072) );
  AOI22_X1 U14016 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14017 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U14018 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11067) );
  AOI22_X1 U14019 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11066) );
  AND3_X1 U14020 ( .A1(n11068), .A2(n11067), .A3(n11066), .ZN(n11070) );
  NAND2_X1 U14021 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11069) );
  NAND4_X1 U14022 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n11073) );
  AOI22_X1 U14023 ( .A1(n11129), .A2(n11073), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U14024 ( .A1(n11436), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U14025 ( .C1(n14670), .C2(n14154), .A(n11075), .B(n11074), .ZN(
        n14325) );
  INV_X1 U14026 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14027 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14028 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11076) );
  OAI211_X1 U14029 ( .C1(n9760), .C2(n11078), .A(n11077), .B(n11076), .ZN(
        n11079) );
  INV_X1 U14030 ( .A(n11079), .ZN(n11083) );
  AOI22_X1 U14031 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14032 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9792), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14033 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11080) );
  NAND4_X1 U14034 ( .A1(n11083), .A2(n11082), .A3(n11081), .A4(n11080), .ZN(
        n11089) );
  AOI22_X1 U14035 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14036 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9761), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14037 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11399), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14038 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11084) );
  NAND4_X1 U14039 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n11084), .ZN(
        n11088) );
  NOR2_X1 U14040 ( .A1(n11089), .A2(n11088), .ZN(n11094) );
  NAND2_X1 U14041 ( .A1(n11436), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11093) );
  XOR2_X1 U14042 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11090), .Z(
        n16241) );
  INV_X1 U14043 ( .A(n16241), .ZN(n11091) );
  AOI22_X1 U14044 ( .A1(n11494), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n10934), .B2(n11091), .ZN(n11092) );
  OAI211_X1 U14045 ( .C1(n11095), .C2(n11094), .A(n11093), .B(n11092), .ZN(
        n14446) );
  NAND2_X1 U14046 ( .A1(n14325), .A2(n14446), .ZN(n11096) );
  XNOR2_X1 U14047 ( .A(n11116), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16159) );
  NAND2_X1 U14048 ( .A1(n16159), .A2(n10934), .ZN(n11115) );
  INV_X1 U14049 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14547) );
  AOI22_X1 U14050 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11404), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14051 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14052 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14053 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11098) );
  AND4_X1 U14054 ( .A1(n11101), .A2(n11100), .A3(n11099), .A4(n11098), .ZN(
        n11108) );
  AOI22_X1 U14055 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U14056 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U14057 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11103) );
  AOI22_X1 U14058 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11102) );
  AND3_X1 U14059 ( .A1(n11104), .A2(n11103), .A3(n11102), .ZN(n11106) );
  NAND2_X1 U14060 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11105) );
  NAND4_X1 U14061 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(
        n11109) );
  NAND2_X1 U14062 ( .A1(n11129), .A2(n11109), .ZN(n11111) );
  NAND2_X1 U14063 ( .A1(n11494), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11110) );
  OAI211_X1 U14064 ( .C1(n11112), .C2(n14547), .A(n11111), .B(n11110), .ZN(
        n11113) );
  INV_X1 U14065 ( .A(n11113), .ZN(n11114) );
  NAND2_X1 U14066 ( .A1(n11115), .A2(n11114), .ZN(n14438) );
  XOR2_X1 U14067 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11132), .Z(
        n16235) );
  AOI22_X1 U14068 ( .A1(n9802), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9790), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14069 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14070 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14071 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11117) );
  AND4_X1 U14072 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(
        n11127) );
  AOI22_X1 U14073 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14074 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14075 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11122) );
  AOI22_X1 U14076 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11121) );
  AND3_X1 U14077 ( .A1(n11123), .A2(n11122), .A3(n11121), .ZN(n11125) );
  NAND2_X1 U14078 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11124) );
  NAND4_X1 U14079 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11128) );
  AOI22_X1 U14080 ( .A1(n11129), .A2(n11128), .B1(n11494), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U14081 ( .A1(n11436), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11130) );
  OAI211_X1 U14082 ( .C1(n16235), .C2(n14154), .A(n11131), .B(n11130), .ZN(
        n14433) );
  NAND2_X1 U14083 ( .A1(n14431), .A2(n14433), .ZN(n14307) );
  XOR2_X1 U14084 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11172), .Z(
        n16220) );
  INV_X1 U14085 ( .A(n16220), .ZN(n11151) );
  INV_X1 U14086 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14087 ( .A1(n11405), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14088 ( .A1(n9790), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11133) );
  OAI211_X1 U14089 ( .C1(n9760), .C2(n11135), .A(n11134), .B(n11133), .ZN(
        n11136) );
  INV_X1 U14090 ( .A(n11136), .ZN(n11140) );
  AOI22_X1 U14091 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14092 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U14093 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11137) );
  NAND4_X1 U14094 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11146) );
  AOI22_X1 U14095 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14096 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14097 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14098 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11141) );
  NAND4_X1 U14099 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  NOR2_X1 U14100 ( .A1(n11146), .A2(n11145), .ZN(n11148) );
  AOI22_X1 U14101 ( .A1(n11436), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n11494), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11147) );
  OAI21_X1 U14102 ( .B1(n11488), .B2(n11148), .A(n11147), .ZN(n11149) );
  AOI21_X1 U14103 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n14422) );
  XNOR2_X1 U14104 ( .A(n11152), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14649) );
  INV_X1 U14105 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U14106 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14107 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11153) );
  OAI211_X1 U14108 ( .C1(n9760), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11156) );
  INV_X1 U14109 ( .A(n11156), .ZN(n11160) );
  AOI22_X1 U14110 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14111 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U14112 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11157) );
  NAND4_X1 U14113 ( .A1(n11160), .A2(n11159), .A3(n11158), .A4(n11157), .ZN(
        n11166) );
  AOI22_X1 U14114 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14115 ( .A1(n9790), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14116 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14117 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11161) );
  NAND4_X1 U14118 ( .A1(n11164), .A2(n11163), .A3(n11162), .A4(n11161), .ZN(
        n11165) );
  NOR2_X1 U14119 ( .A1(n11166), .A2(n11165), .ZN(n11168) );
  AOI22_X1 U14120 ( .A1(n11436), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21030), .ZN(n11167) );
  OAI21_X1 U14121 ( .B1(n11488), .B2(n11168), .A(n11167), .ZN(n11169) );
  AND2_X1 U14122 ( .A1(n11169), .A2(n14154), .ZN(n11170) );
  AOI21_X1 U14123 ( .B1(n14649), .B2(n10934), .A(n11170), .ZN(n14309) );
  OR2_X1 U14124 ( .A1(n14422), .A2(n14309), .ZN(n11171) );
  NAND2_X1 U14125 ( .A1(n11173), .A2(n21335), .ZN(n11175) );
  INV_X1 U14126 ( .A(n11211), .ZN(n11174) );
  NAND2_X1 U14127 ( .A1(n11175), .A2(n11174), .ZN(n16132) );
  INV_X1 U14128 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U14129 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14130 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11176) );
  OAI211_X1 U14131 ( .C1(n9760), .C2(n11347), .A(n11177), .B(n11176), .ZN(
        n11178) );
  INV_X1 U14132 ( .A(n11178), .ZN(n11182) );
  AOI22_X1 U14133 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14134 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U14135 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11179) );
  NAND4_X1 U14136 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        n11188) );
  AOI22_X1 U14137 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14138 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14139 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14140 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11183) );
  NAND4_X1 U14141 ( .A1(n11186), .A2(n11185), .A3(n11184), .A4(n11183), .ZN(
        n11187) );
  NOR2_X1 U14142 ( .A1(n11188), .A2(n11187), .ZN(n11191) );
  AOI21_X1 U14143 ( .B1(n11436), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11189), .ZN(
        n11190) );
  OAI21_X1 U14144 ( .B1(n11488), .B2(n11191), .A(n11190), .ZN(n11192) );
  OAI21_X1 U14145 ( .B1(n16132), .B2(n14154), .A(n11192), .ZN(n14411) );
  NOR2_X4 U14146 ( .A1(n14419), .A2(n14411), .ZN(n14412) );
  INV_X1 U14147 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14148 ( .A1(n11405), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11194) );
  NAND2_X1 U14149 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11193) );
  OAI211_X1 U14150 ( .C1(n9760), .C2(n11368), .A(n11194), .B(n11193), .ZN(
        n11195) );
  INV_X1 U14151 ( .A(n11195), .ZN(n11199) );
  AOI22_X1 U14152 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14153 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U14154 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11196) );
  NAND4_X1 U14155 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11206) );
  AOI22_X1 U14156 ( .A1(n9802), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9790), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14157 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14158 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14159 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11201) );
  NAND4_X1 U14160 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .ZN(
        n11205) );
  NOR2_X1 U14161 ( .A1(n11206), .A2(n11205), .ZN(n11210) );
  NAND2_X1 U14162 ( .A1(n21030), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14163 ( .A1(n14154), .A2(n11207), .ZN(n11208) );
  AOI21_X1 U14164 ( .B1(n11436), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11208), .ZN(
        n11209) );
  OAI21_X1 U14165 ( .B1(n11488), .B2(n11210), .A(n11209), .ZN(n11213) );
  OAI21_X1 U14166 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11211), .A(
        n11253), .ZN(n16219) );
  OR2_X1 U14167 ( .A1(n14154), .A2(n16219), .ZN(n11212) );
  AOI22_X1 U14168 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14169 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11327), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14170 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14171 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9792), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14172 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11227) );
  AOI22_X1 U14173 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U14174 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14175 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14176 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14177 ( .A1(n9786), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11218) );
  AND4_X1 U14178 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11224) );
  NAND2_X1 U14179 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14180 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11222) );
  NAND4_X1 U14181 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11226) );
  NOR2_X1 U14182 ( .A1(n11227), .A2(n11226), .ZN(n11230) );
  AOI21_X1 U14183 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16117), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11228) );
  AOI21_X1 U14184 ( .B1(n11436), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11228), .ZN(
        n11229) );
  OAI21_X1 U14185 ( .B1(n11488), .B2(n11230), .A(n11229), .ZN(n11232) );
  XNOR2_X1 U14186 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11253), .ZN(
        n16107) );
  NAND2_X1 U14187 ( .A1(n11150), .A2(n16107), .ZN(n11231) );
  AOI22_X1 U14188 ( .A1(n9802), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U14189 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11238) );
  NAND2_X1 U14190 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U14191 ( .A1(n9786), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11236) );
  NAND2_X1 U14192 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11235) );
  AND4_X1 U14193 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11241) );
  NAND2_X1 U14194 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11240) );
  NAND2_X1 U14195 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11239) );
  NAND4_X1 U14196 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11248) );
  AOI22_X1 U14197 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9791), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14198 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14199 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14200 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11243) );
  NAND4_X1 U14201 ( .A1(n11246), .A2(n11245), .A3(n11244), .A4(n11243), .ZN(
        n11247) );
  NOR2_X1 U14202 ( .A1(n11248), .A2(n11247), .ZN(n11252) );
  NAND2_X1 U14203 ( .A1(n21030), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14204 ( .A1(n14154), .A2(n11249), .ZN(n11250) );
  AOI21_X1 U14205 ( .B1(n11436), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11250), .ZN(
        n11251) );
  OAI21_X1 U14206 ( .B1(n11488), .B2(n11252), .A(n11251), .ZN(n11256) );
  OAI21_X1 U14207 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11254), .A(
        n11276), .ZN(n16208) );
  OR2_X1 U14208 ( .A1(n14154), .A2(n16208), .ZN(n11255) );
  NAND2_X1 U14209 ( .A1(n11256), .A2(n11255), .ZN(n16101) );
  INV_X1 U14210 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11259) );
  NAND2_X1 U14211 ( .A1(n10661), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11258) );
  NAND2_X1 U14212 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11257) );
  OAI211_X1 U14213 ( .C1(n9760), .C2(n11259), .A(n11258), .B(n11257), .ZN(
        n11260) );
  INV_X1 U14214 ( .A(n11260), .ZN(n11264) );
  AOI22_X1 U14215 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14216 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14217 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11261) );
  NAND4_X1 U14218 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .ZN(
        n11272) );
  AOI22_X1 U14219 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14220 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14221 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14222 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14223 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11271) );
  NOR2_X1 U14224 ( .A1(n11272), .A2(n11271), .ZN(n11275) );
  OAI21_X1 U14225 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21139), .A(n14154), 
        .ZN(n11273) );
  AOI21_X1 U14226 ( .B1(n11436), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11273), .ZN(
        n11274) );
  OAI21_X1 U14227 ( .B1(n11488), .B2(n11275), .A(n11274), .ZN(n11280) );
  INV_X1 U14228 ( .A(n11276), .ZN(n11278) );
  INV_X1 U14229 ( .A(n11314), .ZN(n11277) );
  OAI21_X1 U14230 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11278), .A(
        n11277), .ZN(n16087) );
  OR2_X1 U14231 ( .A1(n14154), .A2(n16087), .ZN(n11279) );
  NAND2_X1 U14232 ( .A1(n11280), .A2(n11279), .ZN(n14396) );
  INV_X1 U14233 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11287) );
  INV_X1 U14234 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14235 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14236 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11473), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11281) );
  OAI211_X1 U14237 ( .C1(n9760), .C2(n11283), .A(n11282), .B(n11281), .ZN(
        n11284) );
  INV_X1 U14238 ( .A(n11284), .ZN(n11286) );
  AOI22_X1 U14239 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11285) );
  OAI211_X1 U14240 ( .C1(n9756), .C2(n11287), .A(n11286), .B(n11285), .ZN(
        n11293) );
  AOI22_X1 U14241 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14242 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14243 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9798), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14244 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11288) );
  NAND4_X1 U14245 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11292) );
  NOR2_X1 U14246 ( .A1(n11293), .A2(n11292), .ZN(n11317) );
  INV_X1 U14247 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11303) );
  INV_X1 U14248 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11294) );
  INV_X1 U14249 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11471) );
  OAI22_X1 U14250 ( .A1(n9757), .A2(n11294), .B1(n9787), .B2(n11471), .ZN(
        n11299) );
  INV_X1 U14251 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11296) );
  INV_X1 U14252 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11295) );
  OAI22_X1 U14253 ( .A1(n11297), .A2(n11296), .B1(n9764), .B2(n11295), .ZN(
        n11298) );
  AOI211_X1 U14254 ( .C1(n11402), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11299), .B(n11298), .ZN(n11302) );
  AOI22_X1 U14255 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11301) );
  OAI211_X1 U14256 ( .C1(n9760), .C2(n11303), .A(n11302), .B(n11301), .ZN(
        n11309) );
  AOI22_X1 U14257 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14258 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14259 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14260 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11304) );
  NAND4_X1 U14261 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11308) );
  NOR2_X1 U14262 ( .A1(n11309), .A2(n11308), .ZN(n11318) );
  XNOR2_X1 U14263 ( .A(n11317), .B(n11318), .ZN(n11313) );
  NAND2_X1 U14264 ( .A1(n21030), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14265 ( .A1(n14154), .A2(n11310), .ZN(n11311) );
  AOI21_X1 U14266 ( .B1(n11436), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11311), .ZN(
        n11312) );
  OAI21_X1 U14267 ( .B1(n11313), .B2(n11488), .A(n11312), .ZN(n11316) );
  OAI21_X1 U14268 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n11314), .A(
        n11339), .ZN(n16203) );
  OR2_X1 U14269 ( .A1(n14154), .A2(n16203), .ZN(n11315) );
  NOR2_X1 U14270 ( .A1(n11318), .A2(n11317), .ZN(n11346) );
  INV_X1 U14271 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U14272 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11320) );
  NAND2_X1 U14273 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11319) );
  OAI211_X1 U14274 ( .C1(n9760), .C2(n11321), .A(n11320), .B(n11319), .ZN(
        n11322) );
  INV_X1 U14275 ( .A(n11322), .ZN(n11326) );
  AOI22_X1 U14276 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14277 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14278 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11323) );
  NAND4_X1 U14279 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11333) );
  AOI22_X1 U14280 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14281 ( .A1(n11404), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14282 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14283 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U14284 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11332) );
  OR2_X1 U14285 ( .A1(n11333), .A2(n11332), .ZN(n11345) );
  XNOR2_X1 U14286 ( .A(n11346), .B(n11345), .ZN(n11336) );
  INV_X1 U14287 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14622) );
  AOI21_X1 U14288 ( .B1(n14622), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11334) );
  AOI21_X1 U14289 ( .B1(n11436), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11334), .ZN(
        n11335) );
  OAI21_X1 U14290 ( .B1(n11336), .B2(n11488), .A(n11335), .ZN(n11338) );
  XNOR2_X1 U14291 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n11339), .ZN(
        n14620) );
  NAND2_X1 U14292 ( .A1(n11150), .A2(n14620), .ZN(n11337) );
  NAND2_X1 U14293 ( .A1(n11338), .A2(n11337), .ZN(n14284) );
  INV_X1 U14294 ( .A(n11341), .ZN(n11343) );
  INV_X1 U14295 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14296 ( .A1(n11343), .A2(n11342), .ZN(n11344) );
  NAND2_X1 U14297 ( .A1(n11389), .A2(n11344), .ZN(n14613) );
  NAND2_X1 U14298 ( .A1(n11346), .A2(n11345), .ZN(n11366) );
  INV_X1 U14299 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11355) );
  INV_X1 U14300 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11348) );
  OAI22_X1 U14301 ( .A1(n9757), .A2(n11348), .B1(n9787), .B2(n11347), .ZN(
        n11352) );
  INV_X1 U14302 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11350) );
  OAI22_X1 U14303 ( .A1(n11373), .A2(n11350), .B1(n9800), .B2(n11349), .ZN(
        n11351) );
  AOI211_X1 U14304 ( .C1(n11402), .C2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11352), .B(n11351), .ZN(n11354) );
  AOI22_X1 U14305 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11353) );
  OAI211_X1 U14306 ( .C1(n9760), .C2(n11355), .A(n11354), .B(n11353), .ZN(
        n11361) );
  AOI22_X1 U14307 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14308 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11404), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14309 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14310 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14311 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  NOR2_X1 U14312 ( .A1(n11361), .A2(n11360), .ZN(n11367) );
  XNOR2_X1 U14313 ( .A(n11366), .B(n11367), .ZN(n11364) );
  INV_X1 U14314 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20894) );
  OAI21_X1 U14315 ( .B1(n20894), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n21030), .ZN(n11363) );
  NAND2_X1 U14316 ( .A1(n11436), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11362) );
  OAI211_X1 U14317 ( .C1(n11364), .C2(n11488), .A(n11363), .B(n11362), .ZN(
        n11365) );
  XNOR2_X1 U14318 ( .A(n11389), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14606) );
  INV_X1 U14319 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U14320 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14602), .A(n14154), 
        .ZN(n11387) );
  NOR2_X1 U14321 ( .A1(n11367), .A2(n11366), .ZN(n11394) );
  INV_X1 U14322 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11370) );
  OAI22_X1 U14323 ( .A1(n9757), .A2(n11370), .B1(n9787), .B2(n11368), .ZN(
        n11376) );
  INV_X1 U14324 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11374) );
  INV_X1 U14325 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11372) );
  OAI22_X1 U14326 ( .A1(n10695), .A2(n11374), .B1(n11373), .B2(n11372), .ZN(
        n11375) );
  AOI211_X1 U14327 ( .C1(n11402), .C2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11376), .B(n11375), .ZN(n11384) );
  INV_X1 U14328 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21303) );
  AOI22_X1 U14329 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14330 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14331 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14332 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11377) );
  AND4_X1 U14333 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n11383) );
  AOI22_X1 U14334 ( .A1(n10661), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U14335 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11381) );
  NAND4_X1 U14336 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11393) );
  XNOR2_X1 U14337 ( .A(n11394), .B(n11393), .ZN(n11385) );
  NOR2_X1 U14338 ( .A1(n11385), .A2(n11488), .ZN(n11386) );
  AOI211_X1 U14339 ( .C1(n11436), .C2(P1_EAX_REG_26__SCAN_IN), .A(n11387), .B(
        n11386), .ZN(n11388) );
  AOI21_X1 U14340 ( .B1(n11150), .B2(n14606), .A(n11388), .ZN(n14258) );
  INV_X1 U14341 ( .A(n11390), .ZN(n11391) );
  INV_X1 U14342 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U14343 ( .A1(n11391), .A2(n14249), .ZN(n11392) );
  NAND2_X1 U14344 ( .A1(n11438), .A2(n11392), .ZN(n14594) );
  NAND2_X1 U14345 ( .A1(n11394), .A2(n11393), .ZN(n11417) );
  INV_X1 U14346 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11403) );
  INV_X1 U14347 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14348 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9802), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14349 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11395) );
  OAI211_X1 U14350 ( .C1(n9760), .C2(n11397), .A(n11396), .B(n11395), .ZN(
        n11398) );
  INV_X1 U14351 ( .A(n11398), .ZN(n11401) );
  AOI22_X1 U14352 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11399), .B1(
        n9761), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11400) );
  OAI211_X1 U14353 ( .C1(n11403), .C2(n9756), .A(n11401), .B(n11400), .ZN(
        n11412) );
  AOI22_X1 U14354 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10746), .B1(
        n11404), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14355 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9809), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14356 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9792), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14357 ( .A1(n9818), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U14358 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11411) );
  NOR2_X1 U14359 ( .A1(n11412), .A2(n11411), .ZN(n11418) );
  XNOR2_X1 U14360 ( .A(n11417), .B(n11418), .ZN(n11415) );
  AOI21_X1 U14361 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21030), .A(
        n11150), .ZN(n11414) );
  NAND2_X1 U14362 ( .A1(n11436), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11413) );
  OAI211_X1 U14363 ( .C1(n11415), .C2(n11488), .A(n11414), .B(n11413), .ZN(
        n11416) );
  OAI21_X1 U14364 ( .B1(n14154), .B2(n14594), .A(n11416), .ZN(n14247) );
  NOR2_X2 U14365 ( .A1(n14246), .A2(n14247), .ZN(n14231) );
  XNOR2_X1 U14366 ( .A(n11438), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14579) );
  INV_X1 U14367 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14577) );
  AOI21_X1 U14368 ( .B1(n14577), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11435) );
  NOR2_X1 U14369 ( .A1(n11418), .A2(n11417), .ZN(n11462) );
  INV_X1 U14370 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11421) );
  NAND2_X1 U14371 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11420) );
  NAND2_X1 U14372 ( .A1(n9790), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11419) );
  OAI211_X1 U14373 ( .C1(n9760), .C2(n11421), .A(n11420), .B(n11419), .ZN(
        n11422) );
  INV_X1 U14374 ( .A(n11422), .ZN(n11426) );
  AOI22_X1 U14375 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14376 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14377 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11423) );
  NAND4_X1 U14378 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11432) );
  AOI22_X1 U14379 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14380 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14381 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14382 ( .A1(n9802), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11427) );
  NAND4_X1 U14383 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11431) );
  OR2_X1 U14384 ( .A1(n11432), .A2(n11431), .ZN(n11461) );
  XNOR2_X1 U14385 ( .A(n11462), .B(n11461), .ZN(n11433) );
  NOR2_X1 U14386 ( .A1(n11433), .A2(n11488), .ZN(n11434) );
  AOI211_X1 U14387 ( .C1(n11436), .C2(P1_EAX_REG_28__SCAN_IN), .A(n11435), .B(
        n11434), .ZN(n11437) );
  AOI21_X1 U14388 ( .B1(n11150), .B2(n14579), .A(n11437), .ZN(n14232) );
  INV_X1 U14389 ( .A(n11438), .ZN(n11439) );
  INV_X1 U14390 ( .A(n11440), .ZN(n11441) );
  INV_X1 U14391 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U14392 ( .A1(n11441), .A2(n14224), .ZN(n11442) );
  NAND2_X1 U14393 ( .A1(n11499), .A2(n11442), .ZN(n14572) );
  INV_X1 U14394 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11443) );
  OAI22_X1 U14395 ( .A1(n9800), .A2(n11445), .B1(n9764), .B2(n11443), .ZN(
        n11447) );
  AOI21_X1 U14396 ( .B1(n11402), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11447), .ZN(n11452) );
  AOI22_X1 U14397 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9798), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14398 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9792), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14399 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11449) );
  NAND4_X1 U14400 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11460) );
  AOI22_X1 U14401 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14402 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14403 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11405), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14404 ( .A1(n10466), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11453), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14405 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11459) );
  NOR2_X1 U14406 ( .A1(n11460), .A2(n11459), .ZN(n11468) );
  NAND2_X1 U14407 ( .A1(n11462), .A2(n11461), .ZN(n11467) );
  XNOR2_X1 U14408 ( .A(n11468), .B(n11467), .ZN(n11465) );
  AOI21_X1 U14409 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21030), .A(
        n11150), .ZN(n11464) );
  NAND2_X1 U14410 ( .A1(n11436), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11463) );
  OAI211_X1 U14411 ( .C1(n11465), .C2(n11488), .A(n11464), .B(n11463), .ZN(
        n11466) );
  OAI21_X1 U14412 ( .B1(n14154), .B2(n14572), .A(n11466), .ZN(n14221) );
  NOR2_X1 U14413 ( .A1(n11468), .A2(n11467), .ZN(n11487) );
  OAI22_X1 U14414 ( .A1(n10656), .A2(n11471), .B1(n11470), .B2(n11469), .ZN(
        n11472) );
  AOI21_X1 U14415 ( .B1(n11402), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11472), .ZN(n11477) );
  AOI22_X1 U14416 ( .A1(n11473), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9786), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14417 ( .A1(n9792), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11475) );
  NAND2_X1 U14418 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11474) );
  NAND4_X1 U14419 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11485) );
  AOI22_X1 U14420 ( .A1(n9795), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11454), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14421 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11327), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14422 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10491), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14423 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9818), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11480) );
  NAND4_X1 U14424 ( .A1(n11483), .A2(n11482), .A3(n11481), .A4(n11480), .ZN(
        n11484) );
  NOR2_X1 U14425 ( .A1(n11485), .A2(n11484), .ZN(n11486) );
  XNOR2_X1 U14426 ( .A(n11487), .B(n11486), .ZN(n11490) );
  INV_X1 U14427 ( .A(n11488), .ZN(n11489) );
  NAND2_X1 U14428 ( .A1(n11490), .A2(n11489), .ZN(n11493) );
  INV_X1 U14429 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14562) );
  AOI21_X1 U14430 ( .B1(n14562), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11491) );
  AOI21_X1 U14431 ( .B1(n11436), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11491), .ZN(
        n11492) );
  XNOR2_X1 U14432 ( .A(n11499), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14564) );
  AOI22_X1 U14433 ( .A1(n11493), .A2(n11492), .B1(n14564), .B2(n10934), .ZN(
        n14206) );
  AOI22_X1 U14434 ( .A1(n11436), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11494), .ZN(n11495) );
  NAND3_X1 U14435 ( .A1(n21027), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16409) );
  INV_X1 U14436 ( .A(n16409), .ZN(n11496) );
  NOR2_X2 U14437 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20826) );
  AND2_X2 U14438 ( .A1(n11496), .A2(n20826), .ZN(n20378) );
  NAND2_X1 U14439 ( .A1(n20958), .A2(n11501), .ZN(n21118) );
  AND2_X1 U14440 ( .A1(n21118), .A2(n21027), .ZN(n11497) );
  NAND2_X1 U14441 ( .A1(n21027), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U14442 ( .A1(n20894), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U14443 ( .A1(n16048), .A2(n11498), .ZN(n20366) );
  INV_X1 U14444 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14174) );
  OR2_X2 U14445 ( .A1(n11501), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20243) );
  INV_X2 U14446 ( .A(n20243), .ZN(n16368) );
  NAND2_X1 U14447 ( .A1(n16368), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U14448 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11502) );
  OAI211_X1 U14449 ( .C1(n16254), .C2(n14214), .A(n14706), .B(n11502), .ZN(
        n11503) );
  OAI21_X1 U14450 ( .B1(n16244), .B2(n14710), .A(n11504), .ZN(P1_U2968) );
  AND2_X2 U14451 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12142) );
  AND2_X4 U14452 ( .A1(n12142), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11752) );
  AND2_X4 U14453 ( .A1(n15661), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11744) );
  AOI22_X1 U14454 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11509) );
  AND2_X4 U14455 ( .A1(n11755), .A2(n16597), .ZN(n11602) );
  AOI22_X1 U14456 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11508) );
  NOR2_X2 U14457 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14458 ( .A1(n11511), .A2(n15689), .ZN(n11517) );
  AOI22_X1 U14459 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14460 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14461 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14462 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11513) );
  NAND4_X1 U14463 ( .A1(n10407), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11516) );
  NAND2_X2 U14464 ( .A1(n11517), .A2(n11516), .ZN(n19476) );
  AOI22_X1 U14465 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11744), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14466 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14467 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14468 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14469 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14470 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14471 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n11602), .ZN(n11524) );
  AOI22_X1 U14472 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9824), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14473 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11529) );
  INV_X4 U14474 ( .A(n12774), .ZN(n12919) );
  AOI22_X1 U14475 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11528) );
  AND3_X1 U14476 ( .A1(n11530), .A2(n11529), .A3(n11528), .ZN(n11532) );
  AOI22_X1 U14477 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11744), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11531) );
  NAND2_X1 U14478 ( .A1(n11532), .A2(n11531), .ZN(n11533) );
  AOI22_X1 U14479 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14480 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14481 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14482 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9829), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14483 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  AOI22_X1 U14484 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9835), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14485 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14486 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14487 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14488 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14489 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14490 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14491 ( .A1(n11638), .A2(n13263), .ZN(n11550) );
  NAND2_X1 U14492 ( .A1(n19476), .A2(n11548), .ZN(n11549) );
  INV_X1 U14493 ( .A(n11625), .ZN(n11574) );
  OR2_X1 U14494 ( .A1(n12799), .A2(n11733), .ZN(n11554) );
  NAND2_X1 U14495 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U14496 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11552) );
  NAND4_X1 U14497 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11561) );
  NAND2_X1 U14498 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11559) );
  OR2_X1 U14499 ( .A1(n12774), .A2(n13899), .ZN(n11558) );
  NAND2_X1 U14500 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11557) );
  NAND2_X1 U14501 ( .A1(n9826), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11556) );
  NAND4_X1 U14502 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11560) );
  NOR2_X1 U14503 ( .A1(n11561), .A2(n11560), .ZN(n11573) );
  NAND2_X1 U14504 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11565) );
  OR2_X1 U14505 ( .A1(n12799), .A2(n11726), .ZN(n11564) );
  NAND2_X1 U14506 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11563) );
  OR2_X1 U14507 ( .A1(n12774), .A2(n11724), .ZN(n11562) );
  NAND4_X1 U14508 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11571) );
  OR2_X1 U14509 ( .A1(n11601), .A2(n11709), .ZN(n11569) );
  NAND2_X1 U14510 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14511 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11567) );
  NAND2_X1 U14512 ( .A1(n9825), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11566) );
  NAND4_X1 U14513 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  NOR2_X1 U14514 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  NAND2_X1 U14515 ( .A1(n11574), .A2(n10421), .ZN(n11635) );
  AOI22_X1 U14516 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9828), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14517 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14518 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14519 ( .A1(n11578), .A2(n11575), .A3(n11576), .A4(n11577), .ZN(
        n11644) );
  AOI22_X1 U14520 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14521 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14522 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14523 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9830), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U14524 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11641) );
  MUX2_X2 U14525 ( .A(n11644), .B(n11641), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12576) );
  AND2_X1 U14526 ( .A1(n19476), .A2(n13287), .ZN(n11609) );
  AOI22_X1 U14527 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14528 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14529 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14530 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(
        n11588) );
  AOI22_X1 U14531 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14532 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14533 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14534 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9832), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11589) );
  NAND4_X1 U14535 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11593) );
  AOI22_X1 U14536 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14537 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14538 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14539 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14540 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11551), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14541 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9829), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14542 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11745), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14543 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14544 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  NAND2_X2 U14545 ( .A1(n11608), .A2(n11607), .ZN(n11623) );
  AND3_X2 U14546 ( .A1(n11628), .A2(n11609), .A3(n11611), .ZN(n12587) );
  NAND2_X1 U14547 ( .A1(n12587), .A2(n12576), .ZN(n12546) );
  NAND3_X1 U14548 ( .A1(n20143), .A2(n19467), .A3(n20141), .ZN(n11613) );
  OAI211_X1 U14549 ( .C1(n11635), .C2(n12576), .A(n12546), .B(n11613), .ZN(
        n11618) );
  NAND2_X1 U14550 ( .A1(n11630), .A2(n19467), .ZN(n11617) );
  AND2_X1 U14551 ( .A1(n11623), .A2(n12629), .ZN(n11614) );
  NAND2_X1 U14552 ( .A1(n11618), .A2(n12606), .ZN(n11619) );
  INV_X1 U14553 ( .A(n12389), .ZN(n12943) );
  NAND2_X1 U14554 ( .A1(n12607), .A2(n12609), .ZN(n11622) );
  NAND2_X1 U14555 ( .A1(n11622), .A2(n11621), .ZN(n11636) );
  INV_X1 U14556 ( .A(n12611), .ZN(n12578) );
  NAND2_X1 U14557 ( .A1(n12602), .A2(n10415), .ZN(n11633) );
  NAND2_X1 U14558 ( .A1(n9813), .A2(n11628), .ZN(n11629) );
  NAND2_X1 U14559 ( .A1(n11629), .A2(n11623), .ZN(n11631) );
  NAND2_X1 U14560 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NOR2_X1 U14561 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11680) );
  NAND2_X1 U14562 ( .A1(n11680), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11634) );
  NAND3_X1 U14563 ( .A1(n11636), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11635), 
        .ZN(n11658) );
  INV_X1 U14564 ( .A(n12955), .ZN(n12953) );
  NOR2_X1 U14565 ( .A1(n12953), .A2(n11638), .ZN(n11639) );
  AOI22_X1 U14566 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n9785), .B1(
        n11644), .B2(n15689), .ZN(n11640) );
  NAND3_X1 U14567 ( .A1(n11661), .A2(n11663), .A3(n11640), .ZN(n11646) );
  INV_X1 U14568 ( .A(n12587), .ZN(n11643) );
  OR2_X1 U14569 ( .A1(n9785), .A2(n15689), .ZN(n11642) );
  OAI211_X1 U14570 ( .C1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n11644), .A(
        n11643), .B(n11642), .ZN(n11645) );
  NAND3_X1 U14571 ( .A1(n11646), .A2(n11645), .A3(n16624), .ZN(n11647) );
  NAND2_X2 U14572 ( .A1(n11647), .A2(n15669), .ZN(n12627) );
  NAND2_X2 U14573 ( .A1(n12627), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12244) );
  INV_X1 U14574 ( .A(n12244), .ZN(n11648) );
  INV_X1 U14575 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11650) );
  INV_X1 U14576 ( .A(n11680), .ZN(n11653) );
  NAND2_X1 U14577 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14578 ( .A1(n11653), .A2(n11652), .ZN(n11654) );
  AOI21_X1 U14579 ( .B1(n14869), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11654), .ZN(
        n11655) );
  NAND2_X1 U14580 ( .A1(n9758), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14581 ( .A1(n14869), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11659) );
  INV_X1 U14582 ( .A(n11661), .ZN(n11662) );
  AND2_X2 U14583 ( .A1(n12574), .A2(n12546), .ZN(n16615) );
  NAND2_X1 U14584 ( .A1(n11663), .A2(n16615), .ZN(n15673) );
  INV_X1 U14585 ( .A(n11664), .ZN(n11666) );
  NAND2_X1 U14586 ( .A1(n11666), .A2(n11665), .ZN(n11667) );
  NAND2_X1 U14587 ( .A1(n9758), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14588 ( .A1(n14869), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11668) );
  INV_X1 U14589 ( .A(n11675), .ZN(n11674) );
  OAI21_X1 U14590 ( .B1(n20121), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15656), 
        .ZN(n11672) );
  INV_X1 U14591 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16594) );
  NAND2_X1 U14592 ( .A1(n14870), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14593 ( .A1(n14869), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11678) );
  INV_X1 U14594 ( .A(n11684), .ZN(n11683) );
  AND2_X1 U14595 ( .A1(n11680), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11681) );
  INV_X1 U14596 ( .A(n11685), .ZN(n11682) );
  NAND2_X1 U14597 ( .A1(n11683), .A2(n11682), .ZN(n11686) );
  NAND2_X1 U14598 ( .A1(n11685), .A2(n11684), .ZN(n12166) );
  INV_X1 U14600 ( .A(n11689), .ZN(n11690) );
  INV_X1 U14601 ( .A(n11695), .ZN(n11691) );
  NOR2_X1 U14602 ( .A1(n11687), .A2(n11691), .ZN(n11730) );
  NAND2_X1 U14603 ( .A1(n9839), .A2(n11730), .ZN(n11702) );
  OR2_X2 U14604 ( .A1(n11702), .A2(n10117), .ZN(n19954) );
  INV_X1 U14605 ( .A(n9783), .ZN(n11698) );
  INV_X1 U14606 ( .A(n11696), .ZN(n11697) );
  NAND2_X1 U14607 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  INV_X1 U14608 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11701) );
  OAI22_X1 U14609 ( .A1(n19973), .A2(n19954), .B1(n19783), .B2(n11701), .ZN(
        n11706) );
  INV_X1 U14610 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11704) );
  NOR2_X1 U14611 ( .A1(n9816), .A2(n11696), .ZN(n11707) );
  NAND2_X1 U14612 ( .A1(n9837), .A2(n11707), .ZN(n11708) );
  INV_X1 U14613 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11703) );
  OAI22_X1 U14614 ( .A1(n11704), .A2(n19876), .B1(n19811), .B2(n11703), .ZN(
        n11705) );
  INV_X1 U14615 ( .A(n11707), .ZN(n11714) );
  INV_X1 U14616 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11711) );
  OR2_X1 U14617 ( .A1(n19754), .A2(n11709), .ZN(n11710) );
  OAI211_X1 U14618 ( .C1(n11943), .C2(n11711), .A(n11710), .B(n20155), .ZN(
        n11712) );
  NOR2_X1 U14619 ( .A1(n11713), .A2(n11712), .ZN(n11743) );
  INV_X1 U14620 ( .A(n12665), .ZN(n13206) );
  NOR2_X2 U14621 ( .A1(n11731), .A2(n11729), .ZN(n13887) );
  OAI22_X1 U14622 ( .A1(n11715), .A2(n19507), .B1(n11979), .B2(n13899), .ZN(
        n11721) );
  NAND2_X1 U14623 ( .A1(n15665), .A2(n9816), .ZN(n11735) );
  OR2_X2 U14624 ( .A1(n11731), .A2(n11735), .ZN(n19536) );
  INV_X1 U14625 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11719) );
  INV_X1 U14626 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11718) );
  INV_X1 U14627 ( .A(n11722), .ZN(n11717) );
  OAI22_X1 U14628 ( .A1(n19536), .A2(n11719), .B1(n11718), .B2(n19916), .ZN(
        n11720) );
  NOR2_X1 U14629 ( .A1(n11721), .A2(n11720), .ZN(n11742) );
  INV_X1 U14630 ( .A(n15665), .ZN(n11723) );
  INV_X1 U14631 ( .A(n11730), .ZN(n11734) );
  NOR2_X2 U14632 ( .A1(n11731), .A2(n11734), .ZN(n19570) );
  INV_X1 U14633 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11732) );
  INV_X1 U14634 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11737) );
  INV_X1 U14635 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11736) );
  OAI22_X1 U14636 ( .A1(n11737), .A2(n11941), .B1(n11936), .B2(n11736), .ZN(
        n11738) );
  NOR2_X1 U14637 ( .A1(n11739), .A2(n11738), .ZN(n11740) );
  NAND4_X1 U14638 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11788) );
  AOI22_X1 U14639 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11750) );
  AND2_X2 U14640 ( .A1(n12926), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11817) );
  AOI22_X1 U14641 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11749) );
  AND2_X2 U14642 ( .A1(n12919), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11887) );
  AND2_X2 U14643 ( .A1(n11579), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11848) );
  AOI22_X1 U14644 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14645 ( .A1(n11752), .A2(n15689), .ZN(n11853) );
  AND2_X2 U14646 ( .A1(n9826), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12363) );
  AOI22_X1 U14647 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U14648 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11761) );
  AOI22_X1 U14649 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11759) );
  AND2_X2 U14650 ( .A1(n9825), .A2(n15689), .ZN(n11751) );
  AOI22_X1 U14651 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14652 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14653 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14654 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  INV_X1 U14655 ( .A(n13203), .ZN(n11877) );
  AOI22_X1 U14656 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12363), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14657 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14658 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14659 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12783), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U14660 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11775) );
  AOI22_X1 U14661 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14662 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11772) );
  INV_X2 U14663 ( .A(n11853), .ZN(n12789) );
  AOI22_X1 U14664 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14665 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11751), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11770) );
  NAND4_X1 U14666 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11774) );
  NOR2_X1 U14667 ( .A1(n11775), .A2(n11774), .ZN(n12388) );
  NOR2_X1 U14668 ( .A1(n11877), .A2(n12388), .ZN(n11776) );
  NAND2_X1 U14669 ( .A1(n16624), .A2(n11776), .ZN(n12282) );
  AOI22_X1 U14670 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14671 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14672 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11887), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11777) );
  NAND4_X1 U14674 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11777), .ZN(
        n11786) );
  AOI22_X1 U14675 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14676 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11751), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11781) );
  NAND4_X1 U14679 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11785) );
  INV_X1 U14680 ( .A(n12394), .ZN(n12281) );
  NAND2_X1 U14681 ( .A1(n12282), .A2(n12281), .ZN(n11787) );
  INV_X1 U14682 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11790) );
  INV_X1 U14683 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11789) );
  OAI22_X1 U14684 ( .A1(n11790), .A2(n11943), .B1(n19536), .B2(n11789), .ZN(
        n11794) );
  INV_X1 U14685 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11792) );
  INV_X1 U14686 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11791) );
  OAI22_X1 U14687 ( .A1(n11792), .A2(n11992), .B1(n19507), .B2(n11791), .ZN(
        n11793) );
  NOR2_X1 U14688 ( .A1(n11794), .A2(n11793), .ZN(n11816) );
  INV_X1 U14689 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11795) );
  OAI22_X1 U14690 ( .A1(n19986), .A2(n19954), .B1(n19754), .B2(n11795), .ZN(
        n11799) );
  INV_X1 U14691 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11797) );
  INV_X1 U14692 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11796) );
  OAI22_X1 U14693 ( .A1(n11797), .A2(n19876), .B1(n19811), .B2(n11796), .ZN(
        n11798) );
  INV_X1 U14694 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11800) );
  NOR2_X1 U14695 ( .A1(n19847), .A2(n11800), .ZN(n11801) );
  NOR2_X1 U14696 ( .A1(n11802), .A2(n11801), .ZN(n11815) );
  INV_X1 U14697 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U14698 ( .A1(n13887), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U14699 ( .A1(n19570), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11803) );
  OAI211_X1 U14700 ( .C1(n19721), .C2(n11805), .A(n11804), .B(n11803), .ZN(
        n11806) );
  INV_X1 U14701 ( .A(n11806), .ZN(n11814) );
  INV_X1 U14702 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11808) );
  INV_X1 U14703 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11807) );
  OAI22_X1 U14704 ( .A1(n11808), .A2(n11941), .B1(n11936), .B2(n11807), .ZN(
        n11812) );
  INV_X1 U14705 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11810) );
  INV_X1 U14706 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11809) );
  OAI22_X1 U14707 ( .A1(n11810), .A2(n19916), .B1(n19783), .B2(n11809), .ZN(
        n11811) );
  NOR2_X1 U14708 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  NAND4_X1 U14709 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11830) );
  AOI22_X1 U14710 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12731), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14711 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12783), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14712 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11892), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14714 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11827) );
  AOI22_X1 U14715 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14716 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11751), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14717 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12500), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14718 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11769), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U14719 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11826) );
  INV_X1 U14720 ( .A(n12402), .ZN(n11828) );
  NAND2_X1 U14721 ( .A1(n11828), .A2(n16624), .ZN(n11829) );
  AOI22_X1 U14722 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14723 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11838) );
  INV_X1 U14724 ( .A(n11832), .ZN(n11834) );
  INV_X1 U14725 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11833) );
  OR2_X1 U14726 ( .A1(n11834), .A2(n11833), .ZN(n11837) );
  INV_X1 U14727 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11835) );
  OR2_X1 U14728 ( .A1(n9880), .A2(n11835), .ZN(n11836) );
  NAND4_X1 U14729 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11843) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19498) );
  INV_X1 U14731 ( .A(n11892), .ZN(n11841) );
  INV_X1 U14732 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11840) );
  OAI22_X1 U14733 ( .A1(n19498), .A2(n11841), .B1(n12368), .B2(n11840), .ZN(
        n11842) );
  NOR2_X1 U14734 ( .A1(n11843), .A2(n11842), .ZN(n11859) );
  NAND2_X1 U14735 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11847) );
  NAND2_X1 U14736 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U14737 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U14738 ( .A1(n11762), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11844) );
  INV_X1 U14739 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11851) );
  INV_X1 U14740 ( .A(n11887), .ZN(n11850) );
  INV_X1 U14741 ( .A(n11848), .ZN(n11849) );
  INV_X1 U14742 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12925) );
  OAI22_X1 U14743 ( .A1(n11851), .A2(n11850), .B1(n11849), .B2(n12925), .ZN(
        n11856) );
  INV_X1 U14744 ( .A(n12363), .ZN(n11854) );
  INV_X1 U14745 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11852) );
  OAI22_X1 U14746 ( .A1(n20018), .A2(n11854), .B1(n11853), .B2(n11852), .ZN(
        n11855) );
  NOR2_X1 U14747 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  AND3_X2 U14748 ( .A1(n11859), .A2(n11858), .A3(n11857), .ZN(n15119) );
  MUX2_X1 U14749 ( .A(n12388), .B(P2_EBX_REG_1__SCAN_IN), .S(n11860), .Z(
        n11861) );
  NOR2_X1 U14750 ( .A1(n13885), .A2(n11650), .ZN(n11879) );
  NAND2_X1 U14751 ( .A1(n20141), .A2(n12394), .ZN(n11867) );
  MUX2_X1 U14752 ( .A(n11863), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12134) );
  NAND2_X1 U14753 ( .A1(n12134), .A2(n12135), .ZN(n11865) );
  NAND2_X1 U14754 ( .A1(n11863), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U14755 ( .A1(n11865), .A2(n11864), .ZN(n11870) );
  XNOR2_X1 U14756 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11869) );
  INV_X1 U14757 ( .A(n11869), .ZN(n11866) );
  XNOR2_X1 U14758 ( .A(n11870), .B(n11866), .ZN(n12260) );
  NAND2_X1 U14759 ( .A1(n9789), .A2(n12260), .ZN(n12262) );
  NAND2_X1 U14760 ( .A1(n11867), .A2(n12262), .ZN(n12147) );
  INV_X1 U14761 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11868) );
  MUX2_X1 U14762 ( .A(n12147), .B(n11868), .S(n11860), .Z(n11883) );
  NAND2_X1 U14763 ( .A1(n11870), .A2(n11869), .ZN(n11872) );
  NAND2_X1 U14764 ( .A1(n20121), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11871) );
  MUX2_X1 U14765 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20114), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11900) );
  XNOR2_X1 U14766 ( .A(n11899), .B(n11900), .ZN(n12132) );
  MUX2_X1 U14767 ( .A(n12402), .B(n12132), .S(n9789), .Z(n12150) );
  INV_X1 U14768 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13798) );
  OAI21_X1 U14769 ( .B1(n11874), .B2(n11873), .A(n11907), .ZN(n13794) );
  INV_X1 U14770 ( .A(n12135), .ZN(n11876) );
  NAND2_X1 U14771 ( .A1(n13861), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U14772 ( .A1(n11876), .A2(n11875), .ZN(n12256) );
  MUX2_X1 U14773 ( .A(n11877), .B(n12256), .S(n9789), .Z(n12149) );
  INV_X1 U14774 ( .A(n11879), .ZN(n11878) );
  OAI21_X1 U14775 ( .B1(n12149), .B2(n11860), .A(n11878), .ZN(n19338) );
  NAND2_X1 U14776 ( .A1(n19338), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13201) );
  INV_X1 U14777 ( .A(n11884), .ZN(n11881) );
  NAND2_X1 U14778 ( .A1(n11879), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U14779 ( .A1(n11881), .A2(n11880), .ZN(n13946) );
  NOR2_X1 U14780 ( .A1(n13201), .A2(n13946), .ZN(n11882) );
  NAND2_X1 U14781 ( .A1(n13201), .A2(n13946), .ZN(n13189) );
  OAI21_X1 U14782 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11882), .A(
        n13189), .ZN(n13186) );
  XNOR2_X1 U14783 ( .A(n11884), .B(n11883), .ZN(n11885) );
  INV_X1 U14784 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12617) );
  XNOR2_X1 U14785 ( .A(n11885), .B(n12617), .ZN(n13185) );
  OR2_X1 U14786 ( .A1(n13186), .A2(n13185), .ZN(n13302) );
  INV_X1 U14787 ( .A(n11885), .ZN(n13919) );
  NAND2_X1 U14788 ( .A1(n13919), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U14789 ( .A1(n13302), .A2(n11886), .ZN(n13636) );
  AOI22_X1 U14790 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14791 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14792 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11887), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14793 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14794 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11898) );
  AOI22_X1 U14795 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14796 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11751), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14797 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14798 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11893) );
  NAND4_X1 U14799 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  NAND3_X1 U14800 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12131), .A3(
        n15830), .ZN(n12133) );
  MUX2_X1 U14801 ( .A(n12407), .B(n12133), .S(n9789), .Z(n11903) );
  INV_X1 U14802 ( .A(n11903), .ZN(n12153) );
  MUX2_X1 U14803 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n12153), .S(n13885), .Z(
        n11906) );
  XNOR2_X1 U14804 ( .A(n11906), .B(n11907), .ZN(n11904) );
  XNOR2_X1 U14805 ( .A(n11904), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13698) );
  INV_X1 U14806 ( .A(n11904), .ZN(n13764) );
  NAND2_X1 U14807 ( .A1(n13764), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11905) );
  INV_X1 U14808 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19323) );
  AOI22_X1 U14809 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14810 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14811 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14812 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14813 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U14814 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14815 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14816 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14817 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U14818 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  MUX2_X1 U14819 ( .A(n19323), .B(n12411), .S(n13885), .Z(n11918) );
  INV_X1 U14820 ( .A(n12019), .ZN(n11920) );
  NAND2_X1 U14821 ( .A1(n10232), .A2(n10235), .ZN(n11919) );
  NAND2_X1 U14822 ( .A1(n11920), .A2(n11919), .ZN(n19320) );
  AND2_X1 U14823 ( .A1(n19320), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11957) );
  INV_X1 U14824 ( .A(n11957), .ZN(n11956) );
  INV_X1 U14825 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12295) );
  AND2_X1 U14826 ( .A1(n15119), .A2(n12295), .ZN(n11958) );
  INV_X1 U14827 ( .A(n11958), .ZN(n11955) );
  INV_X1 U14828 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11922) );
  INV_X1 U14829 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11921) );
  OAI22_X1 U14830 ( .A1(n11922), .A2(n19876), .B1(n19754), .B2(n11921), .ZN(
        n11925) );
  INV_X1 U14831 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11923) );
  OAI22_X1 U14832 ( .A1(n20000), .A2(n19954), .B1(n19811), .B2(n11923), .ZN(
        n11924) );
  OR2_X1 U14833 ( .A1(n11925), .A2(n11924), .ZN(n11928) );
  INV_X1 U14834 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11926) );
  NOR2_X1 U14835 ( .A1(n19721), .A2(n11926), .ZN(n11927) );
  NOR2_X1 U14836 ( .A1(n11928), .A2(n11927), .ZN(n11951) );
  INV_X1 U14837 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11930) );
  INV_X1 U14838 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11929) );
  OAI22_X1 U14839 ( .A1(n11930), .A2(n19507), .B1(n19536), .B2(n11929), .ZN(
        n11934) );
  INV_X1 U14840 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11932) );
  INV_X1 U14841 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11931) );
  OAI22_X1 U14842 ( .A1(n11932), .A2(n19916), .B1(n19783), .B2(n11931), .ZN(
        n11933) );
  NOR2_X1 U14843 ( .A1(n11934), .A2(n11933), .ZN(n11950) );
  INV_X1 U14844 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11935) );
  INV_X1 U14845 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13893) );
  OAI22_X1 U14846 ( .A1(n11935), .A2(n11992), .B1(n11979), .B2(n13893), .ZN(
        n11940) );
  INV_X1 U14847 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11938) );
  INV_X1 U14848 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11937) );
  OAI22_X1 U14849 ( .A1(n11938), .A2(n11936), .B1(n11980), .B2(n11937), .ZN(
        n11939) );
  NOR2_X1 U14850 ( .A1(n11940), .A2(n11939), .ZN(n11949) );
  INV_X1 U14851 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11946) );
  INV_X1 U14852 ( .A(n11941), .ZN(n11942) );
  NAND2_X1 U14853 ( .A1(n11942), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U14854 ( .A1(n19634), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11944) );
  OAI211_X1 U14855 ( .C1(n19847), .C2(n11946), .A(n11945), .B(n11944), .ZN(
        n11947) );
  INV_X1 U14856 ( .A(n11947), .ZN(n11948) );
  NAND4_X1 U14857 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11954) );
  INV_X1 U14858 ( .A(n12411), .ZN(n11952) );
  NAND2_X1 U14859 ( .A1(n11952), .A2(n16624), .ZN(n11953) );
  INV_X2 U14860 ( .A(n11969), .ZN(n11964) );
  MUX2_X1 U14861 ( .A(n11956), .B(n11955), .S(n11964), .Z(n11963) );
  MUX2_X1 U14862 ( .A(n11958), .B(n11957), .S(n11964), .Z(n11959) );
  NAND2_X1 U14863 ( .A1(n11965), .A2(n11959), .ZN(n11962) );
  OAI21_X1 U14864 ( .B1(n15119), .B2(n12295), .A(n19320), .ZN(n11960) );
  OAI21_X1 U14865 ( .B1(n12295), .B2(n19320), .A(n11960), .ZN(n11961) );
  OAI211_X1 U14866 ( .C1(n11965), .C2(n11963), .A(n11962), .B(n11961), .ZN(
        n13835) );
  OAI21_X1 U14867 ( .B1(n12296), .B2(n15120), .A(n19320), .ZN(n11966) );
  NAND2_X1 U14868 ( .A1(n11966), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U14869 ( .A1(n11968), .A2(n11967), .ZN(n15650) );
  NAND2_X1 U14870 ( .A1(n11970), .A2(n11969), .ZN(n12016) );
  INV_X1 U14871 ( .A(n12016), .ZN(n12014) );
  INV_X1 U14872 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U14873 ( .A1(n11971), .A2(n19876), .B1(n19954), .B2(n20007), .ZN(
        n11975) );
  INV_X1 U14874 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11973) );
  INV_X1 U14875 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11972) );
  OAI22_X1 U14876 ( .A1(n11973), .A2(n19754), .B1(n19811), .B2(n11972), .ZN(
        n11974) );
  OR2_X1 U14877 ( .A1(n11975), .A2(n11974), .ZN(n11978) );
  INV_X1 U14878 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11976) );
  NOR2_X1 U14879 ( .A1(n19721), .A2(n11976), .ZN(n11977) );
  NOR2_X1 U14880 ( .A1(n11978), .A2(n11977), .ZN(n12000) );
  INV_X1 U14881 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11981) );
  INV_X1 U14882 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n21331) );
  OAI22_X1 U14883 ( .A1(n11981), .A2(n11980), .B1(n11979), .B2(n21331), .ZN(
        n11985) );
  INV_X1 U14884 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11983) );
  INV_X1 U14885 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11982) );
  OAI22_X1 U14886 ( .A1(n11983), .A2(n19916), .B1(n19783), .B2(n11982), .ZN(
        n11984) );
  NOR2_X1 U14887 ( .A1(n11985), .A2(n11984), .ZN(n11999) );
  INV_X1 U14888 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11987) );
  INV_X1 U14889 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11986) );
  OAI22_X1 U14890 ( .A1(n11987), .A2(n11941), .B1(n11936), .B2(n11986), .ZN(
        n11991) );
  INV_X1 U14891 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11989) );
  INV_X1 U14892 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11988) );
  OAI22_X1 U14893 ( .A1(n11989), .A2(n11943), .B1(n19536), .B2(n11988), .ZN(
        n11990) );
  NOR2_X1 U14894 ( .A1(n11991), .A2(n11990), .ZN(n11998) );
  INV_X1 U14895 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11995) );
  INV_X1 U14896 ( .A(n19507), .ZN(n19502) );
  NAND2_X1 U14897 ( .A1(n19502), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11994) );
  NAND2_X1 U14898 ( .A1(n19603), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11993) );
  OAI211_X1 U14899 ( .C1(n19847), .C2(n11995), .A(n11994), .B(n11993), .ZN(
        n11996) );
  INV_X1 U14900 ( .A(n11996), .ZN(n11997) );
  NAND4_X1 U14901 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12013) );
  AOI22_X1 U14902 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U14903 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U14904 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11887), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U14905 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12789), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12001) );
  NAND4_X1 U14906 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12010) );
  AOI22_X1 U14907 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U14908 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11751), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U14909 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U14910 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U14911 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12009) );
  INV_X1 U14912 ( .A(n12414), .ZN(n12011) );
  NAND2_X1 U14913 ( .A1(n12011), .A2(n16624), .ZN(n12012) );
  INV_X1 U14914 ( .A(n12298), .ZN(n12015) );
  NAND2_X1 U14915 ( .A1(n12016), .A2(n12015), .ZN(n12017) );
  INV_X1 U14916 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19308) );
  MUX2_X1 U14917 ( .A(n19308), .B(n12414), .S(n13885), .Z(n12018) );
  NAND2_X2 U14918 ( .A1(n12019), .A2(n12018), .ZN(n12027) );
  OAI21_X1 U14919 ( .B1(n12019), .B2(n12018), .A(n12027), .ZN(n19307) );
  INV_X1 U14920 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15644) );
  XNOR2_X1 U14921 ( .A(n12020), .B(n15644), .ZN(n15652) );
  NAND2_X1 U14922 ( .A1(n15650), .A2(n15652), .ZN(n12022) );
  NAND2_X1 U14923 ( .A1(n12020), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12021) );
  MUX2_X1 U14924 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n9750), .S(n13885), .Z(n12026) );
  NAND2_X1 U14925 ( .A1(n11860), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12023) );
  OR2_X1 U14926 ( .A1(n12033), .A2(n12023), .ZN(n12024) );
  AND2_X1 U14927 ( .A1(n12032), .A2(n12024), .ZN(n12028) );
  INV_X1 U14928 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16579) );
  NOR2_X1 U14929 ( .A1(n15119), .A2(n16579), .ZN(n12025) );
  NAND2_X1 U14930 ( .A1(n12028), .A2(n12025), .ZN(n16535) );
  XNOR2_X1 U14931 ( .A(n12027), .B(n10253), .ZN(n19297) );
  NAND2_X1 U14932 ( .A1(n19297), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16533) );
  INV_X1 U14933 ( .A(n12028), .ZN(n13787) );
  OAI21_X1 U14934 ( .B1(n13787), .B2(n15119), .A(n16579), .ZN(n16536) );
  INV_X1 U14935 ( .A(n19297), .ZN(n12029) );
  INV_X1 U14936 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16569) );
  NAND2_X1 U14937 ( .A1(n12029), .A2(n16569), .ZN(n15322) );
  AND2_X1 U14938 ( .A1(n16536), .A2(n15322), .ZN(n12030) );
  NAND2_X1 U14939 ( .A1(n11860), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12031) );
  XNOR2_X1 U14940 ( .A(n12032), .B(n12031), .ZN(n19286) );
  AOI21_X1 U14941 ( .B1(n19286), .B2(n15120), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15617) );
  NAND3_X1 U14942 ( .A1(n12039), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n11860), 
        .ZN(n12034) );
  OAI211_X1 U14943 ( .C1(n12039), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12034), .B(
        n12122), .ZN(n19273) );
  OR2_X1 U14944 ( .A1(n19273), .A2(n15119), .ZN(n12035) );
  INV_X1 U14945 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U14946 ( .A1(n12035), .A2(n15610), .ZN(n15607) );
  OR2_X1 U14947 ( .A1(n15119), .A2(n15610), .ZN(n12036) );
  OR2_X1 U14948 ( .A1(n19273), .A2(n12036), .ZN(n15606) );
  INV_X1 U14949 ( .A(n19286), .ZN(n12037) );
  INV_X1 U14950 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15576) );
  OR3_X1 U14951 ( .A1(n12037), .A2(n15119), .A3(n15576), .ZN(n15604) );
  AND2_X1 U14952 ( .A1(n15606), .A2(n15604), .ZN(n12038) );
  INV_X1 U14953 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13669) );
  INV_X1 U14954 ( .A(n12040), .ZN(n12041) );
  NAND2_X1 U14955 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12041), .ZN(n12042) );
  NOR2_X1 U14956 ( .A1(n13885), .A2(n12042), .ZN(n12043) );
  OR2_X1 U14957 ( .A1(n12047), .A2(n12043), .ZN(n19260) );
  OR2_X1 U14958 ( .A1(n19260), .A2(n15119), .ZN(n15310) );
  INV_X1 U14959 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U14960 ( .A1(n11860), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12049) );
  OR2_X1 U14961 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  NAND2_X1 U14962 ( .A1(n12053), .A2(n12050), .ZN(n19251) );
  INV_X1 U14963 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15298) );
  INV_X1 U14964 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12051) );
  NOR2_X1 U14965 ( .A1(n13885), .A2(n12051), .ZN(n12052) );
  NAND2_X1 U14966 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  NAND2_X1 U14967 ( .A1(n12081), .A2(n12054), .ZN(n19239) );
  OR2_X1 U14968 ( .A1(n19239), .A2(n15119), .ZN(n12055) );
  INV_X1 U14969 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21229) );
  NAND2_X1 U14970 ( .A1(n12055), .A2(n21229), .ZN(n15284) );
  OR2_X1 U14971 ( .A1(n19251), .A2(n15119), .ZN(n12056) );
  NAND2_X1 U14972 ( .A1(n12056), .A2(n15298), .ZN(n15295) );
  AND2_X1 U14973 ( .A1(n15284), .A2(n15295), .ZN(n12057) );
  INV_X1 U14974 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12203) );
  NOR2_X1 U14975 ( .A1(n13885), .A2(n12203), .ZN(n12079) );
  NOR2_X2 U14976 ( .A1(n12081), .A2(n12079), .ZN(n12072) );
  NAND2_X1 U14977 ( .A1(n11860), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12070) );
  NAND2_X1 U14978 ( .A1(n12072), .A2(n12070), .ZN(n12085) );
  INV_X1 U14979 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19355) );
  NOR2_X1 U14980 ( .A1(n13885), .A2(n19355), .ZN(n12084) );
  OR2_X2 U14981 ( .A1(n12085), .A2(n12084), .ZN(n12075) );
  INV_X1 U14982 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12058) );
  NOR2_X1 U14983 ( .A1(n13885), .A2(n12058), .ZN(n12074) );
  OR2_X2 U14984 ( .A1(n12075), .A2(n12074), .ZN(n12077) );
  INV_X1 U14985 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12059) );
  NOR2_X1 U14986 ( .A1(n13885), .A2(n12059), .ZN(n12067) );
  OR2_X2 U14987 ( .A1(n12077), .A2(n12067), .ZN(n12069) );
  INV_X1 U14988 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12060) );
  NOR2_X1 U14989 ( .A1(n13885), .A2(n12060), .ZN(n12065) );
  INV_X1 U14990 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12061) );
  AND3_X1 U14991 ( .A1(n12062), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11860), .ZN(
        n12063) );
  NOR2_X1 U14992 ( .A1(n12106), .A2(n12063), .ZN(n12983) );
  NAND2_X1 U14993 ( .A1(n12983), .A2(n15120), .ZN(n12064) );
  INV_X1 U14994 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15442) );
  NAND2_X1 U14995 ( .A1(n12064), .A2(n15442), .ZN(n15205) );
  AND2_X1 U14996 ( .A1(n12069), .A2(n12065), .ZN(n12066) );
  NOR2_X1 U14997 ( .A1(n12089), .A2(n12066), .ZN(n19200) );
  NAND2_X1 U14998 ( .A1(n19200), .A2(n15120), .ZN(n12093) );
  INV_X1 U14999 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15455) );
  NAND2_X1 U15000 ( .A1(n12093), .A2(n15455), .ZN(n15231) );
  NAND2_X1 U15001 ( .A1(n12077), .A2(n12067), .ZN(n12068) );
  NAND2_X1 U15002 ( .A1(n12069), .A2(n12068), .ZN(n12094) );
  INV_X1 U15003 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15246) );
  OAI21_X1 U15004 ( .B1(n12094), .B2(n15119), .A(n15246), .ZN(n15242) );
  INV_X1 U15005 ( .A(n12070), .ZN(n12071) );
  XNOR2_X1 U15006 ( .A(n12072), .B(n12071), .ZN(n19230) );
  NAND2_X1 U15007 ( .A1(n19230), .A2(n15120), .ZN(n12073) );
  INV_X1 U15008 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15525) );
  NAND2_X1 U15009 ( .A1(n12073), .A2(n15525), .ZN(n15274) );
  NAND2_X1 U15010 ( .A1(n12075), .A2(n12074), .ZN(n12076) );
  NAND2_X1 U15011 ( .A1(n12077), .A2(n12076), .ZN(n19206) );
  OR2_X1 U15012 ( .A1(n19206), .A2(n15119), .ZN(n12078) );
  INV_X1 U15013 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15014 ( .A1(n12078), .A2(n12310), .ZN(n15211) );
  INV_X1 U15015 ( .A(n12079), .ZN(n12080) );
  XNOR2_X1 U15016 ( .A(n12081), .B(n12080), .ZN(n13854) );
  NAND2_X1 U15017 ( .A1(n13854), .A2(n15120), .ZN(n12082) );
  INV_X1 U15018 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12097) );
  NAND2_X1 U15019 ( .A1(n12082), .A2(n12097), .ZN(n15536) );
  AND4_X1 U15020 ( .A1(n15242), .A2(n15274), .A3(n15211), .A4(n15536), .ZN(
        n12083) );
  AND2_X1 U15021 ( .A1(n15231), .A2(n12083), .ZN(n12091) );
  INV_X1 U15022 ( .A(n12084), .ZN(n12086) );
  MUX2_X1 U15023 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n12086), .S(n12085), .Z(
        n12087) );
  NAND2_X1 U15024 ( .A1(n12087), .A2(n12122), .ZN(n19219) );
  OR2_X1 U15025 ( .A1(n19219), .A2(n15119), .ZN(n12096) );
  XNOR2_X1 U15026 ( .A(n12096), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15261) );
  NOR2_X1 U15027 ( .A1(n13885), .A2(n12061), .ZN(n12088) );
  XNOR2_X1 U15028 ( .A(n12089), .B(n12088), .ZN(n14931) );
  NAND2_X1 U15029 ( .A1(n14931), .A2(n15120), .ZN(n12090) );
  INV_X1 U15030 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15202) );
  NAND2_X1 U15031 ( .A1(n12090), .A2(n15202), .ZN(n15222) );
  NOR2_X1 U15032 ( .A1(n15119), .A2(n15442), .ZN(n12092) );
  NAND2_X1 U15033 ( .A1(n12983), .A2(n12092), .ZN(n15204) );
  OR2_X1 U15034 ( .A1(n12093), .A2(n15455), .ZN(n15232) );
  INV_X1 U15035 ( .A(n12094), .ZN(n14944) );
  NOR2_X1 U15036 ( .A1(n15119), .A2(n15246), .ZN(n12095) );
  NAND2_X1 U15037 ( .A1(n14944), .A2(n12095), .ZN(n15241) );
  AND2_X1 U15038 ( .A1(n15232), .A2(n15241), .ZN(n15213) );
  INV_X1 U15039 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21194) );
  OR2_X1 U15040 ( .A1(n12096), .A2(n21194), .ZN(n15208) );
  NOR2_X1 U15041 ( .A1(n15119), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U15042 ( .A1(n13854), .A2(n12098), .ZN(n15535) );
  OR2_X1 U15043 ( .A1(n15119), .A2(n21229), .ZN(n12099) );
  AND2_X1 U15044 ( .A1(n15535), .A2(n15283), .ZN(n12103) );
  INV_X1 U15045 ( .A(n19230), .ZN(n12100) );
  INV_X1 U15046 ( .A(n19206), .ZN(n12102) );
  NOR2_X1 U15047 ( .A1(n15119), .A2(n12310), .ZN(n12101) );
  NAND2_X1 U15048 ( .A1(n12102), .A2(n12101), .ZN(n15210) );
  AND4_X1 U15049 ( .A1(n15208), .A2(n12103), .A3(n15273), .A4(n15210), .ZN(
        n12105) );
  NOR2_X1 U15050 ( .A1(n15119), .A2(n15202), .ZN(n12104) );
  NAND2_X1 U15051 ( .A1(n14931), .A2(n12104), .ZN(n15221) );
  NAND2_X1 U15052 ( .A1(n11860), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12107) );
  INV_X1 U15053 ( .A(n12107), .ZN(n12108) );
  NAND2_X1 U15054 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  AND2_X1 U15055 ( .A1(n12115), .A2(n12110), .ZN(n13015) );
  NAND2_X1 U15056 ( .A1(n13015), .A2(n15120), .ZN(n12111) );
  INV_X1 U15057 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15430) );
  AND2_X1 U15058 ( .A1(n12111), .A2(n15430), .ZN(n15425) );
  INV_X1 U15059 ( .A(n12111), .ZN(n12112) );
  NAND2_X1 U15060 ( .A1(n12112), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15426) );
  INV_X1 U15061 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12113) );
  NOR2_X1 U15062 ( .A1(n13885), .A2(n12113), .ZN(n12114) );
  NOR2_X2 U15063 ( .A1(n12115), .A2(n12114), .ZN(n16468) );
  AND2_X1 U15064 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  NOR2_X1 U15065 ( .A1(n16468), .A2(n12116), .ZN(n12997) );
  NAND2_X1 U15066 ( .A1(n12997), .A2(n15120), .ZN(n12117) );
  XNOR2_X1 U15067 ( .A(n12117), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15195) );
  INV_X1 U15068 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12231) );
  NOR2_X1 U15069 ( .A1(n15119), .A2(n12231), .ZN(n12118) );
  INV_X1 U15070 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21149) );
  NAND2_X1 U15071 ( .A1(n12122), .A2(n15120), .ZN(n15181) );
  INV_X1 U15072 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16471) );
  AND2_X2 U15073 ( .A1(n16468), .A2(n16471), .ZN(n12121) );
  INV_X1 U15074 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14982) );
  NOR2_X1 U15075 ( .A1(n12121), .A2(n14982), .ZN(n12119) );
  NAND2_X1 U15076 ( .A1(n11860), .A2(n12119), .ZN(n12120) );
  AOI21_X1 U15077 ( .B1(n14915), .B2(n15120), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U15078 ( .A1(n12121), .A2(n14982), .ZN(n16455) );
  OR2_X2 U15079 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16455), .ZN(n16438) );
  NAND2_X2 U15080 ( .A1(n12122), .A2(n16438), .ZN(n16454) );
  NOR2_X1 U15081 ( .A1(n16454), .A2(n15119), .ZN(n12123) );
  XOR2_X1 U15082 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n12123), .Z(
        n15162) );
  INV_X1 U15083 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15397) );
  AOI21_X1 U15084 ( .B1(n12123), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15170), .ZN(n15111) );
  NAND2_X1 U15085 ( .A1(n11860), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16441) );
  NAND2_X1 U15086 ( .A1(n16439), .A2(n15120), .ZN(n15106) );
  NAND2_X1 U15087 ( .A1(n15154), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15155) );
  INV_X1 U15088 ( .A(n12124), .ZN(n12125) );
  INV_X1 U15089 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12249) );
  NOR2_X1 U15090 ( .A1(n13885), .A2(n12249), .ZN(n12126) );
  NAND2_X1 U15091 ( .A1(n16439), .A2(n12126), .ZN(n12127) );
  NAND2_X1 U15092 ( .A1(n15115), .A2(n12127), .ZN(n14899) );
  XNOR2_X1 U15093 ( .A(n15109), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12128) );
  NOR2_X1 U15094 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16074), .ZN(
        n12130) );
  INV_X1 U15095 ( .A(n12134), .ZN(n12257) );
  XNOR2_X1 U15096 ( .A(n12257), .B(n12135), .ZN(n12254) );
  NAND2_X1 U15097 ( .A1(n12260), .A2(n12254), .ZN(n12136) );
  NOR2_X1 U15098 ( .A1(n12268), .A2(n12136), .ZN(n12137) );
  OR2_X1 U15099 ( .A1(n12271), .A2(n12137), .ZN(n16616) );
  INV_X1 U15100 ( .A(n12256), .ZN(n12138) );
  NAND2_X1 U15101 ( .A1(n12260), .A2(n12138), .ZN(n12139) );
  OAI21_X1 U15102 ( .B1(n12268), .B2(n12139), .A(n15656), .ZN(n12140) );
  OR2_X1 U15103 ( .A1(n16616), .A2(n12140), .ZN(n12146) );
  INV_X1 U15104 ( .A(n12142), .ZN(n15685) );
  NAND2_X1 U15105 ( .A1(n12142), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12143) );
  NAND2_X1 U15106 ( .A1(n12143), .A2(n15830), .ZN(n16623) );
  INV_X1 U15107 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12144) );
  OAI21_X1 U15108 ( .B1(n12141), .B2(n16623), .A(n12144), .ZN(n12145) );
  NAND2_X1 U15109 ( .A1(n12145), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20131) );
  NAND2_X1 U15110 ( .A1(n12146), .A2(n20131), .ZN(n16596) );
  NAND2_X1 U15111 ( .A1(n16596), .A2(n20155), .ZN(n12157) );
  INV_X1 U15112 ( .A(n12147), .ZN(n12148) );
  OAI21_X1 U15113 ( .B1(n12149), .B2(n12257), .A(n12148), .ZN(n12151) );
  NAND2_X1 U15114 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  NOR2_X1 U15115 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  OR2_X1 U15116 ( .A1(n12154), .A2(n12271), .ZN(n20139) );
  INV_X1 U15117 ( .A(n20139), .ZN(n12155) );
  NAND2_X1 U15118 ( .A1(n16624), .A2(n12576), .ZN(n12544) );
  NAND2_X1 U15119 ( .A1(n12155), .A2(n20140), .ZN(n12156) );
  NAND2_X1 U15120 ( .A1(n12157), .A2(n12156), .ZN(n12592) );
  NAND2_X1 U15121 ( .A1(n15656), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12550) );
  NOR2_X1 U15122 ( .A1(n20143), .A2(n13874), .ZN(n12158) );
  NAND2_X1 U15123 ( .A1(n12592), .A2(n12158), .ZN(n12313) );
  INV_X1 U15124 ( .A(n12313), .ZN(n12159) );
  NAND2_X1 U15125 ( .A1(n12599), .A2(n16549), .ZN(n12317) );
  NOR2_X1 U15126 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20021) );
  OR2_X1 U15127 ( .A1(n20102), .A2(n20021), .ZN(n20122) );
  NAND2_X1 U15128 ( .A1(n20122), .A2(n21322), .ZN(n12160) );
  INV_X1 U15129 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20153) );
  NAND2_X1 U15130 ( .A1(n20153), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12161) );
  NAND2_X1 U15131 ( .A1(n12253), .A2(n12161), .ZN(n14079) );
  INV_X1 U15132 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12163) );
  AND2_X2 U15133 ( .A1(n12337), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12351) );
  NOR2_X2 U15134 ( .A1(n12332), .A2(n15215), .ZN(n12331) );
  NAND2_X1 U15135 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n12331), .ZN(
        n12329) );
  INV_X1 U15136 ( .A(n12329), .ZN(n12162) );
  AND2_X2 U15137 ( .A1(n12162), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12330) );
  INV_X1 U15138 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15175) );
  INV_X1 U15139 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21232) );
  AOI21_X1 U15140 ( .B1(n12163), .B2(n12325), .A(n12322), .ZN(n14895) );
  NAND2_X1 U15141 ( .A1(n20102), .A2(n15656), .ZN(n19165) );
  NAND2_X1 U15142 ( .A1(n19326), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12643) );
  OAI21_X1 U15143 ( .B1(n16565), .B2(n12163), .A(n12643), .ZN(n12275) );
  INV_X1 U15144 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12290) );
  OR2_X1 U15145 ( .A1(n12244), .A2(n12290), .ZN(n12170) );
  NAND2_X1 U15146 ( .A1(n14870), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15147 ( .A1(n14869), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12167) );
  AND2_X1 U15148 ( .A1(n12168), .A2(n12167), .ZN(n12169) );
  NAND2_X1 U15149 ( .A1(n12170), .A2(n12169), .ZN(n13700) );
  OR2_X1 U15150 ( .A1(n12244), .A2(n12295), .ZN(n12174) );
  NAND2_X1 U15151 ( .A1(n14870), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15152 ( .A1(n14869), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12171) );
  AND2_X1 U15153 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  OR2_X1 U15154 ( .A1(n14873), .A2(n15644), .ZN(n12179) );
  NAND2_X1 U15155 ( .A1(n14870), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15156 ( .A1(n14869), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12176) );
  AND2_X1 U15157 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U15158 ( .A1(n12179), .A2(n12178), .ZN(n13396) );
  OR2_X1 U15159 ( .A1(n14873), .A2(n16569), .ZN(n12183) );
  NAND2_X1 U15160 ( .A1(n14870), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15161 ( .A1(n14869), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12180) );
  AND2_X1 U15162 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  AOI22_X1 U15163 ( .A1(n14869), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12185) );
  NAND2_X1 U15164 ( .A1(n14870), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12184) );
  OAI211_X1 U15165 ( .C1(n14873), .C2(n16579), .A(n12185), .B(n12184), .ZN(
        n13776) );
  NAND2_X1 U15166 ( .A1(n13775), .A2(n13776), .ZN(n13774) );
  INV_X1 U15167 ( .A(n13774), .ZN(n13522) );
  OR2_X1 U15168 ( .A1(n14873), .A2(n15576), .ZN(n12189) );
  NAND2_X1 U15169 ( .A1(n14870), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15170 ( .A1(n14869), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12186) );
  AND2_X1 U15171 ( .A1(n12187), .A2(n12186), .ZN(n12188) );
  NAND2_X1 U15172 ( .A1(n12189), .A2(n12188), .ZN(n13523) );
  NAND2_X1 U15173 ( .A1(n13522), .A2(n13523), .ZN(n15593) );
  AOI22_X1 U15174 ( .A1(n14869), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12190) );
  OAI21_X1 U15175 ( .B1(n12175), .B2(n10247), .A(n12190), .ZN(n12191) );
  AOI21_X1 U15176 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12191), .ZN(n15592) );
  OR2_X1 U15177 ( .A1(n14873), .A2(n12045), .ZN(n12194) );
  INV_X1 U15178 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15313) );
  OAI22_X1 U15179 ( .A1(n12559), .A2(n15313), .B1(n15656), .B2(n19263), .ZN(
        n12192) );
  AOI21_X1 U15180 ( .B1(n14870), .B2(P2_EBX_REG_11__SCAN_IN), .A(n12192), .ZN(
        n12193) );
  OR2_X1 U15181 ( .A1(n14873), .A2(n15298), .ZN(n12198) );
  INV_X1 U15182 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20066) );
  INV_X1 U15183 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12195) );
  OAI22_X1 U15184 ( .A1(n12559), .A2(n20066), .B1(n15656), .B2(n12195), .ZN(
        n12196) );
  AOI21_X1 U15185 ( .B1(n14870), .B2(P2_EBX_REG_12__SCAN_IN), .A(n12196), .ZN(
        n12197) );
  NAND2_X1 U15186 ( .A1(n12198), .A2(n12197), .ZN(n15299) );
  OR2_X1 U15187 ( .A1(n14873), .A2(n21229), .ZN(n12201) );
  INV_X1 U15188 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15288) );
  INV_X1 U15189 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15289) );
  OAI22_X1 U15190 ( .A1(n12559), .A2(n15288), .B1(n15656), .B2(n15289), .ZN(
        n12199) );
  AOI21_X1 U15191 ( .B1(n14870), .B2(P2_EBX_REG_13__SCAN_IN), .A(n12199), .ZN(
        n12200) );
  AOI22_X1 U15192 ( .A1(n14869), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12202) );
  OAI21_X1 U15193 ( .B1(n12175), .B2(n12203), .A(n12202), .ZN(n12204) );
  AOI21_X1 U15194 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12204), .ZN(n13844) );
  OR2_X1 U15195 ( .A1(n14873), .A2(n15525), .ZN(n12207) );
  INV_X1 U15196 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15279) );
  OAI22_X1 U15197 ( .A1(n12559), .A2(n15279), .B1(n15656), .B2(n15278), .ZN(
        n12205) );
  AOI21_X1 U15198 ( .B1(n14870), .B2(P2_EBX_REG_15__SCAN_IN), .A(n12205), .ZN(
        n12206) );
  NAND2_X1 U15199 ( .A1(n12207), .A2(n12206), .ZN(n13744) );
  OR2_X1 U15200 ( .A1(n14873), .A2(n21194), .ZN(n12210) );
  INV_X1 U15201 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15513) );
  OAI22_X1 U15202 ( .A1(n12559), .A2(n15513), .B1(n15656), .B2(n10301), .ZN(
        n12208) );
  AOI21_X1 U15203 ( .B1(n14870), .B2(P2_EBX_REG_16__SCAN_IN), .A(n12208), .ZN(
        n12209) );
  NAND2_X1 U15204 ( .A1(n12210), .A2(n12209), .ZN(n15263) );
  OR2_X1 U15205 ( .A1(n14873), .A2(n12310), .ZN(n12213) );
  INV_X1 U15206 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20073) );
  OAI22_X1 U15207 ( .A1(n12559), .A2(n20073), .B1(n15656), .B2(n19203), .ZN(
        n12211) );
  AOI21_X1 U15208 ( .B1(n14870), .B2(P2_EBX_REG_17__SCAN_IN), .A(n12211), .ZN(
        n12212) );
  OR2_X1 U15209 ( .A1(n14873), .A2(n15246), .ZN(n12217) );
  INV_X1 U15210 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20075) );
  INV_X1 U15211 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12214) );
  OAI22_X1 U15212 ( .A1(n12559), .A2(n20075), .B1(n15656), .B2(n12214), .ZN(
        n12215) );
  AOI21_X1 U15213 ( .B1(n14870), .B2(P2_EBX_REG_18__SCAN_IN), .A(n12215), .ZN(
        n12216) );
  OR2_X1 U15214 ( .A1(n14873), .A2(n15455), .ZN(n12220) );
  INV_X1 U15215 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21162) );
  OAI22_X1 U15216 ( .A1(n12559), .A2(n21162), .B1(n15656), .B2(n19191), .ZN(
        n12218) );
  AOI21_X1 U15217 ( .B1(n14870), .B2(P2_EBX_REG_19__SCAN_IN), .A(n12218), .ZN(
        n12219) );
  NAND2_X1 U15218 ( .A1(n12220), .A2(n12219), .ZN(n14997) );
  AOI22_X1 U15219 ( .A1(n14869), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12221) );
  OAI21_X1 U15220 ( .B1(n12175), .B2(n12061), .A(n12221), .ZN(n12222) );
  AOI21_X1 U15221 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12222), .ZN(n14917) );
  OR2_X1 U15222 ( .A1(n14873), .A2(n15442), .ZN(n12226) );
  INV_X1 U15223 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n12223) );
  OAI22_X1 U15224 ( .A1(n12559), .A2(n12223), .B1(n15656), .B2(n15215), .ZN(
        n12224) );
  AOI21_X1 U15225 ( .B1(n14870), .B2(P2_EBX_REG_21__SCAN_IN), .A(n12224), .ZN(
        n12225) );
  INV_X1 U15226 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15227 ( .A1(n14869), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12228) );
  OAI21_X1 U15228 ( .B1(n12175), .B2(n12229), .A(n12228), .ZN(n12230) );
  AOI21_X1 U15229 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12230), .ZN(n13017) );
  OR2_X1 U15230 ( .A1(n14873), .A2(n12231), .ZN(n12235) );
  INV_X1 U15231 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n12232) );
  INV_X1 U15232 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15196) );
  OAI22_X1 U15233 ( .A1(n12559), .A2(n12232), .B1(n15656), .B2(n15196), .ZN(
        n12233) );
  AOI21_X1 U15234 ( .B1(n14870), .B2(P2_EBX_REG_23__SCAN_IN), .A(n12233), .ZN(
        n12234) );
  NAND2_X1 U15235 ( .A1(n12235), .A2(n12234), .ZN(n12999) );
  OR2_X1 U15236 ( .A1(n14873), .A2(n21149), .ZN(n12238) );
  INV_X1 U15237 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20082) );
  OAI22_X1 U15238 ( .A1(n12559), .A2(n20082), .B1(n15656), .B2(n10296), .ZN(
        n12236) );
  AOI21_X1 U15239 ( .B1(n14870), .B2(P2_EBX_REG_24__SCAN_IN), .A(n12236), .ZN(
        n12237) );
  NAND2_X1 U15240 ( .A1(n12238), .A2(n12237), .ZN(n14988) );
  AOI22_X1 U15241 ( .A1(n14869), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12239) );
  OAI21_X1 U15242 ( .B1(n12175), .B2(n14982), .A(n12239), .ZN(n12240) );
  AOI21_X1 U15243 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12240), .ZN(n14904) );
  INV_X1 U15244 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15245 ( .A1(n14869), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12241) );
  OAI21_X1 U15246 ( .B1(n12175), .B2(n12242), .A(n12241), .ZN(n12243) );
  AOI21_X1 U15247 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12243), .ZN(n14974) );
  INV_X1 U15248 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15369) );
  OR2_X1 U15249 ( .A1(n14873), .A2(n15369), .ZN(n12247) );
  INV_X1 U15250 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20087) );
  OAI22_X1 U15251 ( .A1(n12559), .A2(n20087), .B1(n15656), .B2(n21232), .ZN(
        n12245) );
  AOI21_X1 U15252 ( .B1(n14870), .B2(P2_EBX_REG_27__SCAN_IN), .A(n12245), .ZN(
        n12246) );
  NAND2_X1 U15253 ( .A1(n12247), .A2(n12246), .ZN(n14968) );
  AOI22_X1 U15254 ( .A1(n14869), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12248) );
  OAI21_X1 U15255 ( .B1(n12175), .B2(n12249), .A(n12248), .ZN(n12250) );
  AOI21_X1 U15256 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12250), .ZN(n12251) );
  NAND2_X1 U15257 ( .A1(n14967), .A2(n12251), .ZN(n12252) );
  NAND2_X1 U15258 ( .A1(n14948), .A2(n12252), .ZN(n14961) );
  NAND2_X1 U15259 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U15260 ( .A1(n16624), .A2(n12256), .ZN(n12255) );
  AOI22_X1 U15261 ( .A1(n12255), .A2(n12254), .B1(n16624), .B2(n12260), .ZN(
        n12259) );
  OAI21_X1 U15262 ( .B1(n12257), .B2(n12256), .A(n20141), .ZN(n12258) );
  OAI21_X1 U15263 ( .B1(n12259), .B2(n12576), .A(n12258), .ZN(n12265) );
  INV_X1 U15264 ( .A(n12260), .ZN(n12261) );
  OAI21_X1 U15265 ( .B1(n20152), .B2(n16624), .A(n12261), .ZN(n12263) );
  NAND2_X1 U15266 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  NAND2_X1 U15267 ( .A1(n12265), .A2(n12264), .ZN(n12267) );
  NAND2_X1 U15268 ( .A1(n12268), .A2(n20141), .ZN(n12266) );
  OAI21_X1 U15269 ( .B1(n12268), .B2(n12267), .A(n12266), .ZN(n12269) );
  OR2_X1 U15270 ( .A1(n12271), .A2(n12269), .ZN(n12270) );
  MUX2_X1 U15271 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12270), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12571) );
  NAND2_X1 U15272 ( .A1(n12271), .A2(n20152), .ZN(n12272) );
  INV_X1 U15273 ( .A(n13882), .ZN(n16561) );
  NOR2_X1 U15274 ( .A1(n14961), .A2(n13882), .ZN(n12274) );
  AOI211_X1 U15275 ( .C1(n16555), .C2(n14895), .A(n12275), .B(n12274), .ZN(
        n12315) );
  INV_X1 U15276 ( .A(n12276), .ZN(n12301) );
  OR2_X1 U15277 ( .A1(n12276), .A2(n13828), .ZN(n12297) );
  NOR2_X1 U15278 ( .A1(n13203), .A2(n13273), .ZN(n13202) );
  NAND2_X1 U15279 ( .A1(n13202), .A2(n12279), .ZN(n12280) );
  INV_X1 U15280 ( .A(n12388), .ZN(n12279) );
  NOR2_X1 U15281 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13203), .ZN(
        n12278) );
  XNOR2_X1 U15282 ( .A(n12279), .B(n12278), .ZN(n13192) );
  NAND2_X1 U15283 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13192), .ZN(
        n13191) );
  NAND2_X1 U15284 ( .A1(n12280), .A2(n13191), .ZN(n12283) );
  XNOR2_X1 U15285 ( .A(n12617), .B(n12283), .ZN(n13180) );
  XNOR2_X1 U15286 ( .A(n12282), .B(n12281), .ZN(n13178) );
  NAND2_X1 U15287 ( .A1(n13180), .A2(n13178), .ZN(n12285) );
  NAND2_X1 U15288 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12283), .ZN(
        n12284) );
  NAND2_X1 U15289 ( .A1(n12285), .A2(n12284), .ZN(n12286) );
  NAND2_X1 U15290 ( .A1(n12286), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12287) );
  XNOR2_X1 U15291 ( .A(n12289), .B(n12288), .ZN(n12291) );
  XNOR2_X1 U15292 ( .A(n12292), .B(n12291), .ZN(n13694) );
  NAND2_X1 U15293 ( .A1(n13694), .A2(n12290), .ZN(n13695) );
  INV_X1 U15294 ( .A(n12291), .ZN(n12293) );
  OR2_X1 U15295 ( .A1(n12293), .A2(n12292), .ZN(n12294) );
  NAND2_X1 U15296 ( .A1(n13695), .A2(n12294), .ZN(n13825) );
  NAND2_X1 U15297 ( .A1(n13829), .A2(n12300), .ZN(n12302) );
  NAND2_X1 U15298 ( .A1(n12302), .A2(n12301), .ZN(n12303) );
  NAND2_X1 U15299 ( .A1(n9772), .A2(n15119), .ZN(n12305) );
  NAND2_X1 U15300 ( .A1(n12306), .A2(n12305), .ZN(n15318) );
  INV_X1 U15301 ( .A(n12306), .ZN(n12307) );
  NAND2_X1 U15302 ( .A1(n12307), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12308) );
  AND3_X1 U15303 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15541) );
  AND3_X1 U15304 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12309) );
  AND2_X1 U15305 ( .A1(n15541), .A2(n12309), .ZN(n15490) );
  NAND2_X1 U15306 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15491) );
  NOR2_X1 U15307 ( .A1(n15491), .A2(n12310), .ZN(n12311) );
  AND2_X1 U15308 ( .A1(n15490), .A2(n12311), .ZN(n15477) );
  NAND2_X1 U15309 ( .A1(n15477), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15456) );
  NAND2_X1 U15310 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12312) );
  NOR2_X1 U15311 ( .A1(n15456), .A2(n12312), .ZN(n15443) );
  AND2_X1 U15312 ( .A1(n15443), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12623) );
  AND2_X1 U15313 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U15314 ( .A1(n15402), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15381) );
  OAI21_X1 U15315 ( .B1(n15152), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15147), .ZN(n12649) );
  NAND2_X1 U15316 ( .A1(n12317), .A2(n12316), .ZN(P2_U2986) );
  NAND2_X1 U15317 ( .A1(n12322), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12321) );
  INV_X1 U15318 ( .A(n12321), .ZN(n12318) );
  NAND2_X1 U15319 ( .A1(n12318), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12320) );
  INV_X1 U15320 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12319) );
  INV_X1 U15321 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15335) );
  OAI21_X1 U15322 ( .B1(n12322), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n12321), .ZN(n12323) );
  INV_X1 U15323 ( .A(n12323), .ZN(n16420) );
  INV_X1 U15324 ( .A(n12325), .ZN(n12326) );
  AOI21_X1 U15325 ( .B1(n21232), .B2(n12324), .A(n12326), .ZN(n16435) );
  OR2_X1 U15326 ( .A1(n9945), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12327) );
  NAND2_X1 U15327 ( .A1(n12324), .A2(n12327), .ZN(n15165) );
  INV_X1 U15328 ( .A(n15165), .ZN(n16452) );
  AOI21_X1 U15329 ( .B1(n15175), .B2(n12328), .A(n9945), .ZN(n15177) );
  OAI21_X1 U15330 ( .B1(n12330), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12328), .ZN(n15187) );
  INV_X1 U15331 ( .A(n15187), .ZN(n16467) );
  AOI21_X1 U15332 ( .B1(n15196), .B2(n12329), .A(n12330), .ZN(n15199) );
  OAI21_X1 U15333 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12333), .A(
        n12329), .ZN(n16514) );
  INV_X1 U15334 ( .A(n16514), .ZN(n13013) );
  AOI21_X1 U15335 ( .B1(n15215), .B2(n12332), .A(n12333), .ZN(n15218) );
  OAI21_X1 U15336 ( .B1(n12334), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12332), .ZN(n15226) );
  INV_X1 U15337 ( .A(n15226), .ZN(n14928) );
  AND2_X1 U15338 ( .A1(n12335), .A2(n19203), .ZN(n12336) );
  OR2_X1 U15339 ( .A1(n12336), .A2(n12353), .ZN(n15255) );
  INV_X1 U15340 ( .A(n15255), .ZN(n19209) );
  AOI21_X1 U15341 ( .B1(n15278), .B2(n12350), .A(n9844), .ZN(n15277) );
  NOR2_X1 U15342 ( .A1(n12337), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12338) );
  AOI21_X1 U15343 ( .B1(n12348), .B2(n19263), .A(n12340), .ZN(n19266) );
  AOI21_X1 U15344 ( .B1(n16532), .B2(n9843), .A(n12341), .ZN(n19284) );
  AOI21_X1 U15345 ( .B1(n21274), .B2(n12346), .A(n12342), .ZN(n19295) );
  AOI21_X1 U15346 ( .B1(n16564), .B2(n12343), .A(n12347), .ZN(n19330) );
  AOI21_X1 U15347 ( .B1(n13793), .B2(n12344), .A(n12345), .ZN(n13791) );
  INV_X1 U15348 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13942) );
  OAI22_X1 U15349 ( .A1(n21322), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13942), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13941) );
  AND2_X1 U15350 ( .A1(n19352), .A2(n13941), .ZN(n13914) );
  OAI21_X1 U15351 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12344), .ZN(n13916) );
  NAND2_X1 U15352 ( .A1(n13914), .A2(n13916), .ZN(n13789) );
  OAI21_X1 U15353 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12345), .A(
        n12343), .ZN(n13756) );
  OAI21_X1 U15354 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12347), .A(
        n12346), .ZN(n19313) );
  NOR2_X1 U15355 ( .A1(n19295), .A2(n19294), .ZN(n13771) );
  OAI21_X1 U15356 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12342), .A(
        n9843), .ZN(n16545) );
  NAND2_X1 U15357 ( .A1(n13771), .A2(n16545), .ZN(n19283) );
  NOR2_X1 U15358 ( .A1(n19284), .A2(n19283), .ZN(n19275) );
  OAI21_X1 U15359 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12341), .A(
        n12348), .ZN(n19277) );
  NAND2_X1 U15360 ( .A1(n19275), .A2(n19277), .ZN(n19265) );
  NOR2_X1 U15361 ( .A1(n12340), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12349) );
  OR2_X1 U15362 ( .A1(n12337), .A2(n12349), .ZN(n19254) );
  OAI21_X1 U15363 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12351), .A(
        n12350), .ZN(n16520) );
  NOR2_X1 U15364 ( .A1(n15277), .A2(n19227), .ZN(n19216) );
  OAI21_X1 U15365 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9844), .A(
        n12335), .ZN(n19217) );
  NAND2_X1 U15366 ( .A1(n19216), .A2(n19217), .ZN(n19208) );
  OR2_X1 U15367 ( .A1(n12353), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12354) );
  NAND2_X1 U15368 ( .A1(n12355), .A2(n12354), .ZN(n15247) );
  AOI21_X1 U15369 ( .B1(n19191), .B2(n12355), .A(n12334), .ZN(n19196) );
  NOR2_X1 U15370 ( .A1(n19197), .A2(n19196), .ZN(n19195) );
  NOR2_X1 U15371 ( .A1(n14928), .A2(n14927), .ZN(n14926) );
  NOR2_X1 U15372 ( .A1(n19312), .A2(n14926), .ZN(n12982) );
  NOR2_X1 U15373 ( .A1(n15218), .A2(n12982), .ZN(n12981) );
  NOR2_X1 U15374 ( .A1(n19312), .A2(n12981), .ZN(n13010) );
  NOR2_X1 U15375 ( .A1(n13013), .A2(n13010), .ZN(n13012) );
  NOR2_X1 U15376 ( .A1(n19312), .A2(n13012), .ZN(n12994) );
  NOR2_X1 U15377 ( .A1(n15199), .A2(n12994), .ZN(n12996) );
  NOR2_X1 U15378 ( .A1(n19312), .A2(n12996), .ZN(n16464) );
  NOR2_X1 U15379 ( .A1(n16452), .A2(n16449), .ZN(n16451) );
  NOR2_X1 U15380 ( .A1(n19312), .A2(n16451), .ZN(n16436) );
  NOR2_X1 U15381 ( .A1(n16435), .A2(n16436), .ZN(n16434) );
  NOR2_X1 U15382 ( .A1(n19312), .A2(n16434), .ZN(n14896) );
  NOR2_X1 U15383 ( .A1(n19312), .A2(n16418), .ZN(n12357) );
  INV_X1 U15384 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12356) );
  XNOR2_X1 U15385 ( .A(n12321), .B(n12356), .ZN(n15139) );
  XNOR2_X1 U15386 ( .A(n12357), .B(n15139), .ZN(n12358) );
  NAND4_X1 U15387 ( .A1(n20132), .A2(n21322), .A3(n20153), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20024) );
  NAND2_X1 U15388 ( .A1(n12358), .A2(n19336), .ZN(n12570) );
  INV_X1 U15389 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n16422) );
  NOR2_X1 U15390 ( .A1(n13885), .A2(n16422), .ZN(n15114) );
  OR2_X2 U15391 ( .A1(n15115), .A2(n15114), .ZN(n14876) );
  NAND2_X1 U15392 ( .A1(n11860), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12359) );
  XNOR2_X1 U15393 ( .A(n14876), .B(n12359), .ZN(n15117) );
  OR2_X1 U15394 ( .A1(n16616), .A2(n13874), .ZN(n13028) );
  NAND2_X1 U15395 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20161) );
  INV_X1 U15396 ( .A(n20161), .ZN(n20150) );
  OR2_X1 U15397 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20150), .ZN(n12564) );
  NAND2_X1 U15398 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12564), .ZN(n12360) );
  NOR2_X1 U15399 ( .A1(n9789), .A2(n12360), .ZN(n12361) );
  NOR2_X1 U15400 ( .A1(n9773), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12384) );
  NOR2_X1 U15401 ( .A1(n13287), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15402 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12377) );
  AND2_X1 U15403 ( .A1(n13287), .A2(n20110), .ZN(n12390) );
  NAND2_X1 U15404 ( .A1(n12534), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12376) );
  AND3_X1 U15405 ( .A1(n9773), .A2(n13885), .A3(n20110), .ZN(n12381) );
  AOI22_X1 U15406 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15407 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12783), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15408 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15409 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11892), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U15410 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n12364), .ZN(
        n12374) );
  AOI22_X1 U15411 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15412 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12789), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15413 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12500), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15414 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11769), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15415 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NAND2_X1 U15416 ( .A1(n9754), .A2(n19360), .ZN(n12375) );
  INV_X1 U15417 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19342) );
  NAND2_X1 U15418 ( .A1(n10266), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12378) );
  OAI211_X1 U15419 ( .C1(n16624), .C2(n13273), .A(n12378), .B(n20110), .ZN(
        n12379) );
  INV_X1 U15420 ( .A(n12379), .ZN(n12380) );
  OAI21_X1 U15421 ( .B1(n14883), .B2(n19342), .A(n12380), .ZN(n13208) );
  AND2_X1 U15422 ( .A1(n21258), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12383) );
  NAND2_X1 U15423 ( .A1(n12384), .A2(n12943), .ZN(n12396) );
  NAND2_X1 U15424 ( .A1(n12381), .A2(n13203), .ZN(n12382) );
  OAI211_X1 U15425 ( .C1(n12390), .C2(n12383), .A(n12396), .B(n12382), .ZN(
        n13207) );
  INV_X1 U15426 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U15427 ( .A1(n12384), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12387) );
  NAND2_X1 U15428 ( .A1(n12385), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n12386) );
  OAI211_X1 U15429 ( .C1(n14883), .C2(n20046), .A(n12387), .B(n12386), .ZN(
        n12393) );
  OR2_X1 U15430 ( .A1(n12388), .A2(n12482), .ZN(n12392) );
  AOI22_X1 U15431 ( .A1(n12389), .A2(n12390), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12391) );
  NAND2_X1 U15432 ( .A1(n12392), .A2(n12391), .ZN(n13276) );
  NAND2_X1 U15433 ( .A1(n9754), .A2(n12394), .ZN(n12395) );
  OAI211_X1 U15434 ( .C1(n20110), .C2(n20121), .A(n12396), .B(n12395), .ZN(
        n12397) );
  AND2_X1 U15435 ( .A1(n12397), .A2(n10423), .ZN(n12398) );
  AND2_X1 U15436 ( .A1(n13279), .A2(n12398), .ZN(n12399) );
  INV_X1 U15437 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20048) );
  INV_X2 U15438 ( .A(n12419), .ZN(n14879) );
  NAND2_X1 U15439 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12401) );
  NAND2_X1 U15440 ( .A1(n14880), .A2(P2_EAX_REG_2__SCAN_IN), .ZN(n12400) );
  OAI211_X1 U15441 ( .C1(n14883), .C2(n20048), .A(n12401), .B(n12400), .ZN(
        n13296) );
  NAND2_X1 U15442 ( .A1(n12534), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15443 ( .A1(n14880), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12405) );
  NAND2_X1 U15444 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12404) );
  NAND2_X1 U15445 ( .A1(n9754), .A2(n12402), .ZN(n12403) );
  NAND4_X1 U15446 ( .A1(n12406), .A2(n12405), .A3(n12404), .A4(n12403), .ZN(
        n13607) );
  NAND2_X1 U15447 ( .A1(n13606), .A2(n13607), .ZN(n13671) );
  AOI22_X1 U15448 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U15449 ( .A1(n12534), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U15450 ( .A1(n9754), .A2(n12407), .ZN(n12408) );
  AOI22_X1 U15451 ( .A1(n12534), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n9754), .B2(
        n12411), .ZN(n12413) );
  AOI22_X1 U15452 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15453 ( .A1(n12413), .A2(n12412), .ZN(n13831) );
  NAND2_X1 U15454 ( .A1(n9754), .A2(n12414), .ZN(n12415) );
  AOI22_X1 U15455 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15456 ( .A1(n12534), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12416) );
  INV_X1 U15457 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19446) );
  INV_X1 U15458 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20057) );
  OAI222_X1 U15459 ( .A1(n16569), .A2(n12419), .B1(n12418), .B2(n19446), .C1(
        n14883), .C2(n20057), .ZN(n13197) );
  AOI22_X1 U15460 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12432) );
  NAND2_X1 U15461 ( .A1(n12534), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15462 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15463 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15464 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15465 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12420) );
  NAND4_X1 U15466 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12429) );
  AOI22_X1 U15467 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15468 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15469 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15470 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12424) );
  NAND4_X1 U15471 ( .A1(n12427), .A2(n12426), .A3(n12425), .A4(n12424), .ZN(
        n12428) );
  NAND2_X1 U15472 ( .A1(n9754), .A2(n19379), .ZN(n12430) );
  INV_X1 U15473 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U15474 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15475 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15476 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15477 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12433) );
  NAND4_X1 U15478 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12442) );
  AOI22_X1 U15479 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15480 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15481 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15482 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12437) );
  NAND4_X1 U15483 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12441) );
  AOI22_X1 U15484 ( .A1(n12534), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n9754), .B2(
        n12686), .ZN(n12444) );
  AOI22_X1 U15485 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U15486 ( .A1(n12444), .A2(n12443), .ZN(n13319) );
  AOI22_X1 U15487 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U15488 ( .A1(n12534), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15489 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15490 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15491 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15492 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11892), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U15493 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12454) );
  AOI22_X1 U15494 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15495 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12789), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15496 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15497 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15498 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12453) );
  NOR2_X1 U15499 ( .A1(n12454), .A2(n12453), .ZN(n19373) );
  INV_X1 U15500 ( .A(n19373), .ZN(n12455) );
  NAND2_X1 U15501 ( .A1(n9754), .A2(n12455), .ZN(n12456) );
  NOR2_X2 U15502 ( .A1(n15589), .A2(n15588), .ZN(n15590) );
  AOI22_X1 U15503 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15504 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15505 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15506 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12459) );
  NAND4_X1 U15507 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12468) );
  AOI22_X1 U15508 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15509 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15511 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U15512 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12467) );
  AOI22_X1 U15513 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U15514 ( .A1(n12534), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12469) );
  OAI211_X1 U15515 ( .C1(n12482), .C2(n13662), .A(n12470), .B(n12469), .ZN(
        n13424) );
  AOI22_X1 U15516 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12141), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15517 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12783), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15518 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15519 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11892), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12471) );
  NAND4_X1 U15520 ( .A1(n12474), .A2(n12473), .A3(n12472), .A4(n12471), .ZN(
        n12480) );
  AOI22_X1 U15521 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15522 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12789), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15523 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12500), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11769), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12475) );
  NAND4_X1 U15525 ( .A1(n12478), .A2(n12477), .A3(n12476), .A4(n12475), .ZN(
        n12479) );
  INV_X1 U15526 ( .A(n12689), .ZN(n19368) );
  AOI22_X1 U15527 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12481) );
  OAI21_X1 U15528 ( .B1(n19368), .B2(n12482), .A(n12481), .ZN(n12483) );
  AOI21_X1 U15529 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n12534), .A(n12483), 
        .ZN(n15568) );
  AOI22_X1 U15530 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15531 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15532 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15533 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15534 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12493) );
  AOI22_X1 U15535 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15536 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15537 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15538 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12488) );
  NAND4_X1 U15539 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12492) );
  AOI22_X1 U15540 ( .A1(n12534), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n9754), 
        .B2(n19361), .ZN(n12495) );
  AOI22_X1 U15541 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15542 ( .A1(n12495), .A2(n12494), .ZN(n13588) );
  AOI22_X1 U15543 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15544 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12783), .B1(
        n12141), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15545 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15546 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15547 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12496) );
  NAND4_X1 U15548 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n12506) );
  AOI22_X1 U15549 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15550 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15551 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15552 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11769), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12501) );
  NAND4_X1 U15553 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12505) );
  NAND2_X1 U15554 ( .A1(n9754), .A2(n9918), .ZN(n12507) );
  OAI211_X1 U15555 ( .C1(n14883), .C2(n15279), .A(n12508), .B(n12507), .ZN(
        n13627) );
  NAND2_X1 U15556 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12510) );
  NAND2_X1 U15557 ( .A1(n14880), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n12509) );
  OAI211_X1 U15558 ( .C1(n14883), .C2(n15513), .A(n12510), .B(n12509), .ZN(
        n15510) );
  NAND2_X1 U15559 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12512) );
  NAND2_X1 U15560 ( .A1(n14880), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n12511) );
  OAI211_X1 U15561 ( .C1(n14883), .C2(n20073), .A(n12512), .B(n12511), .ZN(
        n15097) );
  AOI22_X1 U15562 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U15563 ( .A1(n12534), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15564 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U15565 ( .A1(n12534), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12515) );
  NOR2_X2 U15566 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  INV_X1 U15567 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U15568 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12518) );
  NAND2_X1 U15569 ( .A1(n14880), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n12517) );
  OAI211_X1 U15570 ( .C1(n14883), .C2(n15225), .A(n12518), .B(n12517), .ZN(
        n14920) );
  AND2_X2 U15571 ( .A1(n15087), .A2(n14920), .ZN(n14922) );
  NAND2_X1 U15572 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15573 ( .A1(n14880), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n12519) );
  OAI211_X1 U15574 ( .C1(n14883), .C2(n12223), .A(n12520), .B(n12519), .ZN(
        n12988) );
  AND2_X2 U15575 ( .A1(n14922), .A2(n12988), .ZN(n13002) );
  INV_X1 U15576 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U15577 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12522) );
  NAND2_X1 U15578 ( .A1(n14880), .A2(P2_EAX_REG_22__SCAN_IN), .ZN(n12521) );
  OAI211_X1 U15579 ( .C1(n14883), .C2(n12523), .A(n12522), .B(n12521), .ZN(
        n13022) );
  NAND2_X1 U15580 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U15581 ( .A1(n14880), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n12524) );
  OAI211_X1 U15582 ( .C1(n14883), .C2(n12232), .A(n12525), .B(n12524), .ZN(
        n13001) );
  AOI22_X1 U15583 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15584 ( .A1(n12534), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12526) );
  AND2_X1 U15585 ( .A1(n12527), .A2(n12526), .ZN(n15052) );
  AOI22_X1 U15586 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U15587 ( .A1(n12534), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12528) );
  AND2_X1 U15588 ( .A1(n12529), .A2(n12528), .ZN(n14906) );
  INV_X1 U15589 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16453) );
  NAND2_X1 U15590 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15591 ( .A1(n14880), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n12530) );
  OAI211_X1 U15592 ( .C1(n14883), .C2(n16453), .A(n12531), .B(n12530), .ZN(
        n15038) );
  AOI22_X1 U15593 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12533) );
  NAND2_X1 U15594 ( .A1(n12534), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12532) );
  AND2_X1 U15595 ( .A1(n12533), .A2(n12532), .ZN(n15028) );
  AOI22_X1 U15596 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n14880), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15597 ( .A1(n12534), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12535) );
  AND2_X1 U15598 ( .A1(n12536), .A2(n12535), .ZN(n12633) );
  INV_X1 U15599 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20089) );
  NAND2_X1 U15600 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U15601 ( .A1(n14880), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n12537) );
  OAI211_X1 U15602 ( .C1(n14883), .C2(n20089), .A(n12538), .B(n12537), .ZN(
        n15011) );
  INV_X1 U15603 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U15604 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12540) );
  NAND2_X1 U15605 ( .A1(n14880), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n12539) );
  OAI211_X1 U15606 ( .C1(n14883), .C2(n15138), .A(n12540), .B(n12539), .ZN(
        n12541) );
  INV_X1 U15607 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19163) );
  NOR2_X1 U15608 ( .A1(n19163), .A2(n20045), .ZN(n20037) );
  NOR2_X1 U15609 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20038) );
  NOR3_X1 U15610 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20037), .A3(n20038), 
        .ZN(n20151) );
  NAND2_X1 U15611 ( .A1(n20161), .A2(n20151), .ZN(n13034) );
  NOR2_X1 U15612 ( .A1(n13034), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14887) );
  INV_X1 U15613 ( .A(n14887), .ZN(n12543) );
  NOR2_X1 U15614 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  NAND2_X1 U15615 ( .A1(n12587), .A2(n12545), .ZN(n16635) );
  NOR2_X1 U15616 ( .A1(n13028), .A2(n16635), .ZN(n19337) );
  INV_X2 U15617 ( .A(n19337), .ZN(n19335) );
  OR2_X1 U15618 ( .A1(n14888), .A2(n14887), .ZN(n12549) );
  INV_X1 U15619 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12547) );
  NAND3_X1 U15620 ( .A1(n13040), .A2(n12547), .A3(n12564), .ZN(n12548) );
  NAND2_X1 U15621 ( .A1(n19344), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12554) );
  NOR3_X1 U15622 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12550), .A3(n20110), 
        .ZN(n16633) );
  NOR2_X1 U15623 ( .A1(n19336), .A2(n16633), .ZN(n12551) );
  NAND2_X1 U15624 ( .A1(n19305), .A2(n12551), .ZN(n12552) );
  NAND2_X1 U15625 ( .A1(n19341), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19282) );
  AOI22_X1 U15626 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19349), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19327), .ZN(n12553) );
  OAI211_X1 U15627 ( .C1(n15343), .C2(n19335), .A(n12554), .B(n12553), .ZN(
        n12555) );
  AOI21_X1 U15628 ( .B1(n15117), .B2(n19339), .A(n12555), .ZN(n12568) );
  INV_X1 U15629 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15630 ( .A1(n14869), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12556) );
  OAI21_X1 U15631 ( .B1(n12175), .B2(n12557), .A(n12556), .ZN(n12558) );
  AOI21_X1 U15632 ( .B1(n11671), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12558), .ZN(n12563) );
  INV_X1 U15633 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15357) );
  OR2_X1 U15634 ( .A1(n14873), .A2(n15357), .ZN(n12562) );
  INV_X1 U15635 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16423) );
  OAI22_X1 U15636 ( .A1(n12559), .A2(n20089), .B1(n15656), .B2(n16423), .ZN(
        n12560) );
  AOI21_X1 U15637 ( .B1(n14870), .B2(P2_EBX_REG_29__SCAN_IN), .A(n12560), .ZN(
        n12561) );
  AND2_X1 U15638 ( .A1(n12562), .A2(n12561), .ZN(n14947) );
  AOI21_X1 U15639 ( .B1(n12563), .B2(n14950), .A(n14875), .ZN(n15342) );
  NOR2_X1 U15640 ( .A1(n9789), .A2(n12564), .ZN(n12565) );
  NAND2_X1 U15641 ( .A1(n19166), .A2(n12565), .ZN(n19346) );
  NAND2_X1 U15642 ( .A1(n15342), .A2(n12566), .ZN(n12567) );
  NAND2_X1 U15643 ( .A1(n12570), .A2(n12569), .ZN(P2_U2825) );
  NOR2_X1 U15644 ( .A1(n16614), .A2(n16624), .ZN(n13871) );
  INV_X1 U15645 ( .A(n13034), .ZN(n13870) );
  NAND3_X1 U15646 ( .A1(n13871), .A2(n13870), .A3(n12629), .ZN(n12595) );
  INV_X1 U15647 ( .A(n13871), .ZN(n12573) );
  AOI21_X1 U15648 ( .B1(n12571), .B2(n9812), .A(n19476), .ZN(n12572) );
  NAND2_X1 U15649 ( .A1(n12573), .A2(n12572), .ZN(n12594) );
  INV_X1 U15650 ( .A(n20143), .ZN(n12646) );
  NAND2_X1 U15651 ( .A1(n12587), .A2(n13870), .ZN(n12586) );
  NAND2_X1 U15652 ( .A1(n12389), .A2(n12580), .ZN(n12575) );
  NAND2_X1 U15653 ( .A1(n12575), .A2(n19467), .ZN(n12582) );
  AOI21_X1 U15654 ( .B1(n12580), .B2(n16624), .A(n12576), .ZN(n12577) );
  OAI21_X1 U15655 ( .B1(n12577), .B2(n10266), .A(n19467), .ZN(n12579) );
  OAI211_X1 U15656 ( .C1(n12583), .C2(n12580), .A(n12579), .B(n12578), .ZN(
        n12581) );
  AOI21_X1 U15657 ( .B1(n12574), .B2(n12582), .A(n12581), .ZN(n12585) );
  NAND2_X1 U15658 ( .A1(n12583), .A2(n13287), .ZN(n12584) );
  NAND2_X1 U15659 ( .A1(n12584), .A2(n20140), .ZN(n12608) );
  OAI211_X1 U15660 ( .C1(n16616), .C2(n12586), .A(n12585), .B(n12608), .ZN(
        n13865) );
  MUX2_X1 U15661 ( .A(n12587), .B(n12629), .S(n16624), .Z(n12588) );
  NAND2_X1 U15662 ( .A1(n12588), .A2(n20161), .ZN(n12589) );
  NOR2_X1 U15663 ( .A1(n16616), .A2(n12589), .ZN(n12590) );
  OR2_X1 U15664 ( .A1(n13865), .A2(n12590), .ZN(n12591) );
  AOI21_X1 U15665 ( .B1(n12592), .B2(n12646), .A(n12591), .ZN(n12593) );
  NAND3_X1 U15666 ( .A1(n12595), .A2(n12594), .A3(n12593), .ZN(n12596) );
  INV_X1 U15667 ( .A(n12648), .ZN(n12598) );
  NOR2_X1 U15668 ( .A1(n20143), .A2(n9789), .ZN(n12597) );
  NAND2_X1 U15669 ( .A1(n12599), .A2(n16592), .ZN(n12653) );
  AND3_X1 U15670 ( .A1(n19467), .A2(n16624), .A3(n13885), .ZN(n12601) );
  NAND2_X1 U15671 ( .A1(n12600), .A2(n12601), .ZN(n16620) );
  OAI22_X1 U15672 ( .A1(n12602), .A2(n19476), .B1(n19467), .B2(n9813), .ZN(
        n12603) );
  INV_X1 U15673 ( .A(n12603), .ZN(n12605) );
  NAND2_X1 U15674 ( .A1(n13285), .A2(n12604), .ZN(n12940) );
  AND3_X1 U15675 ( .A1(n12606), .A2(n12605), .A3(n12940), .ZN(n12615) );
  NAND2_X1 U15676 ( .A1(n12607), .A2(n20155), .ZN(n13859) );
  NAND2_X1 U15677 ( .A1(n13859), .A2(n12608), .ZN(n12610) );
  NAND2_X1 U15678 ( .A1(n12610), .A2(n12609), .ZN(n12614) );
  OAI21_X1 U15679 ( .B1(n13285), .B2(n10421), .A(n12602), .ZN(n12612) );
  NAND2_X1 U15680 ( .A1(n12612), .A2(n12611), .ZN(n12613) );
  AND2_X1 U15681 ( .A1(n15660), .A2(n11574), .ZN(n12616) );
  NOR2_X1 U15682 ( .A1(n12648), .A2(n12616), .ZN(n15500) );
  AND2_X1 U15683 ( .A1(n12648), .A2(n19305), .ZN(n13299) );
  NOR2_X1 U15684 ( .A1(n15498), .A2(n13299), .ZN(n15611) );
  AND2_X1 U15685 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U15686 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U15687 ( .A1(n12617), .A2(n13271), .ZN(n13292) );
  INV_X1 U15688 ( .A(n13292), .ZN(n12618) );
  NOR2_X1 U15689 ( .A1(n12617), .A2(n13271), .ZN(n12636) );
  INV_X1 U15690 ( .A(n12636), .ZN(n13293) );
  OAI211_X1 U15691 ( .C1(n15500), .C2(n12618), .A(n15498), .B(n13293), .ZN(
        n12619) );
  INV_X1 U15692 ( .A(n12619), .ZN(n12620) );
  NOR2_X1 U15693 ( .A1(n13299), .A2(n12620), .ZN(n16595) );
  OAI21_X1 U15694 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16583), .A(
        n16595), .ZN(n13839) );
  NAND3_X1 U15695 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12635) );
  AND2_X1 U15696 ( .A1(n15498), .A2(n12635), .ZN(n12621) );
  NOR2_X1 U15697 ( .A1(n13839), .A2(n12621), .ZN(n16580) );
  NAND2_X1 U15698 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16566) );
  NAND2_X1 U15699 ( .A1(n15498), .A2(n16566), .ZN(n12622) );
  NAND2_X1 U15700 ( .A1(n16580), .A2(n12622), .ZN(n15629) );
  INV_X1 U15701 ( .A(n12623), .ZN(n12624) );
  NOR2_X1 U15702 ( .A1(n15629), .A2(n12624), .ZN(n15413) );
  INV_X1 U15703 ( .A(n15413), .ZN(n12626) );
  INV_X1 U15704 ( .A(n15611), .ZN(n12625) );
  OAI21_X1 U15705 ( .B1(n12626), .B2(n15381), .A(n12625), .ZN(n15407) );
  OAI21_X1 U15706 ( .B1(n15611), .B2(n12639), .A(n15407), .ZN(n15375) );
  INV_X1 U15707 ( .A(n12627), .ZN(n12628) );
  NOR2_X1 U15708 ( .A1(n14961), .A2(n15600), .ZN(n12645) );
  NOR2_X1 U15709 ( .A1(n16615), .A2(n16624), .ZN(n12631) );
  NOR2_X1 U15710 ( .A1(n16624), .A2(n12629), .ZN(n12630) );
  AND2_X1 U15711 ( .A1(n12600), .A2(n12630), .ZN(n16618) );
  NOR2_X1 U15712 ( .A1(n12631), .A2(n16618), .ZN(n12632) );
  AND2_X1 U15713 ( .A1(n9872), .A2(n12633), .ZN(n12634) );
  OR2_X1 U15714 ( .A1(n12634), .A2(n15012), .ZN(n15020) );
  INV_X1 U15715 ( .A(n12635), .ZN(n12637) );
  OAI21_X1 U15716 ( .B1(n15494), .B2(n12636), .A(n13292), .ZN(n16582) );
  NAND2_X1 U15717 ( .A1(n12637), .A2(n15645), .ZN(n16567) );
  NOR2_X1 U15718 ( .A1(n16566), .A2(n16567), .ZN(n15539) );
  AND2_X1 U15719 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15539), .ZN(
        n12638) );
  NAND2_X1 U15720 ( .A1(n15443), .A2(n12638), .ZN(n15417) );
  OR2_X1 U15721 ( .A1(n15417), .A2(n15381), .ZN(n15379) );
  INV_X1 U15722 ( .A(n12639), .ZN(n12640) );
  NOR2_X1 U15723 ( .A1(n15379), .A2(n12640), .ZN(n15370) );
  NAND2_X1 U15724 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15358) );
  INV_X1 U15725 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12641) );
  NAND2_X1 U15726 ( .A1(n12641), .A2(n15369), .ZN(n15108) );
  NAND3_X1 U15727 ( .A1(n15370), .A2(n15358), .A3(n15108), .ZN(n12642) );
  OAI211_X1 U15728 ( .C1(n16581), .C2(n15020), .A(n12643), .B(n12642), .ZN(
        n12644) );
  AOI211_X1 U15729 ( .C1(n15375), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12645), .B(n12644), .ZN(n12651) );
  NAND2_X1 U15730 ( .A1(n12646), .A2(n20140), .ZN(n12647) );
  OR2_X1 U15731 ( .A1(n12649), .A2(n16588), .ZN(n12650) );
  NAND2_X1 U15732 ( .A1(n12653), .A2(n12652), .ZN(P2_U3018) );
  NAND2_X1 U15733 ( .A1(n13263), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U15734 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19948) );
  INV_X1 U15735 ( .A(n19948), .ZN(n12656) );
  AND2_X1 U15736 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12656), .ZN(
        n12657) );
  NAND2_X1 U15737 ( .A1(n12657), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19955) );
  INV_X1 U15738 ( .A(n12657), .ZN(n12674) );
  NAND2_X1 U15739 ( .A1(n20114), .A2(n12674), .ZN(n12658) );
  AND3_X1 U15740 ( .A1(n19955), .A2(n20102), .A3(n12658), .ZN(n19843) );
  AOI21_X1 U15741 ( .B1(n12676), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19843), .ZN(n12659) );
  NOR2_X1 U15742 ( .A1(n13263), .A2(n21322), .ZN(n12660) );
  INV_X1 U15743 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12661) );
  NOR2_X1 U15744 ( .A1(n12880), .A2(n12661), .ZN(n12662) );
  NAND2_X1 U15745 ( .A1(n12663), .A2(n12662), .ZN(n12684) );
  AOI22_X1 U15746 ( .A1(n12676), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20102), .B2(n21258), .ZN(n12666) );
  NAND2_X1 U15747 ( .A1(n12676), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12668) );
  NAND2_X1 U15748 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19809) );
  NAND2_X1 U15749 ( .A1(n11863), .A2(n21258), .ZN(n19719) );
  AND2_X1 U15750 ( .A1(n19809), .A2(n19719), .ZN(n19598) );
  NAND2_X1 U15751 ( .A1(n19598), .A2(n20102), .ZN(n19781) );
  NAND2_X1 U15752 ( .A1(n12668), .A2(n19781), .ZN(n12669) );
  NAND2_X1 U15753 ( .A1(n13283), .A2(n13284), .ZN(n12672) );
  INV_X1 U15754 ( .A(n13261), .ZN(n13864) );
  NAND2_X1 U15755 ( .A1(n13864), .A2(n12670), .ZN(n12671) );
  NAND2_X1 U15756 ( .A1(n12672), .A2(n12671), .ZN(n13309) );
  INV_X1 U15757 ( .A(n13309), .ZN(n12679) );
  NAND2_X1 U15758 ( .A1(n19809), .A2(n20121), .ZN(n12675) );
  AND2_X1 U15759 ( .A1(n12675), .A2(n12674), .ZN(n19599) );
  AOI22_X1 U15760 ( .A1(n12676), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20102), .B2(n19599), .ZN(n12677) );
  NAND2_X1 U15761 ( .A1(n12678), .A2(n12677), .ZN(n12681) );
  INV_X1 U15762 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19472) );
  NOR2_X1 U15763 ( .A1(n12880), .A2(n19472), .ZN(n12680) );
  NAND2_X1 U15764 ( .A1(n12679), .A2(n13311), .ZN(n12682) );
  NAND2_X1 U15765 ( .A1(n12681), .A2(n12680), .ZN(n13310) );
  NAND2_X1 U15766 ( .A1(n13350), .A2(n13351), .ZN(n13349) );
  NAND2_X1 U15767 ( .A1(n13263), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12683) );
  AND2_X1 U15768 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  INV_X1 U15769 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19481) );
  NOR2_X1 U15770 ( .A1(n12880), .A2(n19481), .ZN(n13675) );
  NAND2_X1 U15771 ( .A1(n12688), .A2(n12687), .ZN(n13661) );
  NOR2_X2 U15772 ( .A1(n13661), .A2(n13662), .ZN(n13663) );
  AOI22_X1 U15773 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U15774 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15775 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15776 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U15777 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12699) );
  AOI22_X1 U15778 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15779 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15780 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15781 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12694) );
  NAND4_X1 U15782 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12698) );
  AOI22_X1 U15783 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12141), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15784 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15785 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15786 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15787 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12709) );
  AOI22_X1 U15788 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15789 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15791 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12500), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12704) );
  NAND4_X1 U15792 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n12708) );
  AOI22_X1 U15793 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12141), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15794 ( .A1(n11817), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U15797 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12719) );
  AOI22_X1 U15798 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15799 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15800 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15801 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12500), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12714) );
  NAND4_X1 U15802 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12718) );
  NOR2_X1 U15803 ( .A1(n12719), .A2(n12718), .ZN(n16490) );
  AOI22_X1 U15804 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12141), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15805 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15806 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15807 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12721) );
  NAND4_X1 U15808 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12730) );
  AOI22_X1 U15809 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15810 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11751), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15812 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12500), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12725) );
  NAND4_X1 U15813 ( .A1(n12728), .A2(n12727), .A3(n12726), .A4(n12725), .ZN(
        n12729) );
  AOI22_X1 U15814 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12141), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15815 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15816 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15817 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12732) );
  NAND4_X1 U15818 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12742) );
  AOI22_X1 U15819 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12736), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15820 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15821 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15822 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12500), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12737) );
  NAND4_X1 U15823 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12737), .ZN(
        n12741) );
  NOR2_X1 U15824 ( .A1(n12742), .A2(n12741), .ZN(n16487) );
  INV_X1 U15825 ( .A(n16487), .ZN(n12743) );
  AOI22_X1 U15826 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15827 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U15828 ( .A1(n11887), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U15829 ( .A1(n12789), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12363), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12744) );
  NAND4_X1 U15830 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n12753) );
  AOI22_X1 U15831 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12788), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15832 ( .A1(n11751), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15833 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15834 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U15835 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12752) );
  AOI22_X1 U15836 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12141), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15837 ( .A1(n12731), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15838 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11848), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15839 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12363), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U15840 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12763) );
  AOI22_X1 U15841 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15842 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11892), .B1(
        n11751), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15843 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11767), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15844 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12500), .B1(
        n11769), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U15845 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12762) );
  NOR2_X1 U15846 ( .A1(n12763), .A2(n12762), .ZN(n15073) );
  AOI22_X1 U15847 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11744), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15848 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U15849 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12771) );
  AND2_X1 U15850 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12767) );
  OR2_X1 U15851 ( .A1(n12767), .A2(n12766), .ZN(n12929) );
  INV_X1 U15852 ( .A(n12929), .ZN(n12900) );
  NAND2_X1 U15853 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12769) );
  NAND2_X1 U15854 ( .A1(n9830), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12768) );
  AND3_X1 U15855 ( .A1(n12900), .A2(n12769), .A3(n12768), .ZN(n12770) );
  NAND4_X1 U15856 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12782) );
  AOI22_X1 U15857 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U15858 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12776) );
  NAND2_X1 U15859 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12775) );
  AND3_X1 U15860 ( .A1(n12776), .A2(n12929), .A3(n12775), .ZN(n12779) );
  AOI22_X1 U15861 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U15862 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9831), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U15863 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12781) );
  NAND2_X1 U15864 ( .A1(n12782), .A2(n12781), .ZN(n12819) );
  NOR2_X1 U15865 ( .A1(n16624), .A2(n12819), .ZN(n12796) );
  AOI22_X1 U15866 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11817), .B1(
        n11887), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15867 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12783), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15868 ( .A1(n12141), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11762), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15869 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12363), .B1(
        n11892), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12784) );
  NAND4_X1 U15870 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12795) );
  AOI22_X1 U15871 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12788), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U15872 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11751), .B1(
        n12789), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15873 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12500), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U15874 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11769), .B1(
        n11768), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12790) );
  NAND4_X1 U15875 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  NOR2_X1 U15876 ( .A1(n12795), .A2(n12794), .ZN(n12814) );
  XNOR2_X1 U15877 ( .A(n12796), .B(n12814), .ZN(n12821) );
  INV_X1 U15878 ( .A(n12819), .ZN(n12815) );
  AND2_X1 U15879 ( .A1(n16624), .A2(n12815), .ZN(n15062) );
  AOI22_X1 U15880 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U15881 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12801) );
  NAND2_X1 U15882 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12800) );
  AND3_X1 U15883 ( .A1(n12900), .A2(n12801), .A3(n12800), .ZN(n12804) );
  AOI22_X1 U15884 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15885 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12802) );
  NAND4_X1 U15886 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12813) );
  AOI22_X1 U15887 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U15888 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12807) );
  NAND2_X1 U15889 ( .A1(n9832), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12806) );
  AND3_X1 U15890 ( .A1(n12807), .A2(n12929), .A3(n12806), .ZN(n12810) );
  AOI22_X1 U15891 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15892 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12808) );
  NAND4_X1 U15893 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n12812) );
  NAND2_X1 U15894 ( .A1(n12813), .A2(n12812), .ZN(n12822) );
  INV_X1 U15895 ( .A(n12814), .ZN(n12816) );
  NAND2_X1 U15896 ( .A1(n12816), .A2(n12815), .ZN(n12823) );
  XOR2_X1 U15897 ( .A(n12822), .B(n12823), .Z(n12817) );
  INV_X1 U15898 ( .A(n12880), .ZN(n12859) );
  NAND2_X1 U15899 ( .A1(n12817), .A2(n12859), .ZN(n14985) );
  INV_X1 U15900 ( .A(n12822), .ZN(n12818) );
  NAND2_X1 U15901 ( .A1(n16624), .A2(n12818), .ZN(n14987) );
  NOR2_X1 U15902 ( .A1(n14987), .A2(n12819), .ZN(n12820) );
  NOR2_X1 U15903 ( .A1(n12823), .A2(n12822), .ZN(n12838) );
  AOI22_X1 U15904 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U15905 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U15906 ( .A1(n9836), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12824) );
  AND3_X1 U15907 ( .A1(n12900), .A2(n12825), .A3(n12824), .ZN(n12828) );
  AOI22_X1 U15908 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U15909 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12826) );
  NAND4_X1 U15910 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        n12837) );
  AOI22_X1 U15911 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U15912 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12831) );
  NAND2_X1 U15913 ( .A1(n9835), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12830) );
  AND3_X1 U15914 ( .A1(n12831), .A2(n12929), .A3(n12830), .ZN(n12834) );
  AOI22_X1 U15915 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15916 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U15917 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  AND2_X1 U15918 ( .A1(n12837), .A2(n12836), .ZN(n12840) );
  NAND2_X1 U15919 ( .A1(n12838), .A2(n12840), .ZN(n12879) );
  OAI211_X1 U15920 ( .C1(n12838), .C2(n12840), .A(n12859), .B(n12879), .ZN(
        n12842) );
  INV_X1 U15921 ( .A(n12842), .ZN(n12839) );
  INV_X1 U15922 ( .A(n12840), .ZN(n12841) );
  NOR2_X1 U15923 ( .A1(n20155), .A2(n12841), .ZN(n14980) );
  AOI22_X1 U15924 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U15925 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12846) );
  NAND2_X1 U15926 ( .A1(n9828), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12845) );
  AND3_X1 U15927 ( .A1(n12900), .A2(n12846), .A3(n12845), .ZN(n12849) );
  AOI22_X1 U15928 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U15929 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12847) );
  NAND4_X1 U15930 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12858) );
  AOI22_X1 U15931 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12856) );
  NAND2_X1 U15932 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12852) );
  NAND2_X1 U15933 ( .A1(n9829), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12851) );
  AND3_X1 U15934 ( .A1(n12852), .A2(n12929), .A3(n12851), .ZN(n12855) );
  AOI22_X1 U15935 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15936 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12853) );
  NAND4_X1 U15937 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  AND2_X1 U15938 ( .A1(n12858), .A2(n12857), .ZN(n12862) );
  XNOR2_X1 U15939 ( .A(n12879), .B(n12862), .ZN(n12860) );
  NAND2_X1 U15940 ( .A1(n12860), .A2(n12859), .ZN(n12863) );
  INV_X1 U15941 ( .A(n12862), .ZN(n12878) );
  NOR2_X1 U15942 ( .A1(n20155), .A2(n12878), .ZN(n14972) );
  AOI22_X1 U15944 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12869) );
  NAND2_X1 U15945 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12865) );
  NAND2_X1 U15946 ( .A1(n9829), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12864) );
  AND3_X1 U15947 ( .A1(n12900), .A2(n12865), .A3(n12864), .ZN(n12868) );
  AOI22_X1 U15948 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U15949 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12866) );
  NAND4_X1 U15950 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12877) );
  AOI22_X1 U15951 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U15952 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U15953 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12870) );
  AND3_X1 U15954 ( .A1(n12871), .A2(n12929), .A3(n12870), .ZN(n12874) );
  AOI22_X1 U15955 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U15956 ( .A1(n11744), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12872) );
  NAND4_X1 U15957 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12872), .ZN(
        n12876) );
  NAND2_X1 U15958 ( .A1(n12877), .A2(n12876), .ZN(n12883) );
  OR2_X1 U15959 ( .A1(n12879), .A2(n12878), .ZN(n12881) );
  NOR2_X1 U15960 ( .A1(n12881), .A2(n12883), .ZN(n14957) );
  NOR2_X1 U15961 ( .A1(n20155), .A2(n12883), .ZN(n14965) );
  AOI22_X1 U15962 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U15963 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12885) );
  NAND2_X1 U15964 ( .A1(n9826), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12884) );
  AND3_X1 U15965 ( .A1(n12900), .A2(n12885), .A3(n12884), .ZN(n12888) );
  AOI22_X1 U15966 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U15967 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12886) );
  NAND4_X1 U15968 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n12897) );
  AOI22_X1 U15969 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12895) );
  NAND2_X1 U15970 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12891) );
  NAND2_X1 U15971 ( .A1(n9825), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12890) );
  AND3_X1 U15972 ( .A1(n12891), .A2(n12929), .A3(n12890), .ZN(n12894) );
  AOI22_X1 U15973 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U15974 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12892) );
  NAND4_X1 U15975 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12896) );
  NAND2_X1 U15976 ( .A1(n12897), .A2(n12896), .ZN(n14959) );
  AOI21_X1 U15977 ( .B1(n14964), .B2(n14956), .A(n14959), .ZN(n14952) );
  AOI22_X1 U15978 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U15979 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12899) );
  NAND2_X1 U15980 ( .A1(n9831), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12898) );
  AND3_X1 U15981 ( .A1(n12900), .A2(n12899), .A3(n12898), .ZN(n12904) );
  AOI22_X1 U15982 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12903) );
  INV_X1 U15983 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U15984 ( .A1(n11752), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12902) );
  NAND4_X1 U15985 ( .A1(n12905), .A2(n12904), .A3(n12903), .A4(n12902), .ZN(
        n12913) );
  AOI22_X1 U15986 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12911) );
  NAND2_X1 U15987 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12907) );
  NAND2_X1 U15988 ( .A1(n9830), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12906) );
  AND3_X1 U15989 ( .A1(n12907), .A2(n12929), .A3(n12906), .ZN(n12910) );
  AOI22_X1 U15990 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U15991 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12908) );
  NAND4_X1 U15992 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12912) );
  NAND2_X1 U15993 ( .A1(n12913), .A2(n12912), .ZN(n12916) );
  NOR2_X1 U15994 ( .A1(n16624), .A2(n14959), .ZN(n12914) );
  NAND2_X1 U15995 ( .A1(n14957), .A2(n12914), .ZN(n12915) );
  NOR2_X1 U15996 ( .A1(n12915), .A2(n12916), .ZN(n12917) );
  AOI21_X1 U15997 ( .B1(n12916), .B2(n12915), .A(n12917), .ZN(n14951) );
  NAND2_X1 U15998 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  INV_X1 U15999 ( .A(n12917), .ZN(n12918) );
  NAND2_X1 U16000 ( .A1(n14953), .A2(n12918), .ZN(n12939) );
  AOI22_X1 U16001 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12919), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16002 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U16003 ( .A1(n12921), .A2(n12920), .ZN(n12936) );
  AOI21_X1 U16004 ( .B1(n12922), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12929), .ZN(n12924) );
  AOI22_X1 U16005 ( .A1(n11745), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U16006 ( .A1(n12919), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11579), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16007 ( .A1(n12926), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12927) );
  NAND2_X1 U16008 ( .A1(n12928), .A2(n12927), .ZN(n12934) );
  AOI22_X1 U16009 ( .A1(n9774), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11752), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16010 ( .A1(n12922), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12931) );
  NAND2_X1 U16011 ( .A1(n9832), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12930) );
  NAND4_X1 U16012 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12933) );
  OAI22_X1 U16013 ( .A1(n12936), .A2(n12935), .B1(n12934), .B2(n12933), .ZN(
        n12937) );
  INV_X1 U16014 ( .A(n12937), .ZN(n12938) );
  XNOR2_X1 U16015 ( .A(n12939), .B(n12938), .ZN(n14204) );
  OR2_X1 U16016 ( .A1(n16616), .A2(n16615), .ZN(n13037) );
  NAND2_X1 U16017 ( .A1(n12602), .A2(n20161), .ZN(n13035) );
  OAI22_X1 U16018 ( .A1(n16614), .A2(n16620), .B1(n13037), .B2(n13035), .ZN(
        n13869) );
  INV_X1 U16019 ( .A(n12940), .ZN(n12941) );
  NAND2_X1 U16020 ( .A1(n12943), .A2(n15094), .ZN(n19422) );
  NOR4_X1 U16021 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12947) );
  NOR4_X1 U16022 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12946) );
  NOR4_X1 U16023 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12945) );
  NOR4_X1 U16024 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12944) );
  NAND4_X1 U16025 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12952) );
  NOR4_X1 U16026 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12950) );
  NOR4_X1 U16027 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12949) );
  NOR4_X1 U16028 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12948) );
  INV_X1 U16029 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20050) );
  NAND4_X1 U16030 ( .A1(n12950), .A2(n12949), .A3(n12948), .A4(n20050), .ZN(
        n12951) );
  NOR3_X2 U16031 ( .A1(n19419), .A2(n13103), .A3(n12953), .ZN(n19397) );
  INV_X1 U16032 ( .A(n15343), .ZN(n12954) );
  NOR2_X2 U16033 ( .A1(n19419), .A2(n13287), .ZN(n19392) );
  AOI22_X1 U16034 ( .A1(n19397), .A2(BUF1_REG_30__SCAN_IN), .B1(n12954), .B2(
        n19392), .ZN(n12963) );
  NAND2_X1 U16035 ( .A1(n12955), .A2(n13103), .ZN(n12956) );
  NOR2_X2 U16036 ( .A1(n19419), .A2(n12956), .ZN(n19398) );
  NOR2_X1 U16037 ( .A1(n10266), .A2(n13885), .ZN(n12957) );
  NAND2_X1 U16038 ( .A1(n15094), .A2(n12957), .ZN(n15096) );
  INV_X1 U16039 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n12958) );
  NOR2_X1 U16040 ( .A1(n13881), .A2(n12958), .ZN(n12959) );
  AOI21_X1 U16041 ( .B1(BUF1_REG_14__SCAN_IN), .B2(n13881), .A(n12959), .ZN(
        n13112) );
  INV_X1 U16042 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12960) );
  OAI22_X1 U16043 ( .A1(n15096), .A2(n13112), .B1(n15094), .B2(n12960), .ZN(
        n12961) );
  AOI21_X1 U16044 ( .B1(n19398), .B2(BUF2_REG_30__SCAN_IN), .A(n12961), .ZN(
        n12962) );
  AND2_X1 U16045 ( .A1(n12963), .A2(n12962), .ZN(n12964) );
  OAI21_X1 U16046 ( .B1(n14204), .B2(n19422), .A(n12964), .ZN(P2_U2889) );
  NOR2_X1 U16047 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12966) );
  NOR4_X1 U16048 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12965) );
  NAND4_X1 U16049 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(P2_M_IO_N_REG_SCAN_IN), 
        .A3(n12966), .A4(n12965), .ZN(n12980) );
  NOR4_X1 U16050 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12970) );
  NOR4_X1 U16051 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12969) );
  NOR4_X1 U16052 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12968) );
  NOR4_X1 U16053 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12967) );
  AND4_X1 U16054 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n12976) );
  NOR4_X1 U16055 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_11__SCAN_IN), .A4(
        P1_ADDRESS_REG_5__SCAN_IN), .ZN(n12974) );
  NOR4_X1 U16056 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12973) );
  NOR4_X1 U16057 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12972) );
  INV_X1 U16058 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12971) );
  AND4_X1 U16059 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n12975) );
  NAND2_X1 U16060 ( .A1(n12976), .A2(n12975), .ZN(n12977) );
  INV_X1 U16061 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21115) );
  NOR3_X1 U16062 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21115), .ZN(n12979) );
  NOR4_X1 U16063 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12978) );
  NAND4_X1 U16064 ( .A1(n20377), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12979), .A4(
        n12978), .ZN(U214) );
  NOR2_X1 U16065 ( .A1(n13883), .A2(n12980), .ZN(n16727) );
  NAND2_X1 U16066 ( .A1(n16727), .A2(U214), .ZN(U212) );
  AOI211_X1 U16067 ( .C1(n15218), .C2(n12982), .A(n12981), .B(n20024), .ZN(
        n12993) );
  OAI22_X1 U16068 ( .A1(n15215), .A2(n19282), .B1(n12223), .B2(n19341), .ZN(
        n12992) );
  INV_X1 U16069 ( .A(n12983), .ZN(n12984) );
  OAI22_X1 U16070 ( .A1(n12984), .A2(n19306), .B1(n19324), .B2(n10243), .ZN(
        n12991) );
  INV_X1 U16071 ( .A(n12985), .ZN(n14919) );
  NAND2_X1 U16072 ( .A1(n14919), .A2(n12986), .ZN(n12987) );
  NAND2_X1 U16073 ( .A1(n13018), .A2(n12987), .ZN(n15441) );
  OR2_X1 U16074 ( .A1(n14922), .A2(n12988), .ZN(n12989) );
  NAND2_X1 U16075 ( .A1(n12989), .A2(n13021), .ZN(n15446) );
  OAI22_X1 U16076 ( .A1(n15441), .A2(n19346), .B1(n15446), .B2(n19335), .ZN(
        n12990) );
  OR4_X1 U16077 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        P2_U2834) );
  AOI211_X1 U16078 ( .C1(n15199), .C2(n12995), .A(n12996), .B(n20024), .ZN(
        n13009) );
  OAI22_X1 U16079 ( .A1(n15196), .A2(n19282), .B1(n12232), .B2(n19341), .ZN(
        n13008) );
  INV_X1 U16080 ( .A(n12997), .ZN(n12998) );
  OAI22_X1 U16081 ( .A1(n12998), .A2(n19306), .B1(n19324), .B2(n12113), .ZN(
        n13007) );
  NOR2_X1 U16082 ( .A1(n13019), .A2(n12999), .ZN(n13000) );
  OR2_X1 U16083 ( .A1(n14989), .A2(n13000), .ZN(n16481) );
  INV_X1 U16084 ( .A(n13001), .ZN(n13004) );
  NAND2_X1 U16085 ( .A1(n13022), .A2(n13002), .ZN(n13003) );
  NAND2_X1 U16086 ( .A1(n13004), .A2(n13003), .ZN(n13005) );
  AND2_X1 U16087 ( .A1(n13005), .A2(n15053), .ZN(n15420) );
  INV_X1 U16088 ( .A(n15420), .ZN(n15066) );
  OAI22_X1 U16089 ( .A1(n16481), .A2(n19346), .B1(n19335), .B2(n15066), .ZN(
        n13006) );
  OR4_X1 U16090 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        P2_U2832) );
  AOI211_X1 U16091 ( .C1(n13013), .C2(n13011), .A(n13012), .B(n20024), .ZN(
        n13027) );
  AOI22_X1 U16092 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19327), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19349), .ZN(n13014) );
  INV_X1 U16093 ( .A(n13014), .ZN(n13026) );
  INV_X1 U16094 ( .A(n13015), .ZN(n13016) );
  OAI22_X1 U16095 ( .A1(n13016), .A2(n19306), .B1(n19324), .B2(n12229), .ZN(
        n13025) );
  AND2_X1 U16096 ( .A1(n13018), .A2(n13017), .ZN(n13020) );
  OR2_X1 U16097 ( .A1(n13020), .A2(n13019), .ZN(n16510) );
  XNOR2_X1 U16098 ( .A(n13022), .B(n13021), .ZN(n15435) );
  INV_X1 U16099 ( .A(n15435), .ZN(n13023) );
  OAI22_X1 U16100 ( .A1(n16510), .A2(n19346), .B1(n19335), .B2(n13023), .ZN(
        n13024) );
  OR4_X1 U16101 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        P2_U2833) );
  INV_X1 U16102 ( .A(n13028), .ZN(n13029) );
  INV_X1 U16103 ( .A(n12574), .ZN(n16625) );
  NAND2_X1 U16104 ( .A1(n13029), .A2(n16625), .ZN(n13927) );
  INV_X1 U16105 ( .A(n13927), .ZN(n19348) );
  INV_X1 U16106 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13030) );
  INV_X1 U16107 ( .A(n13040), .ZN(n13039) );
  OAI211_X1 U16108 ( .C1(n19348), .C2(n13030), .A(n19165), .B(n13039), .ZN(
        P2_U2814) );
  INV_X1 U16109 ( .A(n12602), .ZN(n13033) );
  INV_X1 U16110 ( .A(n19166), .ZN(n20162) );
  INV_X1 U16111 ( .A(n19165), .ZN(n13031) );
  OAI21_X1 U16112 ( .B1(n13031), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20162), 
        .ZN(n13032) );
  OAI21_X1 U16113 ( .B1(n13033), .B2(n20162), .A(n13032), .ZN(P2_U3612) );
  NAND2_X1 U16114 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NOR2_X1 U16115 ( .A1(n13037), .A2(n13036), .ZN(n16622) );
  NOR2_X1 U16116 ( .A1(n16622), .A2(n13874), .ZN(n20149) );
  OAI21_X1 U16117 ( .B1(n20149), .B2(n12144), .A(n13038), .ZN(P2_U2819) );
  INV_X1 U16118 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13042) );
  OAI21_X1 U16119 ( .B1(n13039), .B2(n20150), .A(n14888), .ZN(n13101) );
  NAND3_X1 U16120 ( .A1(n13040), .A2(n20155), .A3(n20161), .ZN(n13127) );
  AOI22_X1 U16121 ( .A1(n13881), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13883), .ZN(n13630) );
  INV_X1 U16122 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13041) );
  OAI222_X1 U16123 ( .A1(n13042), .A2(n13101), .B1(n13127), .B2(n13630), .C1(
        n14888), .C2(n13041), .ZN(P2_U2982) );
  INV_X1 U16124 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13044) );
  OAI22_X1 U16125 ( .A1(n13103), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13881), .ZN(n19461) );
  INV_X1 U16126 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13043) );
  OAI222_X1 U16127 ( .A1(n13044), .A2(n13101), .B1(n13127), .B2(n19461), .C1(
        n14888), .C2(n13043), .ZN(P2_U2967) );
  INV_X1 U16128 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16129 ( .A1(n13881), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13103), .ZN(n19482) );
  NOR2_X1 U16130 ( .A1(n13127), .A2(n19482), .ZN(n13075) );
  AOI21_X1 U16131 ( .B1(n13098), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13075), .ZN(
        n13045) );
  OAI21_X1 U16132 ( .B1(n13101), .B2(n13046), .A(n13045), .ZN(P2_U2973) );
  INV_X1 U16133 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13048) );
  INV_X1 U16134 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16768) );
  INV_X1 U16135 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18494) );
  AOI22_X1 U16136 ( .A1(n13881), .A2(n16768), .B1(n18494), .B2(n13103), .ZN(
        n16493) );
  INV_X1 U16137 ( .A(n16493), .ZN(n19477) );
  NOR2_X1 U16138 ( .A1(n13127), .A2(n19477), .ZN(n13081) );
  AOI21_X1 U16139 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n13098), .A(n13081), .ZN(
        n13047) );
  OAI21_X1 U16140 ( .B1(n13101), .B2(n13048), .A(n13047), .ZN(P2_U2971) );
  INV_X1 U16141 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13050) );
  OAI22_X1 U16142 ( .A1(n13103), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13881), .ZN(n19468) );
  NOR2_X1 U16143 ( .A1(n13127), .A2(n19468), .ZN(n13069) );
  AOI21_X1 U16144 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n13098), .A(n13069), .ZN(
        n13049) );
  OAI21_X1 U16145 ( .B1(n13101), .B2(n13050), .A(n13049), .ZN(P2_U2969) );
  NOR4_X1 U16146 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13056) );
  NOR2_X1 U16147 ( .A1(n13057), .A2(n13056), .ZN(n13365) );
  NAND2_X1 U16148 ( .A1(n13051), .A2(n13365), .ZN(n13243) );
  INV_X1 U16149 ( .A(n13403), .ZN(n20171) );
  AND2_X1 U16150 ( .A1(n20826), .A2(n21324), .ZN(n13062) );
  NOR2_X1 U16151 ( .A1(n13137), .A2(n20171), .ZN(n13058) );
  INV_X1 U16152 ( .A(n13337), .ZN(n13059) );
  AOI211_X1 U16153 ( .C1(n13061), .C2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13062), 
        .B(n13059), .ZN(n13060) );
  INV_X1 U16154 ( .A(n13060), .ZN(P1_U2801) );
  OAI21_X1 U16155 ( .B1(n13062), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14359), 
        .ZN(n13063) );
  OAI21_X1 U16156 ( .B1(n13064), .B2(n14359), .A(n13063), .ZN(P1_U3487) );
  INV_X1 U16157 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16158 ( .A1(n13881), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13103), .ZN(n19418) );
  NOR2_X1 U16159 ( .A1(n13127), .A2(n19418), .ZN(n13078) );
  AOI21_X1 U16160 ( .B1(n13098), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13078), .ZN(
        n13065) );
  OAI21_X1 U16161 ( .B1(n13126), .B2(n13066), .A(n13065), .ZN(P2_U2972) );
  INV_X1 U16162 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16163 ( .A1(n13881), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13883), .ZN(n15095) );
  NOR2_X1 U16164 ( .A1(n13127), .A2(n15095), .ZN(n13072) );
  AOI21_X1 U16165 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n13098), .A(n13072), .ZN(
        n13067) );
  OAI21_X1 U16166 ( .B1(n13126), .B2(n13068), .A(n13067), .ZN(P2_U2968) );
  INV_X1 U16167 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13071) );
  AOI21_X1 U16168 ( .B1(n13098), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13069), .ZN(
        n13070) );
  OAI21_X1 U16169 ( .B1(n13126), .B2(n13071), .A(n13070), .ZN(P2_U2954) );
  INV_X1 U16170 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13074) );
  AOI21_X1 U16171 ( .B1(n13098), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13072), .ZN(
        n13073) );
  OAI21_X1 U16172 ( .B1(n13126), .B2(n13074), .A(n13073), .ZN(P2_U2953) );
  INV_X1 U16173 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13077) );
  AOI21_X1 U16174 ( .B1(n13098), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13075), .ZN(
        n13076) );
  OAI21_X1 U16175 ( .B1(n13126), .B2(n13077), .A(n13076), .ZN(P2_U2958) );
  INV_X1 U16176 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13080) );
  AOI21_X1 U16177 ( .B1(n13098), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13078), .ZN(
        n13079) );
  OAI21_X1 U16178 ( .B1(n13126), .B2(n13080), .A(n13079), .ZN(P2_U2957) );
  INV_X1 U16179 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13083) );
  AOI21_X1 U16180 ( .B1(n13098), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13081), .ZN(
        n13082) );
  OAI21_X1 U16181 ( .B1(n13126), .B2(n13083), .A(n13082), .ZN(P2_U2956) );
  INV_X1 U16182 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16183 ( .A1(n13881), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13883), .ZN(n19473) );
  NOR2_X1 U16184 ( .A1(n13127), .A2(n19473), .ZN(n13091) );
  AOI21_X1 U16185 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n13098), .A(n13091), .ZN(
        n13084) );
  OAI21_X1 U16186 ( .B1(n13126), .B2(n13085), .A(n13084), .ZN(P2_U2970) );
  INV_X1 U16187 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16188 ( .A1(n13881), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13103), .ZN(n19492) );
  NOR2_X1 U16189 ( .A1(n13127), .A2(n19492), .ZN(n13088) );
  AOI21_X1 U16190 ( .B1(n13098), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13088), .ZN(
        n13086) );
  OAI21_X1 U16191 ( .B1(n13126), .B2(n13087), .A(n13086), .ZN(P2_U2974) );
  INV_X1 U16192 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13090) );
  AOI21_X1 U16193 ( .B1(n13098), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13088), .ZN(
        n13089) );
  OAI21_X1 U16194 ( .B1(n13126), .B2(n13090), .A(n13089), .ZN(P2_U2959) );
  INV_X1 U16195 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13093) );
  AOI21_X1 U16196 ( .B1(n13098), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13091), .ZN(
        n13092) );
  OAI21_X1 U16197 ( .B1(n13126), .B2(n13093), .A(n13092), .ZN(P2_U2955) );
  INV_X1 U16198 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13095) );
  INV_X1 U16199 ( .A(n13127), .ZN(n13116) );
  MUX2_X1 U16200 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n13103), .Z(n15043) );
  NAND2_X1 U16201 ( .A1(n13116), .A2(n15043), .ZN(n13108) );
  NAND2_X1 U16202 ( .A1(n13098), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13094) );
  OAI211_X1 U16203 ( .C1(n13126), .C2(n13095), .A(n13108), .B(n13094), .ZN(
        P2_U2976) );
  INV_X1 U16204 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13097) );
  MUX2_X1 U16205 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n13103), .Z(n15010) );
  NAND2_X1 U16206 ( .A1(n13116), .A2(n15010), .ZN(n13123) );
  NAND2_X1 U16207 ( .A1(n13098), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13096) );
  OAI211_X1 U16208 ( .C1(n13126), .C2(n13097), .A(n13123), .B(n13096), .ZN(
        P2_U2980) );
  INV_X1 U16209 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13100) );
  MUX2_X1 U16210 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n13103), .Z(n15027) );
  NAND2_X1 U16211 ( .A1(n13116), .A2(n15027), .ZN(n13105) );
  NAND2_X1 U16212 ( .A1(n13098), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13099) );
  OAI211_X1 U16213 ( .C1(n13126), .C2(n13100), .A(n13105), .B(n13099), .ZN(
        P2_U2978) );
  INV_X1 U16214 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19436) );
  INV_X1 U16215 ( .A(n13101), .ZN(n13122) );
  NAND2_X1 U16216 ( .A1(n13122), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13104) );
  INV_X1 U16217 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16756) );
  NOR2_X1 U16218 ( .A1(n13103), .A2(n16756), .ZN(n13102) );
  AOI21_X1 U16219 ( .B1(n13103), .B2(BUF2_REG_12__SCAN_IN), .A(n13102), .ZN(
        n15022) );
  INV_X1 U16220 ( .A(n15022), .ZN(n19409) );
  NAND2_X1 U16221 ( .A1(n13116), .A2(n19409), .ZN(n13110) );
  OAI211_X1 U16222 ( .C1(n19436), .C2(n14888), .A(n13104), .B(n13110), .ZN(
        P2_U2979) );
  INV_X1 U16223 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16224 ( .A1(n13122), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13106) );
  OAI211_X1 U16225 ( .C1(n14888), .C2(n13155), .A(n13106), .B(n13105), .ZN(
        P2_U2963) );
  INV_X1 U16226 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U16227 ( .A1(n13122), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13107) );
  MUX2_X1 U16228 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n13103), .Z(n19415) );
  NAND2_X1 U16229 ( .A1(n13116), .A2(n19415), .ZN(n13120) );
  OAI211_X1 U16230 ( .C1(n13151), .C2(n14888), .A(n13107), .B(n13120), .ZN(
        P2_U2960) );
  INV_X1 U16231 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U16232 ( .A1(n13122), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13109) );
  OAI211_X1 U16233 ( .C1(n14888), .C2(n13157), .A(n13109), .B(n13108), .ZN(
        P2_U2961) );
  INV_X1 U16234 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U16235 ( .A1(n13122), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13111) );
  OAI211_X1 U16236 ( .C1(n13149), .C2(n14888), .A(n13111), .B(n13110), .ZN(
        P2_U2964) );
  NAND2_X1 U16237 ( .A1(n13122), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13113) );
  INV_X1 U16238 ( .A(n13112), .ZN(n19406) );
  NAND2_X1 U16239 ( .A1(n13116), .A2(n19406), .ZN(n13114) );
  OAI211_X1 U16240 ( .C1(n12960), .C2(n14888), .A(n13113), .B(n13114), .ZN(
        P2_U2966) );
  INV_X1 U16241 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19432) );
  NAND2_X1 U16242 ( .A1(n13122), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13115) );
  OAI211_X1 U16243 ( .C1(n19432), .C2(n14888), .A(n13115), .B(n13114), .ZN(
        P2_U2981) );
  INV_X1 U16244 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19440) );
  NAND2_X1 U16245 ( .A1(n13122), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13117) );
  MUX2_X1 U16246 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13103), .Z(n19412) );
  NAND2_X1 U16247 ( .A1(n13116), .A2(n19412), .ZN(n13118) );
  OAI211_X1 U16248 ( .C1(n19440), .C2(n14888), .A(n13117), .B(n13118), .ZN(
        P2_U2977) );
  INV_X1 U16249 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U16250 ( .A1(n13122), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13119) );
  OAI211_X1 U16251 ( .C1(n13160), .C2(n14888), .A(n13119), .B(n13118), .ZN(
        P2_U2962) );
  INV_X1 U16252 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19444) );
  NAND2_X1 U16253 ( .A1(n13122), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U16254 ( .C1(n19444), .C2(n14888), .A(n13121), .B(n13120), .ZN(
        P2_U2975) );
  INV_X1 U16255 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15015) );
  NAND2_X1 U16256 ( .A1(n13122), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13124) );
  OAI211_X1 U16257 ( .C1(n14888), .C2(n15015), .A(n13124), .B(n13123), .ZN(
        P2_U2965) );
  INV_X1 U16258 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13413) );
  INV_X1 U16259 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13125) );
  OAI222_X1 U16260 ( .A1(n13127), .A2(n19461), .B1(n14888), .B2(n13413), .C1(
        n13126), .C2(n13125), .ZN(P2_U2952) );
  NAND2_X1 U16261 ( .A1(n13128), .A2(n9765), .ZN(n13369) );
  NOR2_X1 U16262 ( .A1(n13129), .A2(n13369), .ZN(n13240) );
  INV_X1 U16263 ( .A(n13240), .ZN(n13387) );
  NOR2_X1 U16264 ( .A1(n13387), .A2(n16056), .ZN(n13136) );
  OR2_X1 U16265 ( .A1(n13249), .A2(n13130), .ZN(n13374) );
  INV_X1 U16266 ( .A(n13374), .ZN(n13131) );
  AOI21_X1 U16267 ( .B1(n13132), .B2(n13324), .A(n13131), .ZN(n13134) );
  INV_X1 U16268 ( .A(n13051), .ZN(n13133) );
  OAI22_X1 U16269 ( .A1(n13134), .A2(n13368), .B1(n13365), .B2(n13133), .ZN(
        n13135) );
  OAI21_X1 U16270 ( .B1(n13136), .B2(n13135), .A(n20424), .ZN(n16037) );
  INV_X1 U16271 ( .A(n13243), .ZN(n13139) );
  INV_X1 U16272 ( .A(n13137), .ZN(n13138) );
  INV_X1 U16273 ( .A(n13140), .ZN(n13141) );
  NAND2_X1 U16274 ( .A1(n13141), .A2(n21043), .ZN(n16069) );
  INV_X1 U16275 ( .A(n16069), .ZN(n16045) );
  AOI21_X1 U16276 ( .B1(n16044), .B2(n14358), .A(n16045), .ZN(n13142) );
  NAND2_X1 U16277 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21119) );
  INV_X1 U16278 ( .A(n21119), .ZN(n16068) );
  NOR2_X1 U16279 ( .A1(n13142), .A2(n16068), .ZN(n21122) );
  NOR2_X1 U16280 ( .A1(n20172), .A2(n21122), .ZN(n16035) );
  OR2_X1 U16281 ( .A1(n16035), .A2(n20171), .ZN(n20177) );
  INV_X1 U16282 ( .A(n20177), .ZN(n13144) );
  INV_X1 U16283 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13143) );
  OR2_X1 U16284 ( .A1(n13144), .A2(n13143), .ZN(n13145) );
  OAI21_X1 U16285 ( .B1(n16037), .B2(n20177), .A(n13145), .ZN(P1_U3484) );
  NAND3_X1 U16286 ( .A1(n13871), .A2(n16625), .A3(n20165), .ZN(n13146) );
  NAND2_X1 U16287 ( .A1(n13146), .A2(n14888), .ZN(n13147) );
  NAND2_X1 U16288 ( .A1(n19429), .A2(n20152), .ZN(n13423) );
  INV_X2 U16289 ( .A(n16630), .ZN(n13158) );
  NOR2_X4 U16290 ( .A1(n13158), .A2(n19429), .ZN(n19458) );
  AOI22_X1 U16291 ( .A1(n13158), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13148) );
  OAI21_X1 U16292 ( .B1(n13149), .B2(n13423), .A(n13148), .ZN(P2_U2923) );
  AOI22_X1 U16293 ( .A1(n13158), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13150) );
  OAI21_X1 U16294 ( .B1(n13151), .B2(n13423), .A(n13150), .ZN(P2_U2927) );
  AOI22_X1 U16295 ( .A1(n13158), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13152) );
  OAI21_X1 U16296 ( .B1(n15015), .B2(n13423), .A(n13152), .ZN(P2_U2922) );
  AOI22_X1 U16297 ( .A1(n13158), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13153) );
  OAI21_X1 U16298 ( .B1(n12960), .B2(n13423), .A(n13153), .ZN(P2_U2921) );
  AOI22_X1 U16299 ( .A1(n13158), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U16300 ( .B1(n13155), .B2(n13423), .A(n13154), .ZN(P2_U2924) );
  AOI22_X1 U16301 ( .A1(n13158), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U16302 ( .B1(n13157), .B2(n13423), .A(n13156), .ZN(P2_U2926) );
  AOI22_X1 U16303 ( .A1(n13158), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13159) );
  OAI21_X1 U16304 ( .B1(n13160), .B2(n13423), .A(n13159), .ZN(P2_U2925) );
  INV_X1 U16305 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13165) );
  NAND2_X1 U16306 ( .A1(n13051), .A2(n20398), .ZN(n16020) );
  NAND2_X1 U16307 ( .A1(n13246), .A2(n9971), .ZN(n13380) );
  NAND2_X1 U16308 ( .A1(n16020), .A2(n13380), .ZN(n13163) );
  NAND2_X1 U16309 ( .A1(n16045), .A2(n13403), .ZN(n13161) );
  NOR2_X1 U16310 ( .A1(n16056), .A2(n13161), .ZN(n13162) );
  NAND2_X1 U16311 ( .A1(n20306), .A2(n9755), .ZN(n13441) );
  NAND2_X1 U16312 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16416) );
  INV_X1 U16313 ( .A(n16416), .ZN(n16411) );
  NAND2_X1 U16314 ( .A1(n21027), .A2(n16411), .ZN(n20304) );
  NOR2_X4 U16315 ( .A1(n20306), .A2(n20332), .ZN(n20331) );
  AOI22_X1 U16316 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13164) );
  OAI21_X1 U16317 ( .B1(n13165), .B2(n13441), .A(n13164), .ZN(P1_U2906) );
  INV_X1 U16318 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U16319 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13166) );
  OAI21_X1 U16320 ( .B1(n13167), .B2(n13441), .A(n13166), .ZN(P1_U2907) );
  INV_X1 U16321 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U16322 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13168) );
  OAI21_X1 U16323 ( .B1(n13169), .B2(n13441), .A(n13168), .ZN(P1_U2908) );
  INV_X1 U16324 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13171) );
  AOI22_X1 U16325 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13170) );
  OAI21_X1 U16326 ( .B1(n13171), .B2(n13441), .A(n13170), .ZN(P1_U2912) );
  INV_X1 U16327 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U16328 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13172) );
  OAI21_X1 U16329 ( .B1(n13173), .B2(n13441), .A(n13172), .ZN(P1_U2909) );
  INV_X1 U16330 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16331 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13174) );
  OAI21_X1 U16332 ( .B1(n13175), .B2(n13441), .A(n13174), .ZN(P1_U2910) );
  INV_X1 U16333 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16334 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13176) );
  OAI21_X1 U16335 ( .B1(n13177), .B2(n13441), .A(n13176), .ZN(P1_U2911) );
  INV_X1 U16336 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13183) );
  INV_X1 U16337 ( .A(n13916), .ZN(n13917) );
  NAND2_X1 U16338 ( .A1(n16555), .A2(n13917), .ZN(n13182) );
  INV_X1 U16339 ( .A(n13178), .ZN(n13179) );
  XNOR2_X1 U16340 ( .A(n13180), .B(n13179), .ZN(n13300) );
  AOI22_X1 U16341 ( .A1(n16550), .A2(n13300), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n19326), .ZN(n13181) );
  OAI211_X1 U16342 ( .C1(n13183), .C2(n16565), .A(n13182), .B(n13181), .ZN(
        n13184) );
  INV_X1 U16343 ( .A(n13184), .ZN(n13188) );
  NAND2_X1 U16344 ( .A1(n13186), .A2(n13185), .ZN(n13301) );
  NAND3_X1 U16345 ( .A1(n13302), .A2(n16549), .A3(n13301), .ZN(n13187) );
  OAI211_X1 U16346 ( .C1(n13882), .C2(n10117), .A(n13188), .B(n13187), .ZN(
        P2_U3012) );
  OAI21_X1 U16347 ( .B1(n13946), .B2(n13201), .A(n13189), .ZN(n13190) );
  INV_X1 U16348 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15659) );
  XOR2_X1 U16349 ( .A(n13190), .B(n15659), .Z(n13280) );
  OAI21_X1 U16350 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13192), .A(
        n13191), .ZN(n13270) );
  NAND2_X1 U16351 ( .A1(n19326), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13269) );
  OAI21_X1 U16352 ( .B1(n16558), .B2(n13270), .A(n13269), .ZN(n13194) );
  MUX2_X1 U16353 ( .A(n16555), .B(n16546), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13193) );
  AOI211_X1 U16354 ( .C1(n13280), .C2(n16549), .A(n13194), .B(n13193), .ZN(
        n13195) );
  OAI21_X1 U16355 ( .B1(n11723), .B2(n13882), .A(n13195), .ZN(P2_U3013) );
  AND2_X1 U16356 ( .A1(n12389), .A2(n13287), .ZN(n13196) );
  OAI21_X1 U16357 ( .B1(n13198), .B2(n13197), .A(n13778), .ZN(n19300) );
  OAI222_X1 U16358 ( .A1(n13679), .A2(n19492), .B1(n19300), .B2(n19428), .C1(
        n19446), .C2(n15094), .ZN(P2_U2912) );
  XNOR2_X1 U16359 ( .A(n13200), .B(n13199), .ZN(n19319) );
  INV_X1 U16360 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19448) );
  OAI222_X1 U16361 ( .A1(n13679), .A2(n19482), .B1(n19319), .B2(n19428), .C1(
        n19448), .C2(n15094), .ZN(P2_U2913) );
  INV_X1 U16362 ( .A(n15600), .ZN(n16586) );
  NOR2_X1 U16363 ( .A1(n19342), .A2(n19305), .ZN(n14077) );
  OAI21_X1 U16364 ( .B1(n19338), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13201), .ZN(n14075) );
  AOI21_X1 U16365 ( .B1(n13203), .B2(n13273), .A(n13202), .ZN(n14078) );
  INV_X1 U16366 ( .A(n14078), .ZN(n13204) );
  OAI22_X1 U16367 ( .A1(n15632), .A2(n14075), .B1(n16588), .B2(n13204), .ZN(
        n13205) );
  AOI211_X1 U16368 ( .C1(n16586), .C2(n13206), .A(n14077), .B(n13205), .ZN(
        n13212) );
  NOR2_X1 U16369 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  AOI22_X1 U16370 ( .A1(n15602), .A2(n10422), .B1(n13299), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13211) );
  OAI211_X1 U16371 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16583), .A(
        n13212), .B(n13211), .ZN(P2_U3046) );
  AND2_X1 U16372 ( .A1(n13369), .A2(n9755), .ZN(n13213) );
  AND2_X1 U16373 ( .A1(n13214), .A2(n13213), .ZN(n13250) );
  INV_X1 U16374 ( .A(n13250), .ZN(n13222) );
  NAND2_X1 U16375 ( .A1(n9910), .A2(n13233), .ZN(n13218) );
  OAI211_X1 U16376 ( .C1(n13216), .C2(n14358), .A(n13215), .B(n14120), .ZN(
        n13217) );
  AOI21_X1 U16377 ( .B1(n13218), .B2(n20398), .A(n13217), .ZN(n13221) );
  NAND3_X1 U16378 ( .A1(n13222), .A2(n13221), .A3(n13220), .ZN(n13385) );
  INV_X1 U16379 ( .A(n13385), .ZN(n13228) );
  INV_X1 U16380 ( .A(n13383), .ZN(n13223) );
  OR2_X1 U16381 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  NOR2_X1 U16382 ( .A1(n13246), .A2(n13225), .ZN(n13227) );
  NAND3_X1 U16383 ( .A1(n13228), .A2(n13227), .A3(n13226), .ZN(n14861) );
  INV_X1 U16384 ( .A(n14861), .ZN(n13314) );
  OR2_X1 U16385 ( .A1(n13249), .A2(n13229), .ZN(n13241) );
  INV_X1 U16386 ( .A(n13241), .ZN(n13230) );
  OR2_X1 U16387 ( .A1(n13240), .A2(n13230), .ZN(n13570) );
  INV_X1 U16388 ( .A(n13563), .ZN(n13231) );
  INV_X1 U16389 ( .A(n10438), .ZN(n14857) );
  NAND2_X1 U16390 ( .A1(n14857), .A2(n10430), .ZN(n13562) );
  NAND2_X1 U16391 ( .A1(n13231), .A2(n13562), .ZN(n13237) );
  XNOR2_X1 U16392 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13232) );
  NOR2_X1 U16393 ( .A1(n16020), .A2(n13232), .ZN(n13235) );
  NOR3_X1 U16394 ( .A1(n14861), .A2(n13233), .A3(n13237), .ZN(n13234) );
  AOI211_X1 U16395 ( .C1(n13570), .C2(n13237), .A(n13235), .B(n13234), .ZN(
        n13236) );
  OAI21_X1 U16396 ( .B1(n20831), .B2(n13314), .A(n13236), .ZN(n13561) );
  INV_X1 U16397 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13536) );
  OAI22_X1 U16398 ( .A1(n10919), .A2(n13536), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14865) );
  INV_X1 U16399 ( .A(n14865), .ZN(n13239) );
  INV_X1 U16400 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14784) );
  NOR2_X1 U16401 ( .A1(n21324), .A2(n14784), .ZN(n14864) );
  INV_X1 U16402 ( .A(n13237), .ZN(n13238) );
  AOI222_X1 U16403 ( .A1(n13561), .A2(n21102), .B1(n13239), .B2(n14864), .C1(
        n21101), .C2(n13238), .ZN(n13260) );
  NAND2_X1 U16404 ( .A1(n13240), .A2(n16056), .ZN(n13328) );
  NAND2_X1 U16405 ( .A1(n13246), .A2(n21119), .ZN(n16043) );
  OAI21_X1 U16406 ( .B1(n16043), .B2(n14082), .A(n13241), .ZN(n13242) );
  NAND2_X1 U16407 ( .A1(n13242), .A2(n13368), .ZN(n13245) );
  OR3_X1 U16408 ( .A1(n13243), .A2(n16068), .A3(n20398), .ZN(n13244) );
  INV_X1 U16409 ( .A(n13246), .ZN(n13248) );
  NAND3_X1 U16410 ( .A1(n13368), .A2(n16045), .A3(n21119), .ZN(n13247) );
  AOI21_X1 U16411 ( .B1(n16020), .B2(n13248), .A(n13247), .ZN(n13253) );
  NOR2_X1 U16412 ( .A1(n13250), .A2(n13249), .ZN(n13251) );
  OR2_X1 U16413 ( .A1(n13251), .A2(n13051), .ZN(n13367) );
  OAI21_X1 U16414 ( .B1(n14358), .B2(n10063), .A(n13367), .ZN(n13252) );
  NOR2_X1 U16415 ( .A1(n13253), .A2(n13252), .ZN(n13254) );
  AND2_X1 U16416 ( .A1(n13402), .A2(n13254), .ZN(n13255) );
  NOR2_X1 U16417 ( .A1(n21027), .A2(n16416), .ZN(n13582) );
  NAND2_X1 U16418 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13582), .ZN(n13257) );
  NAND2_X1 U16419 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21027), .ZN(n13256) );
  AND2_X1 U16420 ( .A1(n13257), .A2(n13256), .ZN(n13258) );
  OAI21_X1 U16421 ( .B1(n16026), .B2(n20171), .A(n13258), .ZN(n16407) );
  INV_X1 U16422 ( .A(n16407), .ZN(n21105) );
  NAND2_X1 U16423 ( .A1(n21105), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13259) );
  OAI21_X1 U16424 ( .B1(n13260), .B2(n21105), .A(n13259), .ZN(P1_U3472) );
  INV_X1 U16425 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19464) );
  NAND2_X1 U16426 ( .A1(n20110), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13262) );
  NOR2_X1 U16427 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  OAI21_X1 U16428 ( .B1(n16624), .B2(n19464), .A(n13264), .ZN(n13265) );
  INV_X1 U16429 ( .A(n13265), .ZN(n13266) );
  NAND2_X1 U16430 ( .A1(n19501), .A2(n10422), .ZN(n13493) );
  OAI211_X1 U16431 ( .C1(n19501), .C2(n10422), .A(n16501), .B(n13493), .ZN(
        n13268) );
  AOI22_X1 U16432 ( .A1(n19392), .A2(n10422), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19419), .ZN(n13267) );
  OAI211_X1 U16433 ( .C1(n13679), .C2(n19461), .A(n13268), .B(n13267), .ZN(
        P2_U2919) );
  OAI21_X1 U16434 ( .B1(n16588), .B2(n13270), .A(n13269), .ZN(n13275) );
  INV_X1 U16435 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13273) );
  INV_X1 U16436 ( .A(n13271), .ZN(n13272) );
  AOI211_X1 U16437 ( .C1(n13273), .C2(n15659), .A(n13272), .B(n16583), .ZN(
        n13274) );
  AOI211_X1 U16438 ( .C1(n13299), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13275), .B(n13274), .ZN(n13282) );
  NAND2_X1 U16439 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  NAND2_X1 U16440 ( .A1(n13279), .A2(n13278), .ZN(n20129) );
  AOI22_X1 U16441 ( .A1(n15602), .A2(n20129), .B1(n16592), .B2(n13280), .ZN(
        n13281) );
  OAI211_X1 U16442 ( .C1(n11723), .C2(n15600), .A(n13282), .B(n13281), .ZN(
        P2_U3045) );
  NAND2_X1 U16443 ( .A1(n16614), .A2(n16618), .ZN(n13867) );
  NAND2_X1 U16444 ( .A1(n15660), .A2(n13285), .ZN(n15670) );
  NAND2_X1 U16445 ( .A1(n13867), .A2(n15670), .ZN(n13286) );
  NAND2_X1 U16446 ( .A1(n19356), .A2(n13287), .ZN(n19380) );
  INV_X1 U16447 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13288) );
  MUX2_X1 U16448 ( .A(n13288), .B(n11723), .S(n19356), .Z(n13289) );
  OAI21_X1 U16449 ( .B1(n20124), .B2(n19380), .A(n13289), .ZN(P2_U2886) );
  NOR2_X1 U16450 ( .A1(n19385), .A2(n9816), .ZN(n13290) );
  AOI21_X1 U16451 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19385), .A(n13290), .ZN(
        n13291) );
  OAI21_X1 U16452 ( .B1(n19380), .B2(n20133), .A(n13291), .ZN(P2_U2887) );
  NAND2_X1 U16453 ( .A1(n13293), .A2(n13292), .ZN(n13307) );
  INV_X1 U16454 ( .A(n13307), .ZN(n13294) );
  NAND2_X1 U16455 ( .A1(n15500), .A2(n13294), .ZN(n13295) );
  OAI21_X1 U16456 ( .B1(n20048), .B2(n15303), .A(n13295), .ZN(n13306) );
  NAND2_X1 U16457 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  AND2_X1 U16458 ( .A1(n13298), .A2(n9946), .ZN(n13922) );
  AOI22_X1 U16459 ( .A1(n16574), .A2(n13300), .B1(n13299), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13304) );
  NAND3_X1 U16460 ( .A1(n16592), .A2(n13302), .A3(n13301), .ZN(n13303) );
  OAI211_X1 U16461 ( .C1(n13922), .C2(n16581), .A(n13304), .B(n13303), .ZN(
        n13305) );
  AOI211_X1 U16462 ( .C1(n15494), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13308) );
  OAI21_X1 U16463 ( .B1(n10117), .B2(n15600), .A(n13308), .ZN(P2_U3044) );
  NAND2_X1 U16464 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  MUX2_X1 U16465 ( .A(n11868), .B(n10117), .S(n19356), .Z(n13313) );
  OAI21_X1 U16466 ( .B1(n20117), .B2(n19380), .A(n13313), .ZN(P2_U2885) );
  INV_X1 U16467 ( .A(n20496), .ZN(n14374) );
  OAI22_X1 U16468 ( .A1(n14374), .A2(n13314), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10622), .ZN(n16018) );
  OAI22_X1 U16469 ( .A1(n21324), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14862), .ZN(n13315) );
  AOI21_X1 U16470 ( .B1(n16018), .B2(n21102), .A(n13315), .ZN(n13318) );
  INV_X1 U16471 ( .A(n16020), .ZN(n13316) );
  AOI21_X1 U16472 ( .B1(n13316), .B2(n21102), .A(n21105), .ZN(n13317) );
  OAI22_X1 U16473 ( .A1(n13318), .A2(n21105), .B1(n13317), .B2(n10928), .ZN(
        P1_U3474) );
  INV_X1 U16474 ( .A(n15043), .ZN(n13320) );
  INV_X1 U16475 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19442) );
  OAI21_X1 U16476 ( .B1(n13777), .B2(n13319), .A(n15589), .ZN(n19289) );
  OAI222_X1 U16477 ( .A1(n13679), .A2(n13320), .B1(n15094), .B2(n19442), .C1(
        n19428), .C2(n19289), .ZN(P2_U2910) );
  NAND2_X1 U16478 ( .A1(n14135), .A2(n14784), .ZN(n13323) );
  OR2_X1 U16479 ( .A1(n14149), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U16480 ( .A1(n14120), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U16481 ( .A1(n13322), .A2(n13321), .ZN(n13504) );
  AND2_X1 U16482 ( .A1(n13323), .A2(n13504), .ZN(n14371) );
  INV_X1 U16483 ( .A(n14371), .ZN(n13335) );
  AND2_X1 U16484 ( .A1(n13324), .A2(n10625), .ZN(n13326) );
  NOR2_X1 U16485 ( .A1(n9765), .A2(n20424), .ZN(n13325) );
  AND3_X1 U16486 ( .A1(n13564), .A2(n13326), .A3(n13325), .ZN(n13400) );
  NAND2_X1 U16487 ( .A1(n13400), .A2(n14143), .ZN(n13327) );
  NAND2_X1 U16488 ( .A1(n13328), .A2(n13327), .ZN(n13329) );
  INV_X1 U16489 ( .A(n20424), .ZN(n14194) );
  INV_X1 U16490 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13334) );
  INV_X1 U16491 ( .A(n13330), .ZN(n13333) );
  OAI21_X1 U16492 ( .B1(n13333), .B2(n13332), .A(n13331), .ZN(n20374) );
  NAND2_X2 U16493 ( .A1(n20302), .A2(n20424), .ZN(n14452) );
  OAI222_X1 U16494 ( .A1(n13335), .A2(n20288), .B1(n13334), .B2(n20302), .C1(
        n20374), .C2(n14452), .ZN(P1_U2872) );
  AND2_X1 U16495 ( .A1(n16044), .A2(n16068), .ZN(n13336) );
  OR2_X2 U16496 ( .A1(n13337), .A2(n13336), .ZN(n20360) );
  OR2_X1 U16497 ( .A1(n20360), .A2(n20398), .ZN(n13452) );
  INV_X1 U16498 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14544) );
  NOR2_X2 U16499 ( .A1(n20360), .A2(n13338), .ZN(n20348) );
  INV_X1 U16500 ( .A(n20348), .ZN(n13341) );
  INV_X1 U16501 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13339) );
  NOR2_X1 U16502 ( .A1(n20379), .A2(n13339), .ZN(n13340) );
  AOI21_X1 U16503 ( .B1(DATAI_15_), .B2(n20379), .A(n13340), .ZN(n14545) );
  INV_X1 U16504 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20305) );
  OAI222_X1 U16505 ( .A1(n13452), .A2(n14544), .B1(n13341), .B2(n14545), .C1(
        n13453), .C2(n20305), .ZN(P1_U2967) );
  XOR2_X1 U16506 ( .A(n13342), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13348)
         );
  NAND2_X1 U16507 ( .A1(n13343), .A2(n13702), .ZN(n13345) );
  INV_X1 U16508 ( .A(n13395), .ZN(n13344) );
  AND2_X1 U16509 ( .A1(n13345), .A2(n13344), .ZN(n19331) );
  NOR2_X1 U16510 ( .A1(n19356), .A2(n19323), .ZN(n13346) );
  AOI21_X1 U16511 ( .B1(n19331), .B2(n19356), .A(n13346), .ZN(n13347) );
  OAI21_X1 U16512 ( .B1(n13348), .B2(n19380), .A(n13347), .ZN(P2_U2882) );
  NAND2_X1 U16513 ( .A1(n9837), .A2(n19356), .ZN(n13354) );
  NAND2_X1 U16514 ( .A1(n19385), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13353) );
  OAI211_X1 U16515 ( .C1(n19504), .C2(n19380), .A(n13354), .B(n13353), .ZN(
        P2_U2884) );
  INV_X1 U16516 ( .A(n13355), .ZN(n13358) );
  INV_X1 U16517 ( .A(n13356), .ZN(n13357) );
  AOI21_X1 U16518 ( .B1(n13358), .B2(n14784), .A(n13357), .ZN(n20370) );
  INV_X1 U16519 ( .A(n20370), .ZN(n13393) );
  NAND2_X1 U16520 ( .A1(n16043), .A2(n9755), .ZN(n13360) );
  NAND2_X1 U16521 ( .A1(n9971), .A2(n16069), .ZN(n13359) );
  AOI21_X1 U16522 ( .B1(n13360), .B2(n13359), .A(n14197), .ZN(n13363) );
  NAND2_X1 U16523 ( .A1(n13368), .A2(n13361), .ZN(n13362) );
  NAND2_X1 U16524 ( .A1(n20398), .A2(n16069), .ZN(n13364) );
  NAND4_X1 U16525 ( .A1(n13365), .A2(n10063), .A3(n21119), .A4(n13364), .ZN(
        n13366) );
  OAI211_X1 U16526 ( .C1(n13369), .C2(n13368), .A(n13367), .B(n13366), .ZN(
        n13370) );
  INV_X1 U16527 ( .A(n13370), .ZN(n13371) );
  NAND2_X1 U16528 ( .A1(n13372), .A2(n13371), .ZN(n13373) );
  OAI21_X1 U16529 ( .B1(n10625), .B2(n13378), .A(n13374), .ZN(n13375) );
  NOR2_X1 U16530 ( .A1(n9778), .A2(n13375), .ZN(n13377) );
  OR2_X1 U16531 ( .A1(n13378), .A2(n20412), .ZN(n13379) );
  AND2_X1 U16532 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  OAI21_X1 U16533 ( .B1(n13383), .B2(n9755), .A(n13382), .ZN(n13384) );
  NOR2_X1 U16534 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  NAND2_X1 U16535 ( .A1(n14783), .A2(n14769), .ZN(n13513) );
  AND2_X1 U16536 ( .A1(n14784), .A2(n13513), .ZN(n13389) );
  NAND2_X1 U16537 ( .A1(n16368), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20371) );
  INV_X1 U16538 ( .A(n20371), .ZN(n13388) );
  AOI211_X1 U16539 ( .C1(n16395), .C2(n14371), .A(n13389), .B(n13388), .ZN(
        n13392) );
  INV_X1 U16540 ( .A(n14802), .ZN(n13511) );
  NAND2_X1 U16541 ( .A1(n20243), .A2(n13390), .ZN(n13534) );
  INV_X1 U16542 ( .A(n13534), .ZN(n13512) );
  OAI21_X1 U16543 ( .B1(n13511), .B2(n13512), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13391) );
  OAI211_X1 U16544 ( .C1(n13393), .C2(n16319), .A(n13392), .B(n13391), .ZN(
        P1_U3031) );
  NOR2_X1 U16545 ( .A1(n13342), .A2(n13893), .ZN(n13394) );
  OAI211_X1 U16546 ( .C1(n13394), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19386), .B(n13443), .ZN(n13399) );
  OR2_X1 U16547 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  AND2_X1 U16548 ( .A1(n13397), .A2(n13444), .ZN(n19315) );
  NAND2_X1 U16549 ( .A1(n19356), .A2(n19315), .ZN(n13398) );
  OAI211_X1 U16550 ( .C1(n19356), .C2(n19308), .A(n13399), .B(n13398), .ZN(
        P2_U2881) );
  NOR2_X1 U16551 ( .A1(n13409), .A2(n14197), .ZN(n13405) );
  INV_X1 U16552 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13406) );
  OR2_X1 U16553 ( .A1(n20379), .A2(n13406), .ZN(n13408) );
  NAND2_X1 U16554 ( .A1(n20379), .A2(DATAI_0_), .ZN(n13407) );
  NAND2_X1 U16555 ( .A1(n13408), .A2(n13407), .ZN(n20390) );
  INV_X1 U16556 ( .A(n20390), .ZN(n13411) );
  NAND2_X1 U16557 ( .A1(n14546), .A2(n13409), .ZN(n14465) );
  INV_X1 U16558 ( .A(n14197), .ZN(n13410) );
  INV_X1 U16559 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20335) );
  OAI222_X1 U16560 ( .A1(n14553), .A2(n20374), .B1(n13411), .B2(n14548), .C1(
        n14546), .C2(n20335), .ZN(P1_U2904) );
  AOI22_X1 U16561 ( .A1(n13158), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13412) );
  OAI21_X1 U16562 ( .B1(n13413), .B2(n13423), .A(n13412), .ZN(P2_U2935) );
  INV_X1 U16563 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16564 ( .A1(n13158), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13414) );
  OAI21_X1 U16565 ( .B1(n13415), .B2(n13423), .A(n13414), .ZN(P2_U2933) );
  INV_X1 U16566 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U16567 ( .A1(n13158), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13416) );
  OAI21_X1 U16568 ( .B1(n15079), .B2(n13423), .A(n13416), .ZN(P2_U2930) );
  INV_X1 U16569 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U16570 ( .A1(n13158), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U16571 ( .B1(n15065), .B2(n13423), .A(n13417), .ZN(P2_U2928) );
  INV_X1 U16572 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U16573 ( .A1(n13158), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13418) );
  OAI21_X1 U16574 ( .B1(n13419), .B2(n13423), .A(n13418), .ZN(P2_U2931) );
  INV_X1 U16575 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21333) );
  AOI22_X1 U16576 ( .A1(n13158), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13420) );
  OAI21_X1 U16577 ( .B1(n21333), .B2(n13423), .A(n13420), .ZN(P2_U2934) );
  INV_X1 U16578 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15084) );
  AOI22_X1 U16579 ( .A1(n13158), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13421) );
  OAI21_X1 U16580 ( .B1(n15084), .B2(n13423), .A(n13421), .ZN(P2_U2932) );
  INV_X1 U16581 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U16582 ( .A1(n13158), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16583 ( .B1(n15074), .B2(n13423), .A(n13422), .ZN(P2_U2929) );
  INV_X1 U16584 ( .A(n15027), .ZN(n13426) );
  OR2_X1 U16585 ( .A1(n15590), .A2(n13424), .ZN(n13425) );
  NAND2_X1 U16586 ( .A1(n15569), .A2(n13425), .ZN(n19272) );
  INV_X1 U16587 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19438) );
  OAI222_X1 U16588 ( .A1(n13679), .A2(n13426), .B1(n19272), .B2(n19428), .C1(
        n19438), .C2(n15094), .ZN(P2_U2908) );
  INV_X1 U16589 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16590 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16591 ( .B1(n13428), .B2(n13441), .A(n13427), .ZN(P1_U2920) );
  INV_X1 U16592 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21338) );
  AOI22_X1 U16593 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16594 ( .B1(n21338), .B2(n13441), .A(n13429), .ZN(P1_U2915) );
  INV_X1 U16595 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16596 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U16597 ( .B1(n13431), .B2(n13441), .A(n13430), .ZN(P1_U2914) );
  INV_X1 U16598 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U16599 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13432) );
  OAI21_X1 U16600 ( .B1(n13433), .B2(n13441), .A(n13432), .ZN(P1_U2917) );
  INV_X1 U16601 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16602 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U16603 ( .B1(n13435), .B2(n13441), .A(n13434), .ZN(P1_U2916) );
  INV_X1 U16604 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U16605 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U16606 ( .B1(n13437), .B2(n13441), .A(n13436), .ZN(P1_U2918) );
  INV_X1 U16607 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U16608 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13438) );
  OAI21_X1 U16609 ( .B1(n13439), .B2(n13441), .A(n13438), .ZN(P1_U2919) );
  INV_X1 U16610 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U16611 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13440) );
  OAI21_X1 U16612 ( .B1(n13442), .B2(n13441), .A(n13440), .ZN(P1_U2913) );
  XOR2_X1 U16613 ( .A(n13443), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13448)
         );
  INV_X1 U16614 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13446) );
  AOI21_X1 U16615 ( .B1(n13445), .B2(n13444), .A(n13775), .ZN(n15635) );
  INV_X1 U16616 ( .A(n15635), .ZN(n19299) );
  MUX2_X1 U16617 ( .A(n13446), .B(n19299), .S(n19356), .Z(n13447) );
  OAI21_X1 U16618 ( .B1(n13448), .B2(n19380), .A(n13447), .ZN(P2_U2880) );
  OAI21_X1 U16619 ( .B1(n13450), .B2(n13449), .A(n13593), .ZN(n13500) );
  MUX2_X1 U16620 ( .A(BUF1_REG_1__SCAN_IN), .B(DATAI_1_), .S(n20379), .Z(
        n20399) );
  INV_X1 U16621 ( .A(n20399), .ZN(n13451) );
  INV_X1 U16622 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20330) );
  OAI222_X1 U16623 ( .A1(n14553), .A2(n13500), .B1(n13451), .B2(n14548), .C1(
        n14546), .C2(n20330), .ZN(P1_U2903) );
  AOI22_X1 U16624 ( .A1(n20363), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20360), .ZN(n13454) );
  NAND2_X1 U16625 ( .A1(n20348), .A2(n20399), .ZN(n13489) );
  NAND2_X1 U16626 ( .A1(n13454), .A2(n13489), .ZN(P1_U2953) );
  AOI22_X1 U16627 ( .A1(n20363), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20360), .ZN(n13455) );
  MUX2_X1 U16628 ( .A(BUF1_REG_5__SCAN_IN), .B(DATAI_5_), .S(n20379), .Z(
        n20416) );
  NAND2_X1 U16629 ( .A1(n20348), .A2(n20416), .ZN(n13479) );
  NAND2_X1 U16630 ( .A1(n13455), .A2(n13479), .ZN(P1_U2957) );
  AOI22_X1 U16631 ( .A1(n20363), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20360), .ZN(n13458) );
  OR2_X1 U16632 ( .A1(n20379), .A2(n16768), .ZN(n13457) );
  NAND2_X1 U16633 ( .A1(n20379), .A2(DATAI_4_), .ZN(n13456) );
  NAND2_X1 U16634 ( .A1(n13457), .A2(n13456), .ZN(n20413) );
  NAND2_X1 U16635 ( .A1(n20348), .A2(n20413), .ZN(n13481) );
  NAND2_X1 U16636 ( .A1(n13458), .A2(n13481), .ZN(P1_U2956) );
  AOI22_X1 U16637 ( .A1(n20363), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20360), .ZN(n13462) );
  INV_X1 U16638 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13459) );
  OR2_X1 U16639 ( .A1(n20379), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U16640 ( .A1(n20379), .A2(DATAI_6_), .ZN(n13460) );
  NAND2_X1 U16641 ( .A1(n13461), .A2(n13460), .ZN(n20419) );
  NAND2_X1 U16642 ( .A1(n20348), .A2(n20419), .ZN(n13477) );
  NAND2_X1 U16643 ( .A1(n13462), .A2(n13477), .ZN(P1_U2958) );
  AOI22_X1 U16644 ( .A1(n20363), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20360), .ZN(n13466) );
  INV_X1 U16645 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13463) );
  OR2_X1 U16646 ( .A1(n20379), .A2(n13463), .ZN(n13465) );
  NAND2_X1 U16647 ( .A1(n20379), .A2(DATAI_2_), .ZN(n13464) );
  NAND2_X1 U16648 ( .A1(n13465), .A2(n13464), .ZN(n20405) );
  NAND2_X1 U16649 ( .A1(n20348), .A2(n20405), .ZN(n13487) );
  NAND2_X1 U16650 ( .A1(n13466), .A2(n13487), .ZN(P1_U2954) );
  AOI22_X1 U16651 ( .A1(n20363), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20360), .ZN(n13467) );
  NAND2_X1 U16652 ( .A1(n20348), .A2(n20390), .ZN(n13485) );
  NAND2_X1 U16653 ( .A1(n13467), .A2(n13485), .ZN(P1_U2937) );
  AOI22_X1 U16654 ( .A1(n20363), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20360), .ZN(n13471) );
  INV_X1 U16655 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13468) );
  OR2_X1 U16656 ( .A1(n20379), .A2(n13468), .ZN(n13470) );
  NAND2_X1 U16657 ( .A1(n20379), .A2(DATAI_3_), .ZN(n13469) );
  NAND2_X1 U16658 ( .A1(n13470), .A2(n13469), .ZN(n20409) );
  NAND2_X1 U16659 ( .A1(n20348), .A2(n20409), .ZN(n13491) );
  NAND2_X1 U16660 ( .A1(n13471), .A2(n13491), .ZN(P1_U2955) );
  AOI22_X1 U16661 ( .A1(n20363), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20360), .ZN(n13475) );
  INV_X1 U16662 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13472) );
  OR2_X1 U16663 ( .A1(n20379), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U16664 ( .A1(n20379), .A2(DATAI_9_), .ZN(n13473) );
  NAND2_X1 U16665 ( .A1(n13474), .A2(n13473), .ZN(n14497) );
  NAND2_X1 U16666 ( .A1(n20348), .A2(n14497), .ZN(n20352) );
  NAND2_X1 U16667 ( .A1(n13475), .A2(n20352), .ZN(P1_U2946) );
  AOI22_X1 U16668 ( .A1(n20363), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20360), .ZN(n13476) );
  MUX2_X1 U16669 ( .A(BUF1_REG_7__SCAN_IN), .B(DATAI_7_), .S(n20379), .Z(
        n20428) );
  NAND2_X1 U16670 ( .A1(n20348), .A2(n20428), .ZN(n13483) );
  NAND2_X1 U16671 ( .A1(n13476), .A2(n13483), .ZN(P1_U2944) );
  AOI22_X1 U16672 ( .A1(n20363), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20360), .ZN(n13478) );
  NAND2_X1 U16673 ( .A1(n13478), .A2(n13477), .ZN(P1_U2943) );
  AOI22_X1 U16674 ( .A1(n20363), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20360), .ZN(n13480) );
  NAND2_X1 U16675 ( .A1(n13480), .A2(n13479), .ZN(P1_U2942) );
  AOI22_X1 U16676 ( .A1(n20363), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20360), .ZN(n13482) );
  NAND2_X1 U16677 ( .A1(n13482), .A2(n13481), .ZN(P1_U2941) );
  AOI22_X1 U16678 ( .A1(n20363), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20360), .ZN(n13484) );
  NAND2_X1 U16679 ( .A1(n13484), .A2(n13483), .ZN(P1_U2959) );
  AOI22_X1 U16680 ( .A1(n20363), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20360), .ZN(n13486) );
  NAND2_X1 U16681 ( .A1(n13486), .A2(n13485), .ZN(P1_U2952) );
  AOI22_X1 U16682 ( .A1(n20363), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20360), .ZN(n13488) );
  NAND2_X1 U16683 ( .A1(n13488), .A2(n13487), .ZN(P1_U2939) );
  AOI22_X1 U16684 ( .A1(n20363), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20360), .ZN(n13490) );
  NAND2_X1 U16685 ( .A1(n13490), .A2(n13489), .ZN(P1_U2938) );
  AOI22_X1 U16686 ( .A1(n20363), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20360), .ZN(n13492) );
  NAND2_X1 U16687 ( .A1(n13492), .A2(n13491), .ZN(P1_U2940) );
  INV_X1 U16688 ( .A(n20129), .ZN(n13499) );
  NOR2_X1 U16689 ( .A1(n20127), .A2(n20129), .ZN(n13553) );
  AOI21_X1 U16690 ( .B1(n20127), .B2(n20129), .A(n13553), .ZN(n13494) );
  NAND2_X1 U16691 ( .A1(n13494), .A2(n13493), .ZN(n13555) );
  OAI21_X1 U16692 ( .B1(n13494), .B2(n13493), .A(n13555), .ZN(n13495) );
  NAND2_X1 U16693 ( .A1(n13495), .A2(n16501), .ZN(n13498) );
  INV_X1 U16694 ( .A(n13679), .ZN(n19421) );
  INV_X1 U16695 ( .A(n15095), .ZN(n13496) );
  AOI22_X1 U16696 ( .A1(n19421), .A2(n13496), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19419), .ZN(n13497) );
  OAI211_X1 U16697 ( .C1(n13499), .C2(n19400), .A(n13498), .B(n13497), .ZN(
        P2_U2918) );
  INV_X1 U16698 ( .A(n13500), .ZN(n20282) );
  INV_X1 U16699 ( .A(n14452), .ZN(n20299) );
  INV_X1 U16700 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20277) );
  NAND2_X1 U16701 ( .A1(n14103), .A2(n20277), .ZN(n13503) );
  INV_X2 U16702 ( .A(n14082), .ZN(n14143) );
  NAND2_X1 U16703 ( .A1(n14143), .A2(n20277), .ZN(n13501) );
  OAI211_X1 U16704 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n14139), .A(
        n13501), .B(n14208), .ZN(n13502) );
  NAND2_X1 U16705 ( .A1(n13503), .A2(n13502), .ZN(n13539) );
  XNOR2_X1 U16706 ( .A(n13539), .B(n13504), .ZN(n13505) );
  NAND2_X1 U16707 ( .A1(n13505), .A2(n14143), .ZN(n13540) );
  OR2_X1 U16708 ( .A1(n13505), .A2(n14143), .ZN(n13506) );
  NAND2_X1 U16709 ( .A1(n13540), .A2(n13506), .ZN(n13519) );
  INV_X1 U16710 ( .A(n13519), .ZN(n20278) );
  OAI22_X1 U16711 ( .A1(n20288), .A2(n20278), .B1(n20277), .B2(n20302), .ZN(
        n13507) );
  AOI21_X1 U16712 ( .B1(n20282), .B2(n20299), .A(n13507), .ZN(n13508) );
  INV_X1 U16713 ( .A(n13508), .ZN(P1_U2871) );
  XNOR2_X1 U16714 ( .A(n13509), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13530) );
  INV_X1 U16715 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21107) );
  NOR2_X1 U16716 ( .A1(n20243), .A2(n21107), .ZN(n13518) );
  INV_X1 U16717 ( .A(n13513), .ZN(n13510) );
  NOR2_X1 U16718 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13511), .ZN(
        n13538) );
  NOR2_X1 U16719 ( .A1(n16303), .A2(n13538), .ZN(n13516) );
  AOI21_X1 U16720 ( .B1(n14784), .B2(n13513), .A(n13512), .ZN(n13514) );
  INV_X1 U16721 ( .A(n13514), .ZN(n13515) );
  MUX2_X1 U16722 ( .A(n13516), .B(n13515), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13517) );
  AOI211_X1 U16723 ( .C1(n16395), .C2(n13519), .A(n13518), .B(n13517), .ZN(
        n13520) );
  OAI21_X1 U16724 ( .B1(n13530), .B2(n16319), .A(n13520), .ZN(P1_U3030) );
  XNOR2_X1 U16725 ( .A(n13521), .B(n19374), .ZN(n13526) );
  OR2_X1 U16726 ( .A1(n13523), .A2(n13522), .ZN(n13524) );
  AND2_X1 U16727 ( .A1(n13524), .A2(n15593), .ZN(n16529) );
  INV_X1 U16728 ( .A(n16529), .ZN(n19288) );
  MUX2_X1 U16729 ( .A(n10250), .B(n19288), .S(n19356), .Z(n13525) );
  OAI21_X1 U16730 ( .B1(n13526), .B2(n19380), .A(n13525), .ZN(P2_U2878) );
  AOI22_X1 U16731 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13527) );
  OAI21_X1 U16732 ( .B1(n16254), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13527), .ZN(n13528) );
  AOI21_X1 U16733 ( .B1(n20282), .B2(n20378), .A(n13528), .ZN(n13529) );
  OAI21_X1 U16734 ( .B1(n13530), .B2(n16244), .A(n13529), .ZN(P1_U2998) );
  XNOR2_X1 U16735 ( .A(n13532), .B(n13531), .ZN(n13598) );
  NAND2_X1 U16736 ( .A1(n14802), .A2(n14783), .ZN(n13818) );
  NOR2_X1 U16737 ( .A1(n13541), .A2(n13536), .ZN(n14692) );
  INV_X1 U16738 ( .A(n14783), .ZN(n13533) );
  NAND2_X1 U16739 ( .A1(n13533), .A2(n14784), .ZN(n13535) );
  OAI21_X1 U16740 ( .B1(n14844), .B2(n14692), .A(n14842), .ZN(n13647) );
  OAI21_X1 U16741 ( .B1(n14784), .B2(n13536), .A(n13541), .ZN(n13814) );
  NAND2_X1 U16742 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13537) );
  AOI221_X1 U16743 ( .B1(n13541), .B2(n13814), .C1(n13537), .C2(n13814), .A(
        n14769), .ZN(n13550) );
  INV_X1 U16744 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21054) );
  NAND3_X1 U16745 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14695), .A3(
        n13541), .ZN(n13548) );
  NAND2_X1 U16746 ( .A1(n13540), .A2(n13539), .ZN(n13545) );
  MUX2_X1 U16747 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13543) );
  NAND2_X1 U16748 ( .A1(n14082), .A2(n14139), .ZN(n14094) );
  OR2_X1 U16749 ( .A1(n14143), .A2(n13541), .ZN(n13542) );
  AND3_X1 U16750 ( .A1(n13543), .A2(n14094), .A3(n13542), .ZN(n13544) );
  NAND2_X1 U16751 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  AND2_X1 U16752 ( .A1(n13624), .A2(n13546), .ZN(n13600) );
  NAND2_X1 U16753 ( .A1(n16395), .A2(n13600), .ZN(n13547) );
  OAI211_X1 U16754 ( .C1(n21054), .C2(n20243), .A(n13548), .B(n13547), .ZN(
        n13549) );
  AOI211_X1 U16755 ( .C1(n13647), .C2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13550), .B(n13549), .ZN(n13551) );
  OAI21_X1 U16756 ( .B1(n16319), .B2(n13598), .A(n13551), .ZN(P1_U3029) );
  INV_X1 U16757 ( .A(n20117), .ZN(n13552) );
  INV_X1 U16758 ( .A(n13922), .ZN(n20119) );
  NOR2_X1 U16759 ( .A1(n13552), .A2(n20119), .ZN(n13609) );
  AOI21_X1 U16760 ( .B1(n13552), .B2(n20119), .A(n13609), .ZN(n13557) );
  INV_X1 U16761 ( .A(n13553), .ZN(n13554) );
  NAND2_X1 U16762 ( .A1(n13555), .A2(n13554), .ZN(n13556) );
  NAND2_X1 U16763 ( .A1(n13557), .A2(n13556), .ZN(n13611) );
  OAI21_X1 U16764 ( .B1(n13557), .B2(n13556), .A(n13611), .ZN(n13558) );
  NAND2_X1 U16765 ( .A1(n13558), .A2(n16501), .ZN(n13560) );
  AOI22_X1 U16766 ( .A1(n19392), .A2(n20119), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19419), .ZN(n13559) );
  OAI211_X1 U16767 ( .C1(n13679), .C2(n19468), .A(n13560), .B(n13559), .ZN(
        P2_U2917) );
  NOR2_X1 U16768 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21324), .ZN(n13581) );
  MUX2_X1 U16769 ( .A(n13561), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16026), .Z(n16028) );
  AOI22_X1 U16770 ( .A1(n13581), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16028), .B2(n21324), .ZN(n13577) );
  NAND2_X1 U16771 ( .A1(n20680), .A2(n14861), .ZN(n13572) );
  XNOR2_X1 U16772 ( .A(n13562), .B(n21260), .ZN(n13569) );
  OAI21_X1 U16773 ( .B1(n13563), .B2(n21260), .A(n9760), .ZN(n21100) );
  NAND2_X1 U16774 ( .A1(n13564), .A2(n21100), .ZN(n13567) );
  XNOR2_X1 U16775 ( .A(n13565), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13566) );
  OAI22_X1 U16776 ( .A1(n14861), .A2(n13567), .B1(n16020), .B2(n13566), .ZN(
        n13568) );
  AOI21_X1 U16777 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n13571) );
  NAND2_X1 U16778 ( .A1(n13572), .A2(n13571), .ZN(n21103) );
  INV_X1 U16779 ( .A(n16026), .ZN(n13573) );
  NAND2_X1 U16780 ( .A1(n21103), .A2(n13573), .ZN(n13575) );
  NAND2_X1 U16781 ( .A1(n16026), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13574) );
  NAND2_X1 U16782 ( .A1(n13575), .A2(n13574), .ZN(n16033) );
  AOI22_X1 U16783 ( .A1(n16033), .A2(n21324), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13581), .ZN(n13576) );
  OR2_X1 U16784 ( .A1(n13577), .A2(n13576), .ZN(n16040) );
  INV_X1 U16785 ( .A(n20535), .ZN(n20830) );
  XNOR2_X1 U16786 ( .A(n13578), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20242) );
  NOR2_X1 U16787 ( .A1(n20242), .A2(n13226), .ZN(n16404) );
  OAI21_X1 U16788 ( .B1(n16404), .B2(n16026), .A(n21324), .ZN(n13579) );
  AOI21_X1 U16789 ( .B1(n16026), .B2(n16406), .A(n13579), .ZN(n13580) );
  AOI21_X1 U16790 ( .B1(n13581), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13580), .ZN(n16039) );
  OAI21_X1 U16791 ( .B1(n13584), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13582), .ZN(
        n13583) );
  NAND2_X1 U16792 ( .A1(n21324), .A2(n21030), .ZN(n16413) );
  INV_X1 U16793 ( .A(n16413), .ZN(n21123) );
  NAND2_X1 U16794 ( .A1(n13583), .A2(n20544), .ZN(n20375) );
  NOR2_X1 U16795 ( .A1(n13584), .A2(n16416), .ZN(n16051) );
  NAND2_X1 U16796 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20840), .ZN(n13602) );
  INV_X1 U16797 ( .A(n13602), .ZN(n13585) );
  OAI22_X1 U16798 ( .A1(n20381), .A2(n20958), .B1(n14374), .B2(n13585), .ZN(
        n13586) );
  OAI21_X1 U16799 ( .B1(n16051), .B2(n13586), .A(n20375), .ZN(n13587) );
  OAI21_X1 U16800 ( .B1(n20375), .B2(n21321), .A(n13587), .ZN(P1_U3478) );
  INV_X1 U16801 ( .A(n15010), .ZN(n13590) );
  INV_X1 U16802 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19434) );
  OAI21_X1 U16803 ( .B1(n13589), .B2(n13588), .A(n13842), .ZN(n19244) );
  OAI222_X1 U16804 ( .A1(n13679), .A2(n13590), .B1(n15094), .B2(n19434), .C1(
        n19428), .C2(n19244), .ZN(P2_U2906) );
  INV_X1 U16805 ( .A(n13591), .ZN(n13592) );
  AOI21_X1 U16806 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13599) );
  AOI22_X1 U16807 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U16808 ( .B1(n16254), .B2(n14361), .A(n13595), .ZN(n13596) );
  AOI21_X1 U16809 ( .B1(n13599), .B2(n20378), .A(n13596), .ZN(n13597) );
  OAI21_X1 U16810 ( .B1(n16244), .B2(n13598), .A(n13597), .ZN(P1_U2997) );
  INV_X1 U16811 ( .A(n13599), .ZN(n14370) );
  INV_X1 U16812 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21147) );
  INV_X1 U16813 ( .A(n13600), .ZN(n14367) );
  OAI222_X1 U16814 ( .A1(n14370), .A2(n14452), .B1(n20302), .B2(n21147), .C1(
        n14367), .C2(n20288), .ZN(P1_U2870) );
  INV_X1 U16815 ( .A(n20405), .ZN(n13601) );
  INV_X1 U16816 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20328) );
  OAI222_X1 U16817 ( .A1(n14553), .A2(n14370), .B1(n13601), .B2(n14548), .C1(
        n14546), .C2(n20328), .ZN(P1_U2902) );
  NAND2_X1 U16818 ( .A1(n20375), .A2(n13602), .ZN(n14192) );
  NAND2_X1 U16819 ( .A1(n20375), .A2(n20826), .ZN(n14187) );
  NAND2_X1 U16820 ( .A1(n13604), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20793) );
  XNOR2_X1 U16821 ( .A(n13603), .B(n20793), .ZN(n13605) );
  OAI222_X1 U16822 ( .A1(n14192), .A2(n20831), .B1(n20375), .B2(n20679), .C1(
        n14187), .C2(n13605), .ZN(P1_U3476) );
  OR2_X1 U16823 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  NAND2_X1 U16824 ( .A1(n13608), .A2(n13671), .ZN(n20111) );
  XNOR2_X1 U16825 ( .A(n20106), .B(n20111), .ZN(n13613) );
  INV_X1 U16826 ( .A(n13609), .ZN(n13610) );
  NAND2_X1 U16827 ( .A1(n13611), .A2(n13610), .ZN(n13612) );
  NAND2_X1 U16828 ( .A1(n13612), .A2(n13613), .ZN(n13674) );
  OAI21_X1 U16829 ( .B1(n13613), .B2(n13612), .A(n13674), .ZN(n13614) );
  NAND2_X1 U16830 ( .A1(n13614), .A2(n16501), .ZN(n13617) );
  INV_X1 U16831 ( .A(n20111), .ZN(n13615) );
  AOI22_X1 U16832 ( .A1(n19392), .A2(n13615), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19419), .ZN(n13616) );
  OAI211_X1 U16833 ( .C1(n19473), .C2(n13679), .A(n13617), .B(n13616), .ZN(
        P2_U2916) );
  OR2_X1 U16834 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  AND2_X1 U16835 ( .A1(n13618), .A2(n13621), .ZN(n20263) );
  INV_X1 U16836 ( .A(n20263), .ZN(n13646) );
  MUX2_X1 U16837 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13623) );
  NAND2_X1 U16838 ( .A1(n14135), .A2(n13725), .ZN(n13622) );
  NAND2_X1 U16839 ( .A1(n13623), .A2(n13622), .ZN(n13625) );
  INV_X1 U16840 ( .A(n13739), .ZN(n16391) );
  AOI21_X1 U16841 ( .B1(n13625), .B2(n13624), .A(n16391), .ZN(n20259) );
  AOI22_X1 U16842 ( .A1(n20298), .A2(n20259), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14458), .ZN(n13626) );
  OAI21_X1 U16843 ( .B1(n13646), .B2(n14452), .A(n13626), .ZN(P1_U2869) );
  OR2_X1 U16844 ( .A1(n13627), .A2(n9914), .ZN(n13629) );
  INV_X1 U16845 ( .A(n15509), .ZN(n13628) );
  NAND2_X1 U16846 ( .A1(n13629), .A2(n13628), .ZN(n19232) );
  OAI222_X1 U16847 ( .A1(n13679), .A2(n13630), .B1(n19232), .B2(n19428), .C1(
        n13041), .C2(n15094), .ZN(P2_U2904) );
  XNOR2_X1 U16848 ( .A(n13632), .B(n13631), .ZN(n13652) );
  AND2_X1 U16849 ( .A1(n16368), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13649) );
  AOI21_X1 U16850 ( .B1(n20367), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13649), .ZN(n13633) );
  OAI21_X1 U16851 ( .B1(n16254), .B2(n20256), .A(n13633), .ZN(n13634) );
  AOI21_X1 U16852 ( .B1(n20263), .B2(n20378), .A(n13634), .ZN(n13635) );
  OAI21_X1 U16853 ( .B1(n13652), .B2(n16244), .A(n13635), .ZN(P1_U2996) );
  XNOR2_X1 U16854 ( .A(n13636), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13637) );
  XNOR2_X1 U16855 ( .A(n9768), .B(n13637), .ZN(n16591) );
  INV_X1 U16856 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13639) );
  OAI22_X1 U16857 ( .A1(n16565), .A2(n13793), .B1(n13639), .B2(n15303), .ZN(
        n13640) );
  AOI21_X1 U16858 ( .B1(n16555), .B2(n13791), .A(n13640), .ZN(n13642) );
  NAND2_X1 U16859 ( .A1(n9837), .A2(n16561), .ZN(n13641) );
  OAI211_X1 U16860 ( .C1(n16589), .C2(n16558), .A(n13642), .B(n13641), .ZN(
        n13643) );
  AOI21_X1 U16861 ( .B1(n16549), .B2(n16591), .A(n13643), .ZN(n13644) );
  INV_X1 U16862 ( .A(n13644), .ZN(P2_U3011) );
  INV_X1 U16863 ( .A(n20409), .ZN(n13645) );
  INV_X1 U16864 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20326) );
  OAI222_X1 U16865 ( .A1(n14553), .A2(n13646), .B1(n13645), .B2(n14548), .C1(
        n14546), .C2(n20326), .ZN(P1_U2901) );
  INV_X1 U16866 ( .A(n13647), .ZN(n13817) );
  OAI21_X1 U16867 ( .B1(n14769), .B2(n13814), .A(n13817), .ZN(n13722) );
  NAND2_X1 U16868 ( .A1(n14692), .A2(n14695), .ZN(n14848) );
  NAND2_X1 U16869 ( .A1(n14769), .A2(n14848), .ZN(n13819) );
  NAND2_X1 U16870 ( .A1(n13814), .A2(n13819), .ZN(n16398) );
  INV_X1 U16871 ( .A(n16398), .ZN(n13648) );
  AOI22_X1 U16872 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13722), .B1(
        n13648), .B2(n13725), .ZN(n13651) );
  AOI21_X1 U16873 ( .B1(n20259), .B2(n16395), .A(n13649), .ZN(n13650) );
  OAI211_X1 U16874 ( .C1(n16319), .C2(n13652), .A(n13651), .B(n13650), .ZN(
        P1_U3028) );
  INV_X1 U16875 ( .A(n20680), .ZN(n13660) );
  INV_X1 U16876 ( .A(n20380), .ZN(n13657) );
  NOR2_X1 U16877 ( .A1(n13603), .A2(n13653), .ZN(n20888) );
  INV_X1 U16878 ( .A(n13604), .ZN(n14188) );
  NAND2_X1 U16879 ( .A1(n20888), .A2(n14188), .ZN(n20864) );
  NAND3_X1 U16880 ( .A1(n20797), .A2(n20864), .A3(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13658) );
  INV_X1 U16881 ( .A(n20793), .ZN(n20493) );
  INV_X1 U16882 ( .A(n13654), .ZN(n13655) );
  AOI22_X1 U16883 ( .A1(n13658), .A2(n13657), .B1(n20493), .B2(n20637), .ZN(
        n13659) );
  OAI222_X1 U16884 ( .A1(n14192), .A2(n13660), .B1(n20375), .B2(n10574), .C1(
        n14187), .C2(n13659), .ZN(P1_U3475) );
  INV_X1 U16885 ( .A(n13661), .ZN(n19372) );
  INV_X1 U16886 ( .A(n13662), .ZN(n13664) );
  INV_X1 U16887 ( .A(n13663), .ZN(n19367) );
  OAI211_X1 U16888 ( .C1(n19372), .C2(n13664), .A(n19367), .B(n19386), .ZN(
        n13668) );
  AND2_X1 U16889 ( .A1(n9877), .A2(n13665), .ZN(n13666) );
  OR2_X1 U16890 ( .A1(n13666), .A2(n15300), .ZN(n15577) );
  INV_X1 U16891 ( .A(n15577), .ZN(n19268) );
  NAND2_X1 U16892 ( .A1(n19356), .A2(n19268), .ZN(n13667) );
  OAI211_X1 U16893 ( .C1(n19356), .C2(n13669), .A(n13668), .B(n13667), .ZN(
        P2_U2876) );
  NAND2_X1 U16894 ( .A1(n19504), .A2(n20111), .ZN(n13673) );
  AOI21_X1 U16895 ( .B1(n13672), .B2(n13671), .A(n13670), .ZN(n13761) );
  AOI21_X1 U16896 ( .B1(n13674), .B2(n13673), .A(n13761), .ZN(n19424) );
  OR2_X1 U16897 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  NAND2_X1 U16898 ( .A1(n13342), .A2(n13677), .ZN(n19423) );
  XNOR2_X1 U16899 ( .A(n19424), .B(n19423), .ZN(n13682) );
  INV_X1 U16900 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n13678) );
  OAI22_X1 U16901 ( .A1(n13679), .A2(n19477), .B1(n15094), .B2(n13678), .ZN(
        n13680) );
  AOI21_X1 U16902 ( .B1(n19392), .B2(n13761), .A(n13680), .ZN(n13681) );
  OAI21_X1 U16903 ( .B1(n13682), .B2(n19422), .A(n13681), .ZN(P2_U2915) );
  INV_X1 U16904 ( .A(n13683), .ZN(n19366) );
  XNOR2_X1 U16905 ( .A(n19366), .B(n19361), .ZN(n13687) );
  NAND2_X1 U16906 ( .A1(n15302), .A2(n13684), .ZN(n13685) );
  NAND2_X1 U16907 ( .A1(n13845), .A2(n13685), .ZN(n19243) );
  MUX2_X1 U16908 ( .A(n12051), .B(n19243), .S(n19356), .Z(n13686) );
  OAI21_X1 U16909 ( .B1(n13687), .B2(n19380), .A(n13686), .ZN(P2_U2874) );
  INV_X1 U16910 ( .A(n13751), .ZN(n13688) );
  AOI21_X1 U16911 ( .B1(n13689), .B2(n13618), .A(n13688), .ZN(n13719) );
  INV_X1 U16912 ( .A(n13719), .ZN(n20248) );
  INV_X1 U16913 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13692) );
  MUX2_X1 U16914 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13690) );
  OAI211_X1 U16915 ( .C1(n14143), .C2(n13691), .A(n13690), .B(n14094), .ZN(
        n16390) );
  XNOR2_X1 U16916 ( .A(n16391), .B(n16390), .ZN(n20237) );
  OAI222_X1 U16917 ( .A1(n20248), .A2(n14452), .B1(n13692), .B2(n20302), .C1(
        n20288), .C2(n20237), .ZN(P1_U2868) );
  INV_X1 U16918 ( .A(n20413), .ZN(n13693) );
  INV_X1 U16919 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21336) );
  OAI222_X1 U16920 ( .A1(n20248), .A2(n14553), .B1(n13693), .B2(n14548), .C1(
        n21336), .C2(n14546), .ZN(P1_U2900) );
  INV_X1 U16921 ( .A(n13694), .ZN(n13697) );
  INV_X1 U16922 ( .A(n13695), .ZN(n13696) );
  AOI21_X1 U16923 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13697), .A(
        n13696), .ZN(n13714) );
  XOR2_X1 U16924 ( .A(n13699), .B(n13698), .Z(n13712) );
  OR2_X1 U16925 ( .A1(n13701), .A2(n13700), .ZN(n13703) );
  NAND2_X1 U16926 ( .A1(n13703), .A2(n13702), .ZN(n19389) );
  INV_X1 U16927 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20051) );
  OAI22_X1 U16928 ( .A1(n20051), .A2(n15303), .B1(n16554), .B2(n13756), .ZN(
        n13704) );
  AOI21_X1 U16929 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16546), .A(
        n13704), .ZN(n13705) );
  OAI21_X1 U16930 ( .B1(n13882), .B2(n19389), .A(n13705), .ZN(n13706) );
  AOI21_X1 U16931 ( .B1(n13712), .B2(n16549), .A(n13706), .ZN(n13707) );
  OAI21_X1 U16932 ( .B1(n13714), .B2(n16558), .A(n13707), .ZN(P2_U3010) );
  NOR2_X1 U16933 ( .A1(n20051), .A2(n19305), .ZN(n13708) );
  AOI221_X1 U16934 ( .B1(n12290), .B2(n15645), .C1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13839), .A(n13708), .ZN(
        n13710) );
  NAND2_X1 U16935 ( .A1(n15602), .A2(n13761), .ZN(n13709) );
  OAI211_X1 U16936 ( .C1(n15600), .C2(n19389), .A(n13710), .B(n13709), .ZN(
        n13711) );
  AOI21_X1 U16937 ( .B1(n13712), .B2(n16592), .A(n13711), .ZN(n13713) );
  OAI21_X1 U16938 ( .B1(n13714), .B2(n16588), .A(n13713), .ZN(P2_U3042) );
  XOR2_X1 U16939 ( .A(n13715), .B(n13716), .Z(n13728) );
  INV_X1 U16940 ( .A(n13728), .ZN(n13721) );
  INV_X1 U16941 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20246) );
  OR2_X1 U16942 ( .A1(n20243), .A2(n20246), .ZN(n13723) );
  NAND2_X1 U16943 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13717) );
  OAI211_X1 U16944 ( .C1(n16254), .C2(n20244), .A(n13723), .B(n13717), .ZN(
        n13718) );
  AOI21_X1 U16945 ( .B1(n13719), .B2(n20378), .A(n13718), .ZN(n13720) );
  OAI21_X1 U16946 ( .B1(n13721), .B2(n16244), .A(n13720), .ZN(P1_U2995) );
  NAND2_X1 U16947 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13722), .ZN(
        n13724) );
  OAI211_X1 U16948 ( .C1(n20237), .C2(n16383), .A(n13724), .B(n13723), .ZN(
        n13727) );
  NAND2_X1 U16949 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14691) );
  INV_X1 U16950 ( .A(n14691), .ZN(n13815) );
  AOI211_X1 U16951 ( .C1(n13691), .C2(n13725), .A(n13815), .B(n16398), .ZN(
        n13726) );
  AOI211_X1 U16952 ( .C1(n13728), .C2(n16400), .A(n13727), .B(n13726), .ZN(
        n13729) );
  INV_X1 U16953 ( .A(n13729), .ZN(P1_U3027) );
  NOR2_X1 U16954 ( .A1(n13730), .A2(n13731), .ZN(n13732) );
  OR2_X1 U16955 ( .A1(n13803), .A2(n13732), .ZN(n20219) );
  INV_X1 U16956 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13734) );
  MUX2_X1 U16957 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13733) );
  OAI211_X1 U16958 ( .C1(n14143), .C2(n13734), .A(n13733), .B(n14094), .ZN(
        n16376) );
  OR2_X1 U16959 ( .A1(n14134), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n13737) );
  INV_X1 U16960 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21135) );
  NAND2_X1 U16961 ( .A1(n14143), .A2(n21135), .ZN(n13735) );
  OAI211_X1 U16962 ( .C1(n14149), .C2(n10850), .A(n13735), .B(n14120), .ZN(
        n13736) );
  AND2_X1 U16963 ( .A1(n13737), .A2(n13736), .ZN(n16389) );
  NAND2_X1 U16964 ( .A1(n16390), .A2(n16389), .ZN(n13738) );
  NOR2_X2 U16965 ( .A1(n13739), .A2(n13738), .ZN(n16392) );
  XOR2_X1 U16966 ( .A(n16376), .B(n16392), .Z(n20213) );
  AOI22_X1 U16967 ( .A1(n20213), .A2(n20298), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14458), .ZN(n13740) );
  OAI21_X1 U16968 ( .B1(n20219), .B2(n14452), .A(n13740), .ZN(P1_U2866) );
  INV_X1 U16969 ( .A(n20419), .ZN(n13741) );
  OAI222_X1 U16970 ( .A1(n20219), .A2(n14553), .B1(n13741), .B2(n14548), .C1(
        n20322), .C2(n14546), .ZN(P1_U2898) );
  INV_X1 U16971 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13749) );
  INV_X1 U16972 ( .A(n13742), .ZN(n13743) );
  OAI211_X1 U16973 ( .C1(n9845), .C2(n9918), .A(n13743), .B(n19386), .ZN(
        n13748) );
  NOR2_X1 U16974 ( .A1(n13846), .A2(n13744), .ZN(n13745) );
  OR2_X1 U16975 ( .A1(n15264), .A2(n13745), .ZN(n19233) );
  INV_X1 U16976 ( .A(n19233), .ZN(n13746) );
  NAND2_X1 U16977 ( .A1(n13746), .A2(n19356), .ZN(n13747) );
  OAI211_X1 U16978 ( .C1(n19356), .C2(n13749), .A(n13748), .B(n13747), .ZN(
        P2_U2872) );
  AND2_X1 U16979 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  NOR2_X1 U16980 ( .A1(n13730), .A2(n13752), .ZN(n20300) );
  INV_X1 U16981 ( .A(n20300), .ZN(n13755) );
  INV_X1 U16982 ( .A(n20416), .ZN(n13754) );
  OAI222_X1 U16983 ( .A1(n14553), .A2(n13755), .B1(n14548), .B2(n13754), .C1(
        n13753), .C2(n14546), .ZN(P1_U2899) );
  INV_X1 U16984 ( .A(n13756), .ZN(n13760) );
  NOR2_X1 U16985 ( .A1(n19312), .A2(n13757), .ZN(n13759) );
  AOI21_X1 U16986 ( .B1(n13760), .B2(n13759), .A(n20024), .ZN(n13758) );
  OAI21_X1 U16987 ( .B1(n13760), .B2(n13759), .A(n13758), .ZN(n13770) );
  INV_X1 U16988 ( .A(n13761), .ZN(n13762) );
  NOR2_X1 U16989 ( .A1(n19335), .A2(n13762), .ZN(n13763) );
  AOI211_X1 U16990 ( .C1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n19349), .A(
        n19326), .B(n13763), .ZN(n13766) );
  NAND2_X1 U16991 ( .A1(n19339), .A2(n13764), .ZN(n13765) );
  OAI211_X1 U16992 ( .C1(n20051), .C2(n19341), .A(n13766), .B(n13765), .ZN(
        n13768) );
  NOR2_X1 U16993 ( .A1(n19389), .A2(n19346), .ZN(n13767) );
  AOI211_X1 U16994 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19344), .A(n13768), .B(
        n13767), .ZN(n13769) );
  OAI211_X1 U16995 ( .C1(n19423), .C2(n13927), .A(n13770), .B(n13769), .ZN(
        P2_U2851) );
  NOR2_X1 U16996 ( .A1(n19312), .A2(n13771), .ZN(n13772) );
  XNOR2_X1 U16997 ( .A(n13772), .B(n16545), .ZN(n13773) );
  NAND2_X1 U16998 ( .A1(n13773), .A2(n19336), .ZN(n13786) );
  OAI21_X1 U16999 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(n19384) );
  AOI21_X1 U17000 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19349), .A(
        n19326), .ZN(n13781) );
  AOI21_X1 U17001 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n16570) );
  NAND2_X1 U17002 ( .A1(n19337), .A2(n16570), .ZN(n13780) );
  OAI211_X1 U17003 ( .C1(n19346), .C2(n19384), .A(n13781), .B(n13780), .ZN(
        n13784) );
  INV_X1 U17004 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13782) );
  NOR2_X1 U17005 ( .A1(n19324), .A2(n13782), .ZN(n13783) );
  AOI211_X1 U17006 ( .C1(n19327), .C2(P2_REIP_REG_8__SCAN_IN), .A(n13784), .B(
        n13783), .ZN(n13785) );
  OAI211_X1 U17007 ( .C1(n19306), .C2(n13787), .A(n13786), .B(n13785), .ZN(
        P2_U2847) );
  NAND2_X1 U17008 ( .A1(n9751), .A2(n13789), .ZN(n13790) );
  XNOR2_X1 U17009 ( .A(n13791), .B(n13790), .ZN(n13792) );
  NAND2_X1 U17010 ( .A1(n13792), .A2(n19336), .ZN(n13801) );
  OAI22_X1 U17011 ( .A1(n13793), .A2(n19282), .B1(n19335), .B2(n20111), .ZN(
        n13796) );
  NOR2_X1 U17012 ( .A1(n19306), .A2(n13794), .ZN(n13795) );
  AOI211_X1 U17013 ( .C1(n19327), .C2(P2_REIP_REG_3__SCAN_IN), .A(n13796), .B(
        n13795), .ZN(n13797) );
  OAI21_X1 U17014 ( .B1(n19324), .B2(n13798), .A(n13797), .ZN(n13799) );
  AOI21_X1 U17015 ( .B1(n9839), .B2(n12566), .A(n13799), .ZN(n13800) );
  OAI211_X1 U17016 ( .C1(n13927), .C2(n19504), .A(n13801), .B(n13800), .ZN(
        P2_U2852) );
  OR2_X1 U17017 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  AND2_X1 U17018 ( .A1(n13901), .A2(n13804), .ZN(n20294) );
  INV_X1 U17019 ( .A(n20294), .ZN(n13806) );
  INV_X1 U17020 ( .A(n20428), .ZN(n13805) );
  INV_X1 U17021 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20320) );
  OAI222_X1 U17022 ( .A1(n14553), .A2(n13806), .B1(n13805), .B2(n14548), .C1(
        n14546), .C2(n20320), .ZN(P1_U2897) );
  XOR2_X1 U17023 ( .A(n13808), .B(n13807), .Z(n13824) );
  INV_X1 U17024 ( .A(n20378), .ZN(n20373) );
  INV_X1 U17025 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21058) );
  NOR2_X1 U17026 ( .A1(n20243), .A2(n21058), .ZN(n13821) );
  AOI21_X1 U17027 ( .B1(n20367), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13821), .ZN(n13811) );
  INV_X1 U17028 ( .A(n20216), .ZN(n13809) );
  NAND2_X1 U17029 ( .A1(n16265), .A2(n13809), .ZN(n13810) );
  OAI211_X1 U17030 ( .C1(n20219), .C2(n20373), .A(n13811), .B(n13810), .ZN(
        n13812) );
  INV_X1 U17031 ( .A(n13812), .ZN(n13813) );
  OAI21_X1 U17032 ( .B1(n13824), .B2(n16244), .A(n13813), .ZN(P1_U2993) );
  NAND2_X1 U17033 ( .A1(n13815), .A2(n10850), .ZN(n16397) );
  NAND3_X1 U17034 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13815), .A3(
        n13814), .ZN(n16340) );
  NAND2_X1 U17035 ( .A1(n14847), .A2(n16340), .ZN(n13816) );
  NAND2_X1 U17036 ( .A1(n13817), .A2(n13816), .ZN(n16339) );
  AOI21_X1 U17037 ( .B1(n14691), .B2(n13818), .A(n16339), .ZN(n16403) );
  OAI21_X1 U17038 ( .B1(n14848), .B2(n16397), .A(n16403), .ZN(n16363) );
  INV_X1 U17039 ( .A(n13819), .ZN(n13820) );
  AOI22_X1 U17040 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16363), .B1(
        n16366), .B2(n13734), .ZN(n13823) );
  AOI21_X1 U17041 ( .B1(n20213), .B2(n16395), .A(n13821), .ZN(n13822) );
  OAI211_X1 U17042 ( .C1(n13824), .C2(n16319), .A(n13823), .B(n13822), .ZN(
        P1_U3025) );
  OAI21_X1 U17043 ( .B1(n13828), .B2(n13826), .A(n13825), .ZN(n13827) );
  OAI21_X1 U17044 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n16559) );
  OAI21_X1 U17045 ( .B1(n13670), .B2(n13831), .A(n13830), .ZN(n19427) );
  NAND2_X1 U17046 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13832) );
  OAI211_X1 U17047 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15645), .B(n13832), .ZN(n13834) );
  AOI22_X1 U17048 ( .A1(n16586), .A2(n19331), .B1(n19326), .B2(
        P2_REIP_REG_5__SCAN_IN), .ZN(n13833) );
  OAI211_X1 U17049 ( .C1(n19427), .C2(n16581), .A(n13834), .B(n13833), .ZN(
        n13838) );
  XNOR2_X1 U17050 ( .A(n13836), .B(n13835), .ZN(n16556) );
  NOR2_X1 U17051 ( .A1(n16556), .A2(n15632), .ZN(n13837) );
  AOI211_X1 U17052 ( .C1(n13839), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13838), .B(n13837), .ZN(n13840) );
  OAI21_X1 U17053 ( .B1(n16588), .B2(n16559), .A(n13840), .ZN(P2_U3041) );
  AOI21_X1 U17054 ( .B1(n13842), .B2(n13841), .A(n9914), .ZN(n13843) );
  INV_X1 U17055 ( .A(n13843), .ZN(n19408) );
  AND2_X1 U17056 ( .A1(n13845), .A2(n13844), .ZN(n13847) );
  OR2_X1 U17057 ( .A1(n13847), .A2(n13846), .ZN(n19365) );
  AOI22_X1 U17058 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19349), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19327), .ZN(n13848) );
  OAI211_X1 U17059 ( .C1(n19324), .C2(n12203), .A(n13848), .B(n15303), .ZN(
        n13849) );
  INV_X1 U17060 ( .A(n13849), .ZN(n13850) );
  OAI21_X1 U17061 ( .B1(n19365), .B2(n19346), .A(n13850), .ZN(n13853) );
  NOR2_X1 U17062 ( .A1(n19312), .A2(n13855), .ZN(n13851) );
  NOR3_X1 U17063 ( .A1(n13851), .A2(n20024), .A3(n16520), .ZN(n13852) );
  AOI211_X1 U17064 ( .C1(n19339), .C2(n13854), .A(n13853), .B(n13852), .ZN(
        n13857) );
  NOR3_X1 U17065 ( .A1(n19312), .A2(n13855), .A3(n20024), .ZN(n19247) );
  NAND2_X1 U17066 ( .A1(n19247), .A2(n16520), .ZN(n13856) );
  OAI211_X1 U17067 ( .C1(n19408), .C2(n19335), .A(n13857), .B(n13856), .ZN(
        P2_U2841) );
  OAI22_X1 U17068 ( .A1(n9751), .A2(n13273), .B1(n19352), .B2(n19312), .ZN(
        n13858) );
  INV_X1 U17069 ( .A(n13858), .ZN(n15657) );
  OR2_X1 U17070 ( .A1(n9816), .A2(n15660), .ZN(n13863) );
  INV_X1 U17071 ( .A(n15673), .ZN(n15686) );
  INV_X1 U17072 ( .A(n13859), .ZN(n13860) );
  NOR2_X1 U17073 ( .A1(n13860), .A2(n12600), .ZN(n15663) );
  MUX2_X1 U17074 ( .A(n15686), .B(n15663), .S(n13861), .Z(n13862) );
  NAND2_X1 U17075 ( .A1(n13863), .A2(n13862), .ZN(n16599) );
  AOI222_X1 U17076 ( .A1(n15657), .A2(P2_STATE2_REG_1__SCAN_IN), .B1(n13864), 
        .B2(n15655), .C1(n16599), .C2(n20021), .ZN(n13877) );
  NOR3_X1 U17077 ( .A1(n20132), .A2(n21322), .A3(n15656), .ZN(n16073) );
  INV_X1 U17078 ( .A(n13865), .ZN(n13866) );
  NAND2_X1 U17079 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  NOR2_X1 U17080 ( .A1(n13869), .A2(n13868), .ZN(n13873) );
  NAND3_X1 U17081 ( .A1(n13871), .A2(n16625), .A3(n13870), .ZN(n13872) );
  NAND2_X1 U17082 ( .A1(n21322), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16642) );
  OAI21_X1 U17083 ( .B1(n16611), .B2(n13874), .A(n16642), .ZN(n13875) );
  AOI21_X1 U17084 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16073), .A(n13875), .ZN(
        n15826) );
  NAND2_X1 U17085 ( .A1(n15826), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13876) );
  OAI21_X1 U17086 ( .B1(n13877), .B2(n15826), .A(n13876), .ZN(P2_U3601) );
  NAND2_X1 U17087 ( .A1(n19500), .A2(n19661), .ZN(n19532) );
  OAI21_X1 U17088 ( .B1(n20015), .B2(n19524), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13878) );
  NAND2_X1 U17089 ( .A1(n13878), .A2(n20102), .ZN(n13890) );
  INV_X1 U17090 ( .A(n13890), .ZN(n13880) );
  NOR2_X1 U17091 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19563) );
  INV_X1 U17092 ( .A(n19563), .ZN(n19565) );
  NOR2_X1 U17093 ( .A1(n19719), .A2(n19565), .ZN(n19491) );
  INV_X1 U17094 ( .A(n19491), .ZN(n13895) );
  AND2_X1 U17095 ( .A1(n19955), .A2(n13895), .ZN(n13889) );
  AOI22_X1 U17096 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19494), .ZN(n19901) );
  INV_X1 U17097 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16744) );
  INV_X1 U17098 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21230) );
  INV_X1 U17099 ( .A(n19490), .ZN(n13894) );
  NAND2_X1 U17100 ( .A1(n13894), .A2(n13885), .ZN(n19521) );
  OAI22_X1 U17101 ( .A1(n19864), .A2(n19532), .B1(n19521), .B2(n13895), .ZN(
        n13886) );
  AOI21_X1 U17102 ( .B1(n20015), .B2(n19997), .A(n13886), .ZN(n13892) );
  OAI21_X1 U17103 ( .B1(n13887), .B2(n19491), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13888) );
  NOR2_X2 U17104 ( .A1(n19418), .A2(n19917), .ZN(n19995) );
  NAND2_X1 U17105 ( .A1(n19495), .A2(n19995), .ZN(n13891) );
  OAI211_X1 U17106 ( .C1(n19499), .C2(n13893), .A(n13892), .B(n13891), .ZN(
        P2_U3053) );
  AOI22_X1 U17107 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19494), .ZN(n19889) );
  INV_X1 U17108 ( .A(n19889), .ZN(n19969) );
  AOI22_X1 U17109 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19494), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19493), .ZN(n19823) );
  NAND2_X1 U17110 ( .A1(n13894), .A2(n20155), .ZN(n19512) );
  OAI22_X1 U17111 ( .A1(n19823), .A2(n19532), .B1(n19512), .B2(n13895), .ZN(
        n13896) );
  AOI21_X1 U17112 ( .B1(n20015), .B2(n19969), .A(n13896), .ZN(n13898) );
  NOR2_X2 U17113 ( .A1(n15095), .A2(n19917), .ZN(n19968) );
  NAND2_X1 U17114 ( .A1(n19495), .A2(n19968), .ZN(n13897) );
  OAI211_X1 U17115 ( .C1(n19499), .C2(n13899), .A(n13898), .B(n13897), .ZN(
        P2_U3049) );
  AOI21_X1 U17116 ( .B1(n13902), .B2(n13901), .A(n11020), .ZN(n13933) );
  INV_X1 U17117 ( .A(n13933), .ZN(n14356) );
  INV_X1 U17118 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16762) );
  OR2_X1 U17119 ( .A1(n20379), .A2(n16762), .ZN(n13904) );
  NAND2_X1 U17120 ( .A1(n20379), .A2(DATAI_8_), .ZN(n13903) );
  NAND2_X1 U17121 ( .A1(n13904), .A2(n13903), .ZN(n20336) );
  AOI22_X1 U17122 ( .A1(n14555), .A2(n20336), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16190), .ZN(n13905) );
  OAI21_X1 U17123 ( .B1(n14356), .B2(n14553), .A(n13905), .ZN(P1_U2896) );
  INV_X1 U17124 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13913) );
  OR2_X1 U17125 ( .A1(n14134), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n13908) );
  INV_X1 U17126 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20296) );
  NAND2_X1 U17127 ( .A1(n14143), .A2(n20296), .ZN(n13906) );
  OAI211_X1 U17128 ( .C1(n14149), .C2(n16387), .A(n13906), .B(n14120), .ZN(
        n13907) );
  AND2_X1 U17129 ( .A1(n13908), .A2(n13907), .ZN(n16375) );
  AND2_X1 U17130 ( .A1(n16376), .A2(n16375), .ZN(n13909) );
  MUX2_X1 U17131 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13911) );
  INV_X1 U17132 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16374) );
  OR2_X1 U17133 ( .A1(n16374), .A2(n14143), .ZN(n13910) );
  NAND3_X1 U17134 ( .A1(n13911), .A2(n14094), .A3(n13910), .ZN(n13912) );
  NAND2_X1 U17135 ( .A1(n16378), .A2(n13912), .ZN(n16353) );
  OAI21_X1 U17136 ( .B1(n16378), .B2(n13912), .A(n16353), .ZN(n16370) );
  OAI222_X1 U17137 ( .A1(n14356), .A2(n14452), .B1(n20302), .B2(n13913), .C1(
        n16370), .C2(n20288), .ZN(P1_U2864) );
  NOR2_X1 U17138 ( .A1(n19312), .A2(n13914), .ZN(n13940) );
  INV_X1 U17139 ( .A(n13940), .ZN(n13915) );
  AOI221_X1 U17140 ( .B1(n13917), .B2(n13940), .C1(n13916), .C2(n13915), .A(
        n20024), .ZN(n13918) );
  INV_X1 U17141 ( .A(n13918), .ZN(n13926) );
  NAND2_X1 U17142 ( .A1(n19339), .A2(n13919), .ZN(n13921) );
  AOI22_X1 U17143 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19327), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19349), .ZN(n13920) );
  OAI211_X1 U17144 ( .C1(n13922), .C2(n19335), .A(n13921), .B(n13920), .ZN(
        n13924) );
  NOR2_X1 U17145 ( .A1(n10117), .A2(n19346), .ZN(n13923) );
  AOI211_X1 U17146 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n19344), .A(n13924), .B(
        n13923), .ZN(n13925) );
  OAI211_X1 U17147 ( .C1(n20117), .C2(n13927), .A(n13926), .B(n13925), .ZN(
        P2_U2853) );
  NAND2_X1 U17148 ( .A1(n9927), .A2(n13928), .ZN(n13929) );
  XNOR2_X1 U17149 ( .A(n13930), .B(n13929), .ZN(n16365) );
  AOI22_X1 U17150 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13931) );
  OAI21_X1 U17151 ( .B1(n16254), .B2(n14352), .A(n13931), .ZN(n13932) );
  AOI21_X1 U17152 ( .B1(n13933), .B2(n20378), .A(n13932), .ZN(n13934) );
  OAI21_X1 U17153 ( .B1(n16365), .B2(n16244), .A(n13934), .ZN(P1_U2991) );
  NAND2_X1 U17154 ( .A1(n13900), .A2(n13936), .ZN(n13937) );
  NAND2_X1 U17155 ( .A1(n13935), .A2(n13937), .ZN(n20289) );
  INV_X1 U17156 ( .A(n14497), .ZN(n13939) );
  OAI222_X1 U17157 ( .A1(n20289), .A2(n14553), .B1(n13939), .B2(n14548), .C1(
        n13938), .C2(n14546), .ZN(P1_U2895) );
  OAI21_X1 U17158 ( .B1(n19352), .B2(n13941), .A(n13940), .ZN(n15658) );
  NAND2_X1 U17159 ( .A1(n15665), .A2(n12566), .ZN(n13951) );
  NAND2_X1 U17160 ( .A1(n19344), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U17161 ( .A1(n19241), .A2(n13942), .ZN(n13944) );
  AOI22_X1 U17162 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19327), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19349), .ZN(n13943) );
  NAND2_X1 U17163 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  AOI21_X1 U17164 ( .B1(n19337), .B2(n20129), .A(n13945), .ZN(n13949) );
  INV_X1 U17165 ( .A(n13946), .ZN(n13947) );
  NAND2_X1 U17166 ( .A1(n19339), .A2(n13947), .ZN(n13948) );
  NAND4_X1 U17167 ( .A1(n13951), .A2(n13950), .A3(n13949), .A4(n13948), .ZN(
        n13952) );
  AOI21_X1 U17168 ( .B1(n20127), .B2(n19348), .A(n13952), .ZN(n13953) );
  OAI21_X1 U17169 ( .B1(n15658), .B2(n20024), .A(n13953), .ZN(P2_U2854) );
  INV_X1 U17170 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17019) );
  INV_X1 U17171 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17396) );
  INV_X1 U17172 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17393) );
  NOR3_X1 U17173 ( .A1(n17019), .A2(n17396), .A3(n17393), .ZN(n15695) );
  NAND3_X1 U17174 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15824) );
  OR2_X2 U17175 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15824), .ZN(
        n13976) );
  INV_X1 U17176 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15736) );
  AOI22_X1 U17177 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13957) );
  OR2_X2 U17178 ( .A1(n13962), .A2(n13958), .ZN(n13975) );
  AOI22_X1 U17179 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13956) );
  OAI211_X1 U17180 ( .C1(n13976), .C2(n15736), .A(n13957), .B(n13956), .ZN(
        n13971) );
  NAND3_X1 U17181 ( .A1(n19096), .A2(n19108), .A3(n18942), .ZN(n15882) );
  INV_X2 U17182 ( .A(n15882), .ZN(n13988) );
  AOI22_X1 U17183 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13969) );
  AOI22_X1 U17184 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13968) );
  INV_X2 U17185 ( .A(n17449), .ZN(n17470) );
  INV_X1 U17186 ( .A(n13962), .ZN(n13963) );
  AOI22_X1 U17187 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13967) );
  INV_X1 U17188 ( .A(n13964), .ZN(n13965) );
  NAND2_X1 U17189 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13966) );
  NAND4_X1 U17190 ( .A1(n13969), .A2(n13968), .A3(n13967), .A4(n13966), .ZN(
        n13970) );
  INV_X1 U17191 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21223) );
  INV_X1 U17192 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17432) );
  INV_X1 U17193 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17112) );
  INV_X1 U17194 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17493) );
  INV_X1 U17195 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17494) );
  INV_X1 U17196 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U17197 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13974) );
  OAI21_X1 U17198 ( .B1(n17449), .B2(n17451), .A(n13974), .ZN(n13985) );
  INV_X2 U17199 ( .A(n13975), .ZN(n17469) );
  AOI22_X1 U17200 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13983) );
  AOI22_X1 U17201 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13977) );
  OAI21_X1 U17202 ( .B1(n21197), .B2(n17381), .A(n13977), .ZN(n13981) );
  AOI22_X1 U17203 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U17204 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13978) );
  OAI211_X1 U17205 ( .C1(n17427), .C2(n18705), .A(n13979), .B(n13978), .ZN(
        n13980) );
  AOI211_X1 U17206 ( .C1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .C2(n17418), .A(
        n13981), .B(n13980), .ZN(n13982) );
  OAI211_X1 U17207 ( .C1(n21224), .C2(n9873), .A(n13983), .B(n13982), .ZN(
        n13984) );
  INV_X1 U17208 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18702) );
  AOI22_X1 U17209 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13987) );
  AOI22_X1 U17210 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13986) );
  OAI211_X1 U17211 ( .C1(n17427), .C2(n18702), .A(n13987), .B(n13986), .ZN(
        n13994) );
  AOI22_X1 U17212 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17213 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U17214 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U17215 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13989) );
  NAND4_X1 U17216 ( .A1(n13992), .A2(n13991), .A3(n13990), .A4(n13989), .ZN(
        n13993) );
  AOI22_X1 U17217 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17218 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U17219 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13997) );
  OAI211_X1 U17220 ( .C1(n17427), .C2(n21319), .A(n13998), .B(n13997), .ZN(
        n14004) );
  AOI22_X1 U17221 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U17222 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17379), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17223 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14000) );
  NAND2_X1 U17224 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13999) );
  NAND4_X1 U17225 ( .A1(n14002), .A2(n14001), .A3(n14000), .A4(n13999), .ZN(
        n14003) );
  AOI22_X1 U17226 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17227 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U17228 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14014) );
  INV_X1 U17229 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18716) );
  OAI22_X1 U17230 ( .A1(n17427), .A2(n18716), .B1(n9875), .B2(n15773), .ZN(
        n14012) );
  AOI22_X1 U17231 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17232 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17233 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U17234 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14007) );
  NAND4_X1 U17235 ( .A1(n14010), .A2(n14009), .A3(n14008), .A4(n14007), .ZN(
        n14011) );
  NAND2_X1 U17236 ( .A1(n17523), .A2(n18499), .ZN(n15813) );
  AOI22_X1 U17237 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14026) );
  INV_X2 U17238 ( .A(n9875), .ZN(n17453) );
  AOI22_X1 U17239 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14018) );
  AOI22_X1 U17240 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14017) );
  OAI211_X1 U17241 ( .C1(n17473), .C2(n21244), .A(n14018), .B(n14017), .ZN(
        n14024) );
  AOI22_X1 U17242 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17243 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17470), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U17244 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14020) );
  NAND2_X1 U17245 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14019) );
  NAND4_X1 U17246 ( .A1(n14022), .A2(n14021), .A3(n14020), .A4(n14019), .ZN(
        n14023) );
  AOI22_X1 U17247 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14036) );
  AOI22_X1 U17248 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U17249 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14027) );
  OAI211_X1 U17250 ( .C1(n17427), .C2(n18710), .A(n14028), .B(n14027), .ZN(
        n14034) );
  AOI22_X1 U17251 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17252 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17253 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14030) );
  NAND2_X1 U17254 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14029) );
  NAND4_X1 U17255 ( .A1(n14032), .A2(n14031), .A3(n14030), .A4(n14029), .ZN(
        n14033) );
  NOR2_X1 U17256 ( .A1(n14045), .A2(n15803), .ZN(n18933) );
  NAND2_X1 U17257 ( .A1(n14044), .A2(n18933), .ZN(n15794) );
  AOI22_X1 U17258 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14037) );
  OAI21_X1 U17259 ( .B1(n17450), .B2(n17305), .A(n14037), .ZN(n14043) );
  AOI22_X1 U17260 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14042) );
  INV_X1 U17261 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17313) );
  INV_X1 U17262 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17403) );
  OAI22_X1 U17263 ( .A1(n17427), .A2(n17313), .B1(n15882), .B2(n17403), .ZN(
        n14041) );
  AOI22_X1 U17264 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17265 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17266 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14038) );
  INV_X1 U17267 ( .A(n18495), .ZN(n15812) );
  NAND2_X1 U17268 ( .A1(n17527), .A2(n18488), .ZN(n15986) );
  OAI22_X1 U17269 ( .A1(n19114), .A2(n18958), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15807) );
  NAND2_X1 U17270 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14048), .ZN(
        n14050) );
  OAI22_X1 U17271 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18967), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14048), .ZN(n14052) );
  AOI21_X1 U17272 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14050), .A(
        n14052), .ZN(n14049) );
  NOR2_X1 U17273 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18967), .ZN(
        n14051) );
  AOI22_X1 U17274 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14052), .B1(
        n14051), .B2(n14050), .ZN(n14056) );
  OAI21_X1 U17275 ( .B1(n14055), .B2(n14054), .A(n14056), .ZN(n14053) );
  AOI21_X1 U17276 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19121), .A(
        n15806), .ZN(n15981) );
  NAND3_X1 U17277 ( .A1(n15807), .A2(n14056), .A3(n15981), .ZN(n14057) );
  NAND3_X1 U17278 ( .A1(n15808), .A2(n15809), .A3(n14057), .ZN(n16645) );
  NAND4_X1 U17279 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n17502) );
  NAND2_X1 U17280 ( .A1(n18511), .A2(n9907), .ZN(n17392) );
  NOR2_X1 U17281 ( .A1(n17396), .A2(n17393), .ZN(n14059) );
  AOI21_X1 U17282 ( .B1(n9907), .B2(n14059), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n14060) );
  NOR2_X1 U17283 ( .A1(n17363), .A2(n14060), .ZN(n14074) );
  INV_X1 U17284 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21325) );
  INV_X1 U17285 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18724) );
  OAI22_X1 U17286 ( .A1(n17381), .A2(n21325), .B1(n17467), .B2(n18724), .ZN(
        n14071) );
  AOI22_X1 U17287 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U17288 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14068) );
  INV_X1 U17289 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17290 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14061) );
  OAI21_X1 U17291 ( .B1(n17230), .B2(n14062), .A(n14061), .ZN(n14066) );
  AOI22_X1 U17292 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17293 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14063) );
  OAI211_X1 U17294 ( .C1(n13976), .C2(n17490), .A(n14064), .B(n14063), .ZN(
        n14065) );
  AOI211_X1 U17295 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14066), .B(n14065), .ZN(n14067) );
  NAND3_X1 U17296 ( .A1(n14069), .A2(n14068), .A3(n14067), .ZN(n14070) );
  AOI211_X1 U17297 ( .C1(n17349), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14071), .B(n14070), .ZN(n17604) );
  INV_X1 U17298 ( .A(n17604), .ZN(n14073) );
  MUX2_X1 U17299 ( .A(n14074), .B(n14073), .S(n17517), .Z(P3_U2688) );
  NOR2_X1 U17300 ( .A1(n16557), .A2(n14075), .ZN(n14076) );
  AOI211_X1 U17301 ( .C1(n16550), .C2(n14078), .A(n14077), .B(n14076), .ZN(
        n14081) );
  OAI21_X1 U17302 ( .B1(n16546), .B2(n14079), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14080) );
  OAI211_X1 U17303 ( .C1(n13882), .C2(n9816), .A(n14081), .B(n14080), .ZN(
        P2_U3014) );
  AOI22_X1 U17304 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n14082), .B1(
        n14145), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n14151) );
  NAND2_X1 U17305 ( .A1(n14145), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14084) );
  INV_X1 U17306 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14714) );
  OR2_X1 U17307 ( .A1(n14143), .A2(n14714), .ZN(n14083) );
  NAND2_X1 U17308 ( .A1(n14084), .A2(n14083), .ZN(n14209) );
  OR2_X1 U17309 ( .A1(n14134), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n14087) );
  INV_X1 U17310 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20292) );
  NAND2_X1 U17311 ( .A1(n14143), .A2(n20292), .ZN(n14085) );
  OAI211_X1 U17312 ( .C1(n14149), .C2(n16361), .A(n14085), .B(n14120), .ZN(
        n14086) );
  NAND2_X1 U17313 ( .A1(n14087), .A2(n14086), .ZN(n16352) );
  OR2_X1 U17314 ( .A1(n14146), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14090) );
  INV_X1 U17315 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14460) );
  NAND2_X1 U17316 ( .A1(n14143), .A2(n14460), .ZN(n14088) );
  OAI211_X1 U17317 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n14139), .A(
        n14088), .B(n14208), .ZN(n14089) );
  MUX2_X1 U17318 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14091) );
  MUX2_X1 U17319 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14095) );
  OR2_X1 U17320 ( .A1(n14092), .A2(n14143), .ZN(n14093) );
  MUX2_X1 U17321 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14096) );
  OAI21_X1 U17322 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14145), .A(
        n14096), .ZN(n14330) );
  NOR2_X1 U17323 ( .A1(n14450), .A2(n14330), .ZN(n14097) );
  OR2_X1 U17324 ( .A1(n14146), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14101) );
  INV_X1 U17325 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U17326 ( .A1(n14143), .A2(n14098), .ZN(n14099) );
  OAI211_X1 U17327 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n14139), .A(
        n14099), .B(n14208), .ZN(n14100) );
  MUX2_X1 U17328 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14102) );
  OAI21_X1 U17329 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14145), .A(
        n14102), .ZN(n14434) );
  INV_X1 U17330 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U17331 ( .A1(n14103), .A2(n14428), .ZN(n14106) );
  NAND2_X1 U17332 ( .A1(n14143), .A2(n14428), .ZN(n14104) );
  OAI211_X1 U17333 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n14139), .A(
        n14104), .B(n14208), .ZN(n14105) );
  NAND2_X1 U17334 ( .A1(n14106), .A2(n14105), .ZN(n14310) );
  INV_X1 U17335 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14427) );
  MUX2_X1 U17336 ( .A(n14208), .B(n14134), .S(n14427), .Z(n14108) );
  NAND2_X1 U17337 ( .A1(n14135), .A2(n10911), .ZN(n14107) );
  NAND2_X1 U17338 ( .A1(n14108), .A2(n14107), .ZN(n14423) );
  OR2_X1 U17339 ( .A1(n14146), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14111) );
  INV_X1 U17340 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16131) );
  NAND2_X1 U17341 ( .A1(n14143), .A2(n16131), .ZN(n14109) );
  OAI211_X1 U17342 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n14139), .A(
        n14109), .B(n14208), .ZN(n14110) );
  MUX2_X1 U17343 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14113) );
  NAND2_X1 U17344 ( .A1(n14135), .A2(n10912), .ZN(n14112) );
  AND2_X1 U17345 ( .A1(n14113), .A2(n14112), .ZN(n14407) );
  MUX2_X1 U17346 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14116) );
  OR2_X1 U17347 ( .A1(n14143), .A2(n14114), .ZN(n14115) );
  NAND2_X1 U17348 ( .A1(n14116), .A2(n14115), .ZN(n14402) );
  OR2_X1 U17349 ( .A1(n14134), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14119) );
  INV_X1 U17350 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U17351 ( .A1(n14143), .A2(n16189), .ZN(n14117) );
  OAI211_X1 U17352 ( .C1(n14149), .C2(n14795), .A(n14117), .B(n14120), .ZN(
        n14118) );
  NAND2_X1 U17353 ( .A1(n14119), .A2(n14118), .ZN(n14790) );
  MUX2_X1 U17354 ( .A(n14146), .B(n14120), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14122) );
  INV_X1 U17355 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21316) );
  OR2_X1 U17356 ( .A1(n14143), .A2(n21316), .ZN(n14121) );
  AND2_X1 U17357 ( .A1(n14122), .A2(n14121), .ZN(n14397) );
  OR2_X2 U17358 ( .A1(n9879), .A2(n14397), .ZN(n14399) );
  MUX2_X1 U17359 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14124) );
  INV_X1 U17360 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16284) );
  NAND2_X1 U17361 ( .A1(n14135), .A2(n16284), .ZN(n14123) );
  NAND2_X1 U17362 ( .A1(n14124), .A2(n14123), .ZN(n14295) );
  OR2_X1 U17363 ( .A1(n14146), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14127) );
  INV_X1 U17364 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14391) );
  NAND2_X1 U17365 ( .A1(n14143), .A2(n14391), .ZN(n14125) );
  OAI211_X1 U17366 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14139), .A(
        n14125), .B(n14208), .ZN(n14126) );
  NAND2_X1 U17367 ( .A1(n14127), .A2(n14126), .ZN(n14281) );
  MUX2_X1 U17368 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14129) );
  INV_X1 U17369 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14610) );
  NAND2_X1 U17370 ( .A1(n14135), .A2(n14610), .ZN(n14128) );
  NAND2_X1 U17371 ( .A1(n14129), .A2(n14128), .ZN(n14271) );
  OR2_X1 U17372 ( .A1(n14146), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14133) );
  INV_X1 U17373 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14130) );
  NAND2_X1 U17374 ( .A1(n14143), .A2(n14130), .ZN(n14131) );
  OAI211_X1 U17375 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n14139), .A(
        n14131), .B(n14208), .ZN(n14132) );
  MUX2_X1 U17376 ( .A(n14134), .B(n14208), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14137) );
  INV_X1 U17377 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14750) );
  NAND2_X1 U17378 ( .A1(n14135), .A2(n14750), .ZN(n14136) );
  AND2_X1 U17379 ( .A1(n14137), .A2(n14136), .ZN(n14243) );
  OR2_X1 U17380 ( .A1(n14146), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14141) );
  INV_X1 U17381 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14384) );
  NAND2_X1 U17382 ( .A1(n14143), .A2(n14384), .ZN(n14138) );
  OAI211_X1 U17383 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14139), .A(
        n14138), .B(n14208), .ZN(n14140) );
  NAND2_X1 U17384 ( .A1(n14141), .A2(n14140), .ZN(n14233) );
  INV_X1 U17385 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U17386 ( .A1(n14143), .A2(n14142), .ZN(n14144) );
  OAI21_X1 U17387 ( .B1(n14145), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14144), .ZN(n14207) );
  OR2_X1 U17388 ( .A1(n14207), .A2(n14149), .ZN(n14148) );
  OR2_X1 U17389 ( .A1(n14146), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14147) );
  AND2_X1 U17390 ( .A1(n14148), .A2(n14147), .ZN(n14223) );
  NOR2_X2 U17391 ( .A1(n14235), .A2(n14223), .ZN(n14222) );
  MUX2_X1 U17392 ( .A(n14149), .B(n14209), .S(n14222), .Z(n14150) );
  NAND2_X1 U17393 ( .A1(n20398), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14169) );
  AND2_X1 U17394 ( .A1(n21119), .A2(n20894), .ZN(n14160) );
  NOR2_X1 U17395 ( .A1(n14169), .A2(n14160), .ZN(n14153) );
  NAND2_X1 U17396 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21123), .ZN(n16057) );
  NAND2_X1 U17397 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21027), .ZN(n14155) );
  OAI21_X1 U17398 ( .B1(n14155), .B2(n14154), .A(n20243), .ZN(n14156) );
  INV_X1 U17399 ( .A(n14156), .ZN(n14157) );
  OAI21_X1 U17400 ( .B1(n16057), .B2(n21027), .A(n14157), .ZN(n14158) );
  NOR2_X1 U17401 ( .A1(n14214), .A2(n21324), .ZN(n14159) );
  NAND2_X1 U17402 ( .A1(n14196), .A2(n20210), .ZN(n14185) );
  AND2_X1 U17403 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14180) );
  OR2_X1 U17404 ( .A1(n20398), .A2(n16045), .ZN(n14161) );
  AND2_X1 U17405 ( .A1(n14161), .A2(n14160), .ZN(n14171) );
  NAND2_X1 U17406 ( .A1(n20273), .A2(n14363), .ZN(n20224) );
  INV_X1 U17407 ( .A(n20224), .ZN(n16125) );
  INV_X1 U17408 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n16097) );
  INV_X1 U17409 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14163) );
  INV_X1 U17410 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21064) );
  INV_X1 U17411 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14162) );
  INV_X1 U17412 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20196) );
  INV_X1 U17413 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21242) );
  INV_X1 U17414 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20234) );
  NAND4_X1 U17415 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20235)
         );
  NOR2_X1 U17416 ( .A1(n20234), .A2(n20235), .ZN(n20214) );
  NAND2_X1 U17417 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20214), .ZN(n20205) );
  NOR2_X1 U17418 ( .A1(n21242), .A2(n20205), .ZN(n14348) );
  NAND2_X1 U17419 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14348), .ZN(n20197) );
  NOR3_X1 U17420 ( .A1(n14162), .A2(n20196), .A3(n20197), .ZN(n16171) );
  NAND3_X1 U17421 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n16171), .ZN(n14327) );
  NOR3_X1 U17422 ( .A1(n14163), .A2(n21064), .A3(n14327), .ZN(n14312) );
  INV_X1 U17423 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21077) );
  NAND3_X1 U17424 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U17425 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16109) );
  NOR3_X1 U17426 ( .A1(n21077), .A2(n16123), .A3(n16109), .ZN(n16084) );
  NAND2_X1 U17427 ( .A1(n14312), .A2(n16084), .ZN(n16096) );
  NOR2_X1 U17428 ( .A1(n16097), .A2(n16096), .ZN(n14301) );
  AND2_X1 U17429 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14164) );
  AND2_X1 U17430 ( .A1(n14301), .A2(n14164), .ZN(n14286) );
  OR2_X1 U17431 ( .A1(n20273), .A2(n14286), .ZN(n14165) );
  NAND2_X1 U17432 ( .A1(n14165), .A2(n14363), .ZN(n14303) );
  NOR2_X1 U17433 ( .A1(n20273), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14166) );
  NOR2_X1 U17434 ( .A1(n14303), .A2(n14166), .ZN(n14278) );
  AND2_X1 U17435 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14176) );
  OR2_X1 U17436 ( .A1(n20273), .A2(n14176), .ZN(n14167) );
  AND2_X1 U17437 ( .A1(n14278), .A2(n14167), .ZN(n14266) );
  NAND2_X1 U17438 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14178) );
  NAND2_X1 U17439 ( .A1(n20224), .A2(n14178), .ZN(n14168) );
  AND2_X1 U17440 ( .A1(n14266), .A2(n14168), .ZN(n14240) );
  OAI21_X1 U17441 ( .B1(n14180), .B2(n16125), .A(n14240), .ZN(n14212) );
  INV_X1 U17442 ( .A(n14169), .ZN(n14170) );
  NOR2_X1 U17443 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  INV_X1 U17444 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14378) );
  AND2_X2 U17445 ( .A1(n14363), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20271) );
  OAI22_X1 U17446 ( .A1(n20276), .A2(n14378), .B1(n14174), .B2(n20240), .ZN(
        n14183) );
  NAND2_X1 U17447 ( .A1(n14286), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14175) );
  OR2_X1 U17448 ( .A1(n20273), .A2(n14175), .ZN(n14262) );
  INV_X1 U17449 ( .A(n14176), .ZN(n14177) );
  NOR2_X1 U17450 ( .A1(n14262), .A2(n14177), .ZN(n14248) );
  INV_X1 U17451 ( .A(n14178), .ZN(n14179) );
  NAND2_X1 U17452 ( .A1(n14248), .A2(n14179), .ZN(n14225) );
  INV_X1 U17453 ( .A(n14180), .ZN(n14181) );
  NOR3_X1 U17454 ( .A1(n14225), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14181), 
        .ZN(n14182) );
  AOI211_X1 U17455 ( .C1(n14212), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14183), 
        .B(n14182), .ZN(n14184) );
  OAI211_X1 U17456 ( .C1(n14689), .C2(n20279), .A(n14185), .B(n14184), .ZN(
        P1_U2809) );
  INV_X1 U17457 ( .A(n20375), .ZN(n14190) );
  AOI211_X1 U17458 ( .C1(n14188), .C2(n20894), .A(n20493), .B(n14187), .ZN(
        n14189) );
  AOI21_X1 U17459 ( .B1(n14190), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n14189), .ZN(n14191) );
  OAI21_X1 U17460 ( .B1(n14186), .B2(n14192), .A(n14191), .ZN(P1_U3477) );
  INV_X1 U17461 ( .A(DATAI_31_), .ZN(n14201) );
  AND2_X1 U17462 ( .A1(n14546), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U17463 ( .A1(n14196), .A2(n14195), .ZN(n14200) );
  AND2_X1 U17464 ( .A1(n14197), .A2(n20377), .ZN(n14198) );
  NAND2_X1 U17465 ( .A1(n14546), .A2(n14198), .ZN(n16196) );
  AOI22_X1 U17466 ( .A1(n14537), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16190), .ZN(n14199) );
  OAI211_X1 U17467 ( .C1(n14540), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        P1_U2873) );
  NOR2_X1 U17468 ( .A1(n15350), .A2(n19385), .ZN(n14202) );
  AOI21_X1 U17469 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19385), .A(n14202), .ZN(
        n14203) );
  OAI21_X1 U17470 ( .B1(n14204), .B2(n19380), .A(n14203), .ZN(P2_U2857) );
  XNOR2_X2 U17471 ( .A(n14205), .B(n14206), .ZN(n14567) );
  OAI22_X1 U17472 ( .A1(n14222), .A2(n14208), .B1(n14207), .B2(n14235), .ZN(
        n14211) );
  INV_X1 U17473 ( .A(n14209), .ZN(n14210) );
  XNOR2_X1 U17474 ( .A(n14211), .B(n14210), .ZN(n14718) );
  INV_X1 U17475 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14380) );
  INV_X1 U17476 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14570) );
  NOR2_X1 U17477 ( .A1(n14225), .A2(n14570), .ZN(n14213) );
  OAI21_X1 U17478 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14213), .A(n14212), 
        .ZN(n14217) );
  AOI22_X1 U17479 ( .A1(n14564), .A2(n20257), .B1(n20271), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14216) );
  OAI211_X1 U17480 ( .C1(n20276), .C2(n14380), .A(n14217), .B(n14216), .ZN(
        n14218) );
  AOI21_X1 U17481 ( .B1(n14718), .B2(n20260), .A(n14218), .ZN(n14219) );
  OAI21_X1 U17482 ( .B1(n14567), .B2(n20218), .A(n14219), .ZN(P1_U2810) );
  INV_X1 U17483 ( .A(n14574), .ZN(n14382) );
  AOI21_X1 U17484 ( .B1(n14223), .B2(n14235), .A(n14222), .ZN(n14728) );
  OAI22_X1 U17485 ( .A1(n14224), .A2(n20240), .B1(n20285), .B2(n14572), .ZN(
        n14227) );
  NOR2_X1 U17486 ( .A1(n14225), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14226) );
  AOI211_X1 U17487 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n20261), .A(n14227), .B(
        n14226), .ZN(n14228) );
  OAI21_X1 U17488 ( .B1(n14240), .B2(n14570), .A(n14228), .ZN(n14229) );
  AOI21_X1 U17489 ( .B1(n14728), .B2(n20260), .A(n14229), .ZN(n14230) );
  OAI21_X1 U17490 ( .B1(n14382), .B2(n20218), .A(n14230), .ZN(P1_U2811) );
  OAI21_X1 U17491 ( .B1(n14231), .B2(n14232), .A(n14220), .ZN(n14589) );
  OR2_X1 U17492 ( .A1(n14245), .A2(n14233), .ZN(n14234) );
  AOI21_X1 U17493 ( .B1(n14248), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17494 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20271), .B1(
        n20257), .B2(n14579), .ZN(n14236) );
  OAI21_X1 U17495 ( .B1(n20276), .B2(n14384), .A(n14236), .ZN(n14237) );
  INV_X1 U17496 ( .A(n14237), .ZN(n14238) );
  OAI21_X1 U17497 ( .B1(n14240), .B2(n14239), .A(n14238), .ZN(n14241) );
  AOI21_X1 U17498 ( .B1(n14737), .B2(n20260), .A(n14241), .ZN(n14242) );
  OAI21_X1 U17499 ( .B1(n14589), .B2(n20218), .A(n14242), .ZN(P1_U2812) );
  NOR2_X1 U17500 ( .A1(n14261), .A2(n14243), .ZN(n14244) );
  OR2_X1 U17501 ( .A1(n14245), .A2(n14244), .ZN(n14748) );
  AOI21_X1 U17502 ( .B1(n14247), .B2(n14246), .A(n14231), .ZN(n14596) );
  NAND2_X1 U17503 ( .A1(n14596), .A2(n20210), .ZN(n14256) );
  INV_X1 U17504 ( .A(n14266), .ZN(n14254) );
  INV_X1 U17505 ( .A(n14248), .ZN(n14252) );
  OAI22_X1 U17506 ( .A1(n14249), .A2(n20240), .B1(n20285), .B2(n14594), .ZN(
        n14250) );
  AOI21_X1 U17507 ( .B1(n20261), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14250), .ZN(
        n14251) );
  OAI21_X1 U17508 ( .B1(n14252), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14251), 
        .ZN(n14253) );
  AOI21_X1 U17509 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14254), .A(n14253), 
        .ZN(n14255) );
  OAI211_X1 U17510 ( .C1(n20279), .C2(n14748), .A(n14256), .B(n14255), .ZN(
        P1_U2813) );
  AND2_X1 U17511 ( .A1(n9925), .A2(n14259), .ZN(n14260) );
  NOR2_X1 U17512 ( .A1(n14261), .A2(n14260), .ZN(n14760) );
  INV_X1 U17513 ( .A(n14262), .ZN(n14276) );
  AOI21_X1 U17514 ( .B1(n14276), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14265) );
  AOI22_X1 U17515 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20271), .B1(
        n20257), .B2(n14606), .ZN(n14264) );
  NAND2_X1 U17516 ( .A1(n20261), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14263) );
  OAI211_X1 U17517 ( .C1(n14266), .C2(n14265), .A(n14264), .B(n14263), .ZN(
        n14267) );
  AOI21_X1 U17518 ( .B1(n14760), .B2(n20260), .A(n14267), .ZN(n14268) );
  OAI21_X1 U17519 ( .B1(n14603), .B2(n20218), .A(n14268), .ZN(P1_U2814) );
  AOI21_X1 U17520 ( .B1(n14270), .B2(n10358), .A(n14257), .ZN(n14615) );
  INV_X1 U17521 ( .A(n14615), .ZN(n14388) );
  NAND2_X1 U17522 ( .A1(n9922), .A2(n14271), .ZN(n14272) );
  NAND2_X1 U17523 ( .A1(n9925), .A2(n14272), .ZN(n14390) );
  INV_X1 U17524 ( .A(n14390), .ZN(n16274) );
  INV_X1 U17525 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21360) );
  INV_X1 U17526 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14389) );
  INV_X1 U17527 ( .A(n14613), .ZN(n14273) );
  AOI22_X1 U17528 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20271), .B1(
        n20257), .B2(n14273), .ZN(n14274) );
  OAI21_X1 U17529 ( .B1(n20276), .B2(n14389), .A(n14274), .ZN(n14275) );
  AOI21_X1 U17530 ( .B1(n14276), .B2(n21360), .A(n14275), .ZN(n14277) );
  OAI21_X1 U17531 ( .B1(n14278), .B2(n21360), .A(n14277), .ZN(n14279) );
  AOI21_X1 U17532 ( .B1(n16274), .B2(n20260), .A(n14279), .ZN(n14280) );
  OAI21_X1 U17533 ( .B1(n14388), .B2(n20218), .A(n14280), .ZN(P1_U2815) );
  OR2_X1 U17534 ( .A1(n14297), .A2(n14281), .ZN(n14282) );
  NAND2_X1 U17535 ( .A1(n9922), .A2(n14282), .ZN(n14764) );
  AOI21_X1 U17536 ( .B1(n14284), .B2(n14283), .A(n14269), .ZN(n14624) );
  NAND2_X1 U17537 ( .A1(n14624), .A2(n20210), .ZN(n14292) );
  INV_X1 U17538 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U17539 ( .A1(n14286), .A2(n14285), .ZN(n14289) );
  OR2_X1 U17540 ( .A1(n20276), .A2(n14391), .ZN(n14288) );
  AOI22_X1 U17541 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20271), .B1(
        n20257), .B2(n14620), .ZN(n14287) );
  OAI211_X1 U17542 ( .C1(n20273), .C2(n14289), .A(n14288), .B(n14287), .ZN(
        n14290) );
  AOI21_X1 U17543 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14303), .A(n14290), 
        .ZN(n14291) );
  OAI211_X1 U17544 ( .C1(n20279), .C2(n14764), .A(n14292), .B(n14291), .ZN(
        P1_U2816) );
  OAI21_X1 U17545 ( .B1(n14293), .B2(n14294), .A(n14283), .ZN(n16197) );
  AND2_X1 U17546 ( .A1(n14399), .A2(n14295), .ZN(n14296) );
  NOR2_X1 U17547 ( .A1(n14297), .A2(n14296), .ZN(n16280) );
  INV_X1 U17548 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14394) );
  INV_X1 U17549 ( .A(n16203), .ZN(n14298) );
  AOI22_X1 U17550 ( .A1(n14298), .A2(n20257), .B1(n20271), .B2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14299) );
  OAI21_X1 U17551 ( .B1(n20276), .B2(n14394), .A(n14299), .ZN(n14300) );
  AOI21_X1 U17552 ( .B1(n16280), .B2(n20260), .A(n14300), .ZN(n14306) );
  INV_X1 U17553 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n16295) );
  NAND2_X1 U17554 ( .A1(n20236), .A2(n14301), .ZN(n16090) );
  INV_X1 U17555 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14302) );
  OAI21_X1 U17556 ( .B1(n16295), .B2(n16090), .A(n14302), .ZN(n14304) );
  NAND2_X1 U17557 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  OAI211_X1 U17558 ( .C1(n16197), .C2(n20218), .A(n14306), .B(n14305), .ZN(
        P1_U2817) );
  OR2_X1 U17559 ( .A1(n14432), .A2(n14309), .ZN(n14421) );
  INV_X1 U17560 ( .A(n14421), .ZN(n14308) );
  AOI21_X1 U17561 ( .B1(n14309), .B2(n14432), .A(n14308), .ZN(n14651) );
  INV_X1 U17562 ( .A(n14651), .ZN(n14319) );
  INV_X1 U17563 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21070) );
  INV_X1 U17564 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n16315) );
  NOR3_X1 U17565 ( .A1(n20273), .A2(n21064), .A3(n14327), .ZN(n16158) );
  NAND2_X1 U17566 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16158), .ZN(n16157) );
  AOI21_X1 U17567 ( .B1(n21070), .B2(n16315), .A(n16157), .ZN(n14317) );
  NAND2_X1 U17568 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16108) );
  NOR2_X1 U17569 ( .A1(n20285), .A2(n14649), .ZN(n14316) );
  OR2_X1 U17570 ( .A1(n14436), .A2(n14310), .ZN(n14311) );
  NAND2_X1 U17571 ( .A1(n14424), .A2(n14311), .ZN(n16309) );
  NAND2_X1 U17572 ( .A1(n14312), .A2(n14363), .ZN(n16083) );
  NAND2_X1 U17573 ( .A1(n20224), .A2(n16083), .ZN(n16168) );
  OAI22_X1 U17574 ( .A1(n20279), .A2(n16309), .B1(n21070), .B2(n16168), .ZN(
        n14313) );
  AOI211_X1 U17575 ( .C1(n20271), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14313), .B(n16368), .ZN(n14314) );
  OAI21_X1 U17576 ( .B1(n14428), .B2(n20276), .A(n14314), .ZN(n14315) );
  AOI211_X1 U17577 ( .C1(n14317), .C2(n16108), .A(n14316), .B(n14315), .ZN(
        n14318) );
  OAI21_X1 U17578 ( .B1(n14319), .B2(n20218), .A(n14318), .ZN(P1_U2824) );
  OAI21_X1 U17579 ( .B1(n14320), .B2(n14321), .A(n14322), .ZN(n14454) );
  OAI21_X1 U17580 ( .B1(n14454), .B2(n10367), .A(n14322), .ZN(n14445) );
  INV_X1 U17581 ( .A(n14323), .ZN(n14324) );
  INV_X1 U17582 ( .A(n14363), .ZN(n20270) );
  AOI21_X1 U17583 ( .B1(n14327), .B2(n20236), .A(n20270), .ZN(n14326) );
  INV_X1 U17584 ( .A(n14326), .ZN(n16174) );
  NOR2_X1 U17585 ( .A1(n20273), .A2(n14327), .ZN(n14334) );
  INV_X1 U17586 ( .A(n14450), .ZN(n14328) );
  NAND2_X1 U17587 ( .A1(n14456), .A2(n14328), .ZN(n14329) );
  AOI21_X1 U17588 ( .B1(n14330), .B2(n14329), .A(n10206), .ZN(n16325) );
  AOI21_X1 U17589 ( .B1(n16325), .B2(n20260), .A(n16368), .ZN(n14331) );
  OAI21_X1 U17590 ( .B1(n14332), .B2(n20240), .A(n14331), .ZN(n14333) );
  AOI221_X1 U17591 ( .B1(n16174), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n14334), 
        .C2(n21064), .A(n14333), .ZN(n14336) );
  AOI22_X1 U17592 ( .A1(n20261), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n20257), 
        .B2(n14670), .ZN(n14335) );
  OAI211_X1 U17593 ( .C1(n14673), .C2(n20218), .A(n14336), .B(n14335), .ZN(
        P1_U2827) );
  AOI21_X1 U17594 ( .B1(n14337), .B2(n13935), .A(n14320), .ZN(n14681) );
  INV_X1 U17595 ( .A(n14681), .ZN(n14557) );
  OAI21_X1 U17596 ( .B1(n16171), .B2(n20273), .A(n14363), .ZN(n16182) );
  NOR2_X1 U17597 ( .A1(n16171), .A2(n20273), .ZN(n14338) );
  AOI211_X1 U17598 ( .C1(n20236), .C2(n20197), .A(n20270), .B(n20196), .ZN(
        n20195) );
  AOI22_X1 U17599 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n16182), .B1(n14338), 
        .B2(n20195), .ZN(n14345) );
  AND2_X1 U17600 ( .A1(n16355), .A2(n14339), .ZN(n14340) );
  OR2_X1 U17601 ( .A1(n14340), .A2(n14455), .ZN(n16346) );
  INV_X1 U17602 ( .A(n14679), .ZN(n14341) );
  AOI22_X1 U17603 ( .A1(n14341), .A2(n20257), .B1(n20261), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14342) );
  OAI21_X1 U17604 ( .B1(n20279), .B2(n16346), .A(n14342), .ZN(n14343) );
  AOI211_X1 U17605 ( .C1(n20271), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n14343), .B(n16368), .ZN(n14344) );
  OAI211_X1 U17606 ( .C1(n14557), .C2(n20218), .A(n14345), .B(n14344), .ZN(
        P1_U2830) );
  NAND2_X1 U17607 ( .A1(n20236), .A2(n20197), .ZN(n14346) );
  NAND2_X1 U17608 ( .A1(n14363), .A2(n14346), .ZN(n14351) );
  INV_X1 U17609 ( .A(n14346), .ZN(n14347) );
  AOI22_X1 U17610 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20271), .B1(
        n14348), .B2(n14347), .ZN(n14349) );
  OAI211_X1 U17611 ( .C1(n20279), .C2(n16370), .A(n14349), .B(n20243), .ZN(
        n14350) );
  AOI21_X1 U17612 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n14351), .A(n14350), .ZN(
        n14355) );
  INV_X1 U17613 ( .A(n14352), .ZN(n14353) );
  AOI22_X1 U17614 ( .A1(n20261), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n14353), .B2(
        n20257), .ZN(n14354) );
  OAI211_X1 U17615 ( .C1(n14356), .C2(n20218), .A(n14355), .B(n14354), .ZN(
        P1_U2832) );
  NAND2_X1 U17616 ( .A1(n20218), .A2(n14357), .ZN(n20281) );
  INV_X1 U17617 ( .A(n20281), .ZN(n20247) );
  INV_X1 U17618 ( .A(n20831), .ZN(n20387) );
  NOR2_X1 U17619 ( .A1(n14359), .A2(n14358), .ZN(n20275) );
  NOR2_X1 U17620 ( .A1(n20273), .A2(n21107), .ZN(n20265) );
  AOI22_X1 U17621 ( .A1(n20271), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21054), .B2(n20265), .ZN(n14360) );
  OAI21_X1 U17622 ( .B1(n20285), .B2(n14361), .A(n14360), .ZN(n14362) );
  AOI21_X1 U17623 ( .B1(n20261), .B2(P1_EBX_REG_2__SCAN_IN), .A(n14362), .ZN(
        n14366) );
  OR2_X1 U17624 ( .A1(n20273), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14364) );
  NAND2_X1 U17625 ( .A1(n14364), .A2(n14363), .ZN(n20262) );
  NAND2_X1 U17626 ( .A1(n20262), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n14365) );
  OAI211_X1 U17627 ( .C1(n14367), .C2(n20279), .A(n14366), .B(n14365), .ZN(
        n14368) );
  AOI21_X1 U17628 ( .B1(n20387), .B2(n20275), .A(n14368), .ZN(n14369) );
  OAI21_X1 U17629 ( .B1(n14370), .B2(n20247), .A(n14369), .ZN(P1_U2838) );
  NAND2_X1 U17630 ( .A1(n20260), .A2(n14371), .ZN(n14373) );
  OAI21_X1 U17631 ( .B1(n20271), .B2(n20257), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14372) );
  OAI211_X1 U17632 ( .C1(n20276), .C2(n13334), .A(n14373), .B(n14372), .ZN(
        n14376) );
  INV_X1 U17633 ( .A(n20275), .ZN(n20241) );
  NOR2_X1 U17634 ( .A1(n14374), .A2(n20241), .ZN(n14375) );
  AOI211_X1 U17635 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20224), .A(n14376), .B(
        n14375), .ZN(n14377) );
  OAI21_X1 U17636 ( .B1(n20374), .B2(n20247), .A(n14377), .ZN(P1_U2840) );
  OAI22_X1 U17637 ( .A1(n14689), .A2(n20288), .B1(n20302), .B2(n14378), .ZN(
        P1_U2841) );
  INV_X1 U17638 ( .A(n14718), .ZN(n14379) );
  OAI222_X1 U17639 ( .A1(n14452), .A2(n14567), .B1(n14380), .B2(n20302), .C1(
        n14379), .C2(n20288), .ZN(P1_U2842) );
  AOI22_X1 U17640 ( .A1(n14728), .A2(n20298), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14458), .ZN(n14381) );
  OAI21_X1 U17641 ( .B1(n14382), .B2(n14452), .A(n14381), .ZN(P1_U2843) );
  INV_X1 U17642 ( .A(n14737), .ZN(n14383) );
  OAI222_X1 U17643 ( .A1(n14452), .A2(n14589), .B1(n14384), .B2(n20302), .C1(
        n14383), .C2(n20288), .ZN(P1_U2844) );
  INV_X1 U17644 ( .A(n14596), .ZN(n14386) );
  INV_X1 U17645 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14385) );
  OAI222_X1 U17646 ( .A1(n14452), .A2(n14386), .B1(n14385), .B2(n20302), .C1(
        n14748), .C2(n20288), .ZN(P1_U2845) );
  AOI22_X1 U17647 ( .A1(n14760), .A2(n20298), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14458), .ZN(n14387) );
  OAI21_X1 U17648 ( .B1(n14603), .B2(n14452), .A(n14387), .ZN(P1_U2846) );
  OAI222_X1 U17649 ( .A1(n14390), .A2(n20288), .B1(n14389), .B2(n20302), .C1(
        n14388), .C2(n14452), .ZN(P1_U2847) );
  INV_X1 U17650 ( .A(n14624), .ZN(n14392) );
  OAI222_X1 U17651 ( .A1(n14452), .A2(n14392), .B1(n14391), .B2(n20302), .C1(
        n14764), .C2(n20288), .ZN(P1_U2848) );
  INV_X1 U17652 ( .A(n16280), .ZN(n14393) );
  OAI222_X1 U17653 ( .A1(n14452), .A2(n16197), .B1(n14394), .B2(n20302), .C1(
        n14393), .C2(n20288), .ZN(P1_U2849) );
  AOI21_X1 U17654 ( .B1(n14396), .B2(n14395), .A(n14293), .ZN(n14631) );
  INV_X1 U17655 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U17656 ( .A1(n9879), .A2(n14397), .ZN(n14398) );
  NAND2_X1 U17657 ( .A1(n14399), .A2(n14398), .ZN(n16287) );
  OAI222_X1 U17658 ( .A1(n16091), .A2(n14452), .B1(n20302), .B2(n14400), .C1(
        n16287), .C2(n20288), .ZN(P1_U2850) );
  OAI21_X1 U17659 ( .B1(n14406), .B2(n14401), .A(n16102), .ZN(n16111) );
  INV_X1 U17660 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14403) );
  OAI21_X1 U17661 ( .B1(n14409), .B2(n14402), .A(n9926), .ZN(n16110) );
  OAI222_X1 U17662 ( .A1(n16111), .A2(n14452), .B1(n20302), .B2(n14403), .C1(
        n16110), .C2(n20288), .ZN(P1_U2852) );
  NOR2_X1 U17663 ( .A1(n14412), .A2(n14404), .ZN(n14405) );
  OR2_X1 U17664 ( .A1(n14406), .A2(n14405), .ZN(n16120) );
  INV_X1 U17665 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14410) );
  NOR2_X1 U17666 ( .A1(n14415), .A2(n14407), .ZN(n14408) );
  OR2_X1 U17667 ( .A1(n14409), .A2(n14408), .ZN(n16297) );
  OAI222_X1 U17668 ( .A1(n14452), .A2(n16120), .B1(n14410), .B2(n20302), .C1(
        n16297), .C2(n20288), .ZN(P1_U2853) );
  AND2_X1 U17669 ( .A1(n14419), .A2(n14411), .ZN(n14413) );
  OR2_X1 U17670 ( .A1(n14413), .A2(n14412), .ZN(n16140) );
  AND2_X1 U17671 ( .A1(n14426), .A2(n14414), .ZN(n14416) );
  OR2_X1 U17672 ( .A1(n14416), .A2(n14415), .ZN(n16143) );
  OAI22_X1 U17673 ( .A1(n16143), .A2(n20288), .B1(n16131), .B2(n20302), .ZN(
        n14417) );
  INV_X1 U17674 ( .A(n14417), .ZN(n14418) );
  OAI21_X1 U17675 ( .B1(n16140), .B2(n14452), .A(n14418), .ZN(P1_U2854) );
  INV_X1 U17676 ( .A(n14419), .ZN(n14420) );
  AOI21_X1 U17677 ( .B1(n14422), .B2(n14421), .A(n14420), .ZN(n16221) );
  INV_X1 U17678 ( .A(n16221), .ZN(n14536) );
  NAND2_X1 U17679 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  NAND2_X1 U17680 ( .A1(n14426), .A2(n14425), .ZN(n16144) );
  OAI222_X1 U17681 ( .A1(n14536), .A2(n14452), .B1(n14427), .B2(n20302), .C1(
        n16144), .C2(n20288), .ZN(P1_U2855) );
  OAI22_X1 U17682 ( .A1(n16309), .A2(n20288), .B1(n14428), .B2(n20302), .ZN(
        n14429) );
  AOI21_X1 U17683 ( .B1(n14651), .B2(n20299), .A(n14429), .ZN(n14430) );
  INV_X1 U17684 ( .A(n14430), .ZN(P1_U2856) );
  OAI21_X1 U17685 ( .B1(n14431), .B2(n14433), .A(n14432), .ZN(n16234) );
  AND2_X1 U17686 ( .A1(n14440), .A2(n14434), .ZN(n14435) );
  NOR2_X1 U17687 ( .A1(n14436), .A2(n14435), .ZN(n16317) );
  AOI22_X1 U17688 ( .A1(n16317), .A2(n20298), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14458), .ZN(n14437) );
  OAI21_X1 U17689 ( .B1(n16234), .B2(n14452), .A(n14437), .ZN(P1_U2857) );
  NOR2_X1 U17690 ( .A1(n14323), .A2(n14438), .ZN(n14439) );
  OR2_X1 U17691 ( .A1(n14431), .A2(n14439), .ZN(n16162) );
  AOI21_X1 U17692 ( .B1(n14442), .B2(n14441), .A(n10202), .ZN(n16165) );
  AOI22_X1 U17693 ( .A1(n16165), .A2(n20298), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14458), .ZN(n14443) );
  OAI21_X1 U17694 ( .B1(n16162), .B2(n14452), .A(n14443), .ZN(P1_U2858) );
  AOI22_X1 U17695 ( .A1(n16325), .A2(n20298), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14458), .ZN(n14444) );
  OAI21_X1 U17696 ( .B1(n14673), .B2(n14452), .A(n14444), .ZN(P1_U2859) );
  INV_X1 U17697 ( .A(n14445), .ZN(n14449) );
  INV_X1 U17698 ( .A(n14446), .ZN(n14448) );
  INV_X1 U17699 ( .A(n16240), .ZN(n14551) );
  XNOR2_X1 U17700 ( .A(n14456), .B(n14450), .ZN(n16170) );
  AOI22_X1 U17701 ( .A1(n16170), .A2(n20298), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14458), .ZN(n14451) );
  OAI21_X1 U17702 ( .B1(n14551), .B2(n14452), .A(n14451), .ZN(P1_U2860) );
  XNOR2_X1 U17703 ( .A(n14454), .B(n14453), .ZN(n16250) );
  INV_X1 U17704 ( .A(n16250), .ZN(n14554) );
  INV_X1 U17705 ( .A(n14455), .ZN(n14457) );
  AOI21_X1 U17706 ( .B1(n9950), .B2(n14457), .A(n14456), .ZN(n16332) );
  AOI22_X1 U17707 ( .A1(n16332), .A2(n20298), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14458), .ZN(n14459) );
  OAI21_X1 U17708 ( .B1(n14554), .B2(n14452), .A(n14459), .ZN(P1_U2861) );
  OAI22_X1 U17709 ( .A1(n16346), .A2(n20288), .B1(n14460), .B2(n20302), .ZN(
        n14461) );
  AOI21_X1 U17710 ( .B1(n14681), .B2(n20299), .A(n14461), .ZN(n14462) );
  INV_X1 U17711 ( .A(n14462), .ZN(P1_U2862) );
  INV_X1 U17712 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14463) );
  NOR2_X1 U17713 ( .A1(n20379), .A2(n14463), .ZN(n14464) );
  AOI21_X1 U17714 ( .B1(DATAI_14_), .B2(n20379), .A(n14464), .ZN(n20346) );
  OAI22_X1 U17715 ( .A1(n14465), .A2(n20346), .B1(n14546), .B2(n13165), .ZN(
        n14466) );
  AOI21_X1 U17716 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14537), .A(n14466), .ZN(
        n14468) );
  NAND2_X1 U17717 ( .A1(n16192), .A2(DATAI_30_), .ZN(n14467) );
  OAI211_X1 U17718 ( .C1(n14567), .C2(n14553), .A(n14468), .B(n14467), .ZN(
        P1_U2874) );
  OR2_X1 U17719 ( .A1(n20379), .A2(n16754), .ZN(n14470) );
  NAND2_X1 U17720 ( .A1(n20379), .A2(DATAI_13_), .ZN(n14469) );
  NAND2_X1 U17721 ( .A1(n14470), .A2(n14469), .ZN(n20344) );
  AOI22_X1 U17722 ( .A1(n16191), .A2(n20344), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16190), .ZN(n14472) );
  NAND2_X1 U17723 ( .A1(n14537), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14471) );
  OAI211_X1 U17724 ( .C1(n21291), .C2(n14540), .A(n14472), .B(n14471), .ZN(
        n14473) );
  AOI21_X1 U17725 ( .B1(n14574), .B2(n16193), .A(n14473), .ZN(n14474) );
  INV_X1 U17726 ( .A(n14474), .ZN(P1_U2875) );
  INV_X1 U17727 ( .A(DATAI_28_), .ZN(n14479) );
  OR2_X1 U17728 ( .A1(n20379), .A2(n16756), .ZN(n14476) );
  NAND2_X1 U17729 ( .A1(n20379), .A2(DATAI_12_), .ZN(n14475) );
  NAND2_X1 U17730 ( .A1(n14476), .A2(n14475), .ZN(n20342) );
  AOI22_X1 U17731 ( .A1(n16191), .A2(n20342), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16190), .ZN(n14478) );
  NAND2_X1 U17732 ( .A1(n14537), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14477) );
  OAI211_X1 U17733 ( .C1(n14479), .C2(n14540), .A(n14478), .B(n14477), .ZN(
        n14480) );
  INV_X1 U17734 ( .A(n14480), .ZN(n14481) );
  OAI21_X1 U17735 ( .B1(n14589), .B2(n14553), .A(n14481), .ZN(P1_U2876) );
  INV_X1 U17736 ( .A(DATAI_27_), .ZN(n14487) );
  INV_X1 U17737 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14482) );
  OR2_X1 U17738 ( .A1(n20379), .A2(n14482), .ZN(n14484) );
  NAND2_X1 U17739 ( .A1(n20379), .A2(DATAI_11_), .ZN(n14483) );
  NAND2_X1 U17740 ( .A1(n14484), .A2(n14483), .ZN(n20340) );
  AOI22_X1 U17741 ( .A1(n16191), .A2(n20340), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16190), .ZN(n14486) );
  NAND2_X1 U17742 ( .A1(n14537), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14485) );
  OAI211_X1 U17743 ( .C1(n14487), .C2(n14540), .A(n14486), .B(n14485), .ZN(
        n14488) );
  AOI21_X1 U17744 ( .B1(n14596), .B2(n16193), .A(n14488), .ZN(n14489) );
  INV_X1 U17745 ( .A(n14489), .ZN(P1_U2877) );
  INV_X1 U17746 ( .A(DATAI_26_), .ZN(n14494) );
  INV_X1 U17747 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16759) );
  OR2_X1 U17748 ( .A1(n20379), .A2(n16759), .ZN(n14491) );
  NAND2_X1 U17749 ( .A1(n20379), .A2(DATAI_10_), .ZN(n14490) );
  NAND2_X1 U17750 ( .A1(n14491), .A2(n14490), .ZN(n20338) );
  AOI22_X1 U17751 ( .A1(n16191), .A2(n20338), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16190), .ZN(n14493) );
  NAND2_X1 U17752 ( .A1(n14537), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14492) );
  OAI211_X1 U17753 ( .C1(n14494), .C2(n14540), .A(n14493), .B(n14492), .ZN(
        n14495) );
  INV_X1 U17754 ( .A(n14495), .ZN(n14496) );
  OAI21_X1 U17755 ( .B1(n14603), .B2(n14553), .A(n14496), .ZN(P1_U2878) );
  INV_X1 U17756 ( .A(DATAI_25_), .ZN(n14500) );
  AOI22_X1 U17757 ( .A1(n16191), .A2(n14497), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16190), .ZN(n14499) );
  NAND2_X1 U17758 ( .A1(n14537), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14498) );
  OAI211_X1 U17759 ( .C1(n14500), .C2(n14540), .A(n14499), .B(n14498), .ZN(
        n14501) );
  AOI21_X1 U17760 ( .B1(n14615), .B2(n16193), .A(n14501), .ZN(n14502) );
  INV_X1 U17761 ( .A(n14502), .ZN(P1_U2879) );
  INV_X1 U17762 ( .A(DATAI_24_), .ZN(n14505) );
  AOI22_X1 U17763 ( .A1(n16191), .A2(n20336), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16190), .ZN(n14504) );
  NAND2_X1 U17764 ( .A1(n14537), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14503) );
  OAI211_X1 U17765 ( .C1(n14505), .C2(n14540), .A(n14504), .B(n14503), .ZN(
        n14506) );
  AOI21_X1 U17766 ( .B1(n14624), .B2(n16193), .A(n14506), .ZN(n14507) );
  INV_X1 U17767 ( .A(n14507), .ZN(P1_U2880) );
  INV_X1 U17768 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15067) );
  AOI22_X1 U17769 ( .A1(n16191), .A2(n20428), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16190), .ZN(n14508) );
  OAI21_X1 U17770 ( .B1(n16196), .B2(n15067), .A(n14508), .ZN(n14509) );
  AOI21_X1 U17771 ( .B1(n16192), .B2(DATAI_23_), .A(n14509), .ZN(n14510) );
  OAI21_X1 U17772 ( .B1(n16197), .B2(n14553), .A(n14510), .ZN(P1_U2881) );
  INV_X1 U17773 ( .A(DATAI_22_), .ZN(n14513) );
  AOI22_X1 U17774 ( .A1(n16191), .A2(n20419), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16190), .ZN(n14512) );
  NAND2_X1 U17775 ( .A1(n14537), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14511) );
  OAI211_X1 U17776 ( .C1(n14513), .C2(n14540), .A(n14512), .B(n14511), .ZN(
        n14514) );
  AOI21_X1 U17777 ( .B1(n14631), .B2(n16193), .A(n14514), .ZN(n14515) );
  INV_X1 U17778 ( .A(n14515), .ZN(P1_U2882) );
  INV_X1 U17779 ( .A(n16111), .ZN(n14520) );
  INV_X1 U17780 ( .A(DATAI_20_), .ZN(n14518) );
  AOI22_X1 U17781 ( .A1(n16191), .A2(n20413), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16190), .ZN(n14517) );
  NAND2_X1 U17782 ( .A1(n14537), .A2(BUF1_REG_20__SCAN_IN), .ZN(n14516) );
  OAI211_X1 U17783 ( .C1(n14518), .C2(n14540), .A(n14517), .B(n14516), .ZN(
        n14519) );
  AOI21_X1 U17784 ( .B1(n14520), .B2(n16193), .A(n14519), .ZN(n14521) );
  INV_X1 U17785 ( .A(n14521), .ZN(P1_U2884) );
  INV_X1 U17786 ( .A(n16120), .ZN(n16216) );
  INV_X1 U17787 ( .A(DATAI_19_), .ZN(n14524) );
  AOI22_X1 U17788 ( .A1(n16191), .A2(n20409), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16190), .ZN(n14523) );
  NAND2_X1 U17789 ( .A1(n14537), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14522) );
  OAI211_X1 U17790 ( .C1(n14524), .C2(n14540), .A(n14523), .B(n14522), .ZN(
        n14525) );
  AOI21_X1 U17791 ( .B1(n16216), .B2(n16193), .A(n14525), .ZN(n14526) );
  INV_X1 U17792 ( .A(n14526), .ZN(P1_U2885) );
  INV_X1 U17793 ( .A(n16140), .ZN(n14531) );
  INV_X1 U17794 ( .A(DATAI_18_), .ZN(n14529) );
  AOI22_X1 U17795 ( .A1(n16191), .A2(n20405), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16190), .ZN(n14528) );
  NAND2_X1 U17796 ( .A1(n14537), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14527) );
  OAI211_X1 U17797 ( .C1(n14529), .C2(n14540), .A(n14528), .B(n14527), .ZN(
        n14530) );
  AOI21_X1 U17798 ( .B1(n14531), .B2(n16193), .A(n14530), .ZN(n14532) );
  INV_X1 U17799 ( .A(n14532), .ZN(P1_U2886) );
  INV_X1 U17800 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U17801 ( .A1(n16191), .A2(n20399), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16190), .ZN(n14533) );
  OAI21_X1 U17802 ( .B1(n16196), .B2(n15100), .A(n14533), .ZN(n14534) );
  AOI21_X1 U17803 ( .B1(n16192), .B2(DATAI_17_), .A(n14534), .ZN(n14535) );
  OAI21_X1 U17804 ( .B1(n14536), .B2(n14553), .A(n14535), .ZN(P1_U2887) );
  INV_X1 U17805 ( .A(DATAI_16_), .ZN(n14541) );
  AOI22_X1 U17806 ( .A1(n16191), .A2(n20390), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16190), .ZN(n14539) );
  NAND2_X1 U17807 ( .A1(n14537), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14538) );
  OAI211_X1 U17808 ( .C1(n14541), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        n14542) );
  AOI21_X1 U17809 ( .B1(n14651), .B2(n16193), .A(n14542), .ZN(n14543) );
  INV_X1 U17810 ( .A(n14543), .ZN(P1_U2888) );
  OAI222_X1 U17811 ( .A1(n14553), .A2(n16234), .B1(n14548), .B2(n14545), .C1(
        n14546), .C2(n14544), .ZN(P1_U2889) );
  OAI222_X1 U17812 ( .A1(n16162), .A2(n14553), .B1(n20346), .B2(n14548), .C1(
        n14547), .C2(n14546), .ZN(P1_U2890) );
  AOI22_X1 U17813 ( .A1(n14555), .A2(n20344), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16190), .ZN(n14549) );
  OAI21_X1 U17814 ( .B1(n14673), .B2(n14553), .A(n14549), .ZN(P1_U2891) );
  AOI22_X1 U17815 ( .A1(n14555), .A2(n20342), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16190), .ZN(n14550) );
  OAI21_X1 U17816 ( .B1(n14551), .B2(n14553), .A(n14550), .ZN(P1_U2892) );
  AOI22_X1 U17817 ( .A1(n14555), .A2(n20340), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16190), .ZN(n14552) );
  OAI21_X1 U17818 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(P1_U2893) );
  AOI22_X1 U17819 ( .A1(n14555), .A2(n20338), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16190), .ZN(n14556) );
  OAI21_X1 U17820 ( .B1(n14557), .B2(n14553), .A(n14556), .ZN(P1_U2894) );
  INV_X1 U17821 ( .A(n14558), .ZN(n14738) );
  INV_X1 U17822 ( .A(n14559), .ZN(n14600) );
  NAND2_X1 U17823 ( .A1(n14711), .A2(n20369), .ZN(n14566) );
  INV_X1 U17824 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14561) );
  NOR2_X1 U17825 ( .A1(n20243), .A2(n14561), .ZN(n14717) );
  NOR2_X1 U17826 ( .A1(n16268), .A2(n14562), .ZN(n14563) );
  AOI211_X1 U17827 ( .C1(n16265), .C2(n14564), .A(n14717), .B(n14563), .ZN(
        n14565) );
  OAI211_X1 U17828 ( .C1(n20373), .C2(n14567), .A(n14566), .B(n14565), .ZN(
        P1_U2969) );
  XNOR2_X1 U17829 ( .A(n10070), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14568) );
  XNOR2_X1 U17830 ( .A(n14569), .B(n14568), .ZN(n14730) );
  NOR2_X1 U17831 ( .A1(n20243), .A2(n14570), .ZN(n14722) );
  AOI21_X1 U17832 ( .B1(n20367), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14722), .ZN(n14571) );
  OAI21_X1 U17833 ( .B1(n16254), .B2(n14572), .A(n14571), .ZN(n14573) );
  AOI21_X1 U17834 ( .B1(n14574), .B2(n20378), .A(n14573), .ZN(n14575) );
  OAI21_X1 U17835 ( .B1(n16244), .B2(n14730), .A(n14575), .ZN(P1_U2970) );
  INV_X1 U17836 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14576) );
  NOR2_X1 U17837 ( .A1(n20243), .A2(n14576), .ZN(n14733) );
  NOR2_X1 U17838 ( .A1(n16268), .A2(n14577), .ZN(n14578) );
  AOI211_X1 U17839 ( .C1(n16265), .C2(n14579), .A(n14733), .B(n14578), .ZN(
        n14588) );
  NOR2_X1 U17840 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14580) );
  NAND4_X1 U17841 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14750), .ZN(
        n14585) );
  NAND3_X1 U17842 ( .A1(n9753), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14584) );
  INV_X1 U17843 ( .A(n16199), .ZN(n14598) );
  AOI21_X1 U17844 ( .B1(n9753), .B2(n14698), .A(n14598), .ZN(n14583) );
  MUX2_X1 U17845 ( .A(n14585), .B(n14584), .S(n14583), .Z(n14586) );
  XNOR2_X1 U17846 ( .A(n14586), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14731) );
  NAND2_X1 U17847 ( .A1(n14731), .A2(n20369), .ZN(n14587) );
  OAI211_X1 U17848 ( .C1(n14589), .C2(n20373), .A(n14588), .B(n14587), .ZN(
        P1_U2971) );
  MUX2_X1 U17849 ( .A(n10914), .B(n14590), .S(n10070), .Z(n14591) );
  XNOR2_X1 U17850 ( .A(n14591), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14753) );
  INV_X1 U17851 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14592) );
  NOR2_X1 U17852 ( .A1(n20243), .A2(n14592), .ZN(n14744) );
  AOI21_X1 U17853 ( .B1(n20367), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14744), .ZN(n14593) );
  OAI21_X1 U17854 ( .B1(n16254), .B2(n14594), .A(n14593), .ZN(n14595) );
  AOI21_X1 U17855 ( .B1(n14596), .B2(n20378), .A(n14595), .ZN(n14597) );
  OAI21_X1 U17856 ( .B1(n16244), .B2(n14753), .A(n14597), .ZN(P1_U2972) );
  OAI21_X1 U17857 ( .B1(n14598), .B2(n14698), .A(n16212), .ZN(n14599) );
  NAND2_X1 U17858 ( .A1(n14600), .A2(n14599), .ZN(n14601) );
  XOR2_X1 U17859 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14601), .Z(
        n14763) );
  NAND2_X1 U17860 ( .A1(n16368), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14758) );
  OAI21_X1 U17861 ( .B1(n16268), .B2(n14602), .A(n14758), .ZN(n14605) );
  NOR2_X1 U17862 ( .A1(n14603), .A2(n20373), .ZN(n14604) );
  OAI21_X1 U17863 ( .B1(n16244), .B2(n14763), .A(n14607), .ZN(P1_U2973) );
  NOR2_X1 U17864 ( .A1(n14608), .A2(n16284), .ZN(n14618) );
  INV_X1 U17865 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14771) );
  MUX2_X1 U17866 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n9900), .S(
        n10070), .Z(n14609) );
  OAI21_X1 U17867 ( .B1(n14618), .B2(n14771), .A(n14609), .ZN(n14611) );
  XNOR2_X1 U17868 ( .A(n14611), .B(n14610), .ZN(n16270) );
  NOR2_X1 U17869 ( .A1(n20243), .A2(n21360), .ZN(n16272) );
  AOI21_X1 U17870 ( .B1(n20367), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16272), .ZN(n14612) );
  OAI21_X1 U17871 ( .B1(n16254), .B2(n14613), .A(n14612), .ZN(n14614) );
  AOI21_X1 U17872 ( .B1(n14615), .B2(n20378), .A(n14614), .ZN(n14616) );
  OAI21_X1 U17873 ( .B1(n16244), .B2(n16270), .A(n14616), .ZN(P1_U2974) );
  NOR2_X1 U17874 ( .A1(n14618), .A2(n16199), .ZN(n14617) );
  MUX2_X1 U17875 ( .A(n14618), .B(n14617), .S(n10070), .Z(n14619) );
  XNOR2_X1 U17876 ( .A(n14619), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14777) );
  NAND2_X1 U17877 ( .A1(n16265), .A2(n14620), .ZN(n14621) );
  NAND2_X1 U17878 ( .A1(n16368), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14765) );
  OAI211_X1 U17879 ( .C1(n16268), .C2(n14622), .A(n14621), .B(n14765), .ZN(
        n14623) );
  AOI21_X1 U17880 ( .B1(n14624), .B2(n20378), .A(n14623), .ZN(n14625) );
  OAI21_X1 U17881 ( .B1(n16244), .B2(n14777), .A(n14625), .ZN(P1_U2975) );
  NAND2_X1 U17882 ( .A1(n14627), .A2(n14626), .ZN(n14628) );
  XOR2_X1 U17883 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14628), .Z(
        n16286) );
  AOI22_X1 U17884 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14629) );
  OAI21_X1 U17885 ( .B1(n16254), .B2(n16087), .A(n14629), .ZN(n14630) );
  AOI21_X1 U17886 ( .B1(n14631), .B2(n20378), .A(n14630), .ZN(n14632) );
  OAI21_X1 U17887 ( .B1(n16244), .B2(n16286), .A(n14632), .ZN(P1_U2977) );
  NAND2_X1 U17888 ( .A1(n14633), .A2(n10070), .ZN(n14778) );
  AND2_X1 U17889 ( .A1(n9753), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14634) );
  NAND2_X1 U17890 ( .A1(n16213), .A2(n14634), .ZN(n14779) );
  NAND2_X1 U17891 ( .A1(n14778), .A2(n14779), .ZN(n14635) );
  XNOR2_X1 U17892 ( .A(n14635), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14807) );
  NAND2_X1 U17893 ( .A1(n16368), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14797) );
  OAI21_X1 U17894 ( .B1(n16268), .B2(n16117), .A(n14797), .ZN(n14637) );
  NOR2_X1 U17895 ( .A1(n16111), .A2(n20373), .ZN(n14636) );
  AOI211_X1 U17896 ( .C1(n16265), .C2(n16107), .A(n14637), .B(n14636), .ZN(
        n14638) );
  OAI21_X1 U17897 ( .B1(n14807), .B2(n16244), .A(n14638), .ZN(P1_U2979) );
  AND2_X1 U17898 ( .A1(n16368), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14814) );
  NOR2_X1 U17899 ( .A1(n16132), .A2(n16254), .ZN(n14639) );
  AOI211_X1 U17900 ( .C1(n20367), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14814), .B(n14639), .ZN(n14643) );
  OR2_X1 U17901 ( .A1(n14641), .A2(n14640), .ZN(n14811) );
  NAND3_X1 U17902 ( .A1(n9973), .A2(n20369), .A3(n14811), .ZN(n14642) );
  OAI211_X1 U17903 ( .C1(n16140), .C2(n20373), .A(n14643), .B(n14642), .ZN(
        P1_U2981) );
  OR2_X1 U17904 ( .A1(n14644), .A2(n14645), .ZN(n16228) );
  AOI21_X1 U17905 ( .B1(n16228), .B2(n14820), .A(n16230), .ZN(n14646) );
  XOR2_X1 U17906 ( .A(n14647), .B(n14646), .Z(n16305) );
  AOI22_X1 U17907 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14648) );
  OAI21_X1 U17908 ( .B1(n16254), .B2(n14649), .A(n14648), .ZN(n14650) );
  AOI21_X1 U17909 ( .B1(n14651), .B2(n20378), .A(n14650), .ZN(n14652) );
  OAI21_X1 U17910 ( .B1(n16244), .B2(n16305), .A(n14652), .ZN(P1_U2983) );
  INV_X1 U17911 ( .A(n14644), .ZN(n14664) );
  INV_X1 U17912 ( .A(n16225), .ZN(n14653) );
  OAI21_X1 U17913 ( .B1(n14664), .B2(n14653), .A(n9932), .ZN(n14655) );
  NAND2_X1 U17914 ( .A1(n14655), .A2(n14654), .ZN(n14657) );
  MUX2_X1 U17915 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n10907), .S(
        n9753), .Z(n14656) );
  XNOR2_X1 U17916 ( .A(n14657), .B(n14656), .ZN(n14832) );
  NAND2_X1 U17917 ( .A1(n14832), .A2(n20369), .ZN(n14660) );
  NOR2_X1 U17918 ( .A1(n20243), .A2(n14163), .ZN(n14835) );
  NOR2_X1 U17919 ( .A1(n16254), .A2(n16159), .ZN(n14658) );
  AOI211_X1 U17920 ( .C1(n20367), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14835), .B(n14658), .ZN(n14659) );
  OAI211_X1 U17921 ( .C1(n20373), .C2(n16162), .A(n14660), .B(n14659), .ZN(
        P1_U2985) );
  INV_X1 U17922 ( .A(n14661), .ZN(n14662) );
  AOI22_X1 U17923 ( .A1(n14664), .A2(n14663), .B1(n10070), .B2(n14662), .ZN(
        n14840) );
  INV_X1 U17924 ( .A(n14666), .ZN(n14665) );
  AOI21_X1 U17925 ( .B1(n10070), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14665), .ZN(n14839) );
  NAND2_X1 U17926 ( .A1(n14840), .A2(n14839), .ZN(n14838) );
  NAND2_X1 U17927 ( .A1(n14838), .A2(n14666), .ZN(n14667) );
  XOR2_X1 U17928 ( .A(n14668), .B(n14667), .Z(n16327) );
  NAND2_X1 U17929 ( .A1(n16327), .A2(n20369), .ZN(n14672) );
  NOR2_X1 U17930 ( .A1(n20243), .A2(n21064), .ZN(n16324) );
  AND2_X1 U17931 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14669) );
  AOI211_X1 U17932 ( .C1(n14670), .C2(n16265), .A(n16324), .B(n14669), .ZN(
        n14671) );
  OAI211_X1 U17933 ( .C1(n20373), .C2(n14673), .A(n14672), .B(n14671), .ZN(
        P1_U2986) );
  XNOR2_X1 U17934 ( .A(n14644), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14676) );
  AND2_X1 U17935 ( .A1(n14674), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14675) );
  MUX2_X1 U17936 ( .A(n14676), .B(n14675), .S(n10070), .Z(n14677) );
  NOR3_X1 U17937 ( .A1(n14674), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9753), .ZN(n16247) );
  NOR2_X1 U17938 ( .A1(n14677), .A2(n16247), .ZN(n16341) );
  AOI22_X1 U17939 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14678) );
  OAI21_X1 U17940 ( .B1(n16254), .B2(n14679), .A(n14678), .ZN(n14680) );
  AOI21_X1 U17941 ( .B1(n14681), .B2(n20378), .A(n14680), .ZN(n14682) );
  OAI21_X1 U17942 ( .B1(n16341), .B2(n16244), .A(n14682), .ZN(P1_U2989) );
  XNOR2_X1 U17943 ( .A(n9753), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14683) );
  XNOR2_X1 U17944 ( .A(n14684), .B(n14683), .ZN(n16351) );
  INV_X1 U17945 ( .A(n20289), .ZN(n20200) );
  AOI22_X1 U17946 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14685) );
  OAI21_X1 U17947 ( .B1(n16254), .B2(n14686), .A(n14685), .ZN(n14687) );
  AOI21_X1 U17948 ( .B1(n20200), .B2(n20378), .A(n14687), .ZN(n14688) );
  OAI21_X1 U17949 ( .B1(n16351), .B2(n16244), .A(n14688), .ZN(P1_U2990) );
  NOR4_X1 U17950 ( .A1(n21199), .A2(n10907), .A3(n16313), .A4(n10911), .ZN(
        n14812) );
  NAND2_X1 U17951 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14812), .ZN(
        n14701) );
  INV_X1 U17952 ( .A(n14701), .ZN(n14696) );
  INV_X1 U17953 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16350) );
  NAND3_X1 U17954 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16343) );
  NOR3_X1 U17955 ( .A1(n16350), .A2(n16361), .A3(n16343), .ZN(n14849) );
  NAND2_X1 U17956 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14849), .ZN(
        n14846) );
  INV_X1 U17957 ( .A(n14846), .ZN(n14690) );
  NAND2_X1 U17958 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14690), .ZN(
        n14694) );
  NOR2_X1 U17959 ( .A1(n16340), .A2(n14694), .ZN(n14786) );
  NAND2_X1 U17960 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14786), .ZN(
        n14810) );
  NOR2_X1 U17961 ( .A1(n10850), .A2(n14691), .ZN(n14693) );
  NAND2_X1 U17962 ( .A1(n14693), .A2(n14692), .ZN(n14841) );
  NOR2_X1 U17963 ( .A1(n14694), .A2(n14841), .ZN(n14699) );
  INV_X1 U17964 ( .A(n14699), .ZN(n14787) );
  NOR2_X1 U17965 ( .A1(n16330), .A2(n14787), .ZN(n14808) );
  NAND2_X1 U17966 ( .A1(n14695), .A2(n14808), .ZN(n14770) );
  OAI21_X1 U17967 ( .B1(n14810), .B2(n14769), .A(n14770), .ZN(n16306) );
  NAND4_X1 U17968 ( .A1(n14697), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14696), .A4(n16306), .ZN(n16278) );
  NOR2_X1 U17969 ( .A1(n16278), .A2(n14698), .ZN(n14757) );
  INV_X1 U17970 ( .A(n14739), .ZN(n14721) );
  NAND3_X1 U17971 ( .A1(n14751), .A2(n14721), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14715) );
  NOR3_X1 U17972 ( .A1(n14715), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14714), .ZN(n14709) );
  NAND2_X1 U17973 ( .A1(n14842), .A2(n16303), .ZN(n14746) );
  NAND2_X1 U17974 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16291) );
  NOR2_X1 U17975 ( .A1(n16330), .A2(n14701), .ZN(n14788) );
  OAI221_X1 U17976 ( .B1(n14844), .B2(n14699), .C1(n14844), .C2(n14788), .A(
        n14842), .ZN(n14700) );
  INV_X1 U17977 ( .A(n14789), .ZN(n14703) );
  INV_X1 U17978 ( .A(n14746), .ZN(n14702) );
  AOI21_X1 U17979 ( .B1(n14801), .B2(n14703), .A(n14702), .ZN(n16289) );
  AOI21_X1 U17980 ( .B1(n16364), .B2(n16291), .A(n16289), .ZN(n16285) );
  OAI21_X1 U17981 ( .B1(n14768), .B2(n16303), .A(n16285), .ZN(n16275) );
  NOR2_X1 U17982 ( .A1(n14704), .A2(n16275), .ZN(n14755) );
  AND2_X1 U17983 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14755), .ZN(
        n14743) );
  NAND2_X1 U17984 ( .A1(n14721), .A2(n14743), .ZN(n14705) );
  NAND2_X1 U17985 ( .A1(n14746), .A2(n14705), .ZN(n14726) );
  OAI211_X1 U17986 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16303), .A(
        n14726), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14712) );
  NAND3_X1 U17987 ( .A1(n14712), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14746), .ZN(n14707) );
  NAND2_X1 U17988 ( .A1(n14707), .A2(n14706), .ZN(n14708) );
  INV_X1 U17989 ( .A(n14711), .ZN(n14720) );
  INV_X1 U17990 ( .A(n14712), .ZN(n14713) );
  AOI21_X1 U17991 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14716) );
  AOI211_X1 U17992 ( .C1(n14718), .C2(n16395), .A(n14717), .B(n14716), .ZN(
        n14719) );
  OAI21_X1 U17993 ( .B1(n14720), .B2(n16319), .A(n14719), .ZN(P1_U3001) );
  INV_X1 U17994 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14725) );
  NAND3_X1 U17995 ( .A1(n14751), .A2(n14721), .A3(n14725), .ZN(n14724) );
  INV_X1 U17996 ( .A(n14722), .ZN(n14723) );
  OAI211_X1 U17997 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14727) );
  AOI21_X1 U17998 ( .B1(n14728), .B2(n16395), .A(n14727), .ZN(n14729) );
  OAI21_X1 U17999 ( .B1(n14730), .B2(n16319), .A(n14729), .ZN(P1_U3002) );
  INV_X1 U18000 ( .A(n14731), .ZN(n14742) );
  INV_X1 U18001 ( .A(n14743), .ZN(n14732) );
  NAND3_X1 U18002 ( .A1(n14746), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n14732), .ZN(n14735) );
  INV_X1 U18003 ( .A(n14733), .ZN(n14734) );
  NAND2_X1 U18004 ( .A1(n14735), .A2(n14734), .ZN(n14736) );
  AOI21_X1 U18005 ( .B1(n14737), .B2(n16395), .A(n14736), .ZN(n14741) );
  NAND3_X1 U18006 ( .A1(n14751), .A2(n14739), .A3(n14738), .ZN(n14740) );
  OAI211_X1 U18007 ( .C1(n14742), .C2(n16319), .A(n14741), .B(n14740), .ZN(
        P1_U3003) );
  NOR2_X1 U18008 ( .A1(n14743), .A2(n14750), .ZN(n14745) );
  AOI21_X1 U18009 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14747) );
  OAI21_X1 U18010 ( .B1(n14748), .B2(n16383), .A(n14747), .ZN(n14749) );
  AOI21_X1 U18011 ( .B1(n14751), .B2(n14750), .A(n14749), .ZN(n14752) );
  OAI21_X1 U18012 ( .B1(n14753), .B2(n16319), .A(n14752), .ZN(P1_U3004) );
  INV_X1 U18013 ( .A(n14768), .ZN(n14754) );
  NOR3_X1 U18014 ( .A1(n16278), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14754), .ZN(n16271) );
  INV_X1 U18015 ( .A(n14755), .ZN(n14756) );
  OAI22_X1 U18016 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14757), .B1(
        n16271), .B2(n14756), .ZN(n14762) );
  INV_X1 U18017 ( .A(n14758), .ZN(n14759) );
  AOI21_X1 U18018 ( .B1(n14760), .B2(n16395), .A(n14759), .ZN(n14761) );
  OAI211_X1 U18019 ( .C1(n14763), .C2(n16319), .A(n14762), .B(n14761), .ZN(
        P1_U3005) );
  INV_X1 U18020 ( .A(n14764), .ZN(n14767) );
  INV_X1 U18021 ( .A(n14765), .ZN(n14766) );
  AOI21_X1 U18022 ( .B1(n14767), .B2(n16395), .A(n14766), .ZN(n14776) );
  INV_X1 U18023 ( .A(n16285), .ZN(n14774) );
  AOI21_X1 U18024 ( .B1(n14770), .B2(n14769), .A(n14768), .ZN(n14773) );
  OAI21_X1 U18025 ( .B1(n16284), .B2(n16278), .A(n14771), .ZN(n14772) );
  OAI21_X1 U18026 ( .B1(n14774), .B2(n14773), .A(n14772), .ZN(n14775) );
  OAI211_X1 U18027 ( .C1(n14777), .C2(n16319), .A(n14776), .B(n14775), .ZN(
        P1_U3007) );
  INV_X1 U18028 ( .A(n16289), .ZN(n14796) );
  NAND2_X1 U18029 ( .A1(n14778), .A2(n14114), .ZN(n14781) );
  NAND2_X1 U18030 ( .A1(n14779), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14780) );
  NAND2_X1 U18031 ( .A1(n14781), .A2(n14780), .ZN(n14782) );
  XNOR2_X1 U18032 ( .A(n14782), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16205) );
  NAND2_X1 U18033 ( .A1(n16205), .A2(n16400), .ZN(n14794) );
  NOR3_X1 U18034 ( .A1(n14784), .A2(n14783), .A3(n14787), .ZN(n14785) );
  AOI21_X1 U18035 ( .B1(n14786), .B2(n14847), .A(n14785), .ZN(n14803) );
  OAI21_X1 U18036 ( .B1(n14787), .B2(n14802), .A(n14803), .ZN(n16326) );
  NAND2_X1 U18037 ( .A1(n14788), .A2(n16326), .ZN(n16302) );
  NOR2_X1 U18038 ( .A1(n14789), .A2(n16302), .ZN(n16292) );
  NAND2_X1 U18039 ( .A1(n9926), .A2(n14790), .ZN(n14791) );
  NAND2_X1 U18040 ( .A1(n9879), .A2(n14791), .ZN(n16186) );
  OAI22_X1 U18041 ( .A1(n16186), .A2(n16383), .B1(n20243), .B2(n16097), .ZN(
        n14792) );
  AOI21_X1 U18042 ( .B1(n16292), .B2(n14795), .A(n14792), .ZN(n14793) );
  OAI211_X1 U18043 ( .C1(n14796), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        P1_U3010) );
  INV_X1 U18044 ( .A(n16110), .ZN(n14800) );
  INV_X1 U18045 ( .A(n14797), .ZN(n14799) );
  NOR3_X1 U18046 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10912), .A3(
        n16302), .ZN(n14798) );
  AOI211_X1 U18047 ( .C1(n16395), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14806) );
  INV_X1 U18048 ( .A(n14801), .ZN(n16296) );
  AOI21_X1 U18049 ( .B1(n14803), .B2(n14802), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14804) );
  OAI21_X1 U18050 ( .B1(n16296), .B2(n14804), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14805) );
  OAI211_X1 U18051 ( .C1(n14807), .C2(n16319), .A(n14806), .B(n14805), .ZN(
        P1_U3011) );
  OAI21_X1 U18052 ( .B1(n14844), .B2(n14808), .A(n14842), .ZN(n14809) );
  AOI21_X1 U18053 ( .B1(n14847), .B2(n14810), .A(n14809), .ZN(n16331) );
  OAI21_X1 U18054 ( .B1(n16303), .B2(n14812), .A(n16331), .ZN(n14829) );
  INV_X1 U18055 ( .A(n14829), .ZN(n14819) );
  NAND3_X1 U18056 ( .A1(n9973), .A2(n16400), .A3(n14811), .ZN(n14817) );
  INV_X1 U18057 ( .A(n16143), .ZN(n14815) );
  AND3_X1 U18058 ( .A1(n14818), .A2(n16306), .A3(n14812), .ZN(n14813) );
  AOI211_X1 U18059 ( .C1(n16395), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14816) );
  OAI211_X1 U18060 ( .C1(n14819), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        P1_U3013) );
  NOR2_X1 U18061 ( .A1(n16212), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14823) );
  NAND2_X1 U18062 ( .A1(n14821), .A2(n14820), .ZN(n14822) );
  MUX2_X1 U18063 ( .A(n14823), .B(n9753), .S(n14822), .Z(n14824) );
  XNOR2_X1 U18064 ( .A(n14824), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16224) );
  INV_X1 U18065 ( .A(n16306), .ZN(n14826) );
  NAND3_X1 U18066 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14825) );
  OAI21_X1 U18067 ( .B1(n14826), .B2(n14825), .A(n10911), .ZN(n14830) );
  INV_X1 U18068 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14827) );
  OAI22_X1 U18069 ( .A1(n16144), .A2(n16383), .B1(n20243), .B2(n14827), .ZN(
        n14828) );
  AOI21_X1 U18070 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14831) );
  OAI21_X1 U18071 ( .B1(n16224), .B2(n16319), .A(n14831), .ZN(P1_U3014) );
  INV_X1 U18072 ( .A(n14832), .ZN(n14837) );
  INV_X1 U18073 ( .A(n16331), .ZN(n14833) );
  MUX2_X1 U18074 ( .A(n16306), .B(n14833), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n14834) );
  AOI211_X1 U18075 ( .C1(n16395), .C2(n16165), .A(n14835), .B(n14834), .ZN(
        n14836) );
  OAI21_X1 U18076 ( .B1(n14837), .B2(n16319), .A(n14836), .ZN(P1_U3017) );
  OAI21_X1 U18077 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n16239) );
  INV_X1 U18078 ( .A(n16366), .ZN(n16342) );
  NOR3_X1 U18079 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14846), .A3(
        n16342), .ZN(n14855) );
  INV_X1 U18080 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21065) );
  INV_X1 U18081 ( .A(n14841), .ZN(n14843) );
  OAI221_X1 U18082 ( .B1(n14844), .B2(n14843), .C1(n14844), .C2(n14849), .A(
        n14842), .ZN(n14845) );
  AOI221_X1 U18083 ( .B1(n16340), .B2(n14847), .C1(n14846), .C2(n14847), .A(
        n14845), .ZN(n16338) );
  INV_X1 U18084 ( .A(n16338), .ZN(n14851) );
  INV_X1 U18085 ( .A(n14848), .ZN(n14850) );
  INV_X1 U18086 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16337) );
  AND2_X1 U18087 ( .A1(n16337), .A2(n14849), .ZN(n16333) );
  OAI221_X1 U18088 ( .B1(n14851), .B2(n14850), .C1(n14851), .C2(n16333), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U18089 ( .A1(n16170), .A2(n16395), .ZN(n14852) );
  OAI211_X1 U18090 ( .C1(n21065), .C2(n20243), .A(n14853), .B(n14852), .ZN(
        n14854) );
  AOI211_X1 U18091 ( .C1(n16239), .C2(n16400), .A(n14855), .B(n14854), .ZN(
        n14856) );
  INV_X1 U18092 ( .A(n14856), .ZN(P1_U3019) );
  INV_X1 U18093 ( .A(n14186), .ZN(n20896) );
  NAND2_X1 U18094 ( .A1(n14858), .A2(n14857), .ZN(n14859) );
  OAI22_X1 U18095 ( .A1(n16020), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14859), .B2(n10622), .ZN(n14860) );
  AOI21_X1 U18096 ( .B1(n20896), .B2(n14861), .A(n14860), .ZN(n16021) );
  INV_X1 U18097 ( .A(n21102), .ZN(n14867) );
  AOI21_X1 U18098 ( .B1(n14865), .B2(n14864), .A(n14863), .ZN(n14866) );
  OAI21_X1 U18099 ( .B1(n16021), .B2(n14867), .A(n14866), .ZN(n14868) );
  MUX2_X1 U18100 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14868), .S(
        n16407), .Z(P1_U3473) );
  AOI22_X1 U18101 ( .A1(n14869), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14872) );
  NAND2_X1 U18102 ( .A1(n14870), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14871) );
  OAI211_X1 U18103 ( .C1(n12244), .C2(n15335), .A(n14872), .B(n14871), .ZN(
        n14874) );
  XNOR2_X1 U18104 ( .A(n14875), .B(n14874), .ZN(n16480) );
  NAND4_X1 U18105 ( .A1(n16418), .A2(n19336), .A3(n9751), .A4(n15139), .ZN(
        n14893) );
  INV_X1 U18106 ( .A(n16454), .ZN(n14878) );
  NOR2_X1 U18107 ( .A1(n14876), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14877) );
  MUX2_X1 U18108 ( .A(n14878), .B(n14877), .S(n11860), .Z(n15121) );
  INV_X1 U18109 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20093) );
  OAI22_X1 U18110 ( .A1(n20093), .A2(n19341), .B1(n12319), .B2(n19282), .ZN(
        n14891) );
  NAND2_X1 U18111 ( .A1(n14879), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14882) );
  NAND2_X1 U18112 ( .A1(n14880), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n14881) );
  OAI211_X1 U18113 ( .C1(n14883), .C2(n20093), .A(n14882), .B(n14881), .ZN(
        n14884) );
  INV_X1 U18114 ( .A(n14884), .ZN(n14885) );
  OR3_X1 U18115 ( .A1(n14888), .A2(n12547), .A3(n14887), .ZN(n14889) );
  OAI21_X1 U18116 ( .B1(n19390), .B2(n19335), .A(n14889), .ZN(n14890) );
  AOI211_X1 U18117 ( .C1(n15121), .C2(n19339), .A(n14891), .B(n14890), .ZN(
        n14892) );
  OAI211_X1 U18118 ( .C1(n16480), .C2(n19346), .A(n14893), .B(n14892), .ZN(
        P2_U2824) );
  AOI21_X1 U18119 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  NAND2_X1 U18120 ( .A1(n14897), .A2(n19336), .ZN(n14903) );
  AOI22_X1 U18121 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19349), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19327), .ZN(n14898) );
  OAI21_X1 U18122 ( .B1(n19335), .B2(n15020), .A(n14898), .ZN(n14901) );
  NOR2_X1 U18123 ( .A1(n14899), .A2(n19306), .ZN(n14900) );
  AOI211_X1 U18124 ( .C1(P2_EBX_REG_28__SCAN_IN), .C2(n19344), .A(n14901), .B(
        n14900), .ZN(n14902) );
  OAI211_X1 U18125 ( .C1(n19346), .C2(n14961), .A(n14903), .B(n14902), .ZN(
        P2_U2827) );
  NAND2_X1 U18126 ( .A1(n9887), .A2(n14904), .ZN(n14905) );
  NAND2_X1 U18127 ( .A1(n9876), .A2(n14905), .ZN(n15390) );
  AND2_X1 U18128 ( .A1(n15055), .A2(n14906), .ZN(n14907) );
  OR2_X1 U18129 ( .A1(n14907), .A2(n9886), .ZN(n15393) );
  INV_X1 U18130 ( .A(n15393), .ZN(n15044) );
  AOI22_X1 U18131 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19327), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19344), .ZN(n14908) );
  OAI21_X1 U18132 ( .B1(n15175), .B2(n19282), .A(n14908), .ZN(n14909) );
  AOI21_X1 U18133 ( .B1(n19337), .B2(n15044), .A(n14909), .ZN(n14910) );
  OAI21_X1 U18134 ( .B1(n15390), .B2(n19346), .A(n14910), .ZN(n14914) );
  AOI211_X1 U18135 ( .C1(n14912), .C2(n15177), .A(n14911), .B(n20024), .ZN(
        n14913) );
  AOI211_X1 U18136 ( .C1(n19339), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        n14916) );
  INV_X1 U18137 ( .A(n14916), .ZN(P2_U2830) );
  NAND2_X1 U18138 ( .A1(n9923), .A2(n14917), .ZN(n14918) );
  NAND2_X1 U18139 ( .A1(n14919), .A2(n14918), .ZN(n16489) );
  NOR2_X1 U18140 ( .A1(n15087), .A2(n14920), .ZN(n14921) );
  OR2_X1 U18141 ( .A1(n14922), .A2(n14921), .ZN(n15454) );
  AOI22_X1 U18142 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19349), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19327), .ZN(n14923) );
  OAI21_X1 U18143 ( .B1(n19335), .B2(n15454), .A(n14923), .ZN(n14924) );
  AOI21_X1 U18144 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n19344), .A(n14924), .ZN(
        n14925) );
  OAI21_X1 U18145 ( .B1(n16489), .B2(n19346), .A(n14925), .ZN(n14930) );
  AOI211_X1 U18146 ( .C1(n14928), .C2(n14927), .A(n14926), .B(n20024), .ZN(
        n14929) );
  AOI211_X1 U18147 ( .C1(n19339), .C2(n14931), .A(n14930), .B(n14929), .ZN(
        n14932) );
  INV_X1 U18148 ( .A(n14932), .ZN(P2_U2835) );
  NOR3_X1 U18149 ( .A1(n19312), .A2(n14941), .A3(n20024), .ZN(n19212) );
  INV_X1 U18150 ( .A(n19212), .ZN(n14946) );
  AND2_X1 U18151 ( .A1(n15005), .A2(n14933), .ZN(n14934) );
  OR2_X1 U18152 ( .A1(n14998), .A2(n14934), .ZN(n16492) );
  NAND2_X1 U18153 ( .A1(n15099), .A2(n14935), .ZN(n14936) );
  AND2_X1 U18154 ( .A1(n15086), .A2(n14936), .ZN(n16500) );
  INV_X1 U18155 ( .A(n16500), .ZN(n14938) );
  AOI22_X1 U18156 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19327), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19349), .ZN(n14937) );
  OAI211_X1 U18157 ( .C1(n19335), .C2(n14938), .A(n14937), .B(n19305), .ZN(
        n14939) );
  AOI21_X1 U18158 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19344), .A(n14939), .ZN(
        n14940) );
  OAI21_X1 U18159 ( .B1(n16492), .B2(n19346), .A(n14940), .ZN(n14943) );
  AOI211_X1 U18160 ( .C1(n9751), .C2(n10102), .A(n20024), .B(n15247), .ZN(
        n14942) );
  AOI211_X1 U18161 ( .C1(n19339), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14945) );
  OAI21_X1 U18162 ( .B1(n10101), .B2(n14946), .A(n14945), .ZN(P2_U2837) );
  NAND2_X1 U18163 ( .A1(n14948), .A2(n14947), .ZN(n14949) );
  NAND2_X1 U18164 ( .A1(n14950), .A2(n14949), .ZN(n16428) );
  OR2_X1 U18165 ( .A1(n14952), .A2(n14951), .ZN(n15009) );
  NAND3_X1 U18166 ( .A1(n15009), .A2(n14953), .A3(n19386), .ZN(n14955) );
  NAND2_X1 U18167 ( .A1(n19385), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14954) );
  OAI211_X1 U18168 ( .C1(n19385), .C2(n16428), .A(n14955), .B(n14954), .ZN(
        P2_U2858) );
  INV_X1 U18169 ( .A(n14956), .ZN(n14958) );
  NOR2_X1 U18170 ( .A1(n14958), .A2(n14957), .ZN(n14960) );
  XNOR2_X1 U18171 ( .A(n14960), .B(n14959), .ZN(n15026) );
  NOR2_X1 U18172 ( .A1(n14961), .A2(n19385), .ZN(n14962) );
  AOI21_X1 U18173 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19385), .A(n14962), .ZN(
        n14963) );
  OAI21_X1 U18174 ( .B1(n15026), .B2(n19380), .A(n14963), .ZN(P2_U2859) );
  OAI21_X1 U18175 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n15036) );
  OAI21_X1 U18176 ( .B1(n14975), .B2(n14968), .A(n14967), .ZN(n16444) );
  NOR2_X1 U18177 ( .A1(n16444), .A2(n19385), .ZN(n14969) );
  AOI21_X1 U18178 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19385), .A(n14969), .ZN(
        n14970) );
  OAI21_X1 U18179 ( .B1(n15036), .B2(n19380), .A(n14970), .ZN(P2_U2860) );
  OAI21_X1 U18180 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(n15042) );
  AND2_X1 U18181 ( .A1(n9876), .A2(n14974), .ZN(n14976) );
  OR2_X1 U18182 ( .A1(n14976), .A2(n14975), .ZN(n16459) );
  NOR2_X1 U18183 ( .A1(n16459), .A2(n19385), .ZN(n14977) );
  AOI21_X1 U18184 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19385), .A(n14977), .ZN(
        n14978) );
  OAI21_X1 U18185 ( .B1(n15042), .B2(n19380), .A(n14978), .ZN(P2_U2861) );
  OAI21_X1 U18186 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n15051) );
  MUX2_X1 U18187 ( .A(n15390), .B(n14982), .S(n19385), .Z(n14983) );
  OAI21_X1 U18188 ( .B1(n15051), .B2(n19380), .A(n14983), .ZN(P2_U2862) );
  AOI21_X1 U18189 ( .B1(n14984), .B2(n14985), .A(n9849), .ZN(n14986) );
  XOR2_X1 U18190 ( .A(n14987), .B(n14986), .Z(n15060) );
  OAI21_X1 U18191 ( .B1(n14989), .B2(n14988), .A(n9887), .ZN(n16469) );
  MUX2_X1 U18192 ( .A(n16471), .B(n16469), .S(n19356), .Z(n14990) );
  OAI21_X1 U18193 ( .B1(n15060), .B2(n19380), .A(n14990), .ZN(P2_U2863) );
  OAI21_X1 U18194 ( .B1(n14992), .B2(n14994), .A(n14993), .ZN(n15083) );
  NOR2_X1 U18195 ( .A1(n15441), .A2(n19385), .ZN(n14995) );
  AOI21_X1 U18196 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19385), .A(n14995), .ZN(
        n14996) );
  OAI21_X1 U18197 ( .B1(n15083), .B2(n19380), .A(n14996), .ZN(P2_U2866) );
  OAI21_X1 U18198 ( .B1(n9840), .B2(n9955), .A(n9924), .ZN(n15093) );
  OR2_X1 U18199 ( .A1(n14998), .A2(n14997), .ZN(n14999) );
  NAND2_X1 U18200 ( .A1(n9923), .A2(n14999), .ZN(n19194) );
  NOR2_X1 U18201 ( .A1(n19194), .A2(n19385), .ZN(n15000) );
  AOI21_X1 U18202 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19385), .A(n15000), .ZN(
        n15001) );
  OAI21_X1 U18203 ( .B1(n15093), .B2(n19380), .A(n15001), .ZN(P2_U2868) );
  OAI21_X1 U18204 ( .B1(n15002), .B2(n15004), .A(n15003), .ZN(n15105) );
  NAND2_X1 U18205 ( .A1(n19385), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15008) );
  AOI21_X1 U18206 ( .B1(n15006), .B2(n15266), .A(n10220), .ZN(n19210) );
  NAND2_X1 U18207 ( .A1(n19210), .A2(n19356), .ZN(n15007) );
  OAI211_X1 U18208 ( .C1(n15105), .C2(n19380), .A(n15008), .B(n15007), .ZN(
        P2_U2870) );
  NAND3_X1 U18209 ( .A1(n15009), .A2(n14953), .A3(n16501), .ZN(n15019) );
  AOI22_X1 U18210 ( .A1(n19397), .A2(BUF1_REG_29__SCAN_IN), .B1(n19396), .B2(
        n15010), .ZN(n15018) );
  NOR2_X1 U18211 ( .A1(n15012), .A2(n15011), .ZN(n15013) );
  OAI22_X1 U18212 ( .A1(n19400), .A2(n16433), .B1(n15094), .B2(n15015), .ZN(
        n15016) );
  AOI21_X1 U18213 ( .B1(n19398), .B2(BUF2_REG_29__SCAN_IN), .A(n15016), .ZN(
        n15017) );
  NAND3_X1 U18214 ( .A1(n15019), .A2(n15018), .A3(n15017), .ZN(P2_U2890) );
  INV_X1 U18215 ( .A(n15020), .ZN(n15021) );
  AOI22_X1 U18216 ( .A1(n19397), .A2(BUF1_REG_28__SCAN_IN), .B1(n19392), .B2(
        n15021), .ZN(n15025) );
  OAI22_X1 U18217 ( .A1(n15096), .A2(n15022), .B1(n15094), .B2(n13149), .ZN(
        n15023) );
  AOI21_X1 U18218 ( .B1(n19398), .B2(BUF2_REG_28__SCAN_IN), .A(n15023), .ZN(
        n15024) );
  OAI211_X1 U18219 ( .C1(n15026), .C2(n19422), .A(n15025), .B(n15024), .ZN(
        P2_U2891) );
  INV_X1 U18220 ( .A(n19398), .ZN(n15048) );
  INV_X1 U18221 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U18222 ( .A1(n19397), .A2(BUF1_REG_27__SCAN_IN), .B1(n19396), .B2(
        n15027), .ZN(n15032) );
  NAND2_X1 U18223 ( .A1(n15037), .A2(n15028), .ZN(n15029) );
  NAND2_X1 U18224 ( .A1(n9872), .A2(n15029), .ZN(n16448) );
  INV_X1 U18225 ( .A(n16448), .ZN(n15030) );
  AOI22_X1 U18226 ( .A1(n19392), .A2(n15030), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n19419), .ZN(n15031) );
  OAI211_X1 U18227 ( .C1(n15048), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15034) );
  INV_X1 U18228 ( .A(n15034), .ZN(n15035) );
  OAI21_X1 U18229 ( .B1(n15036), .B2(n19422), .A(n15035), .ZN(P2_U2892) );
  AOI22_X1 U18230 ( .A1(n19397), .A2(BUF1_REG_26__SCAN_IN), .B1(n19396), .B2(
        n19412), .ZN(n15041) );
  OAI21_X1 U18231 ( .B1(n9886), .B2(n15038), .A(n15037), .ZN(n15380) );
  OAI22_X1 U18232 ( .A1(n19400), .A2(n15380), .B1(n15094), .B2(n13160), .ZN(
        n15039) );
  AOI21_X1 U18233 ( .B1(n19398), .B2(BUF2_REG_26__SCAN_IN), .A(n15039), .ZN(
        n15040) );
  OAI211_X1 U18234 ( .C1(n15042), .C2(n19422), .A(n15041), .B(n15040), .ZN(
        P2_U2893) );
  INV_X1 U18235 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15047) );
  AOI22_X1 U18236 ( .A1(n19397), .A2(BUF1_REG_25__SCAN_IN), .B1(n19396), .B2(
        n15043), .ZN(n15046) );
  AOI22_X1 U18237 ( .A1(n19392), .A2(n15044), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19419), .ZN(n15045) );
  OAI211_X1 U18238 ( .C1(n15048), .C2(n15047), .A(n15046), .B(n15045), .ZN(
        n15049) );
  INV_X1 U18239 ( .A(n15049), .ZN(n15050) );
  OAI21_X1 U18240 ( .B1(n15051), .B2(n19422), .A(n15050), .ZN(P2_U2894) );
  AOI22_X1 U18241 ( .A1(n19397), .A2(BUF1_REG_24__SCAN_IN), .B1(n19396), .B2(
        n19415), .ZN(n15059) );
  NAND2_X1 U18242 ( .A1(n15053), .A2(n15052), .ZN(n15054) );
  AND2_X1 U18243 ( .A1(n15055), .A2(n15054), .ZN(n16478) );
  INV_X1 U18244 ( .A(n16478), .ZN(n15056) );
  OAI22_X1 U18245 ( .A1(n19400), .A2(n15056), .B1(n15094), .B2(n13151), .ZN(
        n15057) );
  AOI21_X1 U18246 ( .B1(n19398), .B2(BUF2_REG_24__SCAN_IN), .A(n15057), .ZN(
        n15058) );
  OAI211_X1 U18247 ( .C1(n15060), .C2(n19422), .A(n15059), .B(n15058), .ZN(
        P2_U2895) );
  NOR2_X1 U18248 ( .A1(n15061), .A2(n15062), .ZN(n15064) );
  NOR2_X1 U18249 ( .A1(n15064), .A2(n15063), .ZN(n16483) );
  INV_X1 U18250 ( .A(n16483), .ZN(n15071) );
  OAI22_X1 U18251 ( .A1(n15096), .A2(n19492), .B1(n15094), .B2(n15065), .ZN(
        n15069) );
  INV_X1 U18252 ( .A(n19397), .ZN(n15101) );
  OAI22_X1 U18253 ( .A1(n15101), .A2(n15067), .B1(n19400), .B2(n15066), .ZN(
        n15068) );
  AOI211_X1 U18254 ( .C1(n19398), .C2(BUF2_REG_23__SCAN_IN), .A(n15069), .B(
        n15068), .ZN(n15070) );
  OAI21_X1 U18255 ( .B1(n15071), .B2(n19422), .A(n15070), .ZN(P2_U2896) );
  AOI21_X1 U18256 ( .B1(n15073), .B2(n14993), .A(n15072), .ZN(n16485) );
  INV_X1 U18257 ( .A(n16485), .ZN(n15078) );
  AOI22_X1 U18258 ( .A1(n19397), .A2(BUF1_REG_22__SCAN_IN), .B1(n19392), .B2(
        n15435), .ZN(n15077) );
  OAI22_X1 U18259 ( .A1(n15096), .A2(n19482), .B1(n15094), .B2(n15074), .ZN(
        n15075) );
  AOI21_X1 U18260 ( .B1(n19398), .B2(BUF2_REG_22__SCAN_IN), .A(n15075), .ZN(
        n15076) );
  OAI211_X1 U18261 ( .C1(n15078), .C2(n19422), .A(n15077), .B(n15076), .ZN(
        P2_U2897) );
  OAI22_X1 U18262 ( .A1(n15096), .A2(n19418), .B1(n15094), .B2(n15079), .ZN(
        n15081) );
  OAI22_X1 U18263 ( .A1(n15101), .A2(n16744), .B1(n19400), .B2(n15446), .ZN(
        n15080) );
  AOI211_X1 U18264 ( .C1(n19398), .C2(BUF2_REG_21__SCAN_IN), .A(n15081), .B(
        n15080), .ZN(n15082) );
  OAI21_X1 U18265 ( .B1(n15083), .B2(n19422), .A(n15082), .ZN(P2_U2898) );
  OAI22_X1 U18266 ( .A1(n15096), .A2(n19473), .B1(n15094), .B2(n15084), .ZN(
        n15091) );
  INV_X1 U18267 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15089) );
  AND2_X1 U18268 ( .A1(n15086), .A2(n15085), .ZN(n15088) );
  OR2_X1 U18269 ( .A1(n15088), .A2(n15087), .ZN(n19202) );
  OAI22_X1 U18270 ( .A1(n15101), .A2(n15089), .B1(n19400), .B2(n19202), .ZN(
        n15090) );
  AOI211_X1 U18271 ( .C1(n19398), .C2(BUF2_REG_19__SCAN_IN), .A(n15091), .B(
        n15090), .ZN(n15092) );
  OAI21_X1 U18272 ( .B1(n15093), .B2(n19422), .A(n15092), .ZN(P2_U2900) );
  OAI22_X1 U18273 ( .A1(n15096), .A2(n15095), .B1(n15094), .B2(n21333), .ZN(
        n15103) );
  OR2_X1 U18274 ( .A1(n15512), .A2(n15097), .ZN(n15098) );
  NAND2_X1 U18275 ( .A1(n15099), .A2(n15098), .ZN(n19215) );
  OAI22_X1 U18276 ( .A1(n15101), .A2(n15100), .B1(n19400), .B2(n19215), .ZN(
        n15102) );
  AOI211_X1 U18277 ( .C1(n19398), .C2(BUF2_REG_17__SCAN_IN), .A(n15103), .B(
        n15102), .ZN(n15104) );
  OAI21_X1 U18278 ( .B1(n15105), .B2(n19422), .A(n15104), .ZN(P2_U2902) );
  INV_X1 U18279 ( .A(n15106), .ZN(n15107) );
  OAI22_X1 U18280 ( .A1(n15109), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15107), .ZN(n15112) );
  NAND2_X1 U18281 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  OAI211_X1 U18282 ( .C1(n15113), .C2(n15112), .A(n15111), .B(n15110), .ZN(
        n15144) );
  XNOR2_X1 U18283 ( .A(n15115), .B(n15114), .ZN(n15118) );
  OAI21_X1 U18284 ( .B1(n15118), .B2(n15119), .A(n15357), .ZN(n15142) );
  NAND2_X1 U18285 ( .A1(n15144), .A2(n15142), .ZN(n15132) );
  AOI21_X1 U18286 ( .B1(n15117), .B2(n15120), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15135) );
  INV_X1 U18287 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U18288 ( .A1(n15119), .A2(n15333), .ZN(n15116) );
  NAND2_X1 U18289 ( .A1(n15117), .A2(n15116), .ZN(n15133) );
  INV_X1 U18290 ( .A(n15118), .ZN(n16426) );
  NAND3_X1 U18291 ( .A1(n16426), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15120), .ZN(n15143) );
  OAI211_X1 U18292 ( .C1(n15132), .C2(n15135), .A(n15133), .B(n15143), .ZN(
        n15124) );
  NAND2_X1 U18293 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  XNOR2_X1 U18294 ( .A(n15122), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15123) );
  XNOR2_X1 U18295 ( .A(n15124), .B(n15123), .ZN(n15341) );
  XNOR2_X1 U18296 ( .A(n15125), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15338) );
  NOR2_X1 U18297 ( .A1(n19305), .A2(n20093), .ZN(n15329) );
  NOR2_X1 U18298 ( .A1(n16554), .A2(n15126), .ZN(n15127) );
  AOI211_X1 U18299 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16546), .A(
        n15329), .B(n15127), .ZN(n15128) );
  OAI21_X1 U18300 ( .B1(n15341), .B2(n16557), .A(n15131), .ZN(P2_U2983) );
  NAND2_X1 U18301 ( .A1(n15132), .A2(n15143), .ZN(n15137) );
  INV_X1 U18302 ( .A(n15133), .ZN(n15134) );
  NOR2_X1 U18303 ( .A1(n15135), .A2(n15134), .ZN(n15136) );
  XOR2_X1 U18304 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15146), .Z(
        n15352) );
  NOR2_X1 U18305 ( .A1(n19305), .A2(n15138), .ZN(n15346) );
  NOR2_X1 U18306 ( .A1(n16554), .A2(n15139), .ZN(n15140) );
  AOI211_X1 U18307 ( .C1(n16546), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15346), .B(n15140), .ZN(n15141) );
  NAND2_X1 U18308 ( .A1(n15143), .A2(n15142), .ZN(n15145) );
  XOR2_X1 U18309 ( .A(n15145), .B(n15144), .Z(n15367) );
  AOI21_X1 U18310 ( .B1(n15357), .B2(n15147), .A(n15146), .ZN(n15365) );
  NOR2_X1 U18311 ( .A1(n15303), .A2(n20089), .ZN(n15360) );
  NOR2_X1 U18312 ( .A1(n16565), .A2(n16423), .ZN(n15148) );
  AOI211_X1 U18313 ( .C1(n16420), .C2(n16555), .A(n15360), .B(n15148), .ZN(
        n15149) );
  OAI21_X1 U18314 ( .B1(n16428), .B2(n13882), .A(n15149), .ZN(n15150) );
  AOI21_X1 U18315 ( .B1(n15365), .B2(n16550), .A(n15150), .ZN(n15151) );
  OAI21_X1 U18316 ( .B1(n15367), .B2(n16557), .A(n15151), .ZN(P2_U2985) );
  INV_X1 U18317 ( .A(n15152), .ZN(n15153) );
  OAI21_X1 U18318 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15163), .A(
        n15153), .ZN(n15378) );
  OR2_X1 U18319 ( .A1(n15154), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15368) );
  NAND3_X1 U18320 ( .A1(n15368), .A2(n15155), .A3(n16549), .ZN(n15159) );
  OR2_X1 U18321 ( .A1(n15303), .A2(n20087), .ZN(n15372) );
  OAI21_X1 U18322 ( .B1(n16565), .B2(n21232), .A(n15372), .ZN(n15157) );
  NOR2_X1 U18323 ( .A1(n16444), .A2(n13882), .ZN(n15156) );
  AOI211_X1 U18324 ( .C1(n16555), .C2(n16435), .A(n15157), .B(n15156), .ZN(
        n15158) );
  OAI211_X1 U18325 ( .C1(n16558), .C2(n15378), .A(n15159), .B(n15158), .ZN(
        P2_U2987) );
  NOR2_X1 U18326 ( .A1(n15160), .A2(n15170), .ZN(n15161) );
  XOR2_X1 U18327 ( .A(n15162), .B(n15161), .Z(n15389) );
  INV_X1 U18328 ( .A(n15174), .ZN(n15164) );
  AOI21_X1 U18329 ( .B1(n10036), .B2(n15164), .A(n15163), .ZN(n15387) );
  NOR2_X1 U18330 ( .A1(n19305), .A2(n16453), .ZN(n15383) );
  NOR2_X1 U18331 ( .A1(n16554), .A2(n15165), .ZN(n15166) );
  AOI211_X1 U18332 ( .C1(n16546), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15383), .B(n15166), .ZN(n15167) );
  OAI21_X1 U18333 ( .B1(n16459), .B2(n13882), .A(n15167), .ZN(n15168) );
  AOI21_X1 U18334 ( .B1(n15387), .B2(n16550), .A(n15168), .ZN(n15169) );
  OAI21_X1 U18335 ( .B1(n15389), .B2(n16557), .A(n15169), .ZN(P2_U2988) );
  NOR2_X1 U18336 ( .A1(n15171), .A2(n15170), .ZN(n15173) );
  XOR2_X1 U18337 ( .A(n15173), .B(n15172), .Z(n15401) );
  AOI21_X1 U18338 ( .B1(n15397), .B2(n15185), .A(n15174), .ZN(n15399) );
  NAND2_X1 U18339 ( .A1(n19326), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15392) );
  OAI21_X1 U18340 ( .B1(n16565), .B2(n15175), .A(n15392), .ZN(n15176) );
  AOI21_X1 U18341 ( .B1(n16555), .B2(n15177), .A(n15176), .ZN(n15178) );
  OAI21_X1 U18342 ( .B1(n15390), .B2(n13882), .A(n15178), .ZN(n15179) );
  AOI21_X1 U18343 ( .B1(n15399), .B2(n16550), .A(n15179), .ZN(n15180) );
  OAI21_X1 U18344 ( .B1(n15401), .B2(n16557), .A(n15180), .ZN(P2_U2989) );
  XOR2_X1 U18345 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15181), .Z(
        n15182) );
  XNOR2_X1 U18346 ( .A(n15183), .B(n15182), .ZN(n15411) );
  INV_X1 U18347 ( .A(n15424), .ZN(n15184) );
  NAND2_X1 U18348 ( .A1(n15184), .A2(n15402), .ZN(n15192) );
  INV_X1 U18349 ( .A(n15185), .ZN(n15186) );
  AOI21_X1 U18350 ( .B1(n21149), .B2(n15192), .A(n15186), .ZN(n15409) );
  NOR2_X1 U18351 ( .A1(n15303), .A2(n20082), .ZN(n15404) );
  NOR2_X1 U18352 ( .A1(n16554), .A2(n15187), .ZN(n15188) );
  AOI211_X1 U18353 ( .C1(n16546), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15404), .B(n15188), .ZN(n15189) );
  OAI21_X1 U18354 ( .B1(n16469), .B2(n13882), .A(n15189), .ZN(n15190) );
  AOI21_X1 U18355 ( .B1(n15409), .B2(n16550), .A(n15190), .ZN(n15191) );
  OAI21_X1 U18356 ( .B1(n15411), .B2(n16557), .A(n15191), .ZN(P2_U2990) );
  NOR2_X1 U18357 ( .A1(n15424), .A2(n15430), .ZN(n15193) );
  OAI21_X1 U18358 ( .B1(n15193), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15192), .ZN(n15423) );
  XOR2_X1 U18359 ( .A(n15195), .B(n15194), .Z(n15412) );
  NAND2_X1 U18360 ( .A1(n15412), .A2(n16549), .ZN(n15201) );
  OAI22_X1 U18361 ( .A1(n16565), .A2(n15196), .B1(n12232), .B2(n15303), .ZN(
        n15198) );
  NOR2_X1 U18362 ( .A1(n16481), .A2(n13882), .ZN(n15197) );
  AOI211_X1 U18363 ( .C1(n16555), .C2(n15199), .A(n15198), .B(n15197), .ZN(
        n15200) );
  OAI211_X1 U18364 ( .C1(n16558), .C2(n15423), .A(n15201), .B(n15200), .ZN(
        P2_U2991) );
  NAND2_X1 U18365 ( .A1(n15622), .A2(n15477), .ZN(n15257) );
  NAND2_X1 U18366 ( .A1(n15245), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15471) );
  OAI21_X1 U18367 ( .B1(n15471), .B2(n15202), .A(n15442), .ZN(n15203) );
  NAND2_X1 U18368 ( .A1(n15203), .A2(n15424), .ZN(n15452) );
  NAND2_X1 U18369 ( .A1(n15205), .A2(n15204), .ZN(n15214) );
  INV_X1 U18370 ( .A(n15536), .ZN(n15206) );
  INV_X1 U18371 ( .A(n15273), .ZN(n15207) );
  INV_X1 U18372 ( .A(n15261), .ZN(n15209) );
  OAI21_X1 U18373 ( .B1(n15262), .B2(n15209), .A(n15208), .ZN(n15252) );
  NAND2_X1 U18374 ( .A1(n15211), .A2(n15210), .ZN(n15253) );
  INV_X1 U18375 ( .A(n15231), .ZN(n15212) );
  INV_X1 U18376 ( .A(n15242), .ZN(n15233) );
  NAND2_X1 U18377 ( .A1(n15440), .A2(n16549), .ZN(n15220) );
  NAND2_X1 U18378 ( .A1(n19326), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15445) );
  OAI21_X1 U18379 ( .B1(n16565), .B2(n15215), .A(n15445), .ZN(n15217) );
  NOR2_X1 U18380 ( .A1(n15441), .A2(n13882), .ZN(n15216) );
  AOI211_X1 U18381 ( .C1(n16555), .C2(n15218), .A(n15217), .B(n15216), .ZN(
        n15219) );
  OAI211_X1 U18382 ( .C1(n16558), .C2(n15452), .A(n15220), .B(n15219), .ZN(
        P2_U2993) );
  NAND2_X1 U18383 ( .A1(n15222), .A2(n15221), .ZN(n15224) );
  XOR2_X1 U18384 ( .A(n15224), .B(n15223), .Z(n15464) );
  XNOR2_X1 U18385 ( .A(n15471), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15462) );
  NOR2_X1 U18386 ( .A1(n15303), .A2(n15225), .ZN(n15458) );
  NOR2_X1 U18387 ( .A1(n16554), .A2(n15226), .ZN(n15227) );
  AOI211_X1 U18388 ( .C1(n16546), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15458), .B(n15227), .ZN(n15228) );
  OAI21_X1 U18389 ( .B1(n16489), .B2(n13882), .A(n15228), .ZN(n15229) );
  AOI21_X1 U18390 ( .B1(n15462), .B2(n16550), .A(n15229), .ZN(n15230) );
  OAI21_X1 U18391 ( .B1(n15464), .B2(n16557), .A(n15230), .ZN(P2_U2994) );
  NAND2_X1 U18392 ( .A1(n15232), .A2(n15231), .ZN(n15235) );
  AOI21_X1 U18393 ( .B1(n15244), .B2(n15241), .A(n15233), .ZN(n15234) );
  XOR2_X1 U18394 ( .A(n15235), .B(n15234), .Z(n15475) );
  NAND2_X1 U18395 ( .A1(n19326), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15467) );
  OAI21_X1 U18396 ( .B1(n16565), .B2(n19191), .A(n15467), .ZN(n15237) );
  NOR2_X1 U18397 ( .A1(n19194), .A2(n13882), .ZN(n15236) );
  AOI211_X1 U18398 ( .C1(n16555), .C2(n19196), .A(n15237), .B(n15236), .ZN(
        n15240) );
  INV_X1 U18399 ( .A(n15245), .ZN(n15238) );
  NAND2_X1 U18400 ( .A1(n15238), .A2(n15455), .ZN(n15472) );
  NAND3_X1 U18401 ( .A1(n15472), .A2(n16550), .A3(n15471), .ZN(n15239) );
  OAI211_X1 U18402 ( .C1(n15475), .C2(n16557), .A(n15240), .B(n15239), .ZN(
        P2_U2995) );
  NAND2_X1 U18403 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  XNOR2_X1 U18404 ( .A(n15244), .B(n15243), .ZN(n15486) );
  AOI21_X1 U18405 ( .B1(n15246), .B2(n15257), .A(n15245), .ZN(n15484) );
  NOR2_X1 U18406 ( .A1(n15303), .A2(n20075), .ZN(n15480) );
  NOR2_X1 U18407 ( .A1(n16554), .A2(n15247), .ZN(n15248) );
  AOI211_X1 U18408 ( .C1(n16546), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15480), .B(n15248), .ZN(n15249) );
  OAI21_X1 U18409 ( .B1(n16492), .B2(n13882), .A(n15249), .ZN(n15250) );
  AOI21_X1 U18410 ( .B1(n15484), .B2(n16550), .A(n15250), .ZN(n15251) );
  OAI21_X1 U18411 ( .B1(n15486), .B2(n16557), .A(n15251), .ZN(P2_U2996) );
  XOR2_X1 U18412 ( .A(n15253), .B(n15252), .Z(n15507) );
  NOR2_X1 U18413 ( .A1(n15303), .A2(n20073), .ZN(n15487) );
  AOI21_X1 U18414 ( .B1(n16546), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15487), .ZN(n15254) );
  OAI21_X1 U18415 ( .B1(n16554), .B2(n15255), .A(n15254), .ZN(n15256) );
  AOI21_X1 U18416 ( .B1(n19210), .B2(n16561), .A(n15256), .ZN(n15259) );
  NAND2_X1 U18417 ( .A1(n15622), .A2(n15490), .ZN(n15489) );
  NOR2_X1 U18418 ( .A1(n15260), .A2(n21194), .ZN(n15496) );
  OAI211_X1 U18419 ( .C1(n15496), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16550), .B(n15257), .ZN(n15258) );
  OAI211_X1 U18420 ( .C1(n15507), .C2(n16557), .A(n15259), .B(n15258), .ZN(
        P2_U2997) );
  XOR2_X1 U18421 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n15260), .Z(
        n15272) );
  XNOR2_X1 U18422 ( .A(n15262), .B(n15261), .ZN(n15508) );
  NAND2_X1 U18423 ( .A1(n15508), .A2(n16549), .ZN(n15271) );
  OR2_X1 U18424 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  NAND2_X1 U18425 ( .A1(n15266), .A2(n15265), .ZN(n19359) );
  INV_X1 U18426 ( .A(n19359), .ZN(n15269) );
  NOR2_X1 U18427 ( .A1(n15513), .A2(n19305), .ZN(n15268) );
  OAI22_X1 U18428 ( .A1(n16565), .A2(n10301), .B1(n16554), .B2(n19217), .ZN(
        n15267) );
  AOI211_X1 U18429 ( .C1(n16561), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15270) );
  OAI211_X1 U18430 ( .C1(n16558), .C2(n15272), .A(n15271), .B(n15270), .ZN(
        P2_U2998) );
  NAND2_X1 U18431 ( .A1(n15274), .A2(n15273), .ZN(n15276) );
  XOR2_X1 U18432 ( .A(n15276), .B(n15275), .Z(n15532) );
  XNOR2_X1 U18433 ( .A(n15489), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15530) );
  INV_X1 U18434 ( .A(n15277), .ZN(n19228) );
  OAI22_X1 U18435 ( .A1(n16565), .A2(n15278), .B1(n16554), .B2(n19228), .ZN(
        n15281) );
  OAI22_X1 U18436 ( .A1(n19233), .A2(n13882), .B1(n15279), .B2(n15303), .ZN(
        n15280) );
  AOI211_X1 U18437 ( .C1(n15530), .C2(n16550), .A(n15281), .B(n15280), .ZN(
        n15282) );
  OAI21_X1 U18438 ( .B1(n15532), .B2(n16557), .A(n15282), .ZN(P2_U2999) );
  NAND2_X1 U18439 ( .A1(n15587), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15309) );
  XNOR2_X1 U18440 ( .A(n15533), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15563) );
  NAND2_X1 U18441 ( .A1(n15284), .A2(n15283), .ZN(n15287) );
  NAND2_X1 U18442 ( .A1(n15285), .A2(n15295), .ZN(n15286) );
  XOR2_X1 U18443 ( .A(n15287), .B(n15286), .Z(n15560) );
  NOR2_X1 U18444 ( .A1(n15303), .A2(n15288), .ZN(n15551) );
  NOR2_X1 U18445 ( .A1(n16565), .A2(n15289), .ZN(n15290) );
  AOI211_X1 U18446 ( .C1(n9874), .C2(n16555), .A(n15551), .B(n15290), .ZN(
        n15291) );
  OAI21_X1 U18447 ( .B1(n13882), .B2(n19243), .A(n15291), .ZN(n15292) );
  AOI21_X1 U18448 ( .B1(n15560), .B2(n16549), .A(n15292), .ZN(n15293) );
  OAI21_X1 U18449 ( .B1(n15563), .B2(n16558), .A(n15293), .ZN(P2_U3001) );
  NAND2_X1 U18450 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  XNOR2_X1 U18451 ( .A(n15297), .B(n15296), .ZN(n15575) );
  NAND2_X1 U18452 ( .A1(n15309), .A2(n15298), .ZN(n15564) );
  NAND3_X1 U18453 ( .A1(n10034), .A2(n16550), .A3(n15564), .ZN(n15308) );
  INV_X1 U18454 ( .A(n19254), .ZN(n15306) );
  OR2_X1 U18455 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  NAND2_X1 U18456 ( .A1(n15302), .A2(n15301), .ZN(n19371) );
  NOR2_X1 U18457 ( .A1(n15303), .A2(n20066), .ZN(n15566) );
  AOI21_X1 U18458 ( .B1(n16546), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15566), .ZN(n15304) );
  OAI21_X1 U18459 ( .B1(n13882), .B2(n19371), .A(n15304), .ZN(n15305) );
  AOI21_X1 U18460 ( .B1(n16555), .B2(n15306), .A(n15305), .ZN(n15307) );
  OAI211_X1 U18461 ( .C1(n16557), .C2(n15575), .A(n15308), .B(n15307), .ZN(
        P2_U3002) );
  OAI21_X1 U18462 ( .B1(n15587), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15309), .ZN(n15586) );
  XOR2_X1 U18463 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15310), .Z(
        n15311) );
  XNOR2_X1 U18464 ( .A(n15312), .B(n15311), .ZN(n15584) );
  NOR2_X1 U18465 ( .A1(n19305), .A2(n15313), .ZN(n15579) );
  NOR2_X1 U18466 ( .A1(n16565), .A2(n19263), .ZN(n15314) );
  AOI211_X1 U18467 ( .C1(n19266), .C2(n16555), .A(n15579), .B(n15314), .ZN(
        n15315) );
  OAI21_X1 U18468 ( .B1(n13882), .B2(n15577), .A(n15315), .ZN(n15316) );
  AOI21_X1 U18469 ( .B1(n15584), .B2(n16549), .A(n15316), .ZN(n15317) );
  OAI21_X1 U18470 ( .B1(n15586), .B2(n16558), .A(n15317), .ZN(P2_U3003) );
  XNOR2_X1 U18471 ( .A(n15318), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15319) );
  XNOR2_X1 U18472 ( .A(n15320), .B(n15319), .ZN(n15641) );
  NAND2_X1 U18473 ( .A1(n15321), .A2(n15322), .ZN(n16534) );
  INV_X1 U18474 ( .A(n16534), .ZN(n15324) );
  AOI21_X1 U18475 ( .B1(n16533), .B2(n15322), .A(n15321), .ZN(n15323) );
  AOI21_X1 U18476 ( .B1(n15324), .B2(n16533), .A(n15323), .ZN(n15639) );
  OAI22_X1 U18477 ( .A1(n16565), .A2(n21274), .B1(n20057), .B2(n15303), .ZN(
        n15327) );
  INV_X1 U18478 ( .A(n19295), .ZN(n15325) );
  OAI22_X1 U18479 ( .A1(n13882), .A2(n19299), .B1(n16554), .B2(n15325), .ZN(
        n15326) );
  AOI211_X1 U18480 ( .C1(n15639), .C2(n16549), .A(n15327), .B(n15326), .ZN(
        n15328) );
  OAI21_X1 U18481 ( .B1(n15641), .B2(n16558), .A(n15328), .ZN(P2_U3007) );
  INV_X1 U18482 ( .A(n15329), .ZN(n15331) );
  NOR2_X1 U18483 ( .A1(n15357), .A2(n15358), .ZN(n15356) );
  NAND4_X1 U18484 ( .A1(n15370), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15356), .A4(n15335), .ZN(n15330) );
  OAI211_X1 U18485 ( .C1(n16581), .C2(n19390), .A(n15331), .B(n15330), .ZN(
        n15332) );
  INV_X1 U18486 ( .A(n15332), .ZN(n15336) );
  INV_X1 U18487 ( .A(n15356), .ZN(n15334) );
  AOI211_X1 U18488 ( .C1(n15498), .C2(n15334), .A(n15333), .B(n15375), .ZN(
        n15345) );
  INV_X1 U18489 ( .A(n15337), .ZN(n15340) );
  NAND2_X1 U18490 ( .A1(n15338), .A2(n16574), .ZN(n15339) );
  OAI211_X1 U18491 ( .C1(n15341), .C2(n15632), .A(n15340), .B(n15339), .ZN(
        P2_U3015) );
  AOI21_X1 U18492 ( .B1(n15370), .B2(n15356), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15344) );
  OR2_X1 U18493 ( .A1(n15345), .A2(n15344), .ZN(n15348) );
  INV_X1 U18494 ( .A(n15346), .ZN(n15347) );
  AOI21_X1 U18495 ( .B1(n15352), .B2(n16574), .A(n15351), .ZN(n15353) );
  OAI21_X1 U18496 ( .B1(n15354), .B2(n15632), .A(n15353), .ZN(P2_U3016) );
  NAND2_X1 U18497 ( .A1(n15375), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15363) );
  INV_X1 U18498 ( .A(n15370), .ZN(n15355) );
  AOI211_X1 U18499 ( .C1(n15358), .C2(n15357), .A(n15356), .B(n15355), .ZN(
        n15359) );
  AOI211_X1 U18500 ( .C1(n15602), .C2(n15361), .A(n15360), .B(n15359), .ZN(
        n15362) );
  OAI211_X1 U18501 ( .C1(n16428), .C2(n15600), .A(n15363), .B(n15362), .ZN(
        n15364) );
  AOI21_X1 U18502 ( .B1(n15365), .B2(n16574), .A(n15364), .ZN(n15366) );
  OAI21_X1 U18503 ( .B1(n15367), .B2(n15632), .A(n15366), .ZN(P2_U3017) );
  NAND3_X1 U18504 ( .A1(n15368), .A2(n15155), .A3(n16592), .ZN(n15377) );
  NOR2_X1 U18505 ( .A1(n16444), .A2(n15600), .ZN(n15374) );
  NAND2_X1 U18506 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  OAI211_X1 U18507 ( .C1(n16581), .C2(n16448), .A(n15372), .B(n15371), .ZN(
        n15373) );
  AOI211_X1 U18508 ( .C1(n15375), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15374), .B(n15373), .ZN(n15376) );
  OAI211_X1 U18509 ( .C1(n15378), .C2(n16588), .A(n15377), .B(n15376), .ZN(
        P2_U3019) );
  OR2_X1 U18510 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15391) );
  AOI21_X1 U18511 ( .B1(n15407), .B2(n15391), .A(n10036), .ZN(n15386) );
  INV_X1 U18512 ( .A(n15380), .ZN(n16462) );
  NOR4_X1 U18513 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15397), .A4(n15381), .ZN(n15382) );
  AOI211_X1 U18514 ( .C1(n15602), .C2(n16462), .A(n15383), .B(n15382), .ZN(
        n15384) );
  OAI21_X1 U18515 ( .B1(n16459), .B2(n15600), .A(n15384), .ZN(n15385) );
  AOI211_X1 U18516 ( .C1(n15387), .C2(n16574), .A(n15386), .B(n15385), .ZN(
        n15388) );
  OAI21_X1 U18517 ( .B1(n15389), .B2(n15632), .A(n15388), .ZN(P2_U3020) );
  INV_X1 U18518 ( .A(n15390), .ZN(n15395) );
  OAI211_X1 U18519 ( .C1(n16581), .C2(n15393), .A(n15392), .B(n15391), .ZN(
        n15394) );
  AOI21_X1 U18520 ( .B1(n15395), .B2(n16586), .A(n15394), .ZN(n15396) );
  OAI21_X1 U18521 ( .B1(n15407), .B2(n15397), .A(n15396), .ZN(n15398) );
  AOI21_X1 U18522 ( .B1(n15399), .B2(n16574), .A(n15398), .ZN(n15400) );
  OAI21_X1 U18523 ( .B1(n15401), .B2(n15632), .A(n15400), .ZN(P2_U3021) );
  INV_X1 U18524 ( .A(n15417), .ZN(n15431) );
  AOI21_X1 U18525 ( .B1(n15431), .B2(n15402), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15406) );
  NOR2_X1 U18526 ( .A1(n16469), .A2(n15600), .ZN(n15403) );
  AOI211_X1 U18527 ( .C1(n15602), .C2(n16478), .A(n15404), .B(n15403), .ZN(
        n15405) );
  OAI21_X1 U18528 ( .B1(n15407), .B2(n15406), .A(n15405), .ZN(n15408) );
  AOI21_X1 U18529 ( .B1(n15409), .B2(n16574), .A(n15408), .ZN(n15410) );
  OAI21_X1 U18530 ( .B1(n15411), .B2(n15632), .A(n15410), .ZN(P2_U3022) );
  NAND2_X1 U18531 ( .A1(n15412), .A2(n16592), .ZN(n15422) );
  XNOR2_X1 U18532 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15416) );
  NOR2_X1 U18533 ( .A1(n15611), .A2(n15413), .ZN(n15432) );
  NOR2_X1 U18534 ( .A1(n12232), .A2(n19305), .ZN(n15414) );
  AOI21_X1 U18535 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15432), .A(
        n15414), .ZN(n15415) );
  OAI21_X1 U18536 ( .B1(n15417), .B2(n15416), .A(n15415), .ZN(n15419) );
  NOR2_X1 U18537 ( .A1(n16481), .A2(n15600), .ZN(n15418) );
  AOI211_X1 U18538 ( .C1(n15602), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15421) );
  OAI211_X1 U18539 ( .C1(n15423), .C2(n16588), .A(n15422), .B(n15421), .ZN(
        P2_U3023) );
  XNOR2_X1 U18540 ( .A(n15424), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16507) );
  INV_X1 U18541 ( .A(n16507), .ZN(n15439) );
  INV_X1 U18542 ( .A(n15425), .ZN(n15427) );
  AND2_X1 U18543 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  XNOR2_X1 U18544 ( .A(n15429), .B(n15428), .ZN(n16506) );
  NOR2_X1 U18545 ( .A1(n12523), .A2(n19305), .ZN(n15434) );
  MUX2_X1 U18546 ( .A(n15432), .B(n15431), .S(n15430), .Z(n15433) );
  AOI211_X1 U18547 ( .C1(n15602), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        n15436) );
  OAI21_X1 U18548 ( .B1(n16510), .B2(n15600), .A(n15436), .ZN(n15437) );
  AOI21_X1 U18549 ( .B1(n16506), .B2(n16592), .A(n15437), .ZN(n15438) );
  OAI21_X1 U18550 ( .B1(n16588), .B2(n15439), .A(n15438), .ZN(P2_U3024) );
  NAND2_X1 U18551 ( .A1(n15440), .A2(n16592), .ZN(n15451) );
  INV_X1 U18552 ( .A(n15629), .ZN(n15540) );
  OAI21_X1 U18553 ( .B1(n15443), .B2(n16583), .A(n15540), .ZN(n15449) );
  NOR2_X1 U18554 ( .A1(n15441), .A2(n15600), .ZN(n15448) );
  NAND3_X1 U18555 ( .A1(n15443), .A2(n15539), .A3(n15442), .ZN(n15444) );
  OAI211_X1 U18556 ( .C1(n16581), .C2(n15446), .A(n15445), .B(n15444), .ZN(
        n15447) );
  AOI211_X1 U18557 ( .C1(n15449), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15448), .B(n15447), .ZN(n15450) );
  OAI211_X1 U18558 ( .C1(n15452), .C2(n16588), .A(n15451), .B(n15450), .ZN(
        P2_U3025) );
  INV_X1 U18559 ( .A(n15456), .ZN(n15453) );
  OAI21_X1 U18560 ( .B1(n15453), .B2(n16583), .A(n15540), .ZN(n15470) );
  INV_X1 U18561 ( .A(n15539), .ZN(n15623) );
  NOR3_X1 U18562 ( .A1(n15456), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15623), .ZN(n15465) );
  OAI21_X1 U18563 ( .B1(n15470), .B2(n15465), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15460) );
  INV_X1 U18564 ( .A(n15454), .ZN(n16494) );
  NOR4_X1 U18565 ( .A1(n15456), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15455), .A4(n15623), .ZN(n15457) );
  AOI211_X1 U18566 ( .C1(n15602), .C2(n16494), .A(n15458), .B(n15457), .ZN(
        n15459) );
  OAI211_X1 U18567 ( .C1(n16489), .C2(n15600), .A(n15460), .B(n15459), .ZN(
        n15461) );
  AOI21_X1 U18568 ( .B1(n15462), .B2(n16574), .A(n15461), .ZN(n15463) );
  OAI21_X1 U18569 ( .B1(n15464), .B2(n15632), .A(n15463), .ZN(P2_U3026) );
  NOR2_X1 U18570 ( .A1(n19194), .A2(n15600), .ZN(n15469) );
  INV_X1 U18571 ( .A(n15465), .ZN(n15466) );
  OAI211_X1 U18572 ( .C1(n16581), .C2(n19202), .A(n15467), .B(n15466), .ZN(
        n15468) );
  AOI211_X1 U18573 ( .C1(n15470), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15469), .B(n15468), .ZN(n15474) );
  NAND3_X1 U18574 ( .A1(n15472), .A2(n16574), .A3(n15471), .ZN(n15473) );
  OAI211_X1 U18575 ( .C1(n15475), .C2(n15632), .A(n15474), .B(n15473), .ZN(
        P2_U3027) );
  OAI21_X1 U18576 ( .B1(n15477), .B2(n16583), .A(n15540), .ZN(n15476) );
  NAND2_X1 U18577 ( .A1(n15476), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15482) );
  INV_X1 U18578 ( .A(n15477), .ZN(n15478) );
  NOR3_X1 U18579 ( .A1(n15478), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15623), .ZN(n15479) );
  AOI211_X1 U18580 ( .C1(n15602), .C2(n16500), .A(n15480), .B(n15479), .ZN(
        n15481) );
  OAI211_X1 U18581 ( .C1(n16492), .C2(n15600), .A(n15482), .B(n15481), .ZN(
        n15483) );
  AOI21_X1 U18582 ( .B1(n15484), .B2(n16574), .A(n15483), .ZN(n15485) );
  OAI21_X1 U18583 ( .B1(n15486), .B2(n15632), .A(n15485), .ZN(P2_U3028) );
  INV_X1 U18584 ( .A(n15487), .ZN(n15488) );
  OAI21_X1 U18585 ( .B1(n16581), .B2(n19215), .A(n15488), .ZN(n15493) );
  INV_X1 U18586 ( .A(n15489), .ZN(n15534) );
  INV_X1 U18587 ( .A(n15490), .ZN(n15497) );
  NOR2_X1 U18588 ( .A1(n15497), .A2(n15623), .ZN(n15526) );
  AOI21_X1 U18589 ( .B1(n15534), .B2(n16574), .A(n15526), .ZN(n15514) );
  NOR3_X1 U18590 ( .A1(n15514), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15491), .ZN(n15492) );
  AOI211_X1 U18591 ( .C1(n19210), .C2(n16586), .A(n15493), .B(n15492), .ZN(
        n15506) );
  NOR2_X1 U18592 ( .A1(n15494), .A2(n16574), .ZN(n15495) );
  OR2_X1 U18593 ( .A1(n15496), .A2(n15495), .ZN(n15503) );
  AND2_X1 U18594 ( .A1(n15498), .A2(n15497), .ZN(n15499) );
  OR2_X1 U18595 ( .A1(n15629), .A2(n15499), .ZN(n15522) );
  AND2_X1 U18596 ( .A1(n15500), .A2(n15525), .ZN(n15501) );
  NOR2_X1 U18597 ( .A1(n15522), .A2(n15501), .ZN(n15502) );
  NAND2_X1 U18598 ( .A1(n15503), .A2(n15502), .ZN(n15518) );
  NOR2_X1 U18599 ( .A1(n16583), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15504) );
  OAI21_X1 U18600 ( .B1(n15518), .B2(n15504), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15505) );
  OAI211_X1 U18601 ( .C1(n15507), .C2(n15632), .A(n15506), .B(n15505), .ZN(
        P2_U3029) );
  INV_X1 U18602 ( .A(n15508), .ZN(n15521) );
  NOR2_X1 U18603 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  OR2_X1 U18604 ( .A1(n15512), .A2(n15511), .ZN(n19399) );
  INV_X1 U18605 ( .A(n19399), .ZN(n15517) );
  OAI22_X1 U18606 ( .A1(n19359), .A2(n15600), .B1(n15513), .B2(n15303), .ZN(
        n15516) );
  NOR3_X1 U18607 ( .A1(n15514), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15525), .ZN(n15515) );
  AOI211_X1 U18608 ( .C1(n15602), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15520) );
  NAND2_X1 U18609 ( .A1(n15518), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15519) );
  OAI211_X1 U18610 ( .C1(n15521), .C2(n15632), .A(n15520), .B(n15519), .ZN(
        P2_U3030) );
  NAND2_X1 U18611 ( .A1(n15522), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15528) );
  NOR2_X1 U18612 ( .A1(n15279), .A2(n19305), .ZN(n15524) );
  NOR2_X1 U18613 ( .A1(n19233), .A2(n15600), .ZN(n15523) );
  AOI211_X1 U18614 ( .C1(n15526), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        n15527) );
  OAI211_X1 U18615 ( .C1(n16581), .C2(n19232), .A(n15528), .B(n15527), .ZN(
        n15529) );
  AOI21_X1 U18616 ( .B1(n15530), .B2(n16574), .A(n15529), .ZN(n15531) );
  OAI21_X1 U18617 ( .B1(n15532), .B2(n15632), .A(n15531), .ZN(P2_U3031) );
  INV_X1 U18618 ( .A(n16515), .ZN(n15550) );
  AND2_X1 U18619 ( .A1(n15536), .A2(n15535), .ZN(n15537) );
  XNOR2_X1 U18620 ( .A(n15538), .B(n15537), .ZN(n16517) );
  NAND2_X1 U18621 ( .A1(n15541), .A2(n15539), .ZN(n15552) );
  OAI21_X1 U18622 ( .B1(n15541), .B2(n16583), .A(n15540), .ZN(n15572) );
  NOR2_X1 U18623 ( .A1(n15552), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15565) );
  NOR2_X1 U18624 ( .A1(n15572), .A2(n15565), .ZN(n15556) );
  OAI21_X1 U18625 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15552), .A(
        n15556), .ZN(n15546) );
  NAND2_X1 U18626 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15542) );
  NOR3_X1 U18627 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15542), .A3(
        n15552), .ZN(n15545) );
  NAND2_X1 U18628 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19326), .ZN(n15543) );
  OAI21_X1 U18629 ( .B1(n19365), .B2(n15600), .A(n15543), .ZN(n15544) );
  AOI211_X1 U18630 ( .C1(n15546), .C2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15545), .B(n15544), .ZN(n15547) );
  OAI21_X1 U18631 ( .B1(n16581), .B2(n19408), .A(n15547), .ZN(n15548) );
  AOI21_X1 U18632 ( .B1(n16517), .B2(n16592), .A(n15548), .ZN(n15549) );
  OAI21_X1 U18633 ( .B1(n15550), .B2(n16588), .A(n15549), .ZN(P2_U3032) );
  INV_X1 U18634 ( .A(n19244), .ZN(n15559) );
  INV_X1 U18635 ( .A(n15551), .ZN(n15555) );
  INV_X1 U18636 ( .A(n15552), .ZN(n15553) );
  NAND3_X1 U18637 ( .A1(n15553), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n21229), .ZN(n15554) );
  OAI211_X1 U18638 ( .C1(n15600), .C2(n19243), .A(n15555), .B(n15554), .ZN(
        n15558) );
  NOR2_X1 U18639 ( .A1(n15556), .A2(n21229), .ZN(n15557) );
  AOI211_X1 U18640 ( .C1(n15602), .C2(n15559), .A(n15558), .B(n15557), .ZN(
        n15562) );
  NAND2_X1 U18641 ( .A1(n15560), .A2(n16592), .ZN(n15561) );
  OAI211_X1 U18642 ( .C1(n15563), .C2(n16588), .A(n15562), .B(n15561), .ZN(
        P2_U3033) );
  NAND3_X1 U18643 ( .A1(n10034), .A2(n16574), .A3(n15564), .ZN(n15574) );
  NOR2_X1 U18644 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  OAI21_X1 U18645 ( .B1(n15600), .B2(n19371), .A(n15567), .ZN(n15571) );
  XNOR2_X1 U18646 ( .A(n15569), .B(n15568), .ZN(n19411) );
  NOR2_X1 U18647 ( .A1(n19411), .A2(n16581), .ZN(n15570) );
  AOI211_X1 U18648 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15572), .A(
        n15571), .B(n15570), .ZN(n15573) );
  OAI211_X1 U18649 ( .C1(n15575), .C2(n15632), .A(n15574), .B(n15573), .ZN(
        P2_U3034) );
  NOR2_X1 U18650 ( .A1(n15629), .A2(n15576), .ZN(n15612) );
  NOR3_X1 U18651 ( .A1(n15612), .A2(n15611), .A3(n12045), .ZN(n15583) );
  XNOR2_X1 U18652 ( .A(n15610), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15580) );
  NOR2_X1 U18653 ( .A1(n15576), .A2(n15623), .ZN(n15595) );
  NOR2_X1 U18654 ( .A1(n15600), .A2(n15577), .ZN(n15578) );
  AOI211_X1 U18655 ( .C1(n15580), .C2(n15595), .A(n15579), .B(n15578), .ZN(
        n15581) );
  OAI21_X1 U18656 ( .B1(n19272), .B2(n16581), .A(n15581), .ZN(n15582) );
  AOI211_X1 U18657 ( .C1(n15584), .C2(n16592), .A(n15583), .B(n15582), .ZN(
        n15585) );
  OAI21_X1 U18658 ( .B1(n15586), .B2(n16588), .A(n15585), .ZN(P2_U3035) );
  AOI21_X1 U18659 ( .B1(n15610), .B2(n15621), .A(n15587), .ZN(n16521) );
  NAND2_X1 U18660 ( .A1(n16521), .A2(n16574), .ZN(n15616) );
  AND2_X1 U18661 ( .A1(n15589), .A2(n15588), .ZN(n15591) );
  OR2_X1 U18662 ( .A1(n15591), .A2(n15590), .ZN(n19414) );
  INV_X1 U18663 ( .A(n19414), .ZN(n15603) );
  NAND2_X1 U18664 ( .A1(n15593), .A2(n15592), .ZN(n15594) );
  NAND2_X1 U18665 ( .A1(n9877), .A2(n15594), .ZN(n19378) );
  INV_X1 U18666 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20063) );
  NOR2_X1 U18667 ( .A1(n20063), .A2(n19305), .ZN(n15598) );
  INV_X1 U18668 ( .A(n15595), .ZN(n15596) );
  NOR2_X1 U18669 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15596), .ZN(
        n15597) );
  NOR2_X1 U18670 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  OAI21_X1 U18671 ( .B1(n15600), .B2(n19378), .A(n15599), .ZN(n15601) );
  AOI21_X1 U18672 ( .B1(n15603), .B2(n15602), .A(n15601), .ZN(n15615) );
  INV_X1 U18673 ( .A(n15604), .ZN(n15618) );
  OR2_X1 U18674 ( .A1(n15605), .A2(n15618), .ZN(n15609) );
  NAND2_X1 U18675 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  XNOR2_X1 U18676 ( .A(n15609), .B(n15608), .ZN(n16523) );
  NAND2_X1 U18677 ( .A1(n16523), .A2(n16592), .ZN(n15614) );
  OR3_X1 U18678 ( .A1(n15612), .A2(n15611), .A3(n15610), .ZN(n15613) );
  NAND4_X1 U18679 ( .A1(n15616), .A2(n15615), .A3(n15614), .A4(n15613), .ZN(
        P2_U3036) );
  OR2_X1 U18680 ( .A1(n15618), .A2(n15617), .ZN(n15619) );
  XNOR2_X1 U18681 ( .A(n15620), .B(n15619), .ZN(n16526) );
  OAI21_X1 U18682 ( .B1(n15622), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15621), .ZN(n16527) );
  OR2_X1 U18683 ( .A1(n16527), .A2(n16588), .ZN(n15631) );
  INV_X1 U18684 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20061) );
  NOR2_X1 U18685 ( .A1(n20061), .A2(n19305), .ZN(n15625) );
  NOR2_X1 U18686 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15623), .ZN(
        n15624) );
  NOR2_X1 U18687 ( .A1(n15625), .A2(n15624), .ZN(n15627) );
  NAND2_X1 U18688 ( .A1(n16586), .A2(n16529), .ZN(n15626) );
  OAI211_X1 U18689 ( .C1(n19289), .C2(n16581), .A(n15627), .B(n15626), .ZN(
        n15628) );
  AOI21_X1 U18690 ( .B1(n15629), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15628), .ZN(n15630) );
  OAI211_X1 U18691 ( .C1(n16526), .C2(n15632), .A(n15631), .B(n15630), .ZN(
        P2_U3037) );
  NOR2_X1 U18692 ( .A1(n16580), .A2(n16569), .ZN(n15638) );
  NOR2_X1 U18693 ( .A1(n20057), .A2(n19305), .ZN(n15634) );
  NOR2_X1 U18694 ( .A1(n19300), .A2(n16581), .ZN(n15633) );
  AOI211_X1 U18695 ( .C1(n16586), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        n15636) );
  OAI21_X1 U18696 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16567), .A(
        n15636), .ZN(n15637) );
  AOI211_X1 U18697 ( .C1(n15639), .C2(n16592), .A(n15638), .B(n15637), .ZN(
        n15640) );
  OAI21_X1 U18698 ( .B1(n15641), .B2(n16588), .A(n15640), .ZN(P2_U3039) );
  OAI21_X1 U18699 ( .B1(n15643), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15642), .ZN(n16547) );
  INV_X1 U18700 ( .A(n16580), .ZN(n15649) );
  NAND4_X1 U18701 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n15645), .A4(n15644), .ZN(
        n15647) );
  AOI22_X1 U18702 ( .A1(n16586), .A2(n19315), .B1(n19326), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15646) );
  OAI211_X1 U18703 ( .C1(n16581), .C2(n19319), .A(n15647), .B(n15646), .ZN(
        n15648) );
  AOI21_X1 U18704 ( .B1(n15649), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15648), .ZN(n15654) );
  INV_X1 U18705 ( .A(n15650), .ZN(n15651) );
  XNOR2_X1 U18706 ( .A(n15652), .B(n15651), .ZN(n16548) );
  NAND2_X1 U18707 ( .A1(n16548), .A2(n16592), .ZN(n15653) );
  OAI211_X1 U18708 ( .C1(n16547), .C2(n16588), .A(n15654), .B(n15653), .ZN(
        P2_U3040) );
  INV_X1 U18709 ( .A(n15655), .ZN(n16631) );
  OAI21_X1 U18710 ( .B1(n9751), .B2(n15659), .A(n15658), .ZN(n15678) );
  INV_X1 U18711 ( .A(n20021), .ZN(n20104) );
  INV_X1 U18712 ( .A(n15660), .ZN(n15693) );
  NOR2_X1 U18713 ( .A1(n11755), .A2(n15661), .ZN(n15662) );
  OAI22_X1 U18714 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n15686), .B1(
        n15663), .B2(n15662), .ZN(n15664) );
  AOI21_X1 U18715 ( .B1(n15665), .B2(n15693), .A(n15664), .ZN(n16601) );
  OAI222_X1 U18716 ( .A1(n16631), .A2(n20124), .B1(n10414), .B2(n15678), .C1(
        n20104), .C2(n16601), .ZN(n15666) );
  MUX2_X1 U18717 ( .A(n15666), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15826), .Z(P2_U3600) );
  INV_X1 U18718 ( .A(n16618), .ZN(n15667) );
  AND2_X1 U18719 ( .A1(n15667), .A2(n16620), .ZN(n15688) );
  INV_X1 U18720 ( .A(n11753), .ZN(n15668) );
  NAND2_X1 U18721 ( .A1(n15668), .A2(n16597), .ZN(n15684) );
  AND2_X1 U18722 ( .A1(n15681), .A2(n15684), .ZN(n15676) );
  NAND2_X1 U18723 ( .A1(n15670), .A2(n15669), .ZN(n15682) );
  NAND2_X1 U18724 ( .A1(n15682), .A2(n15676), .ZN(n15675) );
  INV_X1 U18725 ( .A(n15671), .ZN(n15672) );
  NAND3_X1 U18726 ( .A1(n15673), .A2(n15672), .A3(n15685), .ZN(n15674) );
  OAI211_X1 U18727 ( .C1(n15688), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        n15677) );
  INV_X1 U18728 ( .A(n15678), .ZN(n15679) );
  OAI222_X1 U18729 ( .A1(n16631), .A2(n20117), .B1(n20104), .B2(n16598), .C1(
        n15679), .C2(n10414), .ZN(n15680) );
  MUX2_X1 U18730 ( .A(n15680), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15826), .Z(P2_U3599) );
  NAND2_X1 U18731 ( .A1(n15682), .A2(n15681), .ZN(n15683) );
  OAI211_X1 U18732 ( .C1(n12142), .C2(n15686), .A(n15683), .B(n15684), .ZN(
        n15691) );
  INV_X1 U18733 ( .A(n15684), .ZN(n15687) );
  OAI22_X1 U18734 ( .A1(n15688), .A2(n15687), .B1(n15686), .B2(n15685), .ZN(
        n15690) );
  MUX2_X1 U18735 ( .A(n15691), .B(n15690), .S(n15689), .Z(n15692) );
  AOI211_X1 U18736 ( .C1(n9839), .C2(n15693), .A(n12789), .B(n15692), .ZN(
        n16605) );
  OAI22_X1 U18737 ( .A1(n19504), .A2(n16631), .B1(n16605), .B2(n20104), .ZN(
        n15694) );
  MUX2_X1 U18738 ( .A(n15694), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15826), .Z(P2_U3596) );
  INV_X1 U18739 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17212) );
  INV_X1 U18740 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17210) );
  INV_X1 U18741 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17213) );
  INV_X1 U18742 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17344) );
  INV_X1 U18743 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17345) );
  NAND2_X1 U18744 ( .A1(n18511), .A2(n17319), .ZN(n17332) );
  NAND2_X1 U18745 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17270), .ZN(n17256) );
  NAND2_X1 U18746 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17261), .ZN(n17248) );
  AOI22_X1 U18747 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15696) );
  OAI21_X1 U18748 ( .B1(n9878), .B2(n21348), .A(n15696), .ZN(n15705) );
  AOI22_X1 U18749 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18750 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15697) );
  OAI21_X1 U18751 ( .B1(n17427), .B2(n18814), .A(n15697), .ZN(n15701) );
  AOI22_X1 U18752 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U18753 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15698) );
  OAI211_X1 U18754 ( .C1(n13976), .C2(n17305), .A(n15699), .B(n15698), .ZN(
        n15700) );
  AOI211_X1 U18755 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15701), .B(n15700), .ZN(n15702) );
  OAI211_X1 U18756 ( .C1(n17230), .C2(n17313), .A(n15703), .B(n15702), .ZN(
        n15704) );
  AOI211_X1 U18757 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15705), .B(n15704), .ZN(n17253) );
  INV_X1 U18758 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15707) );
  AOI22_X1 U18759 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15706) );
  OAI21_X1 U18760 ( .B1(n9875), .B2(n15707), .A(n15706), .ZN(n15716) );
  AOI22_X1 U18761 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15714) );
  INV_X1 U18762 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n21163) );
  OAI22_X1 U18763 ( .A1(n17449), .A2(n21163), .B1(n17381), .B2(n21244), .ZN(
        n15712) );
  AOI22_X1 U18764 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U18765 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18766 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15708) );
  NAND3_X1 U18767 ( .A1(n15710), .A2(n15709), .A3(n15708), .ZN(n15711) );
  AOI211_X1 U18768 ( .C1(n9763), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n15712), .B(n15711), .ZN(n15713) );
  OAI211_X1 U18769 ( .C1(n17483), .C2(n21364), .A(n15714), .B(n15713), .ZN(
        n15715) );
  AOI211_X1 U18770 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15716), .B(n15715), .ZN(n17262) );
  INV_X1 U18771 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21175) );
  AOI22_X1 U18772 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15717) );
  OAI21_X1 U18773 ( .B1(n13975), .B2(n21175), .A(n15717), .ZN(n15727) );
  INV_X1 U18774 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18561) );
  AOI22_X1 U18775 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15725) );
  INV_X1 U18776 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18803) );
  AOI22_X1 U18777 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15719) );
  OAI21_X1 U18778 ( .B1(n17427), .B2(n18803), .A(n15719), .ZN(n15723) );
  INV_X1 U18779 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U18780 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U18781 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15720) );
  OAI211_X1 U18782 ( .C1(n13976), .C2(n17482), .A(n15721), .B(n15720), .ZN(
        n15722) );
  AOI211_X1 U18783 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15723), .B(n15722), .ZN(n15724) );
  OAI211_X1 U18784 ( .C1(n15718), .C2(n18561), .A(n15725), .B(n15724), .ZN(
        n15726) );
  AOI211_X1 U18785 ( .C1(n17349), .C2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n15727), .B(n15726), .ZN(n17272) );
  AOI22_X1 U18786 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15728) );
  OAI21_X1 U18787 ( .B1(n13975), .B2(n18724), .A(n15728), .ZN(n15738) );
  AOI22_X1 U18788 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15735) );
  INV_X1 U18789 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17235) );
  OAI22_X1 U18790 ( .A1(n15718), .A2(n17235), .B1(n17381), .B2(n17490), .ZN(
        n15733) );
  AOI22_X1 U18791 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15731) );
  AOI22_X1 U18792 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U18793 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15729) );
  NAND3_X1 U18794 ( .A1(n15731), .A2(n15730), .A3(n15729), .ZN(n15732) );
  AOI211_X1 U18795 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15733), .B(n15732), .ZN(n15734) );
  OAI211_X1 U18796 ( .C1(n9947), .C2(n15736), .A(n15735), .B(n15734), .ZN(
        n15737) );
  AOI211_X1 U18797 ( .C1(n9763), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15738), .B(n15737), .ZN(n17271) );
  NOR2_X1 U18798 ( .A1(n17272), .A2(n17271), .ZN(n17268) );
  INV_X1 U18799 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U18800 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17468), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n15843), .ZN(n15748) );
  INV_X1 U18801 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15884) );
  AOI22_X1 U18802 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9763), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17417), .ZN(n15740) );
  AOI22_X1 U18803 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n13988), .ZN(n15739) );
  OAI211_X1 U18804 ( .C1(n15884), .C2(n17473), .A(n15740), .B(n15739), .ZN(
        n15746) );
  AOI22_X1 U18805 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U18806 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n15877), .ZN(n15743) );
  AOI22_X1 U18807 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17433), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17453), .ZN(n15742) );
  NAND2_X1 U18808 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15741) );
  NAND4_X1 U18809 ( .A1(n15744), .A2(n15743), .A3(n15742), .A4(n15741), .ZN(
        n15745) );
  AOI211_X1 U18810 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n15746), .B(n15745), .ZN(n15747) );
  OAI211_X1 U18811 ( .C1(n13975), .C2(n17448), .A(n15748), .B(n15747), .ZN(
        n17267) );
  NAND2_X1 U18812 ( .A1(n17268), .A2(n17267), .ZN(n17266) );
  NOR2_X1 U18813 ( .A1(n17262), .A2(n17266), .ZN(n17259) );
  INV_X1 U18814 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U18815 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15758) );
  AOI22_X1 U18816 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18817 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15749) );
  OAI211_X1 U18818 ( .C1(n17427), .C2(n21166), .A(n15750), .B(n15749), .ZN(
        n15756) );
  AOI22_X1 U18819 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15754) );
  AOI22_X1 U18820 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U18821 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15752) );
  NAND2_X1 U18822 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15751) );
  NAND4_X1 U18823 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        n15755) );
  AOI211_X1 U18824 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15756), .B(n15755), .ZN(n15757) );
  OAI211_X1 U18825 ( .C1(n17381), .C2(n17322), .A(n15758), .B(n15757), .ZN(
        n17258) );
  NAND2_X1 U18826 ( .A1(n17259), .A2(n17258), .ZN(n17257) );
  NOR2_X1 U18827 ( .A1(n17253), .A2(n17257), .ZN(n15770) );
  AOI22_X1 U18828 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15768) );
  INV_X1 U18829 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U18830 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U18831 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17470), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15759) );
  OAI211_X1 U18832 ( .C1(n17473), .C2(n17297), .A(n15760), .B(n15759), .ZN(
        n15766) );
  AOI22_X1 U18833 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U18834 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U18835 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15875), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15762) );
  NAND2_X1 U18836 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n15761) );
  NAND4_X1 U18837 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15765) );
  AOI211_X1 U18838 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15766), .B(n15765), .ZN(n15767) );
  OAI211_X1 U18839 ( .C1(n13975), .C2(n15773), .A(n15768), .B(n15767), .ZN(
        n15769) );
  NAND2_X1 U18840 ( .A1(n15770), .A2(n15769), .ZN(n17249) );
  OAI21_X1 U18841 ( .B1(n15770), .B2(n15769), .A(n17249), .ZN(n17540) );
  NAND3_X1 U18842 ( .A1(n17248), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n17511), 
        .ZN(n15771) );
  OAI221_X1 U18843 ( .B1(n17248), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n17511), 
        .C2(n17540), .A(n15771), .ZN(P3_U2675) );
  AOI22_X1 U18844 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15772) );
  OAI21_X1 U18845 ( .B1(n17449), .B2(n15773), .A(n15772), .ZN(n15782) );
  INV_X1 U18846 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n21138) );
  AOI22_X1 U18847 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15780) );
  INV_X1 U18848 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U18849 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15774) );
  OAI21_X1 U18850 ( .B1(n17473), .B2(n17289), .A(n15774), .ZN(n15778) );
  INV_X1 U18851 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U18852 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U18853 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15775) );
  OAI211_X1 U18854 ( .C1(n13976), .C2(n17495), .A(n15776), .B(n15775), .ZN(
        n15777) );
  AOI211_X1 U18855 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15778), .B(n15777), .ZN(n15779) );
  OAI211_X1 U18856 ( .C1(n17230), .C2(n21138), .A(n15780), .B(n15779), .ZN(
        n15781) );
  AOI211_X1 U18857 ( .C1(n17469), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15782), .B(n15781), .ZN(n17611) );
  NOR2_X1 U18858 ( .A1(n17517), .A2(n9907), .ZN(n17378) );
  AOI22_X1 U18859 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17378), .B1(n17411), 
        .B2(n17393), .ZN(n15783) );
  OAI21_X1 U18860 ( .B1(n17611), .B2(n17511), .A(n15783), .ZN(P3_U2690) );
  INV_X1 U18861 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18956) );
  NAND2_X1 U18862 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18956), .ZN(n18465) );
  INV_X1 U18863 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18926) );
  NAND3_X1 U18864 ( .A1(n17381), .A2(n15824), .A3(n18926), .ZN(n18463) );
  NOR2_X1 U18865 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18463), .ZN(n15785) );
  NAND3_X1 U18866 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n19089)
         );
  NAND2_X1 U18867 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18462) );
  NOR2_X1 U18868 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18975) );
  INV_X1 U18869 ( .A(n18975), .ZN(n19145) );
  NAND2_X1 U18870 ( .A1(n18926), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19102) );
  AOI21_X1 U18871 ( .B1(n18462), .B2(n19145), .A(n19115), .ZN(n15784) );
  INV_X1 U18872 ( .A(n15784), .ZN(n18477) );
  OAI21_X1 U18873 ( .B1(n15785), .B2(n19089), .A(n18516), .ZN(n18473) );
  NAND2_X1 U18874 ( .A1(n18465), .A2(n18473), .ZN(n18467) );
  NOR2_X1 U18875 ( .A1(n18958), .A2(n18467), .ZN(n18469) );
  INV_X1 U18876 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19142) );
  INV_X1 U18877 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19091) );
  NAND3_X1 U18878 ( .A1(n19142), .A2(n19091), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18828) );
  INV_X1 U18879 ( .A(n18467), .ZN(n15786) );
  OAI211_X1 U18880 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(
        P3_STATEBS16_REG_SCAN_IN), .A(P3_STATE2_REG_1__SCAN_IN), .B(n19091), 
        .ZN(n18468) );
  AOI21_X1 U18881 ( .B1(n15786), .B2(n18468), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15787) );
  AOI21_X1 U18882 ( .B1(n18469), .B2(n18828), .A(n15787), .ZN(P3_U2864) );
  NOR2_X1 U18883 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19091), .ZN(n18478) );
  INV_X2 U18884 ( .A(n19155), .ZN(n19083) );
  NAND2_X2 U18885 ( .A1(n19083), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19076) );
  OAI211_X1 U18886 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19014), .B(n19076), .ZN(n19005) );
  INV_X1 U18887 ( .A(n19005), .ZN(n19140) );
  INV_X1 U18888 ( .A(n17523), .ZN(n18504) );
  NOR2_X1 U18889 ( .A1(n18504), .A2(n18499), .ZN(n15798) );
  OAI21_X1 U18890 ( .B1(n18511), .B2(n15798), .A(n15812), .ZN(n15789) );
  INV_X1 U18891 ( .A(n15803), .ZN(n18491) );
  NOR2_X1 U18892 ( .A1(n18511), .A2(n17666), .ZN(n15797) );
  NAND4_X1 U18893 ( .A1(n18495), .A2(n18491), .A3(n15798), .A4(n15797), .ZN(
        n15805) );
  INV_X1 U18894 ( .A(n15795), .ZN(n15791) );
  NAND2_X1 U18895 ( .A1(n18484), .A2(n17666), .ZN(n15945) );
  NAND2_X1 U18896 ( .A1(n18484), .A2(n18479), .ZN(n16076) );
  INV_X1 U18897 ( .A(n15797), .ZN(n15801) );
  AOI221_X1 U18898 ( .B1(n18499), .B2(n15815), .C1(n15812), .C2(n15815), .A(
        n15798), .ZN(n15800) );
  AOI211_X1 U18899 ( .C1(n18491), .C2(n15801), .A(n15800), .B(n15799), .ZN(
        n15802) );
  INV_X1 U18900 ( .A(n15802), .ZN(n15817) );
  NAND2_X1 U18901 ( .A1(n17527), .A2(n18504), .ZN(n18949) );
  AOI21_X1 U18902 ( .B1(n17625), .B2(n18949), .A(n15945), .ZN(n15816) );
  AOI21_X1 U18903 ( .B1(n19140), .B2(n17663), .A(n16075), .ZN(n15821) );
  XNOR2_X1 U18904 ( .A(n15807), .B(n15806), .ZN(n15810) );
  INV_X1 U18905 ( .A(n18921), .ZN(n15984) );
  NAND2_X1 U18906 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19151) );
  NAND2_X1 U18907 ( .A1(n15984), .A2(n19151), .ZN(n16078) );
  INV_X1 U18908 ( .A(n15811), .ZN(n15818) );
  AOI21_X1 U18909 ( .B1(n15812), .B2(n18949), .A(n15947), .ZN(n15814) );
  NAND3_X1 U18910 ( .A1(n15815), .A2(n15814), .A3(n15813), .ZN(n15943) );
  AOI211_X1 U18911 ( .C1(n15818), .C2(n15943), .A(n15817), .B(n15816), .ZN(
        n15990) );
  INV_X1 U18912 ( .A(n15819), .ZN(n15820) );
  OAI211_X1 U18913 ( .C1(n15821), .C2(n16078), .A(n15990), .B(n15820), .ZN(
        n18948) );
  INV_X1 U18914 ( .A(n18948), .ZN(n18961) );
  INV_X1 U18915 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18464) );
  OAI22_X1 U18916 ( .A1(n18961), .A2(n18985), .B1(n18464), .B2(n19089), .ZN(
        n15822) );
  INV_X1 U18917 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19100) );
  NAND2_X1 U18918 ( .A1(n19100), .A2(n19091), .ZN(n19103) );
  INV_X1 U18919 ( .A(n19103), .ZN(n19117) );
  AOI21_X1 U18920 ( .B1(n15824), .B2(n18926), .A(n15823), .ZN(n18973) );
  NAND3_X1 U18921 ( .A1(n19119), .A2(n19117), .A3(n18973), .ZN(n15825) );
  OAI21_X1 U18922 ( .B1(n19119), .B2(n18926), .A(n15825), .ZN(P3_U3284) );
  INV_X1 U18923 ( .A(n15826), .ZN(n15831) );
  INV_X1 U18924 ( .A(n16623), .ZN(n15827) );
  NOR4_X1 U18925 ( .A1(n12574), .A2(n15827), .A3(n20155), .A4(n20104), .ZN(
        n15828) );
  NAND2_X1 U18926 ( .A1(n15831), .A2(n15828), .ZN(n15829) );
  OAI21_X1 U18927 ( .B1(n15831), .B2(n15830), .A(n15829), .ZN(P2_U3595) );
  NAND2_X1 U18928 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18247) );
  INV_X1 U18929 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18231) );
  NOR2_X1 U18930 ( .A1(n18242), .A2(n18231), .ZN(n18220) );
  NAND3_X1 U18931 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18220), .ZN(n16001) );
  NOR2_X1 U18932 ( .A1(n18247), .A2(n16001), .ZN(n18203) );
  NAND2_X1 U18933 ( .A1(n18203), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18189) );
  INV_X1 U18934 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18195) );
  NOR2_X1 U18935 ( .A1(n18189), .A2(n18195), .ZN(n17828) );
  NAND2_X1 U18936 ( .A1(n17828), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18165) );
  INV_X1 U18937 ( .A(n18165), .ZN(n18167) );
  INV_X1 U18938 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18164) );
  INV_X1 U18939 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18151) );
  NOR2_X1 U18940 ( .A1(n18164), .A2(n18151), .ZN(n18142) );
  NAND2_X1 U18941 ( .A1(n18167), .A2(n18142), .ZN(n17794) );
  INV_X1 U18942 ( .A(n17794), .ZN(n16670) );
  INV_X1 U18943 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18291) );
  NAND2_X1 U18944 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18000) );
  INV_X1 U18945 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18001) );
  NOR2_X1 U18946 ( .A1(n18000), .A2(n18001), .ZN(n18341) );
  NAND2_X1 U18947 ( .A1(n18341), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17978) );
  AOI22_X1 U18948 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15832) );
  OAI21_X1 U18949 ( .B1(n15718), .B2(n17490), .A(n15832), .ZN(n15841) );
  AOI22_X1 U18950 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U18951 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15833) );
  OAI21_X1 U18952 ( .B1(n17473), .B2(n17235), .A(n15833), .ZN(n15837) );
  AOI22_X1 U18953 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15835) );
  AOI22_X1 U18954 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15834) );
  OAI211_X1 U18955 ( .C1(n13976), .C2(n21325), .A(n15835), .B(n15834), .ZN(
        n15836) );
  AOI211_X1 U18956 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n15837), .B(n15836), .ZN(n15838) );
  OAI211_X1 U18957 ( .C1(n17449), .C2(n18724), .A(n15839), .B(n15838), .ZN(
        n15840) );
  AOI211_X4 U18958 ( .C1(n17436), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15841), .B(n15840), .ZN(n18047) );
  AOI22_X1 U18959 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15842) );
  OAI21_X1 U18960 ( .B1(n15718), .B2(n17495), .A(n15842), .ZN(n15853) );
  INV_X1 U18961 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15851) );
  AOI22_X1 U18962 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15850) );
  OAI22_X1 U18963 ( .A1(n9873), .A2(n17297), .B1(n13975), .B2(n21138), .ZN(
        n15848) );
  AOI22_X1 U18964 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15846) );
  AOI22_X1 U18965 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15914), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U18966 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15844) );
  NAND3_X1 U18967 ( .A1(n15846), .A2(n15845), .A3(n15844), .ZN(n15847) );
  AOI211_X1 U18968 ( .C1(n15875), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n15848), .B(n15847), .ZN(n15849) );
  OAI211_X1 U18969 ( .C1(n17381), .C2(n15851), .A(n15850), .B(n15849), .ZN(
        n15852) );
  AOI211_X2 U18970 ( .C1(n17453), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15853), .B(n15852), .ZN(n15952) );
  AOI22_X1 U18971 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15854) );
  OAI21_X1 U18972 ( .B1(n9878), .B2(n21166), .A(n15854), .ZN(n15863) );
  AOI22_X1 U18973 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15861) );
  INV_X1 U18974 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17415) );
  INV_X1 U18975 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21247) );
  OAI22_X1 U18976 ( .A1(n17427), .A2(n17415), .B1(n9875), .B2(n21247), .ZN(
        n15859) );
  AOI22_X1 U18977 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15857) );
  AOI22_X1 U18978 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15856) );
  AOI22_X1 U18979 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15855) );
  NAND3_X1 U18980 ( .A1(n15857), .A2(n15856), .A3(n15855), .ZN(n15858) );
  AOI211_X1 U18981 ( .C1(n17468), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n15859), .B(n15858), .ZN(n15860) );
  OAI211_X1 U18982 ( .C1(n17483), .C2(n17322), .A(n15861), .B(n15860), .ZN(
        n15862) );
  INV_X1 U18983 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U18984 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15873) );
  INV_X1 U18985 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U18986 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15865) );
  AOI22_X1 U18987 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15864) );
  OAI211_X1 U18988 ( .C1(n17427), .C2(n17334), .A(n15865), .B(n15864), .ZN(
        n15871) );
  AOI22_X1 U18989 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15914), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15869) );
  AOI22_X1 U18990 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15868) );
  AOI22_X1 U18991 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15867) );
  NAND2_X1 U18992 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n15866) );
  NAND4_X1 U18993 ( .A1(n15869), .A2(n15868), .A3(n15867), .A4(n15866), .ZN(
        n15870) );
  AOI22_X1 U18994 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15874), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15876) );
  OAI21_X1 U18995 ( .B1(n9878), .B2(n21197), .A(n15876), .ZN(n15881) );
  AOI22_X1 U18996 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n15877), .ZN(n15879) );
  AOI22_X1 U18997 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17417), .ZN(n15878) );
  OAI211_X1 U18998 ( .C1(n17427), .C2(n17448), .A(n15879), .B(n15878), .ZN(
        n15880) );
  AOI211_X1 U18999 ( .C1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n17418), .A(
        n15881), .B(n15880), .ZN(n15888) );
  AOI22_X1 U19000 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15887) );
  NOR2_X1 U19001 ( .A1(n15882), .A2(n21224), .ZN(n15883) );
  AOI22_X1 U19002 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15898) );
  INV_X1 U19003 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U19004 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15890) );
  AOI22_X1 U19005 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15889) );
  OAI211_X1 U19006 ( .C1(n17427), .C2(n17408), .A(n15890), .B(n15889), .ZN(
        n15896) );
  AOI22_X1 U19007 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15894) );
  AOI22_X1 U19008 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U19009 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15892) );
  NAND2_X1 U19010 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n15891) );
  NAND4_X1 U19011 ( .A1(n15894), .A2(n15893), .A3(n15892), .A4(n15891), .ZN(
        n15895) );
  AOI211_X1 U19012 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15896), .B(n15895), .ZN(n15897) );
  OAI211_X1 U19013 ( .C1(n15718), .C2(n21348), .A(n15898), .B(n15897), .ZN(
        n15951) );
  AOI22_X1 U19014 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15908) );
  INV_X1 U19015 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U19016 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15900) );
  AOI22_X1 U19017 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15899) );
  OAI211_X1 U19018 ( .C1(n13976), .C2(n17380), .A(n15900), .B(n15899), .ZN(
        n15906) );
  AOI22_X1 U19019 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19020 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19021 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15902) );
  NAND2_X1 U19022 ( .A1(n15843), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n15901) );
  NAND4_X1 U19023 ( .A1(n15904), .A2(n15903), .A3(n15902), .A4(n15901), .ZN(
        n15905) );
  AOI211_X1 U19024 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n15906), .B(n15905), .ZN(n15907) );
  OAI211_X1 U19025 ( .C1(n17483), .C2(n21259), .A(n15908), .B(n15907), .ZN(
        n15953) );
  NAND2_X1 U19026 ( .A1(n15935), .A2(n15953), .ZN(n15909) );
  AOI21_X1 U19027 ( .B1(n18047), .B2(n15909), .A(n9788), .ZN(n15938) );
  INV_X1 U19028 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21212) );
  INV_X1 U19029 ( .A(n15952), .ZN(n17640) );
  XNOR2_X1 U19030 ( .A(n17640), .B(n15910), .ZN(n18079) );
  INV_X1 U19031 ( .A(n15951), .ZN(n17644) );
  XNOR2_X1 U19032 ( .A(n17644), .B(n15911), .ZN(n15912) );
  NAND2_X1 U19033 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15912), .ZN(
        n15934) );
  XOR2_X1 U19034 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15912), .Z(
        n18092) );
  NAND2_X1 U19035 ( .A1(n17660), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15928) );
  AOI22_X1 U19036 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15913) );
  OAI21_X1 U19037 ( .B1(n17473), .B2(n17482), .A(n15913), .ZN(n15918) );
  AOI22_X1 U19038 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17379), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U19039 ( .A1(n15914), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15915) );
  OAI211_X1 U19040 ( .C1(n17427), .C2(n21175), .A(n15916), .B(n15915), .ZN(
        n15917) );
  AOI211_X1 U19041 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n15918), .B(n15917), .ZN(n15927) );
  AOI22_X1 U19042 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15919) );
  OAI21_X1 U19043 ( .B1(n9878), .B2(n18803), .A(n15919), .ZN(n15925) );
  AOI22_X1 U19044 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15920) );
  INV_X1 U19045 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15921) );
  NAND2_X1 U19046 ( .A1(n15922), .A2(n10411), .ZN(n15923) );
  INV_X1 U19047 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19118) );
  NOR2_X1 U19048 ( .A1(n18134), .A2(n19118), .ZN(n18133) );
  NAND2_X1 U19049 ( .A1(n15928), .A2(n18124), .ZN(n18113) );
  INV_X1 U19050 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18437) );
  NAND2_X1 U19051 ( .A1(n18113), .A2(n18114), .ZN(n18112) );
  OR2_X1 U19052 ( .A1(n18437), .A2(n15929), .ZN(n15930) );
  NAND2_X1 U19053 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15931), .ZN(
        n15933) );
  INV_X1 U19054 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18422) );
  XOR2_X1 U19055 ( .A(n17648), .B(n15932), .Z(n18105) );
  INV_X1 U19056 ( .A(n15953), .ZN(n17637) );
  XNOR2_X1 U19057 ( .A(n17637), .B(n15935), .ZN(n15936) );
  XOR2_X1 U19058 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15936), .Z(
        n18064) );
  NAND2_X1 U19059 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15936), .ZN(
        n15937) );
  NAND2_X2 U19060 ( .A1(n18063), .A2(n15937), .ZN(n15939) );
  NAND2_X1 U19061 ( .A1(n15938), .A2(n15939), .ZN(n15940) );
  NAND2_X2 U19062 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15994), .ZN(
        n18330) );
  NAND2_X1 U19063 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18307), .ZN(
        n17961) );
  NAND2_X1 U19064 ( .A1(n16670), .A2(n18206), .ZN(n17779) );
  NAND3_X1 U19065 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n18150), .ZN(n16712) );
  NAND2_X1 U19066 ( .A1(n18488), .A2(n19141), .ZN(n15941) );
  NOR2_X1 U19067 ( .A1(n18504), .A2(n15941), .ZN(n15988) );
  INV_X1 U19068 ( .A(n15988), .ZN(n15942) );
  NAND2_X1 U19069 ( .A1(n18047), .A2(n18920), .ZN(n18306) );
  INV_X1 U19070 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17780) );
  INV_X1 U19071 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21361) );
  NOR3_X1 U19072 ( .A1(n17780), .A2(n17794), .A3(n21361), .ZN(n15980) );
  NAND2_X1 U19073 ( .A1(n15945), .A2(n15944), .ZN(n19157) );
  NOR2_X1 U19074 ( .A1(n21226), .A2(n17978), .ZN(n18293) );
  NAND2_X1 U19075 ( .A1(n18293), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18276) );
  INV_X1 U19076 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17944) );
  NOR2_X1 U19077 ( .A1(n18276), .A2(n17944), .ZN(n16718) );
  AOI21_X1 U19078 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18425) );
  INV_X1 U19079 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18410) );
  NOR3_X1 U19080 ( .A1(n21212), .A2(n18422), .A3(n18410), .ZN(n18363) );
  NAND4_X1 U19081 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18363), .ZN(n18254) );
  NOR2_X1 U19082 ( .A1(n18425), .A2(n18254), .ZN(n18334) );
  NAND2_X1 U19083 ( .A1(n16718), .A2(n18334), .ZN(n16012) );
  INV_X1 U19084 ( .A(n18363), .ZN(n18379) );
  NOR3_X1 U19085 ( .A1(n18437), .A2(n10078), .A3(n18379), .ZN(n18365) );
  NAND4_X1 U19086 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18365), .ZN(n18353) );
  NOR2_X1 U19087 ( .A1(n18255), .A2(n18353), .ZN(n18147) );
  INV_X1 U19088 ( .A(n18147), .ZN(n18244) );
  AOI21_X2 U19089 ( .B1(n18933), .B2(n15949), .A(n18932), .ZN(n18929) );
  OR2_X2 U19090 ( .A1(n16075), .A2(n17663), .ZN(n18922) );
  NOR2_X4 U19091 ( .A1(n18922), .A2(n15950), .ZN(n18952) );
  NOR2_X1 U19092 ( .A1(n18458), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18442) );
  INV_X1 U19093 ( .A(n18442), .ZN(n18426) );
  NAND2_X1 U19094 ( .A1(n10005), .A2(n18426), .ZN(n18251) );
  OAI22_X1 U19095 ( .A1(n18923), .A2(n16012), .B1(n18244), .B2(n18251), .ZN(
        n18166) );
  NAND2_X1 U19096 ( .A1(n15980), .A2(n18166), .ZN(n16696) );
  OAI21_X1 U19097 ( .B1(n16712), .B2(n18306), .A(n16696), .ZN(n15991) );
  NOR2_X1 U19098 ( .A1(n15961), .A2(n17652), .ZN(n15959) );
  NOR2_X1 U19099 ( .A1(n15959), .A2(n17648), .ZN(n15958) );
  NAND2_X1 U19100 ( .A1(n15958), .A2(n15951), .ZN(n15956) );
  NOR2_X1 U19101 ( .A1(n15952), .A2(n15956), .ZN(n15955) );
  NAND2_X1 U19102 ( .A1(n15955), .A2(n15953), .ZN(n15954) );
  NOR2_X1 U19103 ( .A1(n18047), .A2(n15954), .ZN(n15978) );
  XOR2_X1 U19104 ( .A(n15954), .B(n18047), .Z(n18054) );
  XNOR2_X1 U19105 ( .A(n15955), .B(n17637), .ZN(n15972) );
  XNOR2_X1 U19106 ( .A(n15956), .B(n17640), .ZN(n15957) );
  NAND2_X1 U19107 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15957), .ZN(
        n15971) );
  XOR2_X1 U19108 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15957), .Z(
        n18077) );
  XNOR2_X1 U19109 ( .A(n15958), .B(n17644), .ZN(n15969) );
  XOR2_X1 U19110 ( .A(n15959), .B(n17648), .Z(n15960) );
  NAND2_X1 U19111 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15960), .ZN(
        n15967) );
  XOR2_X1 U19112 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15960), .Z(
        n18103) );
  OR2_X1 U19113 ( .A1(n18437), .A2(n15962), .ZN(n15966) );
  INV_X1 U19114 ( .A(n18134), .ZN(n16081) );
  AOI21_X1 U19115 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15965), .A(
        n16081), .ZN(n15964) );
  NOR2_X1 U19116 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15965), .ZN(
        n15963) );
  AOI221_X1 U19117 ( .B1(n16081), .B2(n15965), .C1(n15964), .C2(n19118), .A(
        n15963), .ZN(n18116) );
  NAND2_X1 U19118 ( .A1(n18117), .A2(n18116), .ZN(n18115) );
  NAND2_X1 U19119 ( .A1(n15966), .A2(n18115), .ZN(n18102) );
  NAND2_X1 U19120 ( .A1(n18103), .A2(n18102), .ZN(n18101) );
  NAND2_X1 U19121 ( .A1(n15967), .A2(n18101), .ZN(n15968) );
  NAND2_X1 U19122 ( .A1(n15969), .A2(n15968), .ZN(n15970) );
  NAND2_X1 U19123 ( .A1(n15971), .A2(n18075), .ZN(n15973) );
  NAND2_X1 U19124 ( .A1(n15972), .A2(n15973), .ZN(n15974) );
  XOR2_X1 U19125 ( .A(n15973), .B(n15972), .Z(n18070) );
  NAND2_X1 U19126 ( .A1(n18070), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18069) );
  INV_X1 U19127 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18366) );
  NAND2_X1 U19128 ( .A1(n15978), .A2(n15975), .ZN(n15979) );
  NAND2_X1 U19129 ( .A1(n18054), .A2(n18055), .ZN(n18053) );
  NAND2_X1 U19130 ( .A1(n15978), .A2(n15977), .ZN(n15976) );
  OAI211_X1 U19131 ( .C1(n15978), .C2(n15977), .A(n18053), .B(n15976), .ZN(
        n18037) );
  NAND2_X1 U19132 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18037), .ZN(
        n18036) );
  AOI21_X1 U19133 ( .B1(n15982), .B2(n15981), .A(n18921), .ZN(n19134) );
  XOR2_X1 U19134 ( .A(n18488), .B(n19141), .Z(n15983) );
  INV_X1 U19135 ( .A(n19151), .ZN(n19143) );
  AOI21_X1 U19136 ( .B1(n15983), .B2(n19005), .A(n19143), .ZN(n16820) );
  NAND3_X1 U19137 ( .A1(n15986), .A2(n16820), .A3(n15984), .ZN(n15985) );
  OAI21_X1 U19138 ( .B1(n15986), .B2(n16645), .A(n15985), .ZN(n15987) );
  AOI21_X1 U19139 ( .B1(n19134), .B2(n15988), .A(n15987), .ZN(n15989) );
  OAI221_X1 U19140 ( .B1(n15991), .B2(n16714), .C1(n15991), .C2(n18974), .A(
        n18439), .ZN(n16064) );
  INV_X1 U19141 ( .A(n18047), .ZN(n18046) );
  INV_X1 U19142 ( .A(n18920), .ZN(n15992) );
  INV_X1 U19143 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16698) );
  NOR2_X1 U19144 ( .A1(n17780), .A2(n16004), .ZN(n16008) );
  NAND2_X1 U19145 ( .A1(n17903), .A2(n18242), .ZN(n15993) );
  INV_X1 U19146 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17870) );
  NAND2_X1 U19147 ( .A1(n17868), .A2(n17870), .ZN(n17847) );
  INV_X1 U19148 ( .A(n15995), .ZN(n18009) );
  NOR2_X2 U19149 ( .A1(n18255), .A2(n17979), .ZN(n15999) );
  NOR2_X1 U19150 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18014) );
  AND2_X1 U19151 ( .A1(n17944), .A2(n18291), .ZN(n15996) );
  NAND2_X1 U19152 ( .A1(n17952), .A2(n15996), .ZN(n17920) );
  INV_X1 U19153 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15997) );
  INV_X1 U19154 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18250) );
  INV_X1 U19155 ( .A(n15999), .ZN(n16000) );
  INV_X1 U19156 ( .A(n17826), .ZN(n17818) );
  NAND2_X1 U19157 ( .A1(n16004), .A2(n17818), .ZN(n16002) );
  OAI221_X1 U19158 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16004), 
        .C1(n18164), .C2(n16003), .A(n16002), .ZN(n17805) );
  NOR2_X1 U19159 ( .A1(n16004), .A2(n18142), .ZN(n16005) );
  OR2_X1 U19160 ( .A1(n17817), .A2(n16005), .ZN(n16006) );
  NOR2_X1 U19161 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9788), .ZN(
        n16707) );
  AOI22_X1 U19162 ( .A1(n16008), .A2(n16708), .B1(n16707), .B2(n16709), .ZN(
        n16009) );
  NOR2_X1 U19163 ( .A1(n19103), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19159) );
  NAND2_X2 U19164 ( .A1(n19146), .A2(n19159), .ZN(n18407) );
  NAND2_X1 U19165 ( .A1(n18923), .A2(n18952), .ZN(n18346) );
  OAI221_X1 U19166 ( .B1(n18952), .B2(n16670), .C1(n18952), .C2(n18147), .A(
        n18439), .ZN(n16014) );
  INV_X1 U19167 ( .A(n18189), .ZN(n16010) );
  NOR2_X1 U19168 ( .A1(n19118), .A2(n18353), .ZN(n18316) );
  INV_X1 U19169 ( .A(n18316), .ZN(n18335) );
  NOR2_X1 U19170 ( .A1(n18255), .A2(n18335), .ZN(n18266) );
  NAND2_X1 U19171 ( .A1(n16010), .A2(n18266), .ZN(n18146) );
  NAND3_X1 U19172 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18142), .ZN(n18141) );
  NOR2_X1 U19173 ( .A1(n21361), .A2(n18141), .ZN(n17781) );
  INV_X1 U19174 ( .A(n17781), .ZN(n16720) );
  OAI21_X1 U19175 ( .B1(n18146), .B2(n16720), .A(n18950), .ZN(n16011) );
  INV_X1 U19176 ( .A(n16011), .ZN(n16013) );
  NAND2_X1 U19177 ( .A1(n18947), .A2(n16012), .ZN(n18202) );
  OAI21_X1 U19178 ( .B1(n16670), .B2(n18923), .A(n18202), .ZN(n18144) );
  NOR3_X1 U19179 ( .A1(n16014), .A2(n16013), .A3(n18144), .ZN(n16061) );
  OAI21_X1 U19180 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18340), .A(
        n16061), .ZN(n16713) );
  AOI21_X1 U19181 ( .B1(n17780), .B2(n18367), .A(n16713), .ZN(n16015) );
  NAND2_X1 U19182 ( .A1(n18974), .A2(n18439), .ZN(n18431) );
  NAND2_X1 U19183 ( .A1(n16714), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16667) );
  NAND2_X1 U19184 ( .A1(n18047), .A2(n18454), .ZN(n18178) );
  INV_X1 U19185 ( .A(n18178), .ZN(n18374) );
  NOR3_X1 U19186 ( .A1(n17780), .A2(n21361), .A3(n16698), .ZN(n16669) );
  NAND2_X1 U19187 ( .A1(n18150), .A2(n16669), .ZN(n16666) );
  AOI22_X1 U19188 ( .A1(n18456), .A2(n16667), .B1(n18374), .B2(n16666), .ZN(
        n16067) );
  OAI21_X1 U19189 ( .B1(n18446), .B2(n16015), .A(n16067), .ZN(n16016) );
  AOI22_X1 U19190 ( .A1(n18373), .A2(n16688), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16016), .ZN(n16017) );
  NAND2_X1 U19191 ( .A1(n18446), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16685) );
  OAI211_X1 U19192 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16064), .A(
        n16017), .B(n16685), .ZN(P3_U2833) );
  INV_X1 U19193 ( .A(n16018), .ZN(n16019) );
  OAI211_X1 U19194 ( .C1(n10928), .C2(n16020), .A(n16019), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16023) );
  INV_X1 U19195 ( .A(n16021), .ZN(n16022) );
  OAI21_X1 U19196 ( .B1(n16023), .B2(n20957), .A(n16022), .ZN(n16025) );
  NAND2_X1 U19197 ( .A1(n16023), .A2(n20957), .ZN(n16024) );
  OAI21_X1 U19198 ( .B1(n16026), .B2(n16025), .A(n16024), .ZN(n16027) );
  AOI222_X1 U19199 ( .A1(n16028), .A2(n20679), .B1(n16028), .B2(n16027), .C1(
        n20679), .C2(n16027), .ZN(n16030) );
  INV_X1 U19200 ( .A(n16030), .ZN(n16032) );
  INV_X1 U19201 ( .A(n16033), .ZN(n16029) );
  AOI21_X1 U19202 ( .B1(n16030), .B2(n16029), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16031) );
  AOI21_X1 U19203 ( .B1(n16033), .B2(n16032), .A(n16031), .ZN(n16042) );
  INV_X1 U19204 ( .A(n16034), .ZN(n16038) );
  OAI21_X1 U19205 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16035), .ZN(n16036) );
  AND4_X1 U19206 ( .A1(n16039), .A2(n16038), .A3(n16037), .A4(n16036), .ZN(
        n16041) );
  OAI211_X1 U19207 ( .C1(n16042), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16041), .B(n16040), .ZN(n16052) );
  INV_X1 U19208 ( .A(n16043), .ZN(n16046) );
  NOR2_X1 U19209 ( .A1(n16044), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21120) );
  NAND3_X1 U19210 ( .A1(n16046), .A2(n21120), .A3(n16045), .ZN(n16050) );
  OAI21_X1 U19211 ( .B1(n21119), .B2(n16048), .A(n16047), .ZN(n16049) );
  NAND2_X1 U19212 ( .A1(n16050), .A2(n16049), .ZN(n16410) );
  AOI221_X1 U19213 ( .B1(n21027), .B2(n21324), .C1(n16052), .C2(n21324), .A(
        n16410), .ZN(n16415) );
  AOI21_X1 U19214 ( .B1(n16053), .B2(n16052), .A(n16051), .ZN(n16054) );
  OAI211_X1 U19215 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21119), .A(n16054), 
        .B(n16057), .ZN(n16055) );
  NOR2_X1 U19216 ( .A1(n16415), .A2(n16055), .ZN(n16060) );
  OR2_X1 U19217 ( .A1(n16057), .A2(n16056), .ZN(n16058) );
  NAND2_X1 U19218 ( .A1(n21027), .A2(n16058), .ZN(n16059) );
  OAI22_X1 U19219 ( .A1(n16060), .A2(n21027), .B1(n16415), .B2(n16059), .ZN(
        P1_U3161) );
  INV_X1 U19220 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16680) );
  NAND2_X1 U19221 ( .A1(n18439), .A2(n18367), .ZN(n18441) );
  OAI22_X1 U19222 ( .A1(n18441), .A2(n16669), .B1(n18451), .B2(n16061), .ZN(
        n16062) );
  INV_X1 U19223 ( .A(n16062), .ZN(n16695) );
  NAND3_X1 U19224 ( .A1(n16709), .A2(n16707), .A3(n16698), .ZN(n16647) );
  NAND2_X1 U19225 ( .A1(n16649), .A2(n16647), .ZN(n16063) );
  XOR2_X1 U19226 ( .A(n16063), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16678) );
  INV_X1 U19227 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19077) );
  NOR2_X1 U19228 ( .A1(n18407), .A2(n19077), .ZN(n16672) );
  NOR3_X1 U19229 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16698), .A3(
        n16064), .ZN(n16065) );
  AOI211_X1 U19230 ( .C1(n18373), .C2(n16678), .A(n16672), .B(n16065), .ZN(
        n16066) );
  OAI221_X1 U19231 ( .B1(n16680), .B2(n16695), .C1(n16680), .C2(n16067), .A(
        n16066), .ZN(P3_U2832) );
  INV_X1 U19232 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21051) );
  INV_X1 U19233 ( .A(HOLD), .ZN(n21050) );
  NOR2_X1 U19234 ( .A1(n21051), .A2(n21050), .ZN(n21036) );
  AOI22_X1 U19235 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16070) );
  NAND2_X1 U19236 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n16068), .ZN(n21044) );
  OAI211_X1 U19237 ( .C1(n21036), .C2(n16070), .A(n16069), .B(n21044), .ZN(
        P1_U3195) );
  AND2_X1 U19238 ( .A1(n20331), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19239 ( .A1(n20150), .A2(n21322), .ZN(n20020) );
  NAND2_X1 U19240 ( .A1(n20020), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16072) );
  NOR2_X1 U19241 ( .A1(n15656), .A2(n20153), .ZN(n20123) );
  AOI21_X1 U19242 ( .B1(n20123), .B2(n21322), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16071) );
  AOI21_X1 U19243 ( .B1(n16072), .B2(n16071), .A(n16073), .ZN(P2_U3178) );
  INV_X1 U19244 ( .A(n16073), .ZN(n16643) );
  OAI221_X1 U19245 ( .B1(n12144), .B2(n16643), .C1(n16596), .C2(n16643), .A(
        n19917), .ZN(n20137) );
  NOR2_X1 U19246 ( .A1(n16074), .A2(n20137), .ZN(P2_U3047) );
  INV_X1 U19247 ( .A(n18985), .ZN(n19149) );
  INV_X1 U19248 ( .A(n16075), .ZN(n16079) );
  INV_X1 U19249 ( .A(n17521), .ZN(n17657) );
  NAND2_X1 U19250 ( .A1(n18511), .A2(n17657), .ZN(n17632) );
  INV_X1 U19251 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21289) );
  AOI22_X1 U19252 ( .A1(n17654), .A2(BUF2_REG_0__SCAN_IN), .B1(n17653), .B2(
        n16081), .ZN(n16082) );
  OAI221_X1 U19253 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17632), .C1(n21289), 
        .C2(n17657), .A(n16082), .ZN(P3_U2735) );
  INV_X1 U19254 ( .A(n16083), .ZN(n16085) );
  NAND2_X1 U19255 ( .A1(n16085), .A2(n16084), .ZN(n16086) );
  AND2_X1 U19256 ( .A1(n16086), .A2(n20224), .ZN(n16114) );
  INV_X1 U19257 ( .A(n16114), .ZN(n16098) );
  NAND2_X1 U19258 ( .A1(n20236), .A2(n16097), .ZN(n16095) );
  INV_X1 U19259 ( .A(n16087), .ZN(n16088) );
  AOI22_X1 U19260 ( .A1(n20261), .A2(P1_EBX_REG_22__SCAN_IN), .B1(n16088), 
        .B2(n20257), .ZN(n16089) );
  OAI21_X1 U19261 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n16090), .A(n16089), 
        .ZN(n16093) );
  OAI22_X1 U19262 ( .A1(n16091), .A2(n20218), .B1(n20279), .B2(n16287), .ZN(
        n16092) );
  OAI221_X1 U19263 ( .B1(n16295), .B2(n16098), .C1(n16295), .C2(n16095), .A(
        n16094), .ZN(P1_U2818) );
  OAI22_X1 U19264 ( .A1(n16208), .A2(n20285), .B1(n16096), .B2(n16095), .ZN(
        n16100) );
  OAI22_X1 U19265 ( .A1(n16098), .A2(n16097), .B1(n16189), .B2(n20276), .ZN(
        n16099) );
  AOI211_X1 U19266 ( .C1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n20271), .A(
        n16100), .B(n16099), .ZN(n16106) );
  NAND2_X1 U19267 ( .A1(n16102), .A2(n16101), .ZN(n16103) );
  NOR2_X1 U19268 ( .A1(n16186), .A2(n20279), .ZN(n16104) );
  AOI21_X1 U19269 ( .B1(n16204), .B2(n20210), .A(n16104), .ZN(n16105) );
  NAND2_X1 U19270 ( .A1(n16106), .A2(n16105), .ZN(P1_U2819) );
  AOI22_X1 U19271 ( .A1(n20261), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20257), 
        .B2(n16107), .ZN(n16116) );
  NOR2_X1 U19272 ( .A1(n16108), .A2(n16157), .ZN(n16147) );
  NAND2_X1 U19273 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n16147), .ZN(n16122) );
  OAI21_X1 U19274 ( .B1(n16109), .B2(n16122), .A(n21077), .ZN(n16113) );
  OAI22_X1 U19275 ( .A1(n16111), .A2(n20218), .B1(n20279), .B2(n16110), .ZN(
        n16112) );
  AOI21_X1 U19276 ( .B1(n16114), .B2(n16113), .A(n16112), .ZN(n16115) );
  OAI211_X1 U19277 ( .C1(n16117), .C2(n20240), .A(n16116), .B(n16115), .ZN(
        P1_U2820) );
  INV_X1 U19278 ( .A(n16219), .ZN(n16118) );
  AOI22_X1 U19279 ( .A1(n20261), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n16118), 
        .B2(n20257), .ZN(n16129) );
  INV_X1 U19280 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21074) );
  NOR3_X1 U19281 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21074), .A3(n16122), 
        .ZN(n16119) );
  AOI211_X1 U19282 ( .C1(n20271), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16119), .B(n16368), .ZN(n16128) );
  OAI22_X1 U19283 ( .A1(n16120), .A2(n20218), .B1(n16297), .B2(n20279), .ZN(
        n16121) );
  INV_X1 U19284 ( .A(n16121), .ZN(n16127) );
  NOR2_X1 U19285 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n16122), .ZN(n16138) );
  INV_X1 U19286 ( .A(n16123), .ZN(n16124) );
  OAI21_X1 U19287 ( .B1(n16125), .B2(n16124), .A(n16168), .ZN(n16146) );
  OAI21_X1 U19288 ( .B1(n16138), .B2(n16146), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n16126) );
  NAND4_X1 U19289 ( .A1(n16129), .A2(n16128), .A3(n16127), .A4(n16126), .ZN(
        P1_U2821) );
  NAND2_X1 U19290 ( .A1(n16146), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16136) );
  NAND2_X1 U19291 ( .A1(n20271), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16130) );
  OAI211_X1 U19292 ( .C1(n20276), .C2(n16131), .A(n20243), .B(n16130), .ZN(
        n16134) );
  NOR2_X1 U19293 ( .A1(n16132), .A2(n20285), .ZN(n16133) );
  NOR2_X1 U19294 ( .A1(n16134), .A2(n16133), .ZN(n16135) );
  NAND2_X1 U19295 ( .A1(n16136), .A2(n16135), .ZN(n16137) );
  NOR2_X1 U19296 ( .A1(n16138), .A2(n16137), .ZN(n16139) );
  OAI21_X1 U19297 ( .B1(n16140), .B2(n20218), .A(n16139), .ZN(n16141) );
  INV_X1 U19298 ( .A(n16141), .ZN(n16142) );
  OAI21_X1 U19299 ( .B1(n20279), .B2(n16143), .A(n16142), .ZN(P1_U2822) );
  AOI22_X1 U19300 ( .A1(n20261), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20271), .ZN(n16151) );
  AOI21_X1 U19301 ( .B1(n20257), .B2(n16220), .A(n16368), .ZN(n16150) );
  INV_X1 U19302 ( .A(n16144), .ZN(n16145) );
  AOI22_X1 U19303 ( .A1(n16221), .A2(n20210), .B1(n20260), .B2(n16145), .ZN(
        n16149) );
  OAI21_X1 U19304 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16147), .A(n16146), 
        .ZN(n16148) );
  NAND4_X1 U19305 ( .A1(n16151), .A2(n16150), .A3(n16149), .A4(n16148), .ZN(
        P1_U2823) );
  AOI22_X1 U19306 ( .A1(n16235), .A2(n20257), .B1(n20260), .B2(n16317), .ZN(
        n16156) );
  NAND2_X1 U19307 ( .A1(n20271), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16152) );
  OAI211_X1 U19308 ( .C1(n16315), .C2(n16168), .A(n16152), .B(n20243), .ZN(
        n16154) );
  NOR2_X1 U19309 ( .A1(n16234), .A2(n20218), .ZN(n16153) );
  AOI211_X1 U19310 ( .C1(n20261), .C2(P1_EBX_REG_15__SCAN_IN), .A(n16154), .B(
        n16153), .ZN(n16155) );
  OAI211_X1 U19311 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16157), .A(n16156), 
        .B(n16155), .ZN(P1_U2825) );
  NOR2_X1 U19312 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16158), .ZN(n16169) );
  INV_X1 U19313 ( .A(n16159), .ZN(n16160) );
  AOI22_X1 U19314 ( .A1(n20261), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n16160), 
        .B2(n20257), .ZN(n16167) );
  INV_X1 U19315 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16161) );
  OAI21_X1 U19316 ( .B1(n20240), .B2(n16161), .A(n20243), .ZN(n16164) );
  NOR2_X1 U19317 ( .A1(n16162), .A2(n20218), .ZN(n16163) );
  AOI211_X1 U19318 ( .C1(n16165), .C2(n20260), .A(n16164), .B(n16163), .ZN(
        n16166) );
  OAI211_X1 U19319 ( .C1(n16169), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        P1_U2826) );
  AOI22_X1 U19320 ( .A1(n20261), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n16241), 
        .B2(n20257), .ZN(n16177) );
  AOI22_X1 U19321 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20271), .B1(
        n20260), .B2(n16170), .ZN(n16176) );
  INV_X1 U19322 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16172) );
  NAND2_X1 U19323 ( .A1(n20236), .A2(n16171), .ZN(n16180) );
  OAI21_X1 U19324 ( .B1(n16172), .B2(n16180), .A(n21065), .ZN(n16173) );
  AOI22_X1 U19325 ( .A1(n20210), .A2(n16240), .B1(n16174), .B2(n16173), .ZN(
        n16175) );
  NAND4_X1 U19326 ( .A1(n16177), .A2(n16176), .A3(n16175), .A4(n20243), .ZN(
        P1_U2828) );
  INV_X1 U19327 ( .A(n16253), .ZN(n16178) );
  AOI22_X1 U19328 ( .A1(n20261), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n16178), 
        .B2(n20257), .ZN(n16185) );
  OAI22_X1 U19329 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16180), .B1(n16179), 
        .B2(n20240), .ZN(n16181) );
  AOI211_X1 U19330 ( .C1(n16332), .C2(n20260), .A(n16368), .B(n16181), .ZN(
        n16184) );
  AOI22_X1 U19331 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16182), .B1(n20210), 
        .B2(n16250), .ZN(n16183) );
  NAND3_X1 U19332 ( .A1(n16185), .A2(n16184), .A3(n16183), .ZN(P1_U2829) );
  NOR2_X1 U19333 ( .A1(n16186), .A2(n20288), .ZN(n16187) );
  AOI21_X1 U19334 ( .B1(n16204), .B2(n20299), .A(n16187), .ZN(n16188) );
  OAI21_X1 U19335 ( .B1(n20302), .B2(n16189), .A(n16188), .ZN(P1_U2851) );
  AOI22_X1 U19336 ( .A1(n16191), .A2(n20416), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16190), .ZN(n16195) );
  AOI22_X1 U19337 ( .A1(n16204), .A2(n16193), .B1(n16192), .B2(DATAI_21_), 
        .ZN(n16194) );
  OAI211_X1 U19338 ( .C1(n16196), .C2(n16744), .A(n16195), .B(n16194), .ZN(
        P1_U2883) );
  AOI22_X1 U19339 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16202) );
  INV_X1 U19340 ( .A(n16197), .ZN(n16200) );
  XNOR2_X1 U19341 ( .A(n9753), .B(n16284), .ZN(n16198) );
  XNOR2_X1 U19342 ( .A(n16199), .B(n16198), .ZN(n16281) );
  AOI22_X1 U19343 ( .A1(n16200), .A2(n20378), .B1(n20369), .B2(n16281), .ZN(
        n16201) );
  OAI211_X1 U19344 ( .C1(n16254), .C2(n16203), .A(n16202), .B(n16201), .ZN(
        P1_U2976) );
  INV_X1 U19345 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21145) );
  NAND2_X1 U19346 ( .A1(n16204), .A2(n20378), .ZN(n16207) );
  NAND2_X1 U19347 ( .A1(n16205), .A2(n20369), .ZN(n16206) );
  OAI211_X1 U19348 ( .C1(n16254), .C2(n16208), .A(n16207), .B(n16206), .ZN(
        n16209) );
  INV_X1 U19349 ( .A(n16209), .ZN(n16211) );
  NAND2_X1 U19350 ( .A1(n16368), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16210) );
  OAI211_X1 U19351 ( .C1(n21145), .C2(n16268), .A(n16211), .B(n16210), .ZN(
        P1_U2978) );
  AOI22_X1 U19352 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16218) );
  NOR2_X1 U19353 ( .A1(n16212), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16214) );
  MUX2_X1 U19354 ( .A(n16214), .B(n9753), .S(n16213), .Z(n16215) );
  XNOR2_X1 U19355 ( .A(n16215), .B(n10912), .ZN(n16299) );
  AOI22_X1 U19356 ( .A1(n16299), .A2(n20369), .B1(n16216), .B2(n20378), .ZN(
        n16217) );
  OAI211_X1 U19357 ( .C1(n16254), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        P1_U2980) );
  AOI22_X1 U19358 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16223) );
  AOI22_X1 U19359 ( .A1(n16221), .A2(n20378), .B1(n16220), .B2(n16265), .ZN(
        n16222) );
  OAI211_X1 U19360 ( .C1(n16244), .C2(n16224), .A(n16223), .B(n16222), .ZN(
        P1_U2982) );
  AND2_X1 U19361 ( .A1(n16226), .A2(n16225), .ZN(n16227) );
  NAND2_X1 U19362 ( .A1(n16228), .A2(n16227), .ZN(n16233) );
  INV_X1 U19363 ( .A(n16229), .ZN(n16231) );
  NOR2_X1 U19364 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  XNOR2_X1 U19365 ( .A(n16233), .B(n16232), .ZN(n16320) );
  AOI22_X1 U19366 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16238) );
  INV_X1 U19367 ( .A(n16234), .ZN(n16236) );
  AOI22_X1 U19368 ( .A1(n16236), .A2(n20378), .B1(n16235), .B2(n16265), .ZN(
        n16237) );
  OAI211_X1 U19369 ( .C1(n16320), .C2(n16244), .A(n16238), .B(n16237), .ZN(
        P1_U2984) );
  INV_X1 U19370 ( .A(n16239), .ZN(n16245) );
  AOI22_X1 U19371 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16243) );
  AOI22_X1 U19372 ( .A1(n16265), .A2(n16241), .B1(n20378), .B2(n16240), .ZN(
        n16242) );
  OAI211_X1 U19373 ( .C1(n16245), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        P1_U2987) );
  AOI22_X1 U19374 ( .A1(n20367), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16368), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16252) );
  NOR3_X1 U19375 ( .A1(n14644), .A2(n10070), .A3(n16350), .ZN(n16248) );
  NOR2_X1 U19376 ( .A1(n16248), .A2(n16247), .ZN(n16249) );
  XNOR2_X1 U19377 ( .A(n16249), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16334) );
  AOI22_X1 U19378 ( .A1(n20369), .A2(n16334), .B1(n20378), .B2(n16250), .ZN(
        n16251) );
  OAI211_X1 U19379 ( .C1(n16254), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P1_U2988) );
  OAI21_X1 U19380 ( .B1(n16257), .B2(n16256), .A(n9775), .ZN(n16385) );
  INV_X1 U19381 ( .A(n20207), .ZN(n16258) );
  AOI222_X1 U19382 ( .A1(n16385), .A2(n20369), .B1(n16258), .B2(n16265), .C1(
        n20378), .C2(n20294), .ZN(n16260) );
  NOR2_X1 U19383 ( .A1(n20243), .A2(n21242), .ZN(n16380) );
  INV_X1 U19384 ( .A(n16380), .ZN(n16259) );
  OAI211_X1 U19385 ( .C1(n16261), .C2(n16268), .A(n16260), .B(n16259), .ZN(
        P1_U2992) );
  XOR2_X1 U19386 ( .A(n16263), .B(n16262), .Z(n16401) );
  INV_X1 U19387 ( .A(n16264), .ZN(n20226) );
  AOI222_X1 U19388 ( .A1(n16401), .A2(n20369), .B1(n20378), .B2(n20300), .C1(
        n20226), .C2(n16265), .ZN(n16267) );
  NOR2_X1 U19389 ( .A1(n20243), .A2(n20234), .ZN(n16394) );
  INV_X1 U19390 ( .A(n16394), .ZN(n16266) );
  OAI211_X1 U19391 ( .C1(n16269), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        P1_U2994) );
  INV_X1 U19392 ( .A(n16270), .ZN(n16273) );
  AOI211_X1 U19393 ( .C1(n16273), .C2(n16400), .A(n16272), .B(n16271), .ZN(
        n16277) );
  AOI22_X1 U19394 ( .A1(n16275), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n16395), .B2(n16274), .ZN(n16276) );
  NAND2_X1 U19395 ( .A1(n16277), .A2(n16276), .ZN(P1_U3006) );
  INV_X1 U19396 ( .A(n16278), .ZN(n16279) );
  AOI22_X1 U19397 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n16368), .B1(n16279), 
        .B2(n16284), .ZN(n16283) );
  AOI22_X1 U19398 ( .A1(n16281), .A2(n16400), .B1(n16395), .B2(n16280), .ZN(
        n16282) );
  OAI211_X1 U19399 ( .C1(n16285), .C2(n16284), .A(n16283), .B(n16282), .ZN(
        P1_U3008) );
  INV_X1 U19400 ( .A(n16286), .ZN(n16290) );
  INV_X1 U19401 ( .A(n16287), .ZN(n16288) );
  AOI222_X1 U19402 ( .A1(n16290), .A2(n16400), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16289), .C1(n16395), .C2(
        n16288), .ZN(n16294) );
  OAI211_X1 U19403 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16292), .B(n16291), .ZN(
        n16293) );
  OAI211_X1 U19404 ( .C1(n16295), .C2(n20243), .A(n16294), .B(n16293), .ZN(
        P1_U3009) );
  AOI22_X1 U19405 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16296), .B1(
        n16368), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16301) );
  INV_X1 U19406 ( .A(n16297), .ZN(n16298) );
  AOI22_X1 U19407 ( .A1(n16299), .A2(n16400), .B1(n16395), .B2(n16298), .ZN(
        n16300) );
  OAI211_X1 U19408 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16302), .A(
        n16301), .B(n16300), .ZN(P1_U3012) );
  OAI21_X1 U19409 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16303), .A(
        n16331), .ZN(n16304) );
  INV_X1 U19410 ( .A(n16304), .ZN(n16323) );
  INV_X1 U19411 ( .A(n16305), .ZN(n16311) );
  NAND2_X1 U19412 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16306), .ZN(
        n16314) );
  AOI221_X1 U19413 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n21199), .C2(n16313), .A(
        n16314), .ZN(n16307) );
  AOI21_X1 U19414 ( .B1(n16368), .B2(P1_REIP_REG_16__SCAN_IN), .A(n16307), 
        .ZN(n16308) );
  OAI21_X1 U19415 ( .B1(n16309), .B2(n16383), .A(n16308), .ZN(n16310) );
  AOI21_X1 U19416 ( .B1(n16311), .B2(n16400), .A(n16310), .ZN(n16312) );
  OAI21_X1 U19417 ( .B1(n16323), .B2(n16313), .A(n16312), .ZN(P1_U3015) );
  OAI22_X1 U19418 ( .A1(n20243), .A2(n16315), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16314), .ZN(n16316) );
  AOI21_X1 U19419 ( .B1(n16317), .B2(n16395), .A(n16316), .ZN(n16318) );
  OAI21_X1 U19420 ( .B1(n16320), .B2(n16319), .A(n16318), .ZN(n16321) );
  INV_X1 U19421 ( .A(n16321), .ZN(n16322) );
  OAI21_X1 U19422 ( .B1(n16323), .B2(n21199), .A(n16322), .ZN(P1_U3016) );
  AOI21_X1 U19423 ( .B1(n16325), .B2(n16395), .A(n16324), .ZN(n16329) );
  AOI22_X1 U19424 ( .A1(n16327), .A2(n16400), .B1(n16330), .B2(n16326), .ZN(
        n16328) );
  OAI211_X1 U19425 ( .C1(n16331), .C2(n16330), .A(n16329), .B(n16328), .ZN(
        P1_U3018) );
  AOI22_X1 U19426 ( .A1(n16332), .A2(n16395), .B1(n16368), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U19427 ( .A1(n16334), .A2(n16400), .B1(n16333), .B2(n16366), .ZN(
        n16335) );
  OAI211_X1 U19428 ( .C1(n16338), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        P1_U3020) );
  AOI221_X1 U19429 ( .B1(n16340), .B2(n16364), .C1(n16343), .C2(n16364), .A(
        n16339), .ZN(n16362) );
  INV_X1 U19430 ( .A(n16341), .ZN(n16348) );
  OR2_X1 U19431 ( .A1(n16343), .A2(n16342), .ZN(n16357) );
  AOI221_X1 U19432 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16350), .C2(n16361), .A(
        n16357), .ZN(n16344) );
  AOI21_X1 U19433 ( .B1(n16368), .B2(P1_REIP_REG_10__SCAN_IN), .A(n16344), 
        .ZN(n16345) );
  OAI21_X1 U19434 ( .B1(n16346), .B2(n16383), .A(n16345), .ZN(n16347) );
  AOI21_X1 U19435 ( .B1(n16348), .B2(n16400), .A(n16347), .ZN(n16349) );
  OAI21_X1 U19436 ( .B1(n16362), .B2(n16350), .A(n16349), .ZN(P1_U3021) );
  INV_X1 U19437 ( .A(n16351), .ZN(n16359) );
  NAND2_X1 U19438 ( .A1(n16353), .A2(n16352), .ZN(n16354) );
  AND2_X1 U19439 ( .A1(n16355), .A2(n16354), .ZN(n20286) );
  AOI22_X1 U19440 ( .A1(n20286), .A2(n16395), .B1(n16368), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16356) );
  OAI21_X1 U19441 ( .B1(n16357), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16356), .ZN(n16358) );
  AOI21_X1 U19442 ( .B1(n16359), .B2(n16400), .A(n16358), .ZN(n16360) );
  OAI21_X1 U19443 ( .B1(n16362), .B2(n16361), .A(n16360), .ZN(P1_U3022) );
  AOI21_X1 U19444 ( .B1(n13734), .B2(n16364), .A(n16363), .ZN(n16388) );
  INV_X1 U19445 ( .A(n16365), .ZN(n16372) );
  NAND2_X1 U19446 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16366), .ZN(
        n16379) );
  AOI221_X1 U19447 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16374), .C2(n16387), .A(
        n16379), .ZN(n16367) );
  AOI21_X1 U19448 ( .B1(n16368), .B2(P1_REIP_REG_8__SCAN_IN), .A(n16367), .ZN(
        n16369) );
  OAI21_X1 U19449 ( .B1(n16370), .B2(n16383), .A(n16369), .ZN(n16371) );
  AOI21_X1 U19450 ( .B1(n16372), .B2(n16400), .A(n16371), .ZN(n16373) );
  OAI21_X1 U19451 ( .B1(n16388), .B2(n16374), .A(n16373), .ZN(P1_U3023) );
  AOI21_X1 U19452 ( .B1(n16392), .B2(n16376), .A(n16375), .ZN(n16377) );
  OR2_X1 U19453 ( .A1(n16378), .A2(n16377), .ZN(n20204) );
  INV_X1 U19454 ( .A(n16379), .ZN(n16381) );
  AOI21_X1 U19455 ( .B1(n16387), .B2(n16381), .A(n16380), .ZN(n16382) );
  OAI21_X1 U19456 ( .B1(n20204), .B2(n16383), .A(n16382), .ZN(n16384) );
  AOI21_X1 U19457 ( .B1(n16385), .B2(n16400), .A(n16384), .ZN(n16386) );
  OAI21_X1 U19458 ( .B1(n16388), .B2(n16387), .A(n16386), .ZN(P1_U3024) );
  AOI21_X1 U19459 ( .B1(n16391), .B2(n16390), .A(n16389), .ZN(n16393) );
  NOR2_X1 U19460 ( .A1(n16393), .A2(n16392), .ZN(n20297) );
  AOI21_X1 U19461 ( .B1(n20297), .B2(n16395), .A(n16394), .ZN(n16396) );
  OAI21_X1 U19462 ( .B1(n16398), .B2(n16397), .A(n16396), .ZN(n16399) );
  AOI21_X1 U19463 ( .B1(n16401), .B2(n16400), .A(n16399), .ZN(n16402) );
  OAI21_X1 U19464 ( .B1(n16403), .B2(n10850), .A(n16402), .ZN(P1_U3026) );
  NAND3_X1 U19465 ( .A1(n16404), .A2(n21102), .A3(n16407), .ZN(n16405) );
  OAI21_X1 U19466 ( .B1(n16407), .B2(n16406), .A(n16405), .ZN(P1_U3468) );
  NAND4_X1 U19467 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n21030), .A4(n21119), .ZN(n16408) );
  NAND2_X1 U19468 ( .A1(n16409), .A2(n16408), .ZN(n21028) );
  OAI21_X1 U19469 ( .B1(n16411), .B2(n21028), .A(n16410), .ZN(n16412) );
  OAI221_X1 U19470 ( .B1(n16413), .B2(n20840), .C1(n16413), .C2(n21119), .A(
        n16412), .ZN(n16414) );
  AOI221_X1 U19471 ( .B1(n16415), .B2(n21324), .C1(n21027), .C2(n21324), .A(
        n16414), .ZN(P1_U3162) );
  NOR2_X1 U19472 ( .A1(n16415), .A2(n21027), .ZN(n16417) );
  OAI22_X1 U19473 ( .A1(n20840), .A2(n16417), .B1(n16416), .B2(n21027), .ZN(
        P1_U3466) );
  INV_X1 U19474 ( .A(n16418), .ZN(n16431) );
  AOI21_X1 U19475 ( .B1(n16421), .B2(n16420), .A(n16419), .ZN(n16430) );
  NOR2_X1 U19476 ( .A1(n19324), .A2(n16422), .ZN(n16425) );
  OAI22_X1 U19477 ( .A1(n19341), .A2(n20089), .B1(n19282), .B2(n16423), .ZN(
        n16424) );
  AOI211_X1 U19478 ( .C1(n16426), .C2(n19339), .A(n16425), .B(n16424), .ZN(
        n16427) );
  OAI21_X1 U19479 ( .B1(n16428), .B2(n19346), .A(n16427), .ZN(n16429) );
  AOI21_X1 U19480 ( .B1(n16431), .B2(n16430), .A(n16429), .ZN(n16432) );
  OAI21_X1 U19481 ( .B1(n16433), .B2(n19335), .A(n16432), .ZN(P2_U2826) );
  AOI21_X1 U19482 ( .B1(n16436), .B2(n16435), .A(n16434), .ZN(n16446) );
  OAI22_X1 U19483 ( .A1(n19341), .A2(n20087), .B1(n19282), .B2(n21232), .ZN(
        n16437) );
  AOI21_X1 U19484 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19344), .A(n16437), .ZN(
        n16443) );
  INV_X1 U19485 ( .A(n16438), .ZN(n16440) );
  OAI211_X1 U19486 ( .C1(n16441), .C2(n16440), .A(n16439), .B(n19339), .ZN(
        n16442) );
  OAI211_X1 U19487 ( .C1(n16444), .C2(n19346), .A(n16443), .B(n16442), .ZN(
        n16445) );
  AOI21_X1 U19488 ( .B1(n19336), .B2(n16446), .A(n16445), .ZN(n16447) );
  OAI21_X1 U19489 ( .B1(n16448), .B2(n19335), .A(n16447), .ZN(P2_U2828) );
  AOI211_X1 U19490 ( .C1(n16452), .C2(n16450), .A(n16451), .B(n20024), .ZN(
        n16461) );
  OAI22_X1 U19491 ( .A1(n19341), .A2(n16453), .B1(n19282), .B2(n10297), .ZN(
        n16457) );
  AOI211_X1 U19492 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n16455), .A(n19306), .B(
        n16454), .ZN(n16456) );
  AOI211_X1 U19493 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n19344), .A(n16457), .B(
        n16456), .ZN(n16458) );
  OAI21_X1 U19494 ( .B1(n16459), .B2(n19346), .A(n16458), .ZN(n16460) );
  AOI211_X1 U19495 ( .C1(n19337), .C2(n16462), .A(n16461), .B(n16460), .ZN(
        n16463) );
  INV_X1 U19496 ( .A(n16463), .ZN(P2_U2829) );
  AOI211_X1 U19497 ( .C1(n16467), .C2(n16465), .A(n16466), .B(n20024), .ZN(
        n16477) );
  XNOR2_X1 U19498 ( .A(n16468), .B(n16471), .ZN(n16475) );
  INV_X1 U19499 ( .A(n16469), .ZN(n16473) );
  AOI22_X1 U19500 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19327), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19349), .ZN(n16470) );
  OAI21_X1 U19501 ( .B1(n19324), .B2(n16471), .A(n16470), .ZN(n16472) );
  AOI21_X1 U19502 ( .B1(n16473), .B2(n12566), .A(n16472), .ZN(n16474) );
  OAI21_X1 U19503 ( .B1(n16475), .B2(n19306), .A(n16474), .ZN(n16476) );
  AOI211_X1 U19504 ( .C1(n19337), .C2(n16478), .A(n16477), .B(n16476), .ZN(
        n16479) );
  INV_X1 U19505 ( .A(n16479), .ZN(P2_U2831) );
  AOI22_X1 U19506 ( .A1(n19356), .A2(n16480), .B1(n12547), .B2(n19385), .ZN(
        P2_U2856) );
  NOR2_X1 U19507 ( .A1(n16481), .A2(n19385), .ZN(n16482) );
  AOI21_X1 U19508 ( .B1(n16483), .B2(n19386), .A(n16482), .ZN(n16484) );
  OAI21_X1 U19509 ( .B1(n19356), .B2(n12113), .A(n16484), .ZN(P2_U2864) );
  AOI22_X1 U19510 ( .A1(n16485), .A2(n19386), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19385), .ZN(n16486) );
  OAI21_X1 U19511 ( .B1(n19385), .B2(n16510), .A(n16486), .ZN(P2_U2865) );
  AOI21_X1 U19512 ( .B1(n16487), .B2(n9924), .A(n14992), .ZN(n16495) );
  AOI22_X1 U19513 ( .A1(n16495), .A2(n19386), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19385), .ZN(n16488) );
  OAI21_X1 U19514 ( .B1(n19385), .B2(n16489), .A(n16488), .ZN(P2_U2867) );
  AOI21_X1 U19515 ( .B1(n16490), .B2(n15003), .A(n9840), .ZN(n16502) );
  AOI22_X1 U19516 ( .A1(n16502), .A2(n19386), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19385), .ZN(n16491) );
  OAI21_X1 U19517 ( .B1(n19385), .B2(n16492), .A(n16491), .ZN(P2_U2869) );
  AOI22_X1 U19518 ( .A1(n19396), .A2(n16493), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19419), .ZN(n16498) );
  AOI22_X1 U19519 ( .A1(n19398), .A2(BUF2_REG_20__SCAN_IN), .B1(n19397), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U19520 ( .A1(n16495), .A2(n16501), .B1(n19392), .B2(n16494), .ZN(
        n16496) );
  NAND3_X1 U19521 ( .A1(n16498), .A2(n16497), .A3(n16496), .ZN(P2_U2899) );
  INV_X1 U19522 ( .A(n19468), .ZN(n16499) );
  AOI22_X1 U19523 ( .A1(n19396), .A2(n16499), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19419), .ZN(n16505) );
  AOI22_X1 U19524 ( .A1(n19398), .A2(BUF2_REG_18__SCAN_IN), .B1(n19397), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19525 ( .A1(n16502), .A2(n16501), .B1(n19392), .B2(n16500), .ZN(
        n16503) );
  NAND3_X1 U19526 ( .A1(n16505), .A2(n16504), .A3(n16503), .ZN(P2_U2901) );
  AOI22_X1 U19527 ( .A1(n16546), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19326), .ZN(n16513) );
  NAND2_X1 U19528 ( .A1(n16506), .A2(n16549), .ZN(n16509) );
  NAND2_X1 U19529 ( .A1(n16507), .A2(n16550), .ZN(n16508) );
  OAI211_X1 U19530 ( .C1(n13882), .C2(n16510), .A(n16509), .B(n16508), .ZN(
        n16511) );
  INV_X1 U19531 ( .A(n16511), .ZN(n16512) );
  OAI211_X1 U19532 ( .C1(n16554), .C2(n16514), .A(n16513), .B(n16512), .ZN(
        P2_U2992) );
  AOI22_X1 U19533 ( .A1(n16546), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19326), .ZN(n16519) );
  INV_X1 U19534 ( .A(n19365), .ZN(n16516) );
  OAI211_X1 U19535 ( .C1(n16554), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        P2_U3000) );
  AOI22_X1 U19536 ( .A1(n16546), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19326), .ZN(n16525) );
  INV_X1 U19537 ( .A(n19378), .ZN(n16522) );
  AOI222_X1 U19538 ( .A1(n16523), .A2(n16549), .B1(n16561), .B2(n16522), .C1(
        n16550), .C2(n16521), .ZN(n16524) );
  OAI211_X1 U19539 ( .C1(n16554), .C2(n19277), .A(n16525), .B(n16524), .ZN(
        P2_U3004) );
  AOI22_X1 U19540 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19326), .B1(n16555), 
        .B2(n19284), .ZN(n16531) );
  OAI22_X1 U19541 ( .A1(n16527), .A2(n16558), .B1(n16557), .B2(n16526), .ZN(
        n16528) );
  AOI21_X1 U19542 ( .B1(n16561), .B2(n16529), .A(n16528), .ZN(n16530) );
  OAI211_X1 U19543 ( .C1(n16565), .C2(n16532), .A(n16531), .B(n16530), .ZN(
        P2_U3005) );
  AOI22_X1 U19544 ( .A1(n16546), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19326), .ZN(n16544) );
  NAND2_X1 U19545 ( .A1(n16534), .A2(n16533), .ZN(n16538) );
  NAND2_X1 U19546 ( .A1(n16536), .A2(n16535), .ZN(n16537) );
  XNOR2_X1 U19547 ( .A(n16538), .B(n16537), .ZN(n16576) );
  INV_X1 U19548 ( .A(n19384), .ZN(n16575) );
  OAI21_X1 U19549 ( .B1(n16541), .B2(n16540), .A(n16539), .ZN(n16542) );
  INV_X1 U19550 ( .A(n16542), .ZN(n16573) );
  AOI222_X1 U19551 ( .A1(n16576), .A2(n16549), .B1(n16561), .B2(n16575), .C1(
        n16550), .C2(n16573), .ZN(n16543) );
  OAI211_X1 U19552 ( .C1(n16554), .C2(n16545), .A(n16544), .B(n16543), .ZN(
        P2_U3006) );
  AOI22_X1 U19553 ( .A1(n16546), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19326), .ZN(n16553) );
  INV_X1 U19554 ( .A(n16547), .ZN(n16551) );
  AOI222_X1 U19555 ( .A1(n16551), .A2(n16550), .B1(n16549), .B2(n16548), .C1(
        n16561), .C2(n19315), .ZN(n16552) );
  OAI211_X1 U19556 ( .C1(n16554), .C2(n19313), .A(n16553), .B(n16552), .ZN(
        P2_U3008) );
  AOI22_X1 U19557 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19326), .B1(n16555), 
        .B2(n19330), .ZN(n16563) );
  OAI22_X1 U19558 ( .A1(n16559), .A2(n16558), .B1(n16557), .B2(n16556), .ZN(
        n16560) );
  AOI21_X1 U19559 ( .B1(n16561), .B2(n19331), .A(n16560), .ZN(n16562) );
  OAI211_X1 U19560 ( .C1(n16565), .C2(n16564), .A(n16563), .B(n16562), .ZN(
        P2_U3009) );
  INV_X1 U19561 ( .A(n16566), .ZN(n16568) );
  AOI211_X1 U19562 ( .C1(n16579), .C2(n16569), .A(n16568), .B(n16567), .ZN(
        n16572) );
  INV_X1 U19563 ( .A(n16570), .ZN(n19417) );
  INV_X1 U19564 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20059) );
  OAI22_X1 U19565 ( .A1(n16581), .A2(n19417), .B1(n20059), .B2(n19305), .ZN(
        n16571) );
  NOR2_X1 U19566 ( .A1(n16572), .A2(n16571), .ZN(n16578) );
  AOI222_X1 U19567 ( .A1(n16576), .A2(n16592), .B1(n16586), .B2(n16575), .C1(
        n16574), .C2(n16573), .ZN(n16577) );
  OAI211_X1 U19568 ( .C1(n16580), .C2(n16579), .A(n16578), .B(n16577), .ZN(
        P2_U3038) );
  OAI22_X1 U19569 ( .A1(n16581), .A2(n20111), .B1(n13639), .B2(n15303), .ZN(
        n16585) );
  NOR3_X1 U19570 ( .A1(n16583), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n16582), .ZN(n16584) );
  AOI211_X1 U19571 ( .C1(n16586), .C2(n9839), .A(n16585), .B(n16584), .ZN(
        n16587) );
  OAI21_X1 U19572 ( .B1(n16589), .B2(n16588), .A(n16587), .ZN(n16590) );
  AOI21_X1 U19573 ( .B1(n16592), .B2(n16591), .A(n16590), .ZN(n16593) );
  OAI21_X1 U19574 ( .B1(n16595), .B2(n16594), .A(n16593), .ZN(P2_U3043) );
  INV_X1 U19575 ( .A(n16596), .ZN(n20142) );
  NOR2_X1 U19576 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n21322), .ZN(n20022) );
  MUX2_X1 U19577 ( .A(n16598), .B(n16597), .S(n16611), .Z(n16612) );
  OR2_X1 U19578 ( .A1(n16612), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16608) );
  INV_X1 U19579 ( .A(n16601), .ZN(n16603) );
  INV_X1 U19580 ( .A(n16599), .ZN(n16600) );
  OAI211_X1 U19581 ( .C1(n16601), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16600), .ZN(n16602) );
  OAI21_X1 U19582 ( .B1(n16603), .B2(n11863), .A(n16602), .ZN(n16604) );
  AOI211_X1 U19583 ( .C1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n16608), .A(
        n16611), .B(n16604), .ZN(n16607) );
  MUX2_X1 U19584 ( .A(n16605), .B(n15689), .S(n16611), .Z(n16613) );
  INV_X1 U19585 ( .A(n16613), .ZN(n16606) );
  AOI222_X1 U19586 ( .A1(n16607), .A2(n20114), .B1(n16607), .B2(n16606), .C1(
        n20114), .C2(n16606), .ZN(n16609) );
  AOI221_X1 U19587 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16609), 
        .C1(n16608), .C2(n16609), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16610) );
  AOI21_X1 U19588 ( .B1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16611), .A(
        n16610), .ZN(n16638) );
  NOR2_X1 U19589 ( .A1(n16613), .A2(n16612), .ZN(n16629) );
  INV_X1 U19590 ( .A(n16614), .ZN(n16621) );
  INV_X1 U19591 ( .A(n16615), .ZN(n16617) );
  AOI22_X1 U19592 ( .A1(n16621), .A2(n16618), .B1(n16617), .B2(n16616), .ZN(
        n16619) );
  OAI21_X1 U19593 ( .B1(n16621), .B2(n16620), .A(n16619), .ZN(n20145) );
  OAI21_X1 U19594 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16622), .ZN(n16627) );
  NAND3_X1 U19595 ( .A1(n16625), .A2(n16624), .A3(n16623), .ZN(n16626) );
  OAI211_X1 U19596 ( .C1(n9812), .C2(n20143), .A(n16627), .B(n16626), .ZN(
        n16628) );
  NOR3_X1 U19597 ( .A1(n16629), .A2(n20145), .A3(n16628), .ZN(n16636) );
  NAND4_X1 U19598 ( .A1(n16638), .A2(n20165), .A3(n16636), .A4(n16635), .ZN(
        n16644) );
  NAND2_X1 U19599 ( .A1(n16630), .A2(n16644), .ZN(n20025) );
  AOI21_X1 U19600 ( .B1(n21322), .B2(n16631), .A(n20159), .ZN(n16632) );
  AOI21_X1 U19601 ( .B1(n20150), .B2(n20025), .A(n16632), .ZN(n16634) );
  AOI211_X1 U19602 ( .C1(n20150), .C2(n20022), .A(n16634), .B(n16633), .ZN(
        n16641) );
  INV_X1 U19603 ( .A(n16635), .ZN(n16637) );
  NAND3_X1 U19604 ( .A1(n16638), .A2(n16637), .A3(n16636), .ZN(n16639) );
  NAND2_X1 U19605 ( .A1(n16639), .A2(n20165), .ZN(n16640) );
  OAI211_X1 U19606 ( .C1(n20142), .C2(n16643), .A(n16641), .B(n16640), .ZN(
        P2_U3176) );
  OAI211_X1 U19607 ( .C1(n20110), .C2(n16644), .A(n16643), .B(n16642), .ZN(
        P2_U3593) );
  INV_X1 U19608 ( .A(n16645), .ZN(n19132) );
  AOI22_X1 U19609 ( .A1(n18974), .A2(n19132), .B1(n19134), .B2(n18920), .ZN(
        n16646) );
  INV_X1 U19610 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19099) );
  AOI22_X1 U19611 ( .A1(n9788), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n19099), .B2(n16004), .ZN(n16655) );
  NAND2_X1 U19612 ( .A1(n16004), .A2(n16647), .ZN(n16651) );
  OAI211_X1 U19613 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16680), .A(
        n16649), .B(n16651), .ZN(n16648) );
  OAI21_X1 U19614 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16004), .A(
        n16648), .ZN(n16654) );
  AOI21_X1 U19615 ( .B1(n16649), .B2(n9788), .A(n16680), .ZN(n16650) );
  INV_X1 U19616 ( .A(n16650), .ZN(n16652) );
  NAND3_X1 U19617 ( .A1(n16655), .A2(n16652), .A3(n16651), .ZN(n16653) );
  OAI21_X1 U19618 ( .B1(n16655), .B2(n16654), .A(n16653), .ZN(n16706) );
  NAND2_X1 U19619 ( .A1(n19091), .A2(n18462), .ZN(n19148) );
  INV_X1 U19620 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16841) );
  NOR2_X1 U19621 ( .A1(n19100), .A2(n16841), .ZN(n18089) );
  INV_X1 U19622 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21214) );
  INV_X1 U19623 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17800) );
  NAND2_X1 U19624 ( .A1(n18085), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17954) );
  NAND2_X1 U19625 ( .A1(n18041), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17069) );
  NAND3_X1 U19626 ( .A1(n18038), .A2(n17955), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17970) );
  NAND2_X1 U19627 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17972) );
  NAND3_X1 U19628 ( .A1(n17924), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17910) );
  INV_X1 U19629 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17834) );
  INV_X1 U19630 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21355) );
  XNOR2_X2 U19631 ( .A(n16656), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17130) );
  INV_X1 U19632 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19079) );
  NOR2_X1 U19633 ( .A1(n18407), .A2(n19079), .ZN(n16700) );
  NAND2_X1 U19634 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17775), .ZN(
        n16686) );
  INV_X1 U19635 ( .A(n16686), .ZN(n16657) );
  NAND2_X1 U19636 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16657), .ZN(
        n16659) );
  NAND2_X1 U19637 ( .A1(n19146), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18135) );
  AOI21_X1 U19638 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16658), .A(
        n18866), .ZN(n17971) );
  OR2_X1 U19639 ( .A1(n16659), .A2(n17971), .ZN(n16675) );
  XNOR2_X1 U19640 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16660) );
  NOR2_X1 U19641 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17856), .ZN(
        n16683) );
  NAND2_X1 U19642 ( .A1(n18866), .A2(n16659), .ZN(n16687) );
  OAI211_X1 U19643 ( .C1(n9862), .C2(n18135), .A(n18136), .B(n16687), .ZN(
        n16692) );
  NOR2_X1 U19644 ( .A1(n16683), .A2(n16692), .ZN(n16674) );
  OAI22_X1 U19645 ( .A1(n16675), .A2(n16660), .B1(n16674), .B2(n21355), .ZN(
        n16661) );
  AOI211_X1 U19646 ( .C1(n17927), .C2(n17130), .A(n16700), .B(n16661), .ZN(
        n16665) );
  OR2_X1 U19647 ( .A1(n16666), .A2(n16680), .ZN(n16662) );
  XOR2_X1 U19648 ( .A(n16662), .B(n19099), .Z(n16703) );
  NAND3_X1 U19649 ( .A1(n16714), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16663) );
  XOR2_X1 U19650 ( .A(n16663), .B(n19099), .Z(n16702) );
  AOI22_X1 U19651 ( .A1(n17998), .A2(n16703), .B1(n18127), .B2(n16702), .ZN(
        n16664) );
  OAI211_X1 U19652 ( .C1(n17967), .C2(n16706), .A(n16665), .B(n16664), .ZN(
        P3_U2799) );
  NAND2_X1 U19653 ( .A1(n17998), .A2(n16666), .ZN(n16694) );
  NAND2_X1 U19654 ( .A1(n18127), .A2(n16667), .ZN(n16689) );
  NOR2_X2 U19655 ( .A1(n18255), .A2(n18035), .ZN(n17933) );
  AND4_X1 U19656 ( .A1(n16680), .A2(n16670), .A3(n16669), .A4(n17933), .ZN(
        n16677) );
  INV_X1 U19657 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21279) );
  AOI22_X1 U19658 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16671), .B1(
        n16681), .B2(n21279), .ZN(n16860) );
  AOI21_X1 U19659 ( .B1(n17927), .B2(n16860), .A(n16672), .ZN(n16673) );
  OAI221_X1 U19660 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16675), .C1(
        n21279), .C2(n16674), .A(n16673), .ZN(n16676) );
  AOI211_X1 U19661 ( .C1(n18032), .C2(n16678), .A(n16677), .B(n16676), .ZN(
        n16679) );
  OAI221_X1 U19662 ( .B1(n16680), .B2(n16694), .C1(n16680), .C2(n16689), .A(
        n16679), .ZN(P3_U2800) );
  OAI21_X1 U19663 ( .B1(n9862), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16681), .ZN(n16682) );
  INV_X1 U19664 ( .A(n16682), .ZN(n16868) );
  OAI21_X1 U19665 ( .B1(n16683), .B2(n17927), .A(n16868), .ZN(n16684) );
  OAI211_X1 U19666 ( .C1(n16687), .C2(n16686), .A(n16685), .B(n16684), .ZN(
        n16691) );
  NOR2_X1 U19667 ( .A1(n16714), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16690) );
  OAI221_X1 U19668 ( .B1(n16694), .B2(n16712), .C1(n16694), .C2(n16698), .A(
        n16693), .ZN(P3_U2801) );
  OAI21_X1 U19669 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18441), .A(
        n16695), .ZN(n16701) );
  NAND2_X1 U19670 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19099), .ZN(
        n16697) );
  NOR4_X1 U19671 ( .A1(n18457), .A2(n16698), .A3(n16697), .A4(n16696), .ZN(
        n16699) );
  AOI211_X1 U19672 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16701), .A(
        n16700), .B(n16699), .ZN(n16705) );
  AOI22_X1 U19673 ( .A1(n16703), .A2(n18374), .B1(n16702), .B2(n18456), .ZN(
        n16704) );
  OAI211_X1 U19674 ( .C1(n18302), .C2(n16706), .A(n16705), .B(n16704), .ZN(
        P3_U2831) );
  NAND2_X1 U19675 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18446), .ZN(n17777) );
  INV_X1 U19676 ( .A(n18306), .ZN(n18331) );
  AOI21_X1 U19677 ( .B1(n9788), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16707), .ZN(n17784) );
  INV_X1 U19678 ( .A(n16709), .ZN(n16721) );
  NAND2_X1 U19679 ( .A1(n16721), .A2(n16710), .ZN(n17783) );
  INV_X1 U19680 ( .A(n18974), .ZN(n19131) );
  OR2_X1 U19681 ( .A1(n16714), .A2(n19131), .ZN(n16715) );
  OAI22_X1 U19682 ( .A1(n18332), .A2(n19131), .B1(n18306), .B2(n18330), .ZN(
        n18319) );
  AOI21_X1 U19683 ( .B1(n16718), .B2(n18319), .A(n18166), .ZN(n18179) );
  INV_X1 U19684 ( .A(n18203), .ZN(n17851) );
  NOR2_X1 U19685 ( .A1(n18179), .A2(n17851), .ZN(n18209) );
  NAND2_X1 U19686 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18209), .ZN(
        n18196) );
  NAND4_X1 U19687 ( .A1(n17777), .A2(n16724), .A3(n16723), .A4(n16722), .ZN(
        P3_U2834) );
  NOR3_X1 U19688 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16726) );
  NOR4_X1 U19689 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16725) );
  NAND4_X1 U19690 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16726), .A3(n16725), .A4(
        U215), .ZN(U213) );
  INV_X1 U19691 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16809) );
  INV_X2 U19692 ( .A(U214), .ZN(n16774) );
  NOR2_X1 U19693 ( .A1(n16774), .A2(n16727), .ZN(n16771) );
  INV_X2 U19694 ( .A(n16771), .ZN(n16776) );
  INV_X1 U19695 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19489) );
  INV_X1 U19696 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16811) );
  OAI222_X1 U19697 ( .A1(U212), .A2(n16809), .B1(n16776), .B2(n19489), .C1(
        U214), .C2(n16811), .ZN(U216) );
  INV_X1 U19698 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16729) );
  AOI22_X1 U19699 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16773), .ZN(n16728) );
  OAI21_X1 U19700 ( .B1(n16729), .B2(n16776), .A(n16728), .ZN(U217) );
  INV_X1 U19701 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16731) );
  AOI22_X1 U19702 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16773), .ZN(n16730) );
  OAI21_X1 U19703 ( .B1(n16731), .B2(n16776), .A(n16730), .ZN(U218) );
  INV_X1 U19704 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19705 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16773), .ZN(n16732) );
  OAI21_X1 U19706 ( .B1(n16733), .B2(n16776), .A(n16732), .ZN(U219) );
  INV_X1 U19707 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16735) );
  AOI22_X1 U19708 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16773), .ZN(n16734) );
  OAI21_X1 U19709 ( .B1(n16735), .B2(n16776), .A(n16734), .ZN(U220) );
  INV_X1 U19710 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19466) );
  AOI22_X1 U19711 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16773), .ZN(n16736) );
  OAI21_X1 U19712 ( .B1(n19466), .B2(n16776), .A(n16736), .ZN(U221) );
  INV_X1 U19713 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19714 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16773), .ZN(n16737) );
  OAI21_X1 U19715 ( .B1(n16738), .B2(n16776), .A(n16737), .ZN(U222) );
  INV_X1 U19716 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16740) );
  AOI22_X1 U19717 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16773), .ZN(n16739) );
  OAI21_X1 U19718 ( .B1(n16740), .B2(n16776), .A(n16739), .ZN(U223) );
  AOI22_X1 U19719 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16773), .ZN(n16741) );
  OAI21_X1 U19720 ( .B1(n15067), .B2(n16776), .A(n16741), .ZN(U224) );
  INV_X1 U19721 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19484) );
  AOI22_X1 U19722 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16773), .ZN(n16742) );
  OAI21_X1 U19723 ( .B1(n19484), .B2(n16776), .A(n16742), .ZN(U225) );
  AOI22_X1 U19724 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16773), .ZN(n16743) );
  OAI21_X1 U19725 ( .B1(n16744), .B2(n16776), .A(n16743), .ZN(U226) );
  INV_X1 U19726 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21160) );
  AOI22_X1 U19727 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16773), .ZN(n16745) );
  OAI21_X1 U19728 ( .B1(n21160), .B2(n16776), .A(n16745), .ZN(U227) );
  AOI22_X1 U19729 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16773), .ZN(n16746) );
  OAI21_X1 U19730 ( .B1(n15089), .B2(n16776), .A(n16746), .ZN(U228) );
  INV_X1 U19731 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20404) );
  AOI22_X1 U19732 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16773), .ZN(n16747) );
  OAI21_X1 U19733 ( .B1(n20404), .B2(n16776), .A(n16747), .ZN(U229) );
  AOI22_X1 U19734 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16773), .ZN(n16748) );
  OAI21_X1 U19735 ( .B1(n15100), .B2(n16776), .A(n16748), .ZN(U230) );
  INV_X1 U19736 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16750) );
  AOI22_X1 U19737 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16773), .ZN(n16749) );
  OAI21_X1 U19738 ( .B1(n16750), .B2(n16776), .A(n16749), .ZN(U231) );
  AOI22_X1 U19739 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16773), .ZN(n16751) );
  OAI21_X1 U19740 ( .B1(n13339), .B2(n16776), .A(n16751), .ZN(U232) );
  AOI22_X1 U19741 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16773), .ZN(n16752) );
  OAI21_X1 U19742 ( .B1(n14463), .B2(n16776), .A(n16752), .ZN(U233) );
  INV_X1 U19743 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16754) );
  AOI22_X1 U19744 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16773), .ZN(n16753) );
  OAI21_X1 U19745 ( .B1(n16754), .B2(n16776), .A(n16753), .ZN(U234) );
  AOI22_X1 U19746 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16773), .ZN(n16755) );
  OAI21_X1 U19747 ( .B1(n16756), .B2(n16776), .A(n16755), .ZN(U235) );
  AOI22_X1 U19748 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16773), .ZN(n16757) );
  OAI21_X1 U19749 ( .B1(n14482), .B2(n16776), .A(n16757), .ZN(U236) );
  AOI22_X1 U19750 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16773), .ZN(n16758) );
  OAI21_X1 U19751 ( .B1(n16759), .B2(n16776), .A(n16758), .ZN(U237) );
  INV_X1 U19752 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U19753 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16771), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16774), .ZN(n16760) );
  OAI21_X1 U19754 ( .B1(n21266), .B2(U212), .A(n16760), .ZN(U238) );
  AOI22_X1 U19755 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16773), .ZN(n16761) );
  OAI21_X1 U19756 ( .B1(n16762), .B2(n16776), .A(n16761), .ZN(U239) );
  INV_X1 U19757 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U19758 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16773), .ZN(n16763) );
  OAI21_X1 U19759 ( .B1(n16764), .B2(n16776), .A(n16763), .ZN(U240) );
  INV_X1 U19760 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16783) );
  AOI22_X1 U19761 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16771), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16774), .ZN(n16765) );
  OAI21_X1 U19762 ( .B1(n16783), .B2(U212), .A(n16765), .ZN(U241) );
  INV_X1 U19763 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n21358) );
  AOI22_X1 U19764 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16771), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16773), .ZN(n16766) );
  OAI21_X1 U19765 ( .B1(n21358), .B2(U214), .A(n16766), .ZN(U242) );
  AOI22_X1 U19766 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16773), .ZN(n16767) );
  OAI21_X1 U19767 ( .B1(n16768), .B2(n16776), .A(n16767), .ZN(U243) );
  INV_X1 U19768 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U19769 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16771), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16774), .ZN(n16769) );
  OAI21_X1 U19770 ( .B1(n16780), .B2(U212), .A(n16769), .ZN(U244) );
  AOI22_X1 U19771 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16773), .ZN(n16770) );
  OAI21_X1 U19772 ( .B1(n13463), .B2(n16776), .A(n16770), .ZN(U245) );
  INV_X1 U19773 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n21269) );
  AOI22_X1 U19774 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16771), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16773), .ZN(n16772) );
  OAI21_X1 U19775 ( .B1(n21269), .B2(U214), .A(n16772), .ZN(U246) );
  AOI22_X1 U19776 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16773), .ZN(n16775) );
  OAI21_X1 U19777 ( .B1(n13406), .B2(n16776), .A(n16775), .ZN(U247) );
  OAI22_X1 U19778 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16808), .ZN(n16777) );
  INV_X1 U19779 ( .A(n16777), .ZN(U251) );
  OAI22_X1 U19780 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16792), .ZN(n16778) );
  INV_X1 U19781 ( .A(n16778), .ZN(U252) );
  OAI22_X1 U19782 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16792), .ZN(n16779) );
  INV_X1 U19783 ( .A(n16779), .ZN(U253) );
  INV_X1 U19784 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21458) );
  AOI22_X1 U19785 ( .A1(n16808), .A2(n16780), .B1(n21458), .B2(U215), .ZN(U254) );
  OAI22_X1 U19786 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16792), .ZN(n16781) );
  INV_X1 U19787 ( .A(n16781), .ZN(U255) );
  OAI22_X1 U19788 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16792), .ZN(n16782) );
  INV_X1 U19789 ( .A(n16782), .ZN(U256) );
  INV_X1 U19790 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18503) );
  AOI22_X1 U19791 ( .A1(n16808), .A2(n16783), .B1(n18503), .B2(U215), .ZN(U257) );
  OAI22_X1 U19792 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16792), .ZN(n16784) );
  INV_X1 U19793 ( .A(n16784), .ZN(U258) );
  OAI22_X1 U19794 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16792), .ZN(n16785) );
  INV_X1 U19795 ( .A(n16785), .ZN(U259) );
  INV_X1 U19796 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17756) );
  AOI22_X1 U19797 ( .A1(n16808), .A2(n21266), .B1(n17756), .B2(U215), .ZN(U260) );
  OAI22_X1 U19798 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16792), .ZN(n16786) );
  INV_X1 U19799 ( .A(n16786), .ZN(U261) );
  OAI22_X1 U19800 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16808), .ZN(n16787) );
  INV_X1 U19801 ( .A(n16787), .ZN(U262) );
  OAI22_X1 U19802 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16792), .ZN(n16788) );
  INV_X1 U19803 ( .A(n16788), .ZN(U263) );
  OAI22_X1 U19804 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16808), .ZN(n16789) );
  INV_X1 U19805 ( .A(n16789), .ZN(U264) );
  OAI22_X1 U19806 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16792), .ZN(n16790) );
  INV_X1 U19807 ( .A(n16790), .ZN(U265) );
  OAI22_X1 U19808 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16808), .ZN(n16791) );
  INV_X1 U19809 ( .A(n16791), .ZN(U266) );
  OAI22_X1 U19810 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16792), .ZN(n16793) );
  INV_X1 U19811 ( .A(n16793), .ZN(U267) );
  OAI22_X1 U19812 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16808), .ZN(n16794) );
  INV_X1 U19813 ( .A(n16794), .ZN(U268) );
  OAI22_X1 U19814 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16808), .ZN(n16795) );
  INV_X1 U19815 ( .A(n16795), .ZN(U269) );
  OAI22_X1 U19816 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16808), .ZN(n16796) );
  INV_X1 U19817 ( .A(n16796), .ZN(U270) );
  INV_X1 U19818 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16797) );
  INV_X1 U19819 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19478) );
  AOI22_X1 U19820 ( .A1(n16808), .A2(n16797), .B1(n19478), .B2(U215), .ZN(U271) );
  OAI22_X1 U19821 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16808), .ZN(n16798) );
  INV_X1 U19822 ( .A(n16798), .ZN(U272) );
  OAI22_X1 U19823 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16808), .ZN(n16799) );
  INV_X1 U19824 ( .A(n16799), .ZN(U273) );
  OAI22_X1 U19825 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16808), .ZN(n16800) );
  INV_X1 U19826 ( .A(n16800), .ZN(U274) );
  OAI22_X1 U19827 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16808), .ZN(n16801) );
  INV_X1 U19828 ( .A(n16801), .ZN(U275) );
  OAI22_X1 U19829 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16808), .ZN(n16802) );
  INV_X1 U19830 ( .A(n16802), .ZN(U276) );
  INV_X1 U19831 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16803) );
  INV_X1 U19832 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19465) );
  AOI22_X1 U19833 ( .A1(n16808), .A2(n16803), .B1(n19465), .B2(U215), .ZN(U277) );
  OAI22_X1 U19834 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16808), .ZN(n16804) );
  INV_X1 U19835 ( .A(n16804), .ZN(U278) );
  OAI22_X1 U19836 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16808), .ZN(n16805) );
  INV_X1 U19837 ( .A(n16805), .ZN(U279) );
  OAI22_X1 U19838 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16808), .ZN(n16806) );
  INV_X1 U19839 ( .A(n16806), .ZN(U280) );
  OAI22_X1 U19840 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16808), .ZN(n16807) );
  INV_X1 U19841 ( .A(n16807), .ZN(U281) );
  INV_X1 U19842 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n21238) );
  AOI22_X1 U19843 ( .A1(n16808), .A2(n16809), .B1(n21238), .B2(U215), .ZN(U282) );
  INV_X1 U19844 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16810) );
  AOI222_X1 U19845 ( .A1(n16811), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16810), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .C1(n16809), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n16812) );
  INV_X2 U19846 ( .A(n16814), .ZN(n16813) );
  INV_X1 U19847 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19036) );
  INV_X1 U19848 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20064) );
  AOI22_X1 U19849 ( .A1(n16813), .A2(n19036), .B1(n20064), .B2(n16814), .ZN(
        U347) );
  INV_X1 U19850 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19034) );
  INV_X1 U19851 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20062) );
  AOI22_X1 U19852 ( .A1(n16813), .A2(n19034), .B1(n20062), .B2(n16814), .ZN(
        U348) );
  INV_X1 U19853 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19031) );
  INV_X1 U19854 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20060) );
  AOI22_X1 U19855 ( .A1(n16813), .A2(n19031), .B1(n20060), .B2(n16814), .ZN(
        U349) );
  INV_X1 U19856 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19030) );
  INV_X1 U19857 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U19858 ( .A1(n16813), .A2(n19030), .B1(n20058), .B2(n16814), .ZN(
        U350) );
  INV_X1 U19859 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19028) );
  INV_X1 U19860 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20056) );
  AOI22_X1 U19861 ( .A1(n16813), .A2(n19028), .B1(n20056), .B2(n16814), .ZN(
        U351) );
  INV_X1 U19862 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19026) );
  INV_X1 U19863 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20054) );
  AOI22_X1 U19864 ( .A1(n16813), .A2(n19026), .B1(n20054), .B2(n16814), .ZN(
        U352) );
  INV_X1 U19865 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19024) );
  INV_X1 U19866 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U19867 ( .A1(n16813), .A2(n19024), .B1(n20052), .B2(n16814), .ZN(
        U353) );
  INV_X1 U19868 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19022) );
  AOI22_X1 U19869 ( .A1(n16813), .A2(n19022), .B1(n20050), .B2(n16814), .ZN(
        U354) );
  INV_X1 U19870 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19078) );
  INV_X1 U19871 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21261) );
  AOI22_X1 U19872 ( .A1(n16813), .A2(n19078), .B1(n21261), .B2(n16814), .ZN(
        U355) );
  INV_X1 U19873 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19075) );
  INV_X1 U19874 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20090) );
  AOI22_X1 U19875 ( .A1(n16813), .A2(n19075), .B1(n20090), .B2(n16814), .ZN(
        U356) );
  INV_X1 U19876 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19072) );
  INV_X1 U19877 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20088) );
  AOI22_X1 U19878 ( .A1(n16813), .A2(n19072), .B1(n20088), .B2(n16814), .ZN(
        U357) );
  INV_X1 U19879 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19069) );
  INV_X1 U19880 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20086) );
  AOI22_X1 U19881 ( .A1(n16813), .A2(n19069), .B1(n20086), .B2(n16814), .ZN(
        U358) );
  INV_X1 U19882 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19068) );
  INV_X1 U19883 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20085) );
  AOI22_X1 U19884 ( .A1(n16813), .A2(n19068), .B1(n20085), .B2(n16814), .ZN(
        U359) );
  INV_X1 U19885 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19066) );
  INV_X1 U19886 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U19887 ( .A1(n16813), .A2(n19066), .B1(n20084), .B2(n16814), .ZN(
        U360) );
  INV_X1 U19888 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19064) );
  INV_X1 U19889 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20083) );
  AOI22_X1 U19890 ( .A1(n16813), .A2(n19064), .B1(n20083), .B2(n16814), .ZN(
        U361) );
  INV_X1 U19891 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19061) );
  INV_X1 U19892 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20081) );
  AOI22_X1 U19893 ( .A1(n16813), .A2(n19061), .B1(n20081), .B2(n16814), .ZN(
        U362) );
  INV_X1 U19894 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19060) );
  INV_X1 U19895 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20080) );
  AOI22_X1 U19896 ( .A1(n16813), .A2(n19060), .B1(n20080), .B2(n16814), .ZN(
        U363) );
  INV_X1 U19897 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19058) );
  INV_X1 U19898 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20079) );
  AOI22_X1 U19899 ( .A1(n16813), .A2(n19058), .B1(n20079), .B2(n16814), .ZN(
        U364) );
  INV_X1 U19900 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19020) );
  INV_X1 U19901 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20049) );
  AOI22_X1 U19902 ( .A1(n16813), .A2(n19020), .B1(n20049), .B2(n16814), .ZN(
        U365) );
  INV_X1 U19903 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19055) );
  INV_X1 U19904 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20078) );
  AOI22_X1 U19905 ( .A1(n16813), .A2(n19055), .B1(n20078), .B2(n16814), .ZN(
        U366) );
  INV_X1 U19906 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19054) );
  INV_X1 U19907 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20077) );
  AOI22_X1 U19908 ( .A1(n16813), .A2(n19054), .B1(n20077), .B2(n16814), .ZN(
        U367) );
  INV_X1 U19909 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19052) );
  INV_X1 U19910 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20076) );
  AOI22_X1 U19911 ( .A1(n16813), .A2(n19052), .B1(n20076), .B2(n16814), .ZN(
        U368) );
  INV_X1 U19912 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19049) );
  INV_X1 U19913 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20074) );
  AOI22_X1 U19914 ( .A1(n16813), .A2(n19049), .B1(n20074), .B2(n16814), .ZN(
        U369) );
  INV_X1 U19915 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19048) );
  INV_X1 U19916 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20072) );
  AOI22_X1 U19917 ( .A1(n16813), .A2(n19048), .B1(n20072), .B2(n16814), .ZN(
        U370) );
  INV_X1 U19918 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19046) );
  INV_X1 U19919 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20071) );
  AOI22_X1 U19920 ( .A1(n16813), .A2(n19046), .B1(n20071), .B2(n16814), .ZN(
        U371) );
  INV_X1 U19921 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19043) );
  INV_X1 U19922 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20070) );
  AOI22_X1 U19923 ( .A1(n16813), .A2(n19043), .B1(n20070), .B2(n16814), .ZN(
        U372) );
  INV_X1 U19924 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19042) );
  INV_X1 U19925 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20068) );
  AOI22_X1 U19926 ( .A1(n16813), .A2(n19042), .B1(n20068), .B2(n16814), .ZN(
        U373) );
  INV_X1 U19927 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19040) );
  INV_X1 U19928 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20067) );
  AOI22_X1 U19929 ( .A1(n16813), .A2(n19040), .B1(n20067), .B2(n16814), .ZN(
        U374) );
  INV_X1 U19930 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19038) );
  INV_X1 U19931 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U19932 ( .A1(n16813), .A2(n19038), .B1(n20065), .B2(n16814), .ZN(
        U375) );
  INV_X1 U19933 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19017) );
  INV_X1 U19934 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U19935 ( .A1(n16813), .A2(n19017), .B1(n20047), .B2(n16814), .ZN(
        U376) );
  INV_X1 U19936 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18998) );
  NOR2_X1 U19937 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n19014), .ZN(n19001) );
  OAI22_X1 U19938 ( .A1(n18998), .A2(n19001), .B1(n19014), .B2(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18996) );
  INV_X1 U19939 ( .A(n18996), .ZN(n19088) );
  AOI21_X1 U19940 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19088), .ZN(n16815) );
  INV_X1 U19941 ( .A(n16815), .ZN(P3_U2633) );
  INV_X1 U19942 ( .A(n19159), .ZN(n16817) );
  INV_X1 U19943 ( .A(n17724), .ZN(n17665) );
  OAI21_X1 U19944 ( .B1(n16821), .B2(n17665), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16816) );
  OAI21_X1 U19945 ( .B1(n16817), .B2(n19146), .A(n16816), .ZN(P3_U2634) );
  INV_X1 U19946 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19016) );
  AOI21_X1 U19947 ( .B1(n19014), .B2(n19016), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16818) );
  AOI22_X1 U19948 ( .A1(n19083), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16818), 
        .B2(n19155), .ZN(P3_U2635) );
  NOR2_X1 U19949 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16819) );
  OAI21_X1 U19950 ( .B1(n16819), .B2(BS16), .A(n19088), .ZN(n19086) );
  OAI21_X1 U19951 ( .B1(n19088), .B2(n16841), .A(n19086), .ZN(P3_U2636) );
  NOR3_X1 U19952 ( .A1(n16821), .A2(n16820), .A3(n18921), .ZN(n18924) );
  NOR2_X1 U19953 ( .A1(n18924), .A2(n18985), .ZN(n19138) );
  OAI21_X1 U19954 ( .B1(n19138), .B2(n18464), .A(n16822), .ZN(P3_U2637) );
  NOR4_X1 U19955 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16826) );
  NOR4_X1 U19956 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16825) );
  NOR4_X1 U19957 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16824) );
  NOR4_X1 U19958 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16823) );
  NAND4_X1 U19959 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n16823), .ZN(
        n16832) );
  NOR4_X1 U19960 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16830) );
  AOI211_X1 U19961 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16829) );
  NOR4_X1 U19962 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16828) );
  NOR4_X1 U19963 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16827) );
  NAND4_X1 U19964 ( .A1(n16830), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16831) );
  NOR2_X1 U19965 ( .A1(n16832), .A2(n16831), .ZN(n19129) );
  INV_X1 U19966 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16834) );
  NOR3_X1 U19967 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16835) );
  OAI21_X1 U19968 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16835), .A(n19129), .ZN(
        n16833) );
  OAI21_X1 U19969 ( .B1(n19129), .B2(n16834), .A(n16833), .ZN(P3_U2638) );
  INV_X1 U19970 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19018) );
  INV_X1 U19971 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19087) );
  AOI21_X1 U19972 ( .B1(n19018), .B2(n19087), .A(n16835), .ZN(n16837) );
  INV_X1 U19973 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16836) );
  INV_X1 U19974 ( .A(n19129), .ZN(n19126) );
  AOI22_X1 U19975 ( .A1(n19129), .A2(n16837), .B1(n16836), .B2(n19126), .ZN(
        P3_U2639) );
  NAND2_X1 U19976 ( .A1(n19142), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18988) );
  INV_X1 U19977 ( .A(n18988), .ZN(n18982) );
  NAND3_X1 U19978 ( .A1(n19146), .A2(n19142), .A3(n16841), .ZN(n18995) );
  NOR2_X2 U19979 ( .A1(n19100), .A2(n18995), .ZN(n17157) );
  NAND2_X1 U19980 ( .A1(n18407), .A2(n18993), .ZN(n17145) );
  INV_X1 U19981 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19063) );
  INV_X1 U19982 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19041) );
  INV_X1 U19983 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19037) );
  INV_X1 U19984 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19029) );
  INV_X1 U19985 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19025) );
  INV_X1 U19986 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19023) );
  INV_X1 U19987 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19019) );
  NOR2_X1 U19988 ( .A1(n19018), .A2(n19019), .ZN(n17180) );
  NAND2_X1 U19989 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17180), .ZN(n17146) );
  OR2_X1 U19990 ( .A1(n19023), .A2(n17146), .ZN(n17128) );
  NOR2_X1 U19991 ( .A1(n19025), .A2(n17128), .ZN(n17108) );
  NAND2_X1 U19992 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17108), .ZN(n17107) );
  NOR2_X1 U19993 ( .A1(n19029), .A2(n17107), .ZN(n17102) );
  NAND2_X1 U19994 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17102), .ZN(n17101) );
  NAND2_X1 U19995 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17061) );
  NOR3_X1 U19996 ( .A1(n19037), .A2(n17101), .A3(n17061), .ZN(n17051) );
  NAND2_X1 U19997 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17051), .ZN(n17034) );
  NOR2_X1 U19998 ( .A1(n19041), .A2(n17034), .ZN(n17025) );
  NAND2_X1 U19999 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17025), .ZN(n16968) );
  INV_X1 U20000 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19050) );
  NAND2_X1 U20001 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16990) );
  NOR2_X1 U20002 ( .A1(n19050), .A2(n16990), .ZN(n16969) );
  NAND4_X1 U20003 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16969), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16926) );
  NOR2_X1 U20004 ( .A1(n16968), .A2(n16926), .ZN(n16937) );
  NAND4_X1 U20005 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16937), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16917) );
  NOR2_X1 U20006 ( .A1(n19063), .A2(n16917), .ZN(n16912) );
  NAND2_X1 U20007 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16912), .ZN(n16852) );
  NOR2_X1 U20008 ( .A1(n17186), .A2(n16852), .ZN(n16898) );
  NAND3_X1 U20009 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(P3_REIP_REG_26__SCAN_IN), 
        .A3(n16898), .ZN(n16876) );
  NAND2_X1 U20010 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n16838) );
  AOI211_X1 U20011 ( .C1(n18484), .C2(n19005), .A(n19143), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16839) );
  INV_X1 U20012 ( .A(n16839), .ZN(n18977) );
  NOR2_X1 U20013 ( .A1(n17186), .A2(n17160), .ZN(n17027) );
  INV_X1 U20014 ( .A(n17027), .ZN(n17202) );
  OAI21_X1 U20015 ( .B1(n16876), .B2(n16838), .A(n17202), .ZN(n16869) );
  AOI211_X4 U20016 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19141), .A(n16839), .B(
        n19160), .ZN(n17204) );
  AOI22_X1 U20017 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n17171), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17204), .ZN(n16856) );
  NAND2_X1 U20018 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19141), .ZN(n16840) );
  AOI211_X4 U20019 ( .C1(n19151), .C2(n16841), .A(n19160), .B(n16840), .ZN(
        n17203) );
  NOR3_X1 U20020 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17173) );
  INV_X1 U20021 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17501) );
  NAND2_X1 U20022 ( .A1(n17173), .A2(n17501), .ZN(n17166) );
  NOR2_X1 U20023 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17166), .ZN(n17147) );
  NAND2_X1 U20024 ( .A1(n17147), .A2(n17494), .ZN(n17137) );
  NAND2_X1 U20025 ( .A1(n17117), .A2(n17112), .ZN(n17109) );
  INV_X1 U20026 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17090) );
  NAND2_X1 U20027 ( .A1(n17096), .A2(n17090), .ZN(n17089) );
  INV_X1 U20028 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17065) );
  NAND2_X1 U20029 ( .A1(n17073), .A2(n17065), .ZN(n17064) );
  NAND2_X1 U20030 ( .A1(n17047), .A2(n17393), .ZN(n17042) );
  NAND2_X1 U20031 ( .A1(n17029), .A2(n17019), .ZN(n17016) );
  NAND2_X1 U20032 ( .A1(n17004), .A2(n17345), .ZN(n16994) );
  INV_X1 U20033 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16976) );
  NAND2_X1 U20034 ( .A1(n16985), .A2(n16976), .ZN(n16975) );
  INV_X1 U20035 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17301) );
  NAND2_X1 U20036 ( .A1(n16956), .A2(n17301), .ZN(n16952) );
  INV_X1 U20037 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17209) );
  NAND2_X1 U20038 ( .A1(n16940), .A2(n17209), .ZN(n16930) );
  NOR2_X1 U20039 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16930), .ZN(n16921) );
  INV_X1 U20040 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17211) );
  NAND2_X1 U20041 ( .A1(n16921), .A2(n17211), .ZN(n16911) );
  NOR2_X1 U20042 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16911), .ZN(n16899) );
  INV_X1 U20043 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16893) );
  NAND2_X1 U20044 ( .A1(n16899), .A2(n16893), .ZN(n16892) );
  NOR2_X1 U20045 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16892), .ZN(n16879) );
  INV_X1 U20046 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U20047 ( .A1(n16879), .A2(n17214), .ZN(n16857) );
  NOR2_X1 U20048 ( .A1(n17194), .A2(n16857), .ZN(n16864) );
  INV_X1 U20049 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17220) );
  INV_X1 U20050 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17824) );
  NAND2_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17853) );
  INV_X1 U20052 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17899) );
  INV_X1 U20053 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17057) );
  NOR2_X1 U20054 ( .A1(n18128), .A2(n17954), .ZN(n17129) );
  NAND2_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17129), .ZN(
        n17120) );
  NAND2_X1 U20056 ( .A1(n17955), .A2(n17106), .ZN(n17070) );
  NOR2_X1 U20057 ( .A1(n17957), .A2(n17035), .ZN(n17925) );
  NAND2_X1 U20058 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16980), .ZN(
        n16848) );
  NAND2_X1 U20059 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17854), .ZN(
        n16846) );
  NAND2_X1 U20060 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17839), .ZN(
        n16844) );
  NOR2_X1 U20061 ( .A1(n17824), .A2(n16844), .ZN(n16843) );
  NAND2_X1 U20062 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16843), .ZN(
        n17773) );
  NOR2_X1 U20063 ( .A1(n17800), .A2(n17773), .ZN(n16842) );
  OAI21_X1 U20064 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16842), .A(
        n16851), .ZN(n17790) );
  INV_X1 U20065 ( .A(n17790), .ZN(n16887) );
  AOI21_X1 U20066 ( .B1(n17800), .B2(n17773), .A(n16842), .ZN(n17804) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16843), .A(
        n17773), .ZN(n17813) );
  INV_X1 U20068 ( .A(n17813), .ZN(n16908) );
  AOI21_X1 U20069 ( .B1(n17824), .B2(n16844), .A(n16843), .ZN(n17831) );
  OAI21_X1 U20070 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17839), .A(
        n16844), .ZN(n17836) );
  INV_X1 U20071 ( .A(n17836), .ZN(n16929) );
  INV_X1 U20072 ( .A(n16846), .ZN(n16847) );
  NAND2_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16847), .ZN(
        n16845) );
  AOI21_X1 U20074 ( .B1(n10162), .B2(n16845), .A(n17839), .ZN(n17857) );
  OAI22_X1 U20075 ( .A1(n10161), .A2(n16846), .B1(n16847), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17863) );
  INV_X1 U20076 ( .A(n17863), .ZN(n16949) );
  AOI21_X1 U20077 ( .B1(n17876), .B2(n16848), .A(n16847), .ZN(n17879) );
  NOR2_X1 U20078 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17888), .ZN(
        n16979) );
  INV_X1 U20079 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17892) );
  INV_X1 U20080 ( .A(n16980), .ZN(n16850) );
  AOI21_X1 U20081 ( .B1(n17892), .B2(n16850), .A(n17854), .ZN(n17890) );
  NOR2_X1 U20082 ( .A1(n16959), .A2(n17156), .ZN(n16948) );
  NOR2_X1 U20083 ( .A1(n16949), .A2(n16948), .ZN(n16947) );
  NOR2_X1 U20084 ( .A1(n16947), .A2(n17156), .ZN(n16939) );
  NOR2_X1 U20085 ( .A1(n17857), .A2(n16939), .ZN(n16938) );
  NOR2_X1 U20086 ( .A1(n16938), .A2(n17156), .ZN(n16928) );
  NOR2_X1 U20087 ( .A1(n16929), .A2(n16928), .ZN(n16927) );
  NOR2_X1 U20088 ( .A1(n16927), .A2(n17156), .ZN(n16920) );
  NOR2_X1 U20089 ( .A1(n17804), .A2(n16901), .ZN(n16900) );
  NOR2_X1 U20090 ( .A1(n16900), .A2(n17156), .ZN(n16886) );
  NOR2_X1 U20091 ( .A1(n16887), .A2(n16886), .ZN(n16885) );
  NOR2_X1 U20092 ( .A1(n16885), .A2(n17156), .ZN(n16878) );
  AOI21_X1 U20093 ( .B1(n21214), .B2(n16851), .A(n9862), .ZN(n17774) );
  NAND2_X1 U20094 ( .A1(n17130), .A2(n17157), .ZN(n17188) );
  NOR3_X1 U20095 ( .A1(n16860), .A2(n16859), .A3(n17188), .ZN(n16854) );
  INV_X1 U20096 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19070) );
  NOR2_X1 U20097 ( .A1(n17195), .A2(n16852), .ZN(n16897) );
  NAND2_X1 U20098 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16897), .ZN(n16889) );
  NOR2_X1 U20099 ( .A1(n19070), .A2(n16889), .ZN(n16882) );
  NAND3_X1 U20100 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16882), .ZN(n16861) );
  AOI221_X1 U20101 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n19079), .C2(n19077), .A(n16861), .ZN(n16853) );
  AOI211_X1 U20102 ( .C1(n16864), .C2(n17220), .A(n16854), .B(n16853), .ZN(
        n16855) );
  OAI211_X1 U20103 ( .C1(n19079), .C2(n16869), .A(n16856), .B(n16855), .ZN(
        P3_U2640) );
  NAND2_X1 U20104 ( .A1(n17203), .A2(n16857), .ZN(n16874) );
  OAI21_X1 U20105 ( .B1(n16859), .B2(n16860), .A(n17157), .ZN(n16858) );
  AOI21_X1 U20106 ( .B1(n16860), .B2(n16859), .A(n16858), .ZN(n16863) );
  AOI22_X1 U20107 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16869), .B1(n16861), 
        .B2(n19077), .ZN(n16862) );
  OAI21_X1 U20108 ( .B1(n17204), .B2(n16864), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16865) );
  NOR2_X1 U20109 ( .A1(n16879), .A2(n17214), .ZN(n16875) );
  AOI211_X1 U20110 ( .C1(n16868), .C2(n9902), .A(n16867), .B(n18993), .ZN(
        n16871) );
  INV_X1 U20111 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19074) );
  OAI22_X1 U20112 ( .A1(n19074), .A2(n16869), .B1(n17161), .B2(n17214), .ZN(
        n16870) );
  AOI211_X1 U20113 ( .C1(n17171), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16871), .B(n16870), .ZN(n16873) );
  NAND3_X1 U20114 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16882), .A3(n19074), 
        .ZN(n16872) );
  OAI211_X1 U20115 ( .C1(n16875), .C2(n16874), .A(n16873), .B(n16872), .ZN(
        P3_U2642) );
  INV_X1 U20116 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19071) );
  NAND2_X1 U20117 ( .A1(n17202), .A2(n16876), .ZN(n16888) );
  AOI22_X1 U20118 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16884) );
  AOI211_X1 U20119 ( .C1(n17774), .C2(n16878), .A(n16877), .B(n18993), .ZN(
        n16881) );
  AOI211_X1 U20120 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16892), .A(n16879), .B(
        n17194), .ZN(n16880) );
  AOI211_X1 U20121 ( .C1(n16882), .C2(n19071), .A(n16881), .B(n16880), .ZN(
        n16883) );
  OAI211_X1 U20122 ( .C1(n19071), .C2(n16888), .A(n16884), .B(n16883), .ZN(
        P3_U2643) );
  AOI22_X1 U20123 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16896) );
  AOI211_X1 U20124 ( .C1(n16887), .C2(n16886), .A(n16885), .B(n18993), .ZN(
        n16891) );
  AOI21_X1 U20125 ( .B1(n16889), .B2(n19070), .A(n16888), .ZN(n16890) );
  NOR2_X1 U20126 ( .A1(n16891), .A2(n16890), .ZN(n16895) );
  OAI211_X1 U20127 ( .C1(n16899), .C2(n16893), .A(n17203), .B(n16892), .ZN(
        n16894) );
  NAND3_X1 U20128 ( .A1(n16896), .A2(n16895), .A3(n16894), .ZN(P3_U2644) );
  INV_X1 U20129 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19067) );
  AOI22_X1 U20130 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17204), .B1(n16897), 
        .B2(n19067), .ZN(n16905) );
  NOR2_X1 U20131 ( .A1(n17027), .A2(n16898), .ZN(n16910) );
  AOI211_X1 U20132 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16911), .A(n16899), .B(
        n17194), .ZN(n16903) );
  AOI211_X1 U20133 ( .C1(n17804), .C2(n16901), .A(n16900), .B(n18993), .ZN(
        n16902) );
  AOI211_X1 U20134 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16910), .A(n16903), 
        .B(n16902), .ZN(n16904) );
  OAI211_X1 U20135 ( .C1(n17800), .C2(n17187), .A(n16905), .B(n16904), .ZN(
        P3_U2645) );
  AOI22_X1 U20136 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16916) );
  AOI211_X1 U20137 ( .C1(n16908), .C2(n16907), .A(n16906), .B(n18993), .ZN(
        n16909) );
  AOI21_X1 U20138 ( .B1(n16910), .B2(P3_REIP_REG_25__SCAN_IN), .A(n16909), 
        .ZN(n16915) );
  OAI211_X1 U20139 ( .C1(n16921), .C2(n17211), .A(n17203), .B(n16911), .ZN(
        n16914) );
  INV_X1 U20140 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19065) );
  NAND3_X1 U20141 ( .A1(n17160), .A2(n16912), .A3(n19065), .ZN(n16913) );
  NAND4_X1 U20142 ( .A1(n16916), .A2(n16915), .A3(n16914), .A4(n16913), .ZN(
        P3_U2646) );
  AOI21_X1 U20143 ( .B1(n17160), .B2(n16917), .A(n17186), .ZN(n16935) );
  NOR3_X1 U20144 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17195), .A3(n16917), 
        .ZN(n16918) );
  AOI21_X1 U20145 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17204), .A(n16918), .ZN(
        n16925) );
  AOI211_X1 U20146 ( .C1(n17831), .C2(n16920), .A(n16919), .B(n18993), .ZN(
        n16923) );
  AOI211_X1 U20147 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16930), .A(n16921), .B(
        n17194), .ZN(n16922) );
  AOI211_X1 U20148 ( .C1(n17171), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16923), .B(n16922), .ZN(n16924) );
  OAI211_X1 U20149 ( .C1(n16935), .C2(n19063), .A(n16925), .B(n16924), .ZN(
        P3_U2647) );
  NAND3_X1 U20150 ( .A1(n17160), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n17025), 
        .ZN(n17003) );
  NOR2_X1 U20151 ( .A1(n16926), .A2(n17003), .ZN(n16951) );
  NAND3_X1 U20152 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16951), .ZN(n16936) );
  INV_X1 U20153 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19062) );
  AOI211_X1 U20154 ( .C1(n16929), .C2(n16928), .A(n16927), .B(n18993), .ZN(
        n16933) );
  OAI211_X1 U20155 ( .C1(n16940), .C2(n17209), .A(n17203), .B(n16930), .ZN(
        n16931) );
  OAI21_X1 U20156 ( .B1(n17209), .B2(n17161), .A(n16931), .ZN(n16932) );
  AOI211_X1 U20157 ( .C1(n17171), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16933), .B(n16932), .ZN(n16934) );
  OAI221_X1 U20158 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16936), .C1(n19062), 
        .C2(n16935), .A(n16934), .ZN(P3_U2648) );
  NAND2_X1 U20159 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16951), .ZN(n16946) );
  INV_X1 U20160 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19059) );
  INV_X1 U20161 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19057) );
  OAI21_X1 U20162 ( .B1(n16937), .B2(n17195), .A(n17205), .ZN(n16963) );
  AOI21_X1 U20163 ( .B1(n16951), .B2(n19057), .A(n16963), .ZN(n16945) );
  AOI211_X1 U20164 ( .C1(n17857), .C2(n16939), .A(n16938), .B(n18993), .ZN(
        n16943) );
  AOI211_X1 U20165 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16952), .A(n16940), .B(
        n17194), .ZN(n16942) );
  OAI22_X1 U20166 ( .A1(n10162), .A2(n17187), .B1(n17161), .B2(n17213), .ZN(
        n16941) );
  NOR3_X1 U20167 ( .A1(n16943), .A2(n16942), .A3(n16941), .ZN(n16944) );
  OAI221_X1 U20168 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n16946), .C1(n19059), 
        .C2(n16945), .A(n16944), .ZN(P3_U2649) );
  AOI22_X1 U20169 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16955) );
  AOI211_X1 U20170 ( .C1(n16949), .C2(n16948), .A(n16947), .B(n18993), .ZN(
        n16950) );
  AOI221_X1 U20171 ( .B1(n16963), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16951), 
        .C2(n19057), .A(n16950), .ZN(n16954) );
  OAI211_X1 U20172 ( .C1(n16956), .C2(n17301), .A(n17203), .B(n16952), .ZN(
        n16953) );
  NAND3_X1 U20173 ( .A1(n16955), .A2(n16954), .A3(n16953), .ZN(P3_U2650) );
  AOI211_X1 U20174 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16975), .A(n16956), .B(
        n17194), .ZN(n16957) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17204), .A(n16957), .ZN(
        n16965) );
  NAND2_X1 U20176 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16958) );
  INV_X1 U20177 ( .A(n17003), .ZN(n17015) );
  NAND2_X1 U20178 ( .A1(n16969), .A2(n17015), .ZN(n16984) );
  NOR2_X1 U20179 ( .A1(n16958), .A2(n16984), .ZN(n16962) );
  INV_X1 U20180 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19056) );
  AOI211_X1 U20181 ( .C1(n17879), .C2(n16960), .A(n16959), .B(n18993), .ZN(
        n16961) );
  AOI221_X1 U20182 ( .B1(n16963), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16962), 
        .C2(n19056), .A(n16961), .ZN(n16964) );
  OAI211_X1 U20183 ( .C1(n17876), .C2(n17187), .A(n16965), .B(n16964), .ZN(
        P3_U2651) );
  AOI211_X1 U20184 ( .C1(n17890), .C2(n16967), .A(n16966), .B(n18993), .ZN(
        n16974) );
  OAI21_X1 U20185 ( .B1(n17161), .B2(n16976), .A(n18407), .ZN(n16973) );
  INV_X1 U20186 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19051) );
  NOR2_X1 U20187 ( .A1(n19051), .A2(n16984), .ZN(n16971) );
  NOR2_X1 U20188 ( .A1(n17186), .A2(n16968), .ZN(n17026) );
  AOI21_X1 U20189 ( .B1(n16969), .B2(n17026), .A(n17027), .ZN(n16999) );
  AOI21_X1 U20190 ( .B1(n17202), .B2(n19051), .A(n16999), .ZN(n16983) );
  INV_X1 U20191 ( .A(n16983), .ZN(n16970) );
  MUX2_X1 U20192 ( .A(n16971), .B(n16970), .S(P3_REIP_REG_19__SCAN_IN), .Z(
        n16972) );
  NOR3_X1 U20193 ( .A1(n16974), .A2(n16973), .A3(n16972), .ZN(n16978) );
  OAI211_X1 U20194 ( .C1(n16985), .C2(n16976), .A(n17203), .B(n16975), .ZN(
        n16977) );
  OAI211_X1 U20195 ( .C1(n17187), .C2(n17892), .A(n16978), .B(n16977), .ZN(
        P3_U2652) );
  NOR2_X1 U20196 ( .A1(n16979), .A2(n17156), .ZN(n16981) );
  AOI21_X1 U20197 ( .B1(n17899), .B2(n17888), .A(n16980), .ZN(n17902) );
  XOR2_X1 U20198 ( .A(n16981), .B(n17902), .Z(n16982) );
  AOI21_X1 U20199 ( .B1(n16982), .B2(n17157), .A(n18446), .ZN(n16989) );
  AOI21_X1 U20200 ( .B1(n19051), .B2(n16984), .A(n16983), .ZN(n16987) );
  AOI211_X1 U20201 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16994), .A(n16985), .B(
        n17194), .ZN(n16986) );
  AOI211_X1 U20202 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17204), .A(n16987), .B(
        n16986), .ZN(n16988) );
  OAI211_X1 U20203 ( .C1(n17899), .C2(n17187), .A(n16989), .B(n16988), .ZN(
        P3_U2653) );
  OAI21_X1 U20204 ( .B1(n16990), .B2(n17003), .A(n19050), .ZN(n16998) );
  OAI21_X1 U20205 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16991), .A(
        n17888), .ZN(n17911) );
  NAND2_X1 U20206 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17925), .ZN(
        n17011) );
  OAI21_X1 U20207 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17011), .A(
        n17130), .ZN(n17012) );
  INV_X1 U20208 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17922) );
  AOI21_X1 U20209 ( .B1(n17922), .B2(n17011), .A(n16991), .ZN(n17926) );
  INV_X1 U20210 ( .A(n17926), .ZN(n17002) );
  NAND2_X1 U20211 ( .A1(n17012), .A2(n17002), .ZN(n17001) );
  NAND2_X1 U20212 ( .A1(n17130), .A2(n17001), .ZN(n16993) );
  AOI21_X1 U20213 ( .B1(n17911), .B2(n16993), .A(n18993), .ZN(n16992) );
  OAI21_X1 U20214 ( .B1(n17911), .B2(n16993), .A(n16992), .ZN(n16996) );
  OAI211_X1 U20215 ( .C1(n17004), .C2(n17345), .A(n17203), .B(n16994), .ZN(
        n16995) );
  OAI211_X1 U20216 ( .C1(n17187), .C2(n17909), .A(n16996), .B(n16995), .ZN(
        n16997) );
  AOI21_X1 U20217 ( .B1(n16999), .B2(n16998), .A(n16997), .ZN(n17000) );
  OAI211_X1 U20218 ( .C1(n17161), .C2(n17345), .A(n17000), .B(n18407), .ZN(
        P3_U2654) );
  OAI21_X1 U20219 ( .B1(n17012), .B2(n17002), .A(n17001), .ZN(n17010) );
  AOI21_X1 U20220 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17026), .A(n17027), 
        .ZN(n17014) );
  INV_X1 U20221 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19045) );
  NOR3_X1 U20222 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19045), .A3(n17003), 
        .ZN(n17008) );
  AOI211_X1 U20223 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17016), .A(n17004), .B(
        n17194), .ZN(n17005) );
  AOI21_X1 U20224 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17204), .A(n17005), .ZN(
        n17006) );
  OAI21_X1 U20225 ( .B1(n17922), .B2(n17187), .A(n17006), .ZN(n17007) );
  AOI211_X1 U20226 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n17014), .A(n17008), 
        .B(n17007), .ZN(n17009) );
  OAI211_X1 U20227 ( .C1(n18993), .C2(n17010), .A(n17009), .B(n18407), .ZN(
        P3_U2655) );
  INV_X1 U20228 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17938) );
  OAI21_X1 U20229 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17925), .A(
        n17011), .ZN(n17951) );
  INV_X1 U20230 ( .A(n17951), .ZN(n17013) );
  NOR3_X1 U20231 ( .A1(n17013), .A2(n17012), .A3(n18993), .ZN(n17022) );
  INV_X1 U20232 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17189) );
  OAI21_X1 U20233 ( .B1(n17156), .B2(n17189), .A(n17157), .ZN(n17192) );
  AOI211_X1 U20234 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17130), .A(
        n17951), .B(n17192), .ZN(n17021) );
  OAI21_X1 U20235 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17015), .A(n17014), 
        .ZN(n17018) );
  OAI211_X1 U20236 ( .C1(n17029), .C2(n17019), .A(n17203), .B(n17016), .ZN(
        n17017) );
  OAI211_X1 U20237 ( .C1(n17019), .C2(n17161), .A(n17018), .B(n17017), .ZN(
        n17020) );
  NOR4_X1 U20238 ( .A1(n18446), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17023) );
  OAI21_X1 U20239 ( .B1(n17938), .B2(n17187), .A(n17023), .ZN(P3_U2656) );
  AOI21_X1 U20240 ( .B1(n17957), .B2(n17035), .A(n17925), .ZN(n17959) );
  OAI21_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17035), .A(
        n17130), .ZN(n17037) );
  XNOR2_X1 U20242 ( .A(n17959), .B(n17037), .ZN(n17024) );
  AOI21_X1 U20243 ( .B1(n17157), .B2(n17024), .A(n18446), .ZN(n17033) );
  INV_X1 U20244 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19044) );
  NAND2_X1 U20245 ( .A1(n17160), .A2(n17025), .ZN(n17028) );
  AOI211_X1 U20246 ( .C1(n19044), .C2(n17028), .A(n17027), .B(n17026), .ZN(
        n17031) );
  AOI211_X1 U20247 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17042), .A(n17029), .B(
        n17194), .ZN(n17030) );
  AOI211_X1 U20248 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17204), .A(n17031), .B(
        n17030), .ZN(n17032) );
  OAI211_X1 U20249 ( .C1(n17957), .C2(n17187), .A(n17033), .B(n17032), .ZN(
        P3_U2657) );
  AOI22_X1 U20250 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17046) );
  NOR3_X1 U20251 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17195), .A3(n17034), 
        .ZN(n17041) );
  INV_X1 U20252 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17987) );
  NOR2_X1 U20253 ( .A1(n17987), .A2(n17055), .ZN(n17036) );
  OAI21_X1 U20254 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17036), .A(
        n17035), .ZN(n17975) );
  INV_X1 U20255 ( .A(n17975), .ZN(n17038) );
  NOR3_X1 U20256 ( .A1(n17038), .A2(n18993), .A3(n17037), .ZN(n17040) );
  AOI211_X1 U20257 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17130), .A(
        n17975), .B(n17192), .ZN(n17039) );
  NOR4_X1 U20258 ( .A1(n18446), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17045) );
  OAI21_X1 U20259 ( .B1(n17051), .B2(n17195), .A(n17205), .ZN(n17063) );
  NOR2_X1 U20260 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17195), .ZN(n17050) );
  OAI21_X1 U20261 ( .B1(n17063), .B2(n17050), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n17044) );
  OAI211_X1 U20262 ( .C1(n17047), .C2(n17393), .A(n17203), .B(n17042), .ZN(
        n17043) );
  NAND4_X1 U20263 ( .A1(n17046), .A2(n17045), .A3(n17044), .A4(n17043), .ZN(
        P3_U2658) );
  AOI211_X1 U20264 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17064), .A(n17047), .B(
        n17194), .ZN(n17048) );
  AOI21_X1 U20265 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17204), .A(n17048), .ZN(
        n17054) );
  OAI21_X1 U20266 ( .B1(n17055), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17130), .ZN(n17059) );
  AOI22_X1 U20267 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17055), .B1(
        n17969), .B2(n17987), .ZN(n17984) );
  XOR2_X1 U20268 ( .A(n17059), .B(n17984), .Z(n17049) );
  AOI22_X1 U20269 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17171), .B1(
        n17157), .B2(n17049), .ZN(n17053) );
  AOI22_X1 U20270 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17063), .B1(n17051), 
        .B2(n17050), .ZN(n17052) );
  NAND4_X1 U20271 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n18407), .ZN(
        P3_U2659) );
  INV_X1 U20272 ( .A(n17070), .ZN(n17056) );
  OAI21_X1 U20273 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17056), .A(
        n17055), .ZN(n18005) );
  NOR2_X1 U20274 ( .A1(n18993), .A2(n17130), .ZN(n17179) );
  INV_X1 U20275 ( .A(n17179), .ZN(n17148) );
  OAI221_X1 U20276 ( .B1(n18005), .B2(n17057), .C1(n18005), .C2(n17189), .A(
        n17157), .ZN(n17058) );
  AOI22_X1 U20277 ( .A1(n18005), .A2(n17059), .B1(n17148), .B2(n17058), .ZN(
        n17060) );
  AOI211_X1 U20278 ( .C1(n17204), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18446), .B(
        n17060), .ZN(n17068) );
  OR2_X1 U20279 ( .A1(n17195), .A2(n17101), .ZN(n17087) );
  OAI21_X1 U20280 ( .B1(n17061), .B2(n17087), .A(n19037), .ZN(n17062) );
  AOI22_X1 U20281 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17171), .B1(
        n17063), .B2(n17062), .ZN(n17067) );
  OAI211_X1 U20282 ( .C1(n17073), .C2(n17065), .A(n17203), .B(n17064), .ZN(
        n17066) );
  NAND3_X1 U20283 ( .A1(n17068), .A2(n17067), .A3(n17066), .ZN(P3_U2660) );
  NOR2_X1 U20284 ( .A1(n17069), .A2(n17120), .ZN(n17080) );
  OAI21_X1 U20285 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17080), .A(
        n17070), .ZN(n18021) );
  NAND2_X1 U20286 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17106), .ZN(
        n17105) );
  NOR3_X1 U20287 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21294), .A3(
        n17105), .ZN(n17082) );
  AOI21_X1 U20288 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17082), .A(
        n17156), .ZN(n17071) );
  INV_X1 U20289 ( .A(n17071), .ZN(n17084) );
  XOR2_X1 U20290 ( .A(n18021), .B(n17084), .Z(n17072) );
  AOI21_X1 U20291 ( .B1(n17072), .B2(n17157), .A(n18446), .ZN(n17079) );
  AOI211_X1 U20292 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17089), .A(n17073), .B(
        n17194), .ZN(n17077) );
  INV_X1 U20293 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19033) );
  NOR2_X1 U20294 ( .A1(n19033), .A2(n17087), .ZN(n17075) );
  AOI221_X1 U20295 ( .B1(n17101), .B2(n17160), .C1(n19033), .C2(n17160), .A(
        n17186), .ZN(n17086) );
  INV_X1 U20296 ( .A(n17086), .ZN(n17074) );
  MUX2_X1 U20297 ( .A(n17075), .B(n17074), .S(P3_REIP_REG_10__SCAN_IN), .Z(
        n17076) );
  AOI211_X1 U20298 ( .C1(n17171), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17077), .B(n17076), .ZN(n17078) );
  OAI211_X1 U20299 ( .C1(n17161), .C2(n17432), .A(n17079), .B(n17078), .ZN(
        P3_U2661) );
  AND2_X1 U20300 ( .A1(n18041), .A2(n17106), .ZN(n17094) );
  INV_X1 U20301 ( .A(n17080), .ZN(n17081) );
  OAI21_X1 U20302 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17094), .A(
        n17081), .ZN(n18027) );
  OAI21_X1 U20303 ( .B1(n17082), .B2(n18027), .A(n17157), .ZN(n17083) );
  AOI22_X1 U20304 ( .A1(n18027), .A2(n17084), .B1(n17148), .B2(n17083), .ZN(
        n17085) );
  AOI211_X1 U20305 ( .C1(n17204), .C2(P3_EBX_REG_9__SCAN_IN), .A(n18446), .B(
        n17085), .ZN(n17093) );
  AOI21_X1 U20306 ( .B1(n19033), .B2(n17087), .A(n17086), .ZN(n17088) );
  AOI21_X1 U20307 ( .B1(n17171), .B2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17088), .ZN(n17092) );
  OAI211_X1 U20308 ( .C1(n17096), .C2(n17090), .A(n17203), .B(n17089), .ZN(
        n17091) );
  NAND3_X1 U20309 ( .A1(n17093), .A2(n17092), .A3(n17091), .ZN(P3_U2662) );
  AOI21_X1 U20310 ( .B1(n21294), .B2(n17105), .A(n17094), .ZN(n18043) );
  OAI21_X1 U20311 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17105), .A(
        n17130), .ZN(n17095) );
  XNOR2_X1 U20312 ( .A(n18043), .B(n17095), .ZN(n17100) );
  AOI211_X1 U20313 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17109), .A(n17096), .B(
        n17194), .ZN(n17099) );
  INV_X1 U20314 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19032) );
  AOI22_X1 U20315 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n17097) );
  OAI211_X1 U20316 ( .C1(n17205), .C2(n19032), .A(n17097), .B(n18407), .ZN(
        n17098) );
  AOI211_X1 U20317 ( .C1(n17157), .C2(n17100), .A(n17099), .B(n17098), .ZN(
        n17104) );
  OAI211_X1 U20318 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n17102), .A(n17160), .B(
        n17101), .ZN(n17103) );
  NAND2_X1 U20319 ( .A1(n17104), .A2(n17103), .ZN(P3_U2663) );
  OAI21_X1 U20320 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17106), .A(
        n17105), .ZN(n18057) );
  INV_X1 U20321 ( .A(n18038), .ZN(n18039) );
  NAND2_X1 U20322 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17189), .ZN(
        n17175) );
  OAI21_X1 U20323 ( .B1(n18039), .B2(n17175), .A(n17130), .ZN(n17119) );
  XNOR2_X1 U20324 ( .A(n18057), .B(n17119), .ZN(n17116) );
  NOR3_X1 U20325 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17195), .A3(n17107), .ZN(
        n17114) );
  INV_X1 U20326 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19027) );
  AND3_X1 U20327 ( .A1(n19027), .A2(n17160), .A3(n17108), .ZN(n17122) );
  OAI21_X1 U20328 ( .B1(n17108), .B2(n17195), .A(n17205), .ZN(n17136) );
  OAI21_X1 U20329 ( .B1(n17122), .B2(n17136), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n17111) );
  OAI211_X1 U20330 ( .C1(n17117), .C2(n17112), .A(n17203), .B(n17109), .ZN(
        n17110) );
  OAI211_X1 U20331 ( .C1(n17112), .C2(n17161), .A(n17111), .B(n17110), .ZN(
        n17113) );
  AOI211_X1 U20332 ( .C1(n17171), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17114), .B(n17113), .ZN(n17115) );
  OAI211_X1 U20333 ( .C1(n18993), .C2(n17116), .A(n17115), .B(n18407), .ZN(
        P3_U2664) );
  AOI211_X1 U20334 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17137), .A(n17117), .B(
        n17194), .ZN(n17118) );
  AOI21_X1 U20335 ( .B1(n17171), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17118), .ZN(n17127) );
  NOR2_X1 U20336 ( .A1(n18993), .A2(n17119), .ZN(n17124) );
  OAI21_X1 U20337 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17129), .A(
        n17120), .ZN(n18071) );
  INV_X1 U20338 ( .A(n17129), .ZN(n17121) );
  AOI211_X1 U20339 ( .C1(n17130), .C2(n17121), .A(n18071), .B(n17192), .ZN(
        n17123) );
  AOI211_X1 U20340 ( .C1(n17124), .C2(n18071), .A(n17123), .B(n17122), .ZN(
        n17126) );
  AOI22_X1 U20341 ( .A1(n17204), .A2(P3_EBX_REG_6__SCAN_IN), .B1(
        P3_REIP_REG_6__SCAN_IN), .B2(n17136), .ZN(n17125) );
  NAND4_X1 U20342 ( .A1(n17127), .A2(n17126), .A3(n17125), .A4(n18407), .ZN(
        P3_U2665) );
  INV_X1 U20343 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17140) );
  OAI21_X1 U20344 ( .B1(n17195), .B2(n17128), .A(n19025), .ZN(n17135) );
  NAND2_X1 U20345 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18085), .ZN(
        n17141) );
  AOI21_X1 U20346 ( .B1(n17140), .B2(n17141), .A(n17129), .ZN(n18083) );
  OAI21_X1 U20347 ( .B1(n17141), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17130), .ZN(n17131) );
  INV_X1 U20348 ( .A(n17131), .ZN(n17142) );
  INV_X1 U20349 ( .A(n18083), .ZN(n17132) );
  OAI221_X1 U20350 ( .B1(n18083), .B2(n17142), .C1(n17132), .C2(n17131), .A(
        n17157), .ZN(n17133) );
  OAI211_X1 U20351 ( .C1(n17161), .C2(n17494), .A(n18407), .B(n17133), .ZN(
        n17134) );
  AOI21_X1 U20352 ( .B1(n17136), .B2(n17135), .A(n17134), .ZN(n17139) );
  OAI211_X1 U20353 ( .C1(n17147), .C2(n17494), .A(n17203), .B(n17137), .ZN(
        n17138) );
  OAI211_X1 U20354 ( .C1(n17187), .C2(n17140), .A(n17139), .B(n17138), .ZN(
        P3_U2666) );
  AOI21_X1 U20355 ( .B1(n17160), .B2(n17146), .A(n17186), .ZN(n17162) );
  OR2_X1 U20356 ( .A1(n18088), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18093) );
  NOR2_X1 U20357 ( .A1(n18128), .A2(n18088), .ZN(n17155) );
  OAI21_X1 U20358 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17155), .A(
        n17141), .ZN(n18096) );
  AOI21_X1 U20359 ( .B1(n17142), .B2(n18096), .A(n18446), .ZN(n17143) );
  OAI21_X1 U20360 ( .B1(n18093), .B2(n17175), .A(n17143), .ZN(n17144) );
  AOI22_X1 U20361 ( .A1(n17204), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n17145), .B2(
        n17144), .ZN(n17154) );
  NOR3_X1 U20362 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17195), .A3(n17146), .ZN(
        n17152) );
  AOI211_X1 U20363 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17166), .A(n17147), .B(
        n17194), .ZN(n17151) );
  NOR2_X1 U20364 ( .A1(n17666), .A2(n19158), .ZN(n17201) );
  INV_X1 U20365 ( .A(n17201), .ZN(n17191) );
  AOI21_X1 U20366 ( .B1(n15718), .B2(n18926), .A(n17191), .ZN(n17150) );
  OAI22_X1 U20367 ( .A1(n18100), .A2(n17187), .B1(n18096), .B2(n17148), .ZN(
        n17149) );
  NOR4_X1 U20368 ( .A1(n17152), .A2(n17151), .A3(n17150), .A4(n17149), .ZN(
        n17153) );
  OAI211_X1 U20369 ( .C1(n19023), .C2(n17162), .A(n17154), .B(n17153), .ZN(
        P3_U2667) );
  INV_X1 U20370 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17169) );
  NOR2_X1 U20371 ( .A1(n19114), .A2(n19108), .ZN(n18944) );
  NAND2_X1 U20372 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18944), .ZN(
        n18935) );
  AOI21_X1 U20373 ( .B1(n19096), .B2(n18935), .A(n17379), .ZN(n19092) );
  NAND2_X1 U20374 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17172) );
  AOI21_X1 U20375 ( .B1(n17169), .B2(n17172), .A(n17155), .ZN(n18110) );
  NOR2_X1 U20376 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17172), .ZN(
        n17174) );
  NOR2_X1 U20377 ( .A1(n17156), .A2(n17174), .ZN(n17159) );
  OAI21_X1 U20378 ( .B1(n18110), .B2(n17159), .A(n17157), .ZN(n17158) );
  AOI21_X1 U20379 ( .B1(n18110), .B2(n17159), .A(n17158), .ZN(n17165) );
  AOI21_X1 U20380 ( .B1(n17160), .B2(n17180), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n17163) );
  OAI22_X1 U20381 ( .A1(n17163), .A2(n17162), .B1(n17161), .B2(n17501), .ZN(
        n17164) );
  AOI211_X1 U20382 ( .C1(n17201), .C2(n19092), .A(n17165), .B(n17164), .ZN(
        n17168) );
  OAI211_X1 U20383 ( .C1(n17173), .C2(n17501), .A(n17203), .B(n17166), .ZN(
        n17167) );
  OAI211_X1 U20384 ( .C1(n17187), .C2(n17169), .A(n17168), .B(n17167), .ZN(
        P3_U2668) );
  NAND2_X1 U20385 ( .A1(n18939), .A2(n19108), .ZN(n18930) );
  NAND2_X1 U20386 ( .A1(n18935), .A2(n18930), .ZN(n19101) );
  OAI22_X1 U20387 ( .A1(n17205), .A2(n19019), .B1(n19101), .B2(n17191), .ZN(
        n17170) );
  INV_X1 U20388 ( .A(n17170), .ZN(n17185) );
  AOI22_X1 U20389 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17171), .B1(
        n17204), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20390 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17172), .ZN(n18118) );
  INV_X1 U20391 ( .A(n18118), .ZN(n17178) );
  INV_X1 U20392 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17519) );
  INV_X1 U20393 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17513) );
  NAND2_X1 U20394 ( .A1(n17519), .A2(n17513), .ZN(n17193) );
  AOI211_X1 U20395 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17193), .A(n17173), .B(
        n17194), .ZN(n17177) );
  AOI211_X1 U20396 ( .C1(n17178), .C2(n17175), .A(n17174), .B(n17188), .ZN(
        n17176) );
  AOI211_X1 U20397 ( .C1(n17179), .C2(n17178), .A(n17177), .B(n17176), .ZN(
        n17183) );
  AOI211_X1 U20398 ( .C1(n19018), .C2(n19019), .A(n17195), .B(n17180), .ZN(
        n17181) );
  INV_X1 U20399 ( .A(n17181), .ZN(n17182) );
  NAND4_X1 U20400 ( .A1(n17185), .A2(n17184), .A3(n17183), .A4(n17182), .ZN(
        P3_U2669) );
  AOI22_X1 U20401 ( .A1(n17204), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17186), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17200) );
  OAI21_X1 U20402 ( .B1(n17189), .B2(n17188), .A(n17187), .ZN(n17198) );
  NOR2_X1 U20403 ( .A1(n18942), .A2(n17190), .ZN(n19111) );
  INV_X1 U20404 ( .A(n19111), .ZN(n18954) );
  OAI22_X1 U20405 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17192), .B1(
        n17191), .B2(n18954), .ZN(n17197) );
  NAND2_X1 U20406 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17506) );
  NAND2_X1 U20407 ( .A1(n17193), .A2(n17506), .ZN(n17514) );
  OAI22_X1 U20408 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17195), .B1(n17194), 
        .B2(n17514), .ZN(n17196) );
  AOI211_X1 U20409 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17198), .A(
        n17197), .B(n17196), .ZN(n17199) );
  NAND2_X1 U20410 ( .A1(n17200), .A2(n17199), .ZN(P3_U2670) );
  AOI22_X1 U20411 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17202), .B1(n17201), 
        .B2(n19121), .ZN(n17208) );
  OAI21_X1 U20412 ( .B1(n17204), .B2(n17203), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17207) );
  NAND3_X1 U20413 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19103), .A3(
        n17205), .ZN(n17206) );
  NAND3_X1 U20414 ( .A1(n17208), .A2(n17207), .A3(n17206), .ZN(P3_U2671) );
  NOR4_X1 U20415 ( .A1(n17212), .A2(n17211), .A3(n17210), .A4(n17209), .ZN(
        n17216) );
  NAND3_X1 U20416 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17319), .ZN(n17300) );
  NOR4_X1 U20417 ( .A1(n17214), .A2(n17213), .A3(n17301), .A4(n17300), .ZN(
        n17215) );
  NAND4_X1 U20418 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17216), .A4(n17215), .ZN(n17219) );
  NAND2_X1 U20419 ( .A1(n17511), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17218) );
  NAND2_X1 U20420 ( .A1(n17247), .A2(n18511), .ZN(n17217) );
  OAI22_X1 U20421 ( .A1(n17247), .A2(n17218), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17217), .ZN(P3_U2672) );
  NAND2_X1 U20422 ( .A1(n17220), .A2(n17219), .ZN(n17221) );
  NAND2_X1 U20423 ( .A1(n17221), .A2(n17511), .ZN(n17246) );
  AOI22_X1 U20424 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17222) );
  OAI21_X1 U20425 ( .B1(n9947), .B2(n17380), .A(n17222), .ZN(n17232) );
  AOI22_X1 U20426 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17229) );
  INV_X1 U20427 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18821) );
  OAI22_X1 U20428 ( .A1(n17381), .A2(n21259), .B1(n17427), .B2(n18821), .ZN(
        n17227) );
  AOI22_X1 U20429 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20430 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20431 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17223) );
  NAND3_X1 U20432 ( .A1(n17225), .A2(n17224), .A3(n17223), .ZN(n17226) );
  AOI211_X1 U20433 ( .C1(n13961), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17227), .B(n17226), .ZN(n17228) );
  OAI211_X1 U20434 ( .C1(n17230), .C2(n21319), .A(n17229), .B(n17228), .ZN(
        n17231) );
  AOI211_X1 U20435 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17232), .B(n17231), .ZN(n17250) );
  NOR2_X1 U20436 ( .A1(n17250), .A2(n17249), .ZN(n17245) );
  AOI22_X1 U20437 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20438 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20439 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17233) );
  OAI211_X1 U20440 ( .C1(n13976), .C2(n17235), .A(n17234), .B(n17233), .ZN(
        n17241) );
  AOI22_X1 U20441 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20442 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20443 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U20444 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n17236) );
  NAND4_X1 U20445 ( .A1(n17239), .A2(n17238), .A3(n17237), .A4(n17236), .ZN(
        n17240) );
  AOI211_X1 U20446 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17241), .B(n17240), .ZN(n17242) );
  OAI211_X1 U20447 ( .C1(n9947), .C2(n21325), .A(n17243), .B(n17242), .ZN(
        n17244) );
  XNOR2_X1 U20448 ( .A(n17245), .B(n17244), .ZN(n17528) );
  OAI22_X1 U20449 ( .A1(n17247), .A2(n17246), .B1(n17528), .B2(n17511), .ZN(
        P3_U2673) );
  INV_X1 U20450 ( .A(n17248), .ZN(n17255) );
  NAND2_X1 U20451 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17255), .ZN(n17252) );
  XNOR2_X1 U20452 ( .A(n17250), .B(n17249), .ZN(n17536) );
  NAND3_X1 U20453 ( .A1(n17252), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17511), 
        .ZN(n17251) );
  OAI221_X1 U20454 ( .B1(n17252), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17511), 
        .C2(n17536), .A(n17251), .ZN(P3_U2674) );
  AOI21_X1 U20455 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17511), .A(n17261), .ZN(
        n17254) );
  XNOR2_X1 U20456 ( .A(n17253), .B(n17257), .ZN(n17545) );
  OAI22_X1 U20457 ( .A1(n17255), .A2(n17254), .B1(n17511), .B2(n17545), .ZN(
        P3_U2676) );
  INV_X1 U20458 ( .A(n17256), .ZN(n17264) );
  AOI21_X1 U20459 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17511), .A(n17264), .ZN(
        n17260) );
  OAI21_X1 U20460 ( .B1(n17259), .B2(n17258), .A(n17257), .ZN(n17549) );
  OAI22_X1 U20461 ( .A1(n17261), .A2(n17260), .B1(n17511), .B2(n17549), .ZN(
        P3_U2677) );
  AOI21_X1 U20462 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17511), .A(n17270), .ZN(
        n17263) );
  XNOR2_X1 U20463 ( .A(n17262), .B(n17266), .ZN(n17553) );
  OAI22_X1 U20464 ( .A1(n17264), .A2(n17263), .B1(n17511), .B2(n17553), .ZN(
        P3_U2678) );
  INV_X1 U20465 ( .A(n17265), .ZN(n17274) );
  AOI21_X1 U20466 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17511), .A(n17274), .ZN(
        n17269) );
  OAI21_X1 U20467 ( .B1(n17268), .B2(n17267), .A(n17266), .ZN(n17558) );
  OAI22_X1 U20468 ( .A1(n17270), .A2(n17269), .B1(n17511), .B2(n17558), .ZN(
        P3_U2679) );
  AOI21_X1 U20469 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17511), .A(n9929), .ZN(
        n17273) );
  XNOR2_X1 U20470 ( .A(n17272), .B(n17271), .ZN(n17563) );
  OAI22_X1 U20471 ( .A1(n17274), .A2(n17273), .B1(n17511), .B2(n17563), .ZN(
        P3_U2680) );
  AOI22_X1 U20472 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U20473 ( .B1(n9875), .B2(n18821), .A(n17275), .ZN(n17285) );
  AOI22_X1 U20474 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17283) );
  INV_X1 U20475 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20476 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15875), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20477 ( .B1(n17473), .B2(n17277), .A(n17276), .ZN(n17281) );
  AOI22_X1 U20478 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U20479 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17278) );
  OAI211_X1 U20480 ( .C1(n13976), .C2(n21259), .A(n17279), .B(n17278), .ZN(
        n17280) );
  AOI211_X1 U20481 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17281), .B(n17280), .ZN(n17282) );
  OAI211_X1 U20482 ( .C1(n13975), .C2(n21319), .A(n17283), .B(n17282), .ZN(
        n17284) );
  AOI211_X1 U20483 ( .C1(n17349), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17285), .B(n17284), .ZN(n17565) );
  NAND3_X1 U20484 ( .A1(n17287), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17511), 
        .ZN(n17286) );
  OAI221_X1 U20485 ( .B1(n17287), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17511), 
        .C2(n17565), .A(n17286), .ZN(P3_U2681) );
  AOI22_X1 U20486 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17288) );
  OAI21_X1 U20487 ( .B1(n17483), .B2(n17289), .A(n17288), .ZN(n17299) );
  AOI22_X1 U20488 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17296) );
  OAI22_X1 U20489 ( .A1(n13975), .A2(n18716), .B1(n17381), .B2(n17495), .ZN(
        n17294) );
  AOI22_X1 U20490 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20491 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20492 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17290) );
  NAND3_X1 U20493 ( .A1(n17292), .A2(n17291), .A3(n17290), .ZN(n17293) );
  AOI211_X1 U20494 ( .C1(n17418), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17294), .B(n17293), .ZN(n17295) );
  OAI211_X1 U20495 ( .C1(n17450), .C2(n17297), .A(n17296), .B(n17295), .ZN(
        n17298) );
  AOI211_X1 U20496 ( .C1(n17436), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n17299), .B(n17298), .ZN(n17570) );
  AND2_X1 U20497 ( .A1(n17511), .A2(n17300), .ZN(n17316) );
  AOI22_X1 U20498 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17316), .B1(n17302), 
        .B2(n17301), .ZN(n17303) );
  OAI21_X1 U20499 ( .B1(n17570), .B2(n17511), .A(n17303), .ZN(P3_U2682) );
  AOI22_X1 U20500 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20501 ( .B1(n15718), .B2(n17305), .A(n17304), .ZN(n17315) );
  AOI22_X1 U20502 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17312) );
  OAI22_X1 U20503 ( .A1(n17381), .A2(n21348), .B1(n9875), .B2(n18814), .ZN(
        n17310) );
  AOI22_X1 U20504 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20505 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20506 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17306) );
  NAND3_X1 U20507 ( .A1(n17308), .A2(n17307), .A3(n17306), .ZN(n17309) );
  AOI211_X1 U20508 ( .C1(n17365), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17310), .B(n17309), .ZN(n17311) );
  OAI211_X1 U20509 ( .C1(n13975), .C2(n17313), .A(n17312), .B(n17311), .ZN(
        n17314) );
  AOI211_X1 U20510 ( .C1(n17436), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17315), .B(n17314), .ZN(n17577) );
  OAI221_X1 U20511 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17317), .A(n17316), .ZN(n17318) );
  OAI21_X1 U20512 ( .B1(n17577), .B2(n17511), .A(n17318), .ZN(P3_U2683) );
  NOR2_X1 U20513 ( .A1(n17517), .A2(n17319), .ZN(n17346) );
  AOI22_X1 U20514 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15874), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20515 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20516 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17320) );
  OAI211_X1 U20517 ( .C1(n13976), .C2(n17322), .A(n17321), .B(n17320), .ZN(
        n17328) );
  AOI22_X1 U20518 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20519 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20520 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17324) );
  NAND2_X1 U20521 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n17323) );
  NAND4_X1 U20522 ( .A1(n17326), .A2(n17325), .A3(n17324), .A4(n17323), .ZN(
        n17327) );
  AOI211_X1 U20523 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17328), .B(n17327), .ZN(n17329) );
  OAI211_X1 U20524 ( .C1(n13975), .C2(n18710), .A(n17330), .B(n17329), .ZN(
        n17578) );
  AOI22_X1 U20525 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17346), .B1(n17517), 
        .B2(n17578), .ZN(n17331) );
  OAI21_X1 U20526 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17332), .A(n17331), .ZN(
        P3_U2684) );
  AOI22_X1 U20527 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17333) );
  OAI21_X1 U20528 ( .B1(n17467), .B2(n17334), .A(n17333), .ZN(n17343) );
  AOI22_X1 U20529 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17341) );
  AOI22_X1 U20530 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17335) );
  OAI21_X1 U20531 ( .B1(n17473), .B2(n21364), .A(n17335), .ZN(n17339) );
  AOI22_X1 U20532 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20533 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17336) );
  OAI211_X1 U20534 ( .C1(n13976), .C2(n21244), .A(n17337), .B(n17336), .ZN(
        n17338) );
  AOI211_X1 U20535 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17339), .B(n17338), .ZN(n17340) );
  OAI211_X1 U20536 ( .C1(n17381), .C2(n17509), .A(n17341), .B(n17340), .ZN(
        n17342) );
  AOI211_X1 U20537 ( .C1(n17365), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17343), .B(n17342), .ZN(n17587) );
  NAND2_X1 U20538 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17363), .ZN(n17362) );
  OAI21_X1 U20539 ( .B1(n17345), .B2(n17362), .A(n17344), .ZN(n17347) );
  NAND2_X1 U20540 ( .A1(n17347), .A2(n17346), .ZN(n17348) );
  OAI21_X1 U20541 ( .B1(n17587), .B2(n17511), .A(n17348), .ZN(P3_U2685) );
  AOI22_X1 U20542 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17349), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20543 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17417), .ZN(n17358) );
  AOI22_X1 U20544 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15843), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17418), .ZN(n17357) );
  OAI22_X1 U20545 ( .A1(n21224), .A2(n17473), .B1(n21197), .B2(n9875), .ZN(
        n17355) );
  AOI22_X1 U20546 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17365), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n15877), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20548 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13988), .ZN(n17351) );
  NAND2_X1 U20549 ( .A1(n17468), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n17350) );
  NAND4_X1 U20550 ( .A1(n17353), .A2(n17352), .A3(n17351), .A4(n17350), .ZN(
        n17354) );
  AOI211_X1 U20551 ( .C1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .C2(n15875), .A(
        n17355), .B(n17354), .ZN(n17356) );
  NAND4_X1 U20552 ( .A1(n17359), .A2(n17358), .A3(n17357), .A4(n17356), .ZN(
        n17588) );
  OAI222_X1 U20553 ( .A1(n17517), .A2(P3_EBX_REG_17__SCAN_IN), .B1(n17517), 
        .B2(n17360), .C1(n17511), .C2(n17588), .ZN(n17361) );
  OAI21_X1 U20554 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17362), .A(n17361), .ZN(
        P3_U2686) );
  INV_X1 U20555 ( .A(n17362), .ZN(n17377) );
  AOI21_X1 U20556 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17511), .A(n17363), .ZN(
        n17376) );
  AOI22_X1 U20557 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20558 ( .B1(n15718), .B2(n17482), .A(n17364), .ZN(n17375) );
  AOI22_X1 U20559 ( .A1(n17365), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U20560 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15843), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17366) );
  INV_X1 U20561 ( .A(n17366), .ZN(n17371) );
  AOI22_X1 U20562 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20563 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20564 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17367) );
  NAND3_X1 U20565 ( .A1(n17369), .A2(n17368), .A3(n17367), .ZN(n17370) );
  AOI211_X1 U20566 ( .C1(n15875), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17371), .B(n17370), .ZN(n17372) );
  OAI211_X1 U20567 ( .C1(n17381), .C2(n17477), .A(n17373), .B(n17372), .ZN(
        n17374) );
  AOI211_X1 U20568 ( .C1(n17436), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17375), .B(n17374), .ZN(n17600) );
  OAI22_X1 U20569 ( .A1(n17377), .A2(n17376), .B1(n17600), .B2(n17511), .ZN(
        P3_U2687) );
  NAND2_X1 U20570 ( .A1(n18511), .A2(n17520), .ZN(n17515) );
  INV_X1 U20571 ( .A(n17515), .ZN(n17516) );
  AOI21_X1 U20572 ( .B1(n17516), .B2(n17393), .A(n17378), .ZN(n17397) );
  AOI22_X1 U20573 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20574 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20575 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17389) );
  OAI22_X1 U20576 ( .A1(n9947), .A2(n18821), .B1(n17381), .B2(n17380), .ZN(
        n17387) );
  AOI22_X1 U20577 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20578 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20579 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15875), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17383) );
  NAND2_X1 U20580 ( .A1(n15843), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n17382) );
  NAND4_X1 U20581 ( .A1(n17385), .A2(n17384), .A3(n17383), .A4(n17382), .ZN(
        n17386) );
  AOI211_X1 U20582 ( .C1(n17349), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17387), .B(n17386), .ZN(n17388) );
  NAND4_X1 U20583 ( .A1(n17391), .A2(n17390), .A3(n17389), .A4(n17388), .ZN(
        n17605) );
  NOR3_X1 U20584 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17393), .A3(n17392), .ZN(
        n17394) );
  AOI21_X1 U20585 ( .B1(n17517), .B2(n17605), .A(n17394), .ZN(n17395) );
  OAI21_X1 U20586 ( .B1(n17397), .B2(n17396), .A(n17395), .ZN(P3_U2689) );
  INV_X1 U20587 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20588 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20589 ( .B1(n9878), .B2(n17399), .A(n17398), .ZN(n17410) );
  AOI22_X1 U20590 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20591 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20592 ( .B1(n13976), .B2(n21348), .A(n17400), .ZN(n17405) );
  AOI22_X1 U20593 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20594 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17401) );
  OAI211_X1 U20595 ( .C1(n17473), .C2(n17403), .A(n17402), .B(n17401), .ZN(
        n17404) );
  AOI211_X1 U20596 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17405), .B(n17404), .ZN(n17406) );
  OAI211_X1 U20597 ( .C1(n17449), .C2(n17408), .A(n17407), .B(n17406), .ZN(
        n17409) );
  AOI211_X1 U20598 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17410), .B(n17409), .ZN(n17615) );
  AOI21_X1 U20599 ( .B1(n21223), .B2(n17428), .A(n17411), .ZN(n17412) );
  INV_X1 U20600 ( .A(n17412), .ZN(n17413) );
  AOI22_X1 U20601 ( .A1(n17517), .A2(n17615), .B1(n17413), .B2(n17511), .ZN(
        P3_U2691) );
  AOI22_X1 U20602 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20603 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20604 ( .B1(n17449), .B2(n17415), .A(n17414), .ZN(n17424) );
  OAI22_X1 U20605 ( .A1(n9947), .A2(n21166), .B1(n17467), .B2(n18710), .ZN(
        n17416) );
  AOI21_X1 U20606 ( .B1(n17468), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n17416), .ZN(n17422) );
  AOI22_X1 U20607 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20608 ( .A1(n13988), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20609 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17418), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17419) );
  NAND4_X1 U20610 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17423) );
  AOI211_X1 U20611 ( .C1(n17379), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17424), .B(n17423), .ZN(n17425) );
  OAI211_X1 U20612 ( .C1(n17427), .C2(n21247), .A(n17426), .B(n17425), .ZN(
        n17618) );
  INV_X1 U20613 ( .A(n17618), .ZN(n17430) );
  OAI21_X1 U20614 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17431), .A(n17428), .ZN(
        n17429) );
  AOI22_X1 U20615 ( .A1(n17517), .A2(n17430), .B1(n17429), .B2(n17511), .ZN(
        P3_U2692) );
  INV_X1 U20616 ( .A(n17431), .ZN(n17446) );
  AOI21_X1 U20617 ( .B1(n17432), .B2(n17464), .A(n17517), .ZN(n17445) );
  AOI22_X1 U20618 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20619 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20620 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17434) );
  OAI211_X1 U20621 ( .C1(n13976), .C2(n17509), .A(n17435), .B(n17434), .ZN(
        n17442) );
  AOI22_X1 U20622 ( .A1(n17469), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20623 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20624 ( .A1(n17436), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17438) );
  NAND2_X1 U20625 ( .A1(n15874), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n17437) );
  NAND4_X1 U20626 ( .A1(n17440), .A2(n17439), .A3(n17438), .A4(n17437), .ZN(
        n17441) );
  AOI211_X1 U20627 ( .C1(n15843), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17442), .B(n17441), .ZN(n17443) );
  OAI211_X1 U20628 ( .C1(n15718), .C2(n21244), .A(n17444), .B(n17443), .ZN(
        n17621) );
  AOI22_X1 U20629 ( .A1(n17446), .A2(n17445), .B1(n17621), .B2(n17517), .ZN(
        n17447) );
  INV_X1 U20630 ( .A(n17447), .ZN(P3_U2693) );
  OAI22_X1 U20631 ( .A1(n17449), .A2(n17448), .B1(n17467), .B2(n18705), .ZN(
        n17463) );
  OAI22_X1 U20632 ( .A1(n17451), .A2(n13975), .B1(n21224), .B2(n17450), .ZN(
        n17462) );
  INV_X1 U20633 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20634 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15875), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20635 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n15843), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17468), .ZN(n17452) );
  OAI21_X1 U20636 ( .B1(n9947), .B2(n21197), .A(n17452), .ZN(n17457) );
  INV_X1 U20637 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20638 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13988), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20639 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17453), .B1(
        n9763), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17454) );
  OAI211_X1 U20640 ( .C1(n13976), .C2(n17512), .A(n17455), .B(n17454), .ZN(
        n17456) );
  AOI211_X1 U20641 ( .C1(n15874), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17457), .B(n17456), .ZN(n17458) );
  OAI211_X1 U20642 ( .C1(n15718), .C2(n17460), .A(n17459), .B(n17458), .ZN(
        n17461) );
  NOR3_X1 U20643 ( .A1(n17463), .A2(n17462), .A3(n17461), .ZN(n17626) );
  OAI21_X1 U20644 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17486), .A(n17464), .ZN(
        n17465) );
  AOI22_X1 U20645 ( .A1(n17517), .A2(n17626), .B1(n17465), .B2(n17511), .ZN(
        P3_U2694) );
  OAI21_X1 U20646 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17487), .A(n17511), .ZN(
        n17485) );
  AOI22_X1 U20647 ( .A1(n15875), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15877), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U20648 ( .A1(n9763), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17453), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20649 ( .B1(n17467), .B2(n18702), .A(n17466), .ZN(n17479) );
  AOI22_X1 U20650 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17468), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20651 ( .A1(n17379), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17469), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20652 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13988), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17471) );
  OAI211_X1 U20653 ( .C1(n17473), .C2(n18561), .A(n17472), .B(n17471), .ZN(
        n17474) );
  AOI21_X1 U20654 ( .B1(n15843), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17474), .ZN(n17475) );
  OAI211_X1 U20655 ( .C1(n13976), .C2(n17477), .A(n17476), .B(n17475), .ZN(
        n17478) );
  AOI211_X1 U20656 ( .C1(n17436), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n17479), .B(n17478), .ZN(n17480) );
  OAI211_X1 U20657 ( .C1(n17483), .C2(n17482), .A(n17481), .B(n17480), .ZN(
        n17629) );
  INV_X1 U20658 ( .A(n17629), .ZN(n17484) );
  OAI22_X1 U20659 ( .A1(n17486), .A2(n17485), .B1(n17484), .B2(n17511), .ZN(
        P3_U2695) );
  NOR2_X1 U20660 ( .A1(n17625), .A2(n9909), .ZN(n17491) );
  INV_X1 U20661 ( .A(n17487), .ZN(n17488) );
  OAI221_X1 U20662 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(P3_EBX_REG_6__SCAN_IN), 
        .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17491), .A(n17488), .ZN(n17489) );
  AOI22_X1 U20663 ( .A1(n17517), .A2(n17490), .B1(n17489), .B2(n17511), .ZN(
        P3_U2696) );
  NAND2_X1 U20664 ( .A1(n17511), .A2(n9909), .ZN(n17496) );
  AOI22_X1 U20665 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17517), .B1(
        n17491), .B2(n17493), .ZN(n17492) );
  OAI21_X1 U20666 ( .B1(n17493), .B2(n17496), .A(n17492), .ZN(P3_U2697) );
  AND2_X1 U20667 ( .A1(n17494), .A2(n17498), .ZN(n17497) );
  OAI22_X1 U20668 ( .A1(n17497), .A2(n17496), .B1(n17495), .B2(n17511), .ZN(
        P3_U2698) );
  OAI21_X1 U20669 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17499), .A(n17498), .ZN(
        n17500) );
  AOI22_X1 U20670 ( .A1(n17517), .A2(n21348), .B1(n17500), .B2(n17511), .ZN(
        P3_U2699) );
  INV_X1 U20671 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17505) );
  INV_X1 U20672 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n21304) );
  NOR3_X1 U20673 ( .A1(n21304), .A2(n17506), .A3(n17515), .ZN(n17508) );
  NOR2_X1 U20674 ( .A1(n17517), .A2(n17501), .ZN(n17503) );
  OAI22_X1 U20675 ( .A1(n17508), .A2(n17503), .B1(n17502), .B2(n17515), .ZN(
        n17504) );
  OAI21_X1 U20676 ( .B1(n17511), .B2(n17505), .A(n17504), .ZN(P3_U2700) );
  INV_X1 U20677 ( .A(n17506), .ZN(n17507) );
  AOI21_X1 U20678 ( .B1(n17520), .B2(n17507), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17510) );
  AOI221_X1 U20679 ( .B1(n17510), .B2(n17511), .C1(n17509), .C2(n17517), .A(
        n17508), .ZN(P3_U2701) );
  OAI222_X1 U20680 ( .A1(n17515), .A2(n17514), .B1(n17513), .B2(n17520), .C1(
        n17512), .C2(n17511), .ZN(P3_U2702) );
  AOI22_X1 U20681 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17517), .B1(
        n17516), .B2(n17519), .ZN(n17518) );
  OAI21_X1 U20682 ( .B1(n17520), .B2(n17519), .A(n17518), .ZN(P3_U2703) );
  INV_X1 U20683 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17673) );
  INV_X1 U20684 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17676) );
  INV_X1 U20685 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17681) );
  INV_X1 U20686 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17692) );
  NAND4_X1 U20687 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17522)
         );
  NAND2_X1 U20688 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n17633) );
  NAND2_X1 U20689 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17634) );
  INV_X1 U20690 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21456) );
  INV_X1 U20691 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17684) );
  INV_X1 U20692 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17687) );
  INV_X1 U20693 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17689) );
  NOR4_X1 U20694 ( .A1(n21456), .A2(n17684), .A3(n17687), .A4(n17689), .ZN(
        n17569) );
  NAND3_X1 U20695 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17596), .A3(n17569), 
        .ZN(n17564) );
  NAND2_X1 U20696 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17560), .ZN(n17559) );
  NAND2_X1 U20697 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17541), .ZN(n17537) );
  NAND2_X1 U20698 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17533), .ZN(n17532) );
  INV_X1 U20699 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17741) );
  OR2_X1 U20700 ( .A1(n17532), .A2(n17741), .ZN(n17526) );
  NAND2_X1 U20701 ( .A1(n17523), .A2(n17607), .ZN(n17593) );
  NAND2_X1 U20702 ( .A1(n17651), .A2(n17532), .ZN(n17531) );
  OAI21_X1 U20703 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17632), .A(n17531), .ZN(
        n17524) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17594), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17524), .ZN(n17525) );
  OAI21_X1 U20705 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17526), .A(n17525), .ZN(
        P3_U2704) );
  NOR2_X2 U20706 ( .A1(n17527), .A2(n17651), .ZN(n17595) );
  INV_X1 U20707 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18502) );
  OAI22_X1 U20708 ( .A1(n17528), .A2(n17661), .B1(n18502), .B2(n17593), .ZN(
        n17529) );
  AOI21_X1 U20709 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17595), .A(n17529), .ZN(
        n17530) );
  OAI221_X1 U20710 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17532), .C1(n17741), 
        .C2(n17531), .A(n17530), .ZN(P3_U2705) );
  AOI22_X1 U20711 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17594), .ZN(n17535) );
  OAI211_X1 U20712 ( .C1(n17533), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17651), .B(
        n17532), .ZN(n17534) );
  OAI211_X1 U20713 ( .C1(n17536), .C2(n17661), .A(n17535), .B(n17534), .ZN(
        P3_U2706) );
  AOI22_X1 U20714 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17594), .ZN(n17539) );
  OAI211_X1 U20715 ( .C1(n17541), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17651), .B(
        n17537), .ZN(n17538) );
  OAI211_X1 U20716 ( .C1(n17540), .C2(n17661), .A(n17539), .B(n17538), .ZN(
        P3_U2707) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17594), .ZN(n17544) );
  AOI211_X1 U20718 ( .C1(n17673), .C2(n17546), .A(n17541), .B(n17607), .ZN(
        n17542) );
  INV_X1 U20719 ( .A(n17542), .ZN(n17543) );
  OAI211_X1 U20720 ( .C1(n17545), .C2(n17661), .A(n17544), .B(n17543), .ZN(
        P3_U2708) );
  AOI22_X1 U20721 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17594), .ZN(n17548) );
  OAI211_X1 U20722 ( .C1(n9911), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17651), .B(
        n17546), .ZN(n17547) );
  OAI211_X1 U20723 ( .C1(n17549), .C2(n17661), .A(n17548), .B(n17547), .ZN(
        P3_U2709) );
  AOI22_X1 U20724 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17594), .ZN(n17552) );
  AOI211_X1 U20725 ( .C1(n17676), .C2(n17554), .A(n9911), .B(n17607), .ZN(
        n17550) );
  INV_X1 U20726 ( .A(n17550), .ZN(n17551) );
  OAI211_X1 U20727 ( .C1(n17553), .C2(n17661), .A(n17552), .B(n17551), .ZN(
        P3_U2710) );
  AOI22_X1 U20728 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17594), .ZN(n17557) );
  OAI211_X1 U20729 ( .C1(n17555), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17651), .B(
        n17554), .ZN(n17556) );
  OAI211_X1 U20730 ( .C1(n17558), .C2(n17661), .A(n17557), .B(n17556), .ZN(
        P3_U2711) );
  AOI22_X1 U20731 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17594), .ZN(n17562) );
  OAI211_X1 U20732 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17560), .A(n17651), .B(
        n17559), .ZN(n17561) );
  OAI211_X1 U20733 ( .C1(n17563), .C2(n17661), .A(n17562), .B(n17561), .ZN(
        P3_U2712) );
  OR2_X1 U20734 ( .A1(n17625), .A2(n17564), .ZN(n17568) );
  NAND2_X1 U20735 ( .A1(n17651), .A2(n17564), .ZN(n17573) );
  INV_X1 U20736 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19483) );
  OAI22_X1 U20737 ( .A1(n17565), .A2(n17661), .B1(n19483), .B2(n17593), .ZN(
        n17566) );
  AOI21_X1 U20738 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17595), .A(n17566), .ZN(
        n17567) );
  OAI221_X1 U20739 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17568), .C1(n17681), 
        .C2(n17573), .A(n17567), .ZN(P3_U2713) );
  AND2_X1 U20740 ( .A1(n18511), .A2(n17596), .ZN(n17590) );
  NAND2_X1 U20741 ( .A1(n17569), .A2(n17590), .ZN(n17574) );
  INV_X1 U20742 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17731) );
  OAI22_X1 U20743 ( .A1(n17570), .A2(n17661), .B1(n21230), .B2(n17593), .ZN(
        n17571) );
  AOI21_X1 U20744 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17595), .A(n17571), .ZN(
        n17572) );
  OAI221_X1 U20745 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17574), .C1(n17731), 
        .C2(n17573), .A(n17572), .ZN(P3_U2714) );
  AOI22_X1 U20746 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17594), .ZN(n17576) );
  NAND3_X1 U20747 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n17590), .ZN(n17583) );
  NOR2_X1 U20748 ( .A1(n21456), .A2(n17583), .ZN(n17579) );
  OAI211_X1 U20749 ( .C1(n17579), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17651), .B(
        n17574), .ZN(n17575) );
  OAI211_X1 U20750 ( .C1(n17577), .C2(n17661), .A(n17576), .B(n17575), .ZN(
        P3_U2715) );
  INV_X1 U20751 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n21181) );
  AOI22_X1 U20752 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17595), .B1(n17653), .B2(
        n17578), .ZN(n17582) );
  AOI211_X1 U20753 ( .C1(n21456), .C2(n17583), .A(n17579), .B(n17607), .ZN(
        n17580) );
  INV_X1 U20754 ( .A(n17580), .ZN(n17581) );
  OAI211_X1 U20755 ( .C1(n17593), .C2(n21181), .A(n17582), .B(n17581), .ZN(
        P3_U2716) );
  AOI22_X1 U20756 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17594), .ZN(n17586) );
  NAND2_X1 U20757 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17590), .ZN(n17589) );
  INV_X1 U20758 ( .A(n17589), .ZN(n17584) );
  OAI211_X1 U20759 ( .C1(n17584), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17651), .B(
        n17583), .ZN(n17585) );
  OAI211_X1 U20760 ( .C1(n17587), .C2(n17661), .A(n17586), .B(n17585), .ZN(
        P3_U2717) );
  INV_X1 U20761 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18482) );
  AOI22_X1 U20762 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17595), .B1(n17653), .B2(
        n17588), .ZN(n17592) );
  OAI211_X1 U20763 ( .C1(n17590), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17651), .B(
        n17589), .ZN(n17591) );
  OAI211_X1 U20764 ( .C1(n17593), .C2(n18482), .A(n17592), .B(n17591), .ZN(
        P3_U2718) );
  AOI22_X1 U20765 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17595), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17594), .ZN(n17599) );
  AOI211_X1 U20766 ( .C1(n17692), .C2(n17601), .A(n17607), .B(n17596), .ZN(
        n17597) );
  INV_X1 U20767 ( .A(n17597), .ZN(n17598) );
  OAI211_X1 U20768 ( .C1(n17600), .C2(n17661), .A(n17599), .B(n17598), .ZN(
        P3_U2719) );
  OAI211_X1 U20769 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17606), .A(n17651), .B(
        n17601), .ZN(n17603) );
  NAND2_X1 U20770 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17654), .ZN(n17602) );
  OAI211_X1 U20771 ( .C1(n17604), .C2(n17661), .A(n17603), .B(n17602), .ZN(
        P3_U2720) );
  INV_X1 U20772 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17700) );
  INV_X1 U20773 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17704) );
  INV_X1 U20774 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17706) );
  NAND2_X1 U20775 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17628), .ZN(n17620) );
  NOR2_X1 U20776 ( .A1(n17700), .A2(n17620), .ZN(n17614) );
  NAND2_X1 U20777 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17617), .ZN(n17610) );
  AOI22_X1 U20778 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17654), .B1(n17653), .B2(
        n17605), .ZN(n17609) );
  INV_X1 U20779 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17766) );
  OR3_X1 U20780 ( .A1(n17766), .A2(n17607), .A3(n17606), .ZN(n17608) );
  OAI211_X1 U20781 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17610), .A(n17609), .B(
        n17608), .ZN(P3_U2721) );
  INV_X1 U20782 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17764) );
  INV_X1 U20783 ( .A(n17610), .ZN(n17613) );
  AOI21_X1 U20784 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17651), .A(n17617), .ZN(
        n17612) );
  OAI222_X1 U20785 ( .A1(n17662), .A2(n17764), .B1(n17613), .B2(n17612), .C1(
        n17661), .C2(n17611), .ZN(P3_U2722) );
  INV_X1 U20786 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21209) );
  AOI21_X1 U20787 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17651), .A(n17614), .ZN(
        n17616) );
  OAI222_X1 U20788 ( .A1(n17662), .A2(n21209), .B1(n17617), .B2(n17616), .C1(
        n17661), .C2(n17615), .ZN(P3_U2723) );
  NAND2_X1 U20789 ( .A1(n17651), .A2(n17620), .ZN(n17624) );
  AOI22_X1 U20790 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17654), .B1(n17653), .B2(
        n17618), .ZN(n17619) );
  OAI221_X1 U20791 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17620), .C1(n17700), 
        .C2(n17624), .A(n17619), .ZN(P3_U2724) );
  INV_X1 U20792 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17702) );
  INV_X1 U20793 ( .A(n17628), .ZN(n17623) );
  AOI22_X1 U20794 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17654), .B1(n17653), .B2(
        n17621), .ZN(n17622) );
  OAI221_X1 U20795 ( .B1(n17624), .B2(n17702), .C1(n17624), .C2(n17623), .A(
        n17622), .ZN(P3_U2725) );
  NOR2_X1 U20796 ( .A1(n17625), .A2(n9854), .ZN(n17636) );
  AOI22_X1 U20797 ( .A1(n17636), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17651), .ZN(n17627) );
  OAI222_X1 U20798 ( .A1(n17662), .A2(n17756), .B1(n17628), .B2(n17627), .C1(
        n17661), .C2(n17626), .ZN(P3_U2726) );
  INV_X1 U20799 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U20800 ( .A1(n17653), .A2(n17629), .B1(n17636), .B2(n17706), .ZN(
        n17631) );
  NAND3_X1 U20801 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17651), .A3(n9854), .ZN(
        n17630) );
  OAI211_X1 U20802 ( .C1(n17662), .C2(n17754), .A(n17631), .B(n17630), .ZN(
        P3_U2727) );
  INV_X1 U20803 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18508) );
  INV_X1 U20804 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21131) );
  NOR2_X1 U20805 ( .A1(n21131), .A2(n17656), .ZN(n17647) );
  NAND2_X1 U20806 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17650), .ZN(n17643) );
  NOR2_X1 U20807 ( .A1(n17634), .A2(n17643), .ZN(n17639) );
  AOI21_X1 U20808 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17651), .A(n17639), .ZN(
        n17635) );
  OAI222_X1 U20809 ( .A1(n17662), .A2(n18508), .B1(n17636), .B2(n17635), .C1(
        n17661), .C2(n18047), .ZN(P3_U2728) );
  INV_X1 U20810 ( .A(n17643), .ZN(n17646) );
  AOI22_X1 U20811 ( .A1(n17646), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17651), .ZN(n17638) );
  OAI222_X1 U20812 ( .A1(n18503), .A2(n17662), .B1(n17639), .B2(n17638), .C1(
        n17661), .C2(n17637), .ZN(P3_U2729) );
  NAND3_X1 U20813 ( .A1(n17651), .A2(P3_EAX_REG_5__SCAN_IN), .A3(n17643), .ZN(
        n17642) );
  AOI22_X1 U20814 ( .A1(n17654), .A2(BUF2_REG_5__SCAN_IN), .B1(n17653), .B2(
        n17640), .ZN(n17641) );
  OAI211_X1 U20815 ( .C1(P3_EAX_REG_5__SCAN_IN), .C2(n17643), .A(n17642), .B(
        n17641), .ZN(P3_U2730) );
  AOI21_X1 U20816 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17651), .A(n17650), .ZN(
        n17645) );
  OAI222_X1 U20817 ( .A1(n18494), .A2(n17662), .B1(n17646), .B2(n17645), .C1(
        n17661), .C2(n17644), .ZN(P3_U2731) );
  AOI21_X1 U20818 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17651), .A(n17647), .ZN(
        n17649) );
  OAI222_X1 U20819 ( .A1(n21458), .A2(n17662), .B1(n17650), .B2(n17649), .C1(
        n17661), .C2(n17648), .ZN(P3_U2732) );
  NAND2_X1 U20820 ( .A1(n17651), .A2(n17656), .ZN(n17659) );
  AOI22_X1 U20821 ( .A1(n17654), .A2(BUF2_REG_2__SCAN_IN), .B1(n17653), .B2(
        n17652), .ZN(n17655) );
  OAI221_X1 U20822 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17656), .C1(n21131), 
        .C2(n17659), .A(n17655), .ZN(P3_U2733) );
  INV_X1 U20823 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18483) );
  AOI21_X1 U20824 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17657), .A(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17658) );
  OAI222_X1 U20825 ( .A1(n17662), .A2(n18483), .B1(n17661), .B2(n17660), .C1(
        n17659), .C2(n17658), .ZN(P3_U2734) );
  NOR2_X2 U20826 ( .A1(n19100), .A2(n18135), .ZN(n19152) );
  NOR2_X4 U20827 ( .A1(n19152), .A2(n17693), .ZN(n17709) );
  AND2_X1 U20828 ( .A1(n17709), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20829 ( .A1(n19152), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17667) );
  OAI21_X1 U20830 ( .B1(n17741), .B2(n17691), .A(n17667), .ZN(P3_U2737) );
  INV_X1 U20831 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17669) );
  AOI22_X1 U20832 ( .A1(n19152), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17668) );
  OAI21_X1 U20833 ( .B1(n17669), .B2(n17691), .A(n17668), .ZN(P3_U2738) );
  INV_X1 U20834 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17671) );
  AOI22_X1 U20835 ( .A1(n19152), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17670) );
  OAI21_X1 U20836 ( .B1(n17671), .B2(n17691), .A(n17670), .ZN(P3_U2739) );
  AOI22_X1 U20837 ( .A1(n19152), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17672) );
  OAI21_X1 U20838 ( .B1(n17673), .B2(n17691), .A(n17672), .ZN(P3_U2740) );
  AOI22_X1 U20839 ( .A1(n19152), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17674) );
  OAI21_X1 U20840 ( .B1(n10169), .B2(n17691), .A(n17674), .ZN(P3_U2741) );
  AOI22_X1 U20841 ( .A1(n19152), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17675) );
  OAI21_X1 U20842 ( .B1(n17676), .B2(n17691), .A(n17675), .ZN(P3_U2742) );
  AOI22_X1 U20843 ( .A1(n19152), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U20844 ( .B1(n10168), .B2(n17691), .A(n17677), .ZN(P3_U2743) );
  INV_X1 U20845 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17679) );
  CLKBUF_X1 U20846 ( .A(n19152), .Z(n17720) );
  AOI22_X1 U20847 ( .A1(n17720), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17678) );
  OAI21_X1 U20848 ( .B1(n17679), .B2(n17691), .A(n17678), .ZN(P3_U2744) );
  AOI22_X1 U20849 ( .A1(n17720), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17680) );
  OAI21_X1 U20850 ( .B1(n17681), .B2(n17691), .A(n17680), .ZN(P3_U2745) );
  AOI22_X1 U20851 ( .A1(n17720), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17682) );
  OAI21_X1 U20852 ( .B1(n17731), .B2(n17691), .A(n17682), .ZN(P3_U2746) );
  AOI22_X1 U20853 ( .A1(n17720), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17683) );
  OAI21_X1 U20854 ( .B1(n17684), .B2(n17691), .A(n17683), .ZN(P3_U2747) );
  AOI22_X1 U20855 ( .A1(n17720), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U20856 ( .B1(n21456), .B2(n17691), .A(n17685), .ZN(P3_U2748) );
  AOI22_X1 U20857 ( .A1(n17720), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17686) );
  OAI21_X1 U20858 ( .B1(n17687), .B2(n17691), .A(n17686), .ZN(P3_U2749) );
  AOI22_X1 U20859 ( .A1(n17720), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17688) );
  OAI21_X1 U20860 ( .B1(n17689), .B2(n17691), .A(n17688), .ZN(P3_U2750) );
  AOI22_X1 U20861 ( .A1(n17720), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17690) );
  OAI21_X1 U20862 ( .B1(n17692), .B2(n17691), .A(n17690), .ZN(P3_U2751) );
  INV_X1 U20863 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U20864 ( .A1(n17720), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U20865 ( .B1(n17769), .B2(n17722), .A(n17694), .ZN(P3_U2752) );
  AOI22_X1 U20866 ( .A1(n17720), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20867 ( .B1(n17766), .B2(n17722), .A(n17695), .ZN(P3_U2753) );
  INV_X1 U20868 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17697) );
  AOI22_X1 U20869 ( .A1(n17720), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17696) );
  OAI21_X1 U20870 ( .B1(n17697), .B2(n17722), .A(n17696), .ZN(P3_U2754) );
  INV_X1 U20871 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21215) );
  AOI22_X1 U20872 ( .A1(n17720), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17698) );
  OAI21_X1 U20873 ( .B1(n21215), .B2(n17722), .A(n17698), .ZN(P3_U2755) );
  AOI22_X1 U20874 ( .A1(n17720), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17699) );
  OAI21_X1 U20875 ( .B1(n17700), .B2(n17722), .A(n17699), .ZN(P3_U2756) );
  AOI22_X1 U20876 ( .A1(n17720), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17701) );
  OAI21_X1 U20877 ( .B1(n17702), .B2(n17722), .A(n17701), .ZN(P3_U2757) );
  AOI22_X1 U20878 ( .A1(n17720), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17703) );
  OAI21_X1 U20879 ( .B1(n17704), .B2(n17722), .A(n17703), .ZN(P3_U2758) );
  AOI22_X1 U20880 ( .A1(n17720), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17705) );
  OAI21_X1 U20881 ( .B1(n17706), .B2(n17722), .A(n17705), .ZN(P3_U2759) );
  INV_X1 U20882 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U20883 ( .A1(n17720), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U20884 ( .B1(n17708), .B2(n17722), .A(n17707), .ZN(P3_U2760) );
  INV_X1 U20885 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U20886 ( .A1(n17720), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17710) );
  OAI21_X1 U20887 ( .B1(n17711), .B2(n17722), .A(n17710), .ZN(P3_U2761) );
  INV_X1 U20888 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20889 ( .A1(n17720), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17712) );
  OAI21_X1 U20890 ( .B1(n17749), .B2(n17722), .A(n17712), .ZN(P3_U2762) );
  INV_X1 U20891 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17714) );
  AOI22_X1 U20892 ( .A1(n17720), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17713) );
  OAI21_X1 U20893 ( .B1(n17714), .B2(n17722), .A(n17713), .ZN(P3_U2763) );
  INV_X1 U20894 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U20895 ( .A1(n17720), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U20896 ( .B1(n17716), .B2(n17722), .A(n17715), .ZN(P3_U2764) );
  AOI22_X1 U20897 ( .A1(n17720), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U20898 ( .B1(n21131), .B2(n17722), .A(n17717), .ZN(P3_U2765) );
  INV_X1 U20899 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17719) );
  AOI22_X1 U20900 ( .A1(n17720), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17718) );
  OAI21_X1 U20901 ( .B1(n17719), .B2(n17722), .A(n17718), .ZN(P3_U2766) );
  AOI22_X1 U20902 ( .A1(n17720), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17709), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17721) );
  OAI21_X1 U20903 ( .B1(n21289), .B2(n17722), .A(n17721), .ZN(P3_U2767) );
  INV_X1 U20904 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18475) );
  AOI22_X1 U20905 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17762), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17752), .ZN(n17726) );
  OAI21_X1 U20906 ( .B1(n18475), .B2(n21457), .A(n17726), .ZN(P3_U2768) );
  AOI22_X1 U20907 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17762), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17752), .ZN(n17727) );
  OAI21_X1 U20908 ( .B1(n18483), .B2(n21457), .A(n17727), .ZN(P3_U2769) );
  INV_X1 U20909 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U20910 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17752), .ZN(n17728) );
  OAI21_X1 U20911 ( .B1(n18487), .B2(n21457), .A(n17728), .ZN(P3_U2770) );
  AOI22_X1 U20912 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17752), .ZN(n17729) );
  OAI21_X1 U20913 ( .B1(n18494), .B2(n21457), .A(n17729), .ZN(P3_U2772) );
  AOI22_X1 U20914 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17767), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17752), .ZN(n17730) );
  OAI21_X1 U20915 ( .B1(n17731), .B2(n21455), .A(n17730), .ZN(P3_U2773) );
  AOI22_X1 U20916 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17752), .ZN(n17732) );
  OAI21_X1 U20917 ( .B1(n18503), .B2(n21457), .A(n17732), .ZN(P3_U2774) );
  AOI22_X1 U20918 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17752), .ZN(n17733) );
  OAI21_X1 U20919 ( .B1(n18508), .B2(n21457), .A(n17733), .ZN(P3_U2775) );
  AOI22_X1 U20920 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17752), .ZN(n17734) );
  OAI21_X1 U20921 ( .B1(n17754), .B2(n17744), .A(n17734), .ZN(P3_U2776) );
  AOI22_X1 U20922 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17752), .ZN(n17735) );
  OAI21_X1 U20923 ( .B1(n17756), .B2(n17744), .A(n17735), .ZN(P3_U2777) );
  INV_X1 U20924 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17758) );
  AOI22_X1 U20925 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17752), .ZN(n17736) );
  OAI21_X1 U20926 ( .B1(n17758), .B2(n17744), .A(n17736), .ZN(P3_U2778) );
  INV_X1 U20927 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21201) );
  AOI22_X1 U20928 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17752), .ZN(n17737) );
  OAI21_X1 U20929 ( .B1(n21201), .B2(n17744), .A(n17737), .ZN(P3_U2779) );
  AOI22_X1 U20930 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17752), .ZN(n17738) );
  OAI21_X1 U20931 ( .B1(n21209), .B2(n17744), .A(n17738), .ZN(P3_U2780) );
  AOI22_X1 U20932 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17760), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17752), .ZN(n17739) );
  OAI21_X1 U20933 ( .B1(n17764), .B2(n17744), .A(n17739), .ZN(P3_U2781) );
  AOI22_X1 U20934 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17767), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17752), .ZN(n17740) );
  OAI21_X1 U20935 ( .B1(n17741), .B2(n21455), .A(n17740), .ZN(P3_U2782) );
  AOI22_X1 U20936 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17752), .ZN(n17742) );
  OAI21_X1 U20937 ( .B1(n18475), .B2(n17744), .A(n17742), .ZN(P3_U2783) );
  AOI22_X1 U20938 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17752), .ZN(n17743) );
  OAI21_X1 U20939 ( .B1(n18483), .B2(n17744), .A(n17743), .ZN(P3_U2784) );
  AOI22_X1 U20940 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17752), .ZN(n17745) );
  OAI21_X1 U20941 ( .B1(n18487), .B2(n21457), .A(n17745), .ZN(P3_U2785) );
  AOI22_X1 U20942 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17752), .ZN(n17746) );
  OAI21_X1 U20943 ( .B1(n21458), .B2(n21457), .A(n17746), .ZN(P3_U2786) );
  AOI22_X1 U20944 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17752), .ZN(n17747) );
  OAI21_X1 U20945 ( .B1(n18494), .B2(n21457), .A(n17747), .ZN(P3_U2787) );
  AOI22_X1 U20946 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17767), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17752), .ZN(n17748) );
  OAI21_X1 U20947 ( .B1(n17749), .B2(n21455), .A(n17748), .ZN(P3_U2788) );
  AOI22_X1 U20948 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17752), .ZN(n17750) );
  OAI21_X1 U20949 ( .B1(n18503), .B2(n21457), .A(n17750), .ZN(P3_U2789) );
  AOI22_X1 U20950 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17752), .ZN(n17751) );
  OAI21_X1 U20951 ( .B1(n18508), .B2(n21457), .A(n17751), .ZN(P3_U2790) );
  AOI22_X1 U20952 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17752), .ZN(n17753) );
  OAI21_X1 U20953 ( .B1(n17754), .B2(n21457), .A(n17753), .ZN(P3_U2791) );
  AOI22_X1 U20954 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17752), .ZN(n17755) );
  OAI21_X1 U20955 ( .B1(n17756), .B2(n21457), .A(n17755), .ZN(P3_U2792) );
  AOI22_X1 U20956 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17752), .ZN(n17757) );
  OAI21_X1 U20957 ( .B1(n17758), .B2(n21457), .A(n17757), .ZN(P3_U2793) );
  AOI22_X1 U20958 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17752), .ZN(n17759) );
  OAI21_X1 U20959 ( .B1(n21201), .B2(n21457), .A(n17759), .ZN(P3_U2794) );
  AOI22_X1 U20960 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17760), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17752), .ZN(n17761) );
  OAI21_X1 U20961 ( .B1(n21209), .B2(n21457), .A(n17761), .ZN(P3_U2795) );
  AOI22_X1 U20962 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17762), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17752), .ZN(n17763) );
  OAI21_X1 U20963 ( .B1(n17764), .B2(n21457), .A(n17763), .ZN(P3_U2796) );
  AOI22_X1 U20964 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17767), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17752), .ZN(n17765) );
  OAI21_X1 U20965 ( .B1(n17766), .B2(n21455), .A(n17765), .ZN(P3_U2797) );
  AOI22_X1 U20966 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17767), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17752), .ZN(n17768) );
  OAI21_X1 U20967 ( .B1(n17769), .B2(n21455), .A(n17768), .ZN(P3_U2798) );
  INV_X1 U20968 ( .A(n17771), .ZN(n17770) );
  NOR3_X1 U20969 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17971), .A3(
        n17770), .ZN(n17792) );
  INV_X1 U20970 ( .A(n18135), .ZN(n17889) );
  INV_X1 U20971 ( .A(n18089), .ZN(n17886) );
  OAI21_X1 U20972 ( .B1(n17771), .B2(n17886), .A(n18136), .ZN(n17772) );
  AOI21_X1 U20973 ( .B1(n17889), .B2(n17773), .A(n17772), .ZN(n17799) );
  OAI21_X1 U20974 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17856), .A(
        n17799), .ZN(n17793) );
  INV_X1 U20975 ( .A(n17971), .ZN(n17923) );
  NAND3_X1 U20976 ( .A1(n17775), .A2(n21214), .A3(n17923), .ZN(n17776) );
  OAI211_X1 U20977 ( .C1(n17985), .C2(n10154), .A(n17777), .B(n17776), .ZN(
        n17778) );
  AOI221_X1 U20978 ( .B1(n17792), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n17793), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17778), .ZN(
        n17788) );
  NOR2_X1 U20979 ( .A1(n18275), .A2(n18165), .ZN(n17816) );
  NAND2_X1 U20980 ( .A1(n18142), .A2(n17816), .ZN(n18145) );
  AOI22_X1 U20981 ( .A1(n18127), .A2(n18145), .B1(n17998), .B2(n17779), .ZN(
        n17808) );
  NAND2_X1 U20982 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17808), .ZN(
        n17795) );
  OAI211_X1 U20983 ( .C1(n17998), .C2(n18127), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17795), .ZN(n17787) );
  INV_X1 U20984 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18211) );
  NAND3_X1 U20985 ( .A1(n17781), .A2(n17844), .A3(n17780), .ZN(n17786) );
  OAI211_X1 U20986 ( .C1(n17784), .C2(n17783), .A(n18032), .B(n17782), .ZN(
        n17785) );
  NAND4_X1 U20987 ( .A1(n17788), .A2(n17787), .A3(n17786), .A4(n17785), .ZN(
        P3_U2802) );
  XOR2_X1 U20988 ( .A(n17789), .B(n9788), .Z(n18156) );
  OAI22_X1 U20989 ( .A1(n18407), .A2(n19070), .B1(n17985), .B2(n17790), .ZN(
        n17791) );
  AOI211_X1 U20990 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17793), .A(
        n17792), .B(n17791), .ZN(n17798) );
  NOR2_X1 U20991 ( .A1(n17794), .A2(n17850), .ZN(n17796) );
  OAI21_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17796), .A(
        n17795), .ZN(n17797) );
  OAI211_X1 U20993 ( .C1(n18156), .C2(n17967), .A(n17798), .B(n17797), .ZN(
        P3_U2803) );
  NAND2_X1 U20994 ( .A1(n18451), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18161) );
  INV_X1 U20995 ( .A(n18161), .ZN(n17803) );
  AOI221_X1 U20996 ( .B1(n17801), .B2(n17800), .C1(n18798), .C2(n17800), .A(
        n17799), .ZN(n17802) );
  AOI211_X1 U20997 ( .C1(n17804), .C2(n18129), .A(n17803), .B(n17802), .ZN(
        n17807) );
  XOR2_X1 U20998 ( .A(n18151), .B(n17805), .Z(n18160) );
  NAND2_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18148) );
  NOR3_X1 U21000 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18164), .A3(
        n18148), .ZN(n18157) );
  AOI22_X1 U21001 ( .A1(n18032), .A2(n18160), .B1(n17844), .B2(n18157), .ZN(
        n17806) );
  OAI211_X1 U21002 ( .C1(n17808), .C2(n18151), .A(n17807), .B(n17806), .ZN(
        P3_U2804) );
  NOR2_X1 U21003 ( .A1(n18278), .A2(n18165), .ZN(n17809) );
  XOR2_X1 U21004 ( .A(n17809), .B(n18164), .Z(n18177) );
  OAI22_X1 U21005 ( .A1(n17811), .A2(n18798), .B1(n17839), .B2(n18135), .ZN(
        n17810) );
  NOR2_X1 U21006 ( .A1(n18122), .A2(n17810), .ZN(n17833) );
  OAI21_X1 U21007 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17856), .A(
        n17833), .ZN(n17822) );
  INV_X1 U21008 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17812) );
  NAND2_X1 U21009 ( .A1(n17811), .A2(n17923), .ZN(n17825) );
  AOI221_X1 U21010 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n17824), .C2(n17812), .A(
        n17825), .ZN(n17815) );
  OAI22_X1 U21011 ( .A1(n18407), .A2(n19065), .B1(n17985), .B2(n17813), .ZN(
        n17814) );
  AOI211_X1 U21012 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17822), .A(
        n17815), .B(n17814), .ZN(n17821) );
  XOR2_X1 U21013 ( .A(n17816), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18173) );
  AOI21_X1 U21014 ( .B1(n17818), .B2(n16004), .A(n17817), .ZN(n17819) );
  XOR2_X1 U21015 ( .A(n17819), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18174) );
  AOI22_X1 U21016 ( .A1(n18127), .A2(n18173), .B1(n18032), .B2(n18174), .ZN(
        n17820) );
  OAI211_X1 U21017 ( .C1(n17977), .C2(n18177), .A(n17821), .B(n17820), .ZN(
        P3_U2805) );
  NAND2_X1 U21018 ( .A1(n17828), .A2(n18206), .ZN(n18186) );
  NAND2_X1 U21019 ( .A1(n18207), .A2(n17828), .ZN(n18184) );
  AOI22_X1 U21020 ( .A1(n17998), .A2(n18186), .B1(n18127), .B2(n18184), .ZN(
        n17846) );
  INV_X1 U21021 ( .A(n17822), .ZN(n17823) );
  NAND2_X1 U21022 ( .A1(n18446), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18193) );
  OAI221_X1 U21023 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17825), .C1(
        n17824), .C2(n17823), .A(n18193), .ZN(n17830) );
  AOI21_X1 U21024 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17827), .A(
        n17826), .ZN(n18182) );
  NAND2_X1 U21025 ( .A1(n17828), .A2(n10140), .ZN(n18180) );
  OAI22_X1 U21026 ( .A1(n18182), .A2(n17967), .B1(n17850), .B2(n18180), .ZN(
        n17829) );
  AOI211_X1 U21027 ( .C1(n17927), .C2(n17831), .A(n17830), .B(n17829), .ZN(
        n17832) );
  OAI21_X1 U21028 ( .B1(n17846), .B2(n10140), .A(n17832), .ZN(P3_U2806) );
  NOR2_X1 U21029 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17856), .ZN(
        n17840) );
  AOI221_X1 U21030 ( .B1(n17835), .B2(n17834), .C1(n18798), .C2(n17834), .A(
        n17833), .ZN(n17838) );
  OAI22_X1 U21031 ( .A1(n18407), .A2(n19062), .B1(n17985), .B2(n17836), .ZN(
        n17837) );
  AOI211_X1 U21032 ( .C1(n17840), .C2(n17839), .A(n17838), .B(n17837), .ZN(
        n17845) );
  AOI22_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16004), .B1(
        n17841), .B2(n17847), .ZN(n17842) );
  NAND2_X1 U21034 ( .A1(n17880), .A2(n17842), .ZN(n17843) );
  XOR2_X1 U21035 ( .A(n17843), .B(n18195), .Z(n18199) );
  INV_X1 U21036 ( .A(n17847), .ZN(n17848) );
  OAI21_X1 U21037 ( .B1(n9903), .B2(n17848), .A(n17880), .ZN(n17849) );
  XOR2_X1 U21038 ( .A(n17849), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n18210) );
  NOR2_X1 U21039 ( .A1(n17851), .A2(n17850), .ZN(n17861) );
  NAND2_X1 U21040 ( .A1(n17977), .A2(n18140), .ZN(n17874) );
  OAI22_X1 U21041 ( .A1(n17977), .A2(n18206), .B1(n18140), .B2(n18207), .ZN(
        n17932) );
  AOI21_X1 U21042 ( .B1(n17851), .B2(n17874), .A(n17932), .ZN(n17852) );
  INV_X1 U21043 ( .A(n17852), .ZN(n17871) );
  NAND2_X1 U21044 ( .A1(n9948), .A2(n17923), .ZN(n17864) );
  OAI21_X1 U21045 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17853), .ZN(n17859) );
  OAI22_X1 U21046 ( .A1(n9948), .A2(n17886), .B1(n17854), .B2(n18135), .ZN(
        n17855) );
  NOR2_X1 U21047 ( .A1(n18122), .A2(n17855), .ZN(n17875) );
  OAI21_X1 U21048 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17856), .A(
        n17875), .ZN(n17866) );
  AOI22_X1 U21049 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17866), .B1(
        n17927), .B2(n17857), .ZN(n17858) );
  NAND2_X1 U21050 ( .A1(n18451), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18213) );
  OAI211_X1 U21051 ( .C1(n17864), .C2(n17859), .A(n17858), .B(n18213), .ZN(
        n17860) );
  AOI221_X1 U21052 ( .B1(n17861), .B2(n18211), .C1(n17871), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17860), .ZN(n17862) );
  OAI21_X1 U21053 ( .B1(n17967), .B2(n18210), .A(n17862), .ZN(P3_U2808) );
  NAND2_X1 U21054 ( .A1(n18220), .A2(n17870), .ZN(n18224) );
  INV_X1 U21055 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17908) );
  NOR2_X1 U21056 ( .A1(n18247), .A2(n17908), .ZN(n18218) );
  NAND2_X1 U21057 ( .A1(n17933), .A2(n18218), .ZN(n17897) );
  NOR2_X1 U21058 ( .A1(n18407), .A2(n19057), .ZN(n18216) );
  OAI22_X1 U21059 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17864), .B1(
        n17863), .B2(n17985), .ZN(n17865) );
  AOI211_X1 U21060 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17866), .A(
        n18216), .B(n17865), .ZN(n17873) );
  AND3_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9788), .A3(
        n17867), .ZN(n17884) );
  AOI22_X1 U21062 ( .A1(n18220), .A2(n17884), .B1(n17905), .B2(n17868), .ZN(
        n17869) );
  XOR2_X1 U21063 ( .A(n17870), .B(n17869), .Z(n18217) );
  AOI22_X1 U21064 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17871), .B1(
        n18032), .B2(n18217), .ZN(n17872) );
  OAI211_X1 U21065 ( .C1(n18224), .C2(n17897), .A(n17873), .B(n17872), .ZN(
        P3_U2809) );
  NAND2_X1 U21066 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18218), .ZN(
        n18229) );
  AOI21_X1 U21067 ( .B1(n17874), .B2(n18229), .A(n17932), .ZN(n17896) );
  AOI221_X1 U21068 ( .B1(n17877), .B2(n17876), .C1(n18798), .C2(n17876), .A(
        n17875), .ZN(n17878) );
  NOR2_X1 U21069 ( .A1(n18407), .A2(n19056), .ZN(n18234) );
  AOI211_X1 U21070 ( .C1(n17879), .C2(n18129), .A(n17878), .B(n18234), .ZN(
        n17883) );
  OAI221_X1 U21071 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17903), 
        .C1(n18242), .C2(n17884), .A(n17880), .ZN(n17881) );
  XOR2_X1 U21072 ( .A(n18231), .B(n17881), .Z(n18225) );
  NOR2_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18229), .ZN(
        n18236) );
  AOI22_X1 U21074 ( .A1(n18032), .A2(n18225), .B1(n17933), .B2(n18236), .ZN(
        n17882) );
  OAI211_X1 U21075 ( .C1(n17896), .C2(n18231), .A(n17883), .B(n17882), .ZN(
        P3_U2810) );
  AOI21_X1 U21076 ( .B1(n17903), .B2(n17905), .A(n17884), .ZN(n17885) );
  XOR2_X1 U21077 ( .A(n18242), .B(n17885), .Z(n18239) );
  NAND2_X1 U21078 ( .A1(n17887), .A2(n17923), .ZN(n17900) );
  AOI221_X1 U21079 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17899), .C2(n17892), .A(
        n17900), .ZN(n17894) );
  OAI21_X1 U21080 ( .B1(n17887), .B2(n17886), .A(n18136), .ZN(n17914) );
  AOI21_X1 U21081 ( .B1(n17889), .B2(n17888), .A(n17914), .ZN(n17898) );
  AOI22_X1 U21082 ( .A1(n18451), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n17927), 
        .B2(n17890), .ZN(n17891) );
  OAI21_X1 U21083 ( .B1(n17898), .B2(n17892), .A(n17891), .ZN(n17893) );
  AOI211_X1 U21084 ( .C1(n18032), .C2(n18239), .A(n17894), .B(n17893), .ZN(
        n17895) );
  OAI221_X1 U21085 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17897), 
        .C1(n18242), .C2(n17896), .A(n17895), .ZN(P3_U2811) );
  AOI21_X1 U21086 ( .B1(n17933), .B2(n18247), .A(n17932), .ZN(n17919) );
  NAND2_X1 U21087 ( .A1(n18446), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18258) );
  OAI221_X1 U21088 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17900), .C1(
        n17899), .C2(n17898), .A(n18258), .ZN(n17901) );
  AOI21_X1 U21089 ( .B1(n17927), .B2(n17902), .A(n17901), .ZN(n17907) );
  AOI21_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n9788), .A(
        n17903), .ZN(n17904) );
  XOR2_X1 U21091 ( .A(n17905), .B(n17904), .Z(n18257) );
  NOR2_X1 U21092 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18247), .ZN(
        n18256) );
  AOI22_X1 U21093 ( .A1(n18032), .A2(n18257), .B1(n17933), .B2(n18256), .ZN(
        n17906) );
  OAI211_X1 U21094 ( .C1(n17919), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2812) );
  OAI21_X1 U21095 ( .B1(n17910), .B2(n18798), .A(n17909), .ZN(n17913) );
  OAI22_X1 U21096 ( .A1(n18119), .A2(n17911), .B1(n18407), .B2(n19050), .ZN(
        n17912) );
  AOI21_X1 U21097 ( .B1(n17914), .B2(n17913), .A(n17912), .ZN(n17918) );
  OAI21_X1 U21098 ( .B1(n17916), .B2(n18250), .A(n17915), .ZN(n18263) );
  NOR2_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15997), .ZN(
        n18262) );
  AOI22_X1 U21100 ( .A1(n18032), .A2(n18263), .B1(n17933), .B2(n18262), .ZN(
        n17917) );
  OAI211_X1 U21101 ( .C1(n17919), .C2(n18250), .A(n17918), .B(n17917), .ZN(
        P3_U2813) );
  INV_X1 U21102 ( .A(n18023), .ZN(n17996) );
  OAI21_X1 U21103 ( .B1(n18255), .B2(n17996), .A(n17920), .ZN(n17921) );
  XOR2_X1 U21104 ( .A(n17921), .B(n15997), .Z(n18274) );
  NOR2_X1 U21105 ( .A1(n17938), .A2(n17922), .ZN(n17930) );
  OAI211_X1 U21106 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17924), .B(n17923), .ZN(n17929) );
  INV_X1 U21107 ( .A(n17924), .ZN(n17935) );
  AOI21_X1 U21108 ( .B1(n18089), .B2(n17935), .A(n18122), .ZN(n17956) );
  OAI21_X1 U21109 ( .B1(n17925), .B2(n18135), .A(n17956), .ZN(n17937) );
  AOI22_X1 U21110 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17937), .B1(
        n17927), .B2(n17926), .ZN(n17928) );
  NAND2_X1 U21111 ( .A1(n18446), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18272) );
  OAI211_X1 U21112 ( .C1(n17930), .C2(n17929), .A(n17928), .B(n18272), .ZN(
        n17931) );
  AOI221_X1 U21113 ( .B1(n17933), .B2(n15997), .C1(n17932), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17931), .ZN(n17934) );
  OAI21_X1 U21114 ( .B1(n18274), .B2(n17967), .A(n17934), .ZN(P3_U2814) );
  NOR2_X1 U21115 ( .A1(n17971), .A2(n17935), .ZN(n17939) );
  NOR2_X1 U21116 ( .A1(n18407), .A2(n19045), .ZN(n17936) );
  AOI221_X1 U21117 ( .B1(n17939), .B2(n17938), .C1(n17937), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17936), .ZN(n17950) );
  INV_X1 U21118 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18328) );
  NAND3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18341), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17941) );
  OAI21_X1 U21120 ( .B1(n17979), .B2(n17941), .A(n17940), .ZN(n17942) );
  OAI221_X1 U21121 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18291), 
        .C1(n18328), .C2(n9788), .A(n17942), .ZN(n17943) );
  XOR2_X1 U21122 ( .A(n17944), .B(n17943), .Z(n18283) );
  NOR2_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17960), .ZN(
        n18280) );
  NAND2_X1 U21124 ( .A1(n17998), .A2(n18278), .ZN(n17947) );
  INV_X1 U21125 ( .A(n18293), .ZN(n17945) );
  NOR3_X1 U21126 ( .A1(n18332), .A2(n17945), .A3(n18291), .ZN(n17963) );
  NOR2_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17963), .ZN(
        n18288) );
  NAND2_X1 U21128 ( .A1(n18127), .A2(n18275), .ZN(n17946) );
  OAI22_X1 U21129 ( .A1(n18280), .A2(n17947), .B1(n18288), .B2(n17946), .ZN(
        n17948) );
  AOI21_X1 U21130 ( .B1(n18032), .B2(n18283), .A(n17948), .ZN(n17949) );
  OAI211_X1 U21131 ( .C1(n17985), .C2(n17951), .A(n17950), .B(n17949), .ZN(
        P3_U2815) );
  AOI21_X1 U21132 ( .B1(n18023), .B2(n18293), .A(n17952), .ZN(n17953) );
  XOR2_X1 U21133 ( .A(n17953), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18303) );
  NOR2_X1 U21134 ( .A1(n17954), .A2(n18798), .ZN(n18067) );
  NAND2_X1 U21135 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18067), .ZN(
        n18052) );
  INV_X1 U21136 ( .A(n18052), .ZN(n18026) );
  AND2_X1 U21137 ( .A1(n17955), .A2(n18026), .ZN(n18012) );
  NAND2_X1 U21138 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18012), .ZN(
        n18002) );
  AOI221_X1 U21139 ( .B1(n17972), .B2(n17957), .C1(n18002), .C2(n17957), .A(
        n17956), .ZN(n17958) );
  NOR2_X1 U21140 ( .A1(n18407), .A2(n19044), .ZN(n18297) );
  AOI211_X1 U21141 ( .C1(n17959), .C2(n18129), .A(n17958), .B(n18297), .ZN(
        n17966) );
  AOI21_X1 U21142 ( .B1(n18291), .B2(n17961), .A(n17960), .ZN(n18299) );
  NAND2_X1 U21143 ( .A1(n18293), .A2(n17962), .ZN(n17964) );
  AOI21_X1 U21144 ( .B1(n18291), .B2(n17964), .A(n17963), .ZN(n18298) );
  AOI22_X1 U21145 ( .A1(n17998), .A2(n18299), .B1(n18127), .B2(n18298), .ZN(
        n17965) );
  OAI211_X1 U21146 ( .C1(n18303), .C2(n17967), .A(n17966), .B(n17965), .ZN(
        P3_U2816) );
  INV_X1 U21147 ( .A(n17978), .ZN(n18317) );
  NAND2_X1 U21148 ( .A1(n18317), .A2(n21226), .ZN(n18315) );
  NAND2_X1 U21149 ( .A1(n18089), .A2(n17970), .ZN(n17968) );
  OAI211_X1 U21150 ( .C1(n17969), .C2(n18135), .A(n17968), .B(n18136), .ZN(
        n17989) );
  NOR2_X1 U21151 ( .A1(n17971), .A2(n17970), .ZN(n17988) );
  OAI211_X1 U21152 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17988), .B(n17972), .ZN(n17974) );
  NAND2_X1 U21153 ( .A1(n18451), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17973) );
  OAI211_X1 U21154 ( .C1(n17985), .C2(n17975), .A(n17974), .B(n17973), .ZN(
        n17976) );
  AOI21_X1 U21155 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17989), .A(
        n17976), .ZN(n17983) );
  NOR2_X1 U21156 ( .A1(n18332), .A2(n17978), .ZN(n18305) );
  OAI22_X1 U21157 ( .A1(n18307), .A2(n17977), .B1(n18305), .B2(n18140), .ZN(
        n17991) );
  OAI22_X1 U21158 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n9788), .B1(
        n17979), .B2(n17978), .ZN(n17980) );
  OAI21_X1 U21159 ( .B1(n9788), .B2(n9912), .A(n17980), .ZN(n17981) );
  XOR2_X1 U21160 ( .A(n17981), .B(n21226), .Z(n18304) );
  AOI22_X1 U21161 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17991), .B1(
        n18032), .B2(n18304), .ZN(n17982) );
  OAI211_X1 U21162 ( .C1(n18035), .C2(n18315), .A(n17983), .B(n17982), .ZN(
        P3_U2817) );
  NAND2_X1 U21163 ( .A1(n18451), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U21164 ( .B1(n17985), .B2(n17984), .A(n18326), .ZN(n17986) );
  AOI221_X1 U21165 ( .B1(n17989), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C1(
        n17988), .C2(n17987), .A(n17986), .ZN(n17994) );
  AOI21_X1 U21166 ( .B1(n18341), .B2(n18023), .A(n9912), .ZN(n17990) );
  XOR2_X1 U21167 ( .A(n17990), .B(n18328), .Z(n18324) );
  AOI22_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17991), .B1(
        n18032), .B2(n18324), .ZN(n17993) );
  INV_X1 U21169 ( .A(n18035), .ZN(n17999) );
  NAND3_X1 U21170 ( .A1(n18341), .A2(n18328), .A3(n17999), .ZN(n17992) );
  NAND3_X1 U21171 ( .A1(n17994), .A2(n17993), .A3(n17992), .ZN(P3_U2818) );
  INV_X1 U21172 ( .A(n18000), .ZN(n18339) );
  NAND2_X1 U21173 ( .A1(n18339), .A2(n18001), .ZN(n18345) );
  OAI21_X1 U21174 ( .B1(n18000), .B2(n17996), .A(n17995), .ZN(n17997) );
  XNOR2_X1 U21175 ( .A(n18001), .B(n17997), .ZN(n18329) );
  AOI22_X1 U21176 ( .A1(n18332), .A2(n18127), .B1(n17998), .B2(n18330), .ZN(
        n18034) );
  NAND2_X1 U21177 ( .A1(n18000), .A2(n17999), .ZN(n18016) );
  AOI21_X1 U21178 ( .B1(n18034), .B2(n18016), .A(n18001), .ZN(n18007) );
  INV_X1 U21179 ( .A(n18068), .ZN(n18130) );
  OAI211_X1 U21180 ( .C1(n18012), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n18130), .B(n18002), .ZN(n18004) );
  NAND2_X1 U21181 ( .A1(n18446), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18003) );
  OAI211_X1 U21182 ( .C1(n18119), .C2(n18005), .A(n18004), .B(n18003), .ZN(
        n18006) );
  AOI211_X1 U21183 ( .C1(n18032), .C2(n18329), .A(n18007), .B(n18006), .ZN(
        n18008) );
  OAI21_X1 U21184 ( .B1(n18035), .B2(n18345), .A(n18008), .ZN(P3_U2819) );
  INV_X1 U21185 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18015) );
  NOR4_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n9788), .A3(
        n18015), .A4(n18009), .ZN(n18011) );
  INV_X1 U21187 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18360) );
  AOI221_X1 U21188 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18023), .C1(
        n18360), .C2(n18022), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18010) );
  AOI211_X1 U21189 ( .C1(n18023), .C2(n18339), .A(n18011), .B(n18010), .ZN(
        n18350) );
  NAND3_X1 U21190 ( .A1(n18041), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18026), .ZN(n18025) );
  AOI211_X1 U21191 ( .C1(n18025), .C2(n18013), .A(n18068), .B(n18012), .ZN(
        n18018) );
  AOI221_X1 U21192 ( .B1(n18034), .B2(n18016), .C1(n18015), .C2(n18016), .A(
        n18014), .ZN(n18017) );
  AOI211_X1 U21193 ( .C1(n18350), .C2(n18032), .A(n18018), .B(n18017), .ZN(
        n18020) );
  NAND2_X1 U21194 ( .A1(n18451), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18019) );
  OAI211_X1 U21195 ( .C1(n18119), .C2(n18021), .A(n18020), .B(n18019), .ZN(
        P3_U2820) );
  NOR2_X1 U21196 ( .A1(n18023), .A2(n18022), .ZN(n18024) );
  XOR2_X1 U21197 ( .A(n18024), .B(n18360), .Z(n18357) );
  NOR2_X1 U21198 ( .A1(n18407), .A2(n19033), .ZN(n18031) );
  INV_X1 U21199 ( .A(n18025), .ZN(n18029) );
  AOI22_X1 U21200 ( .A1(n18041), .A2(n18026), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18130), .ZN(n18028) );
  OAI22_X1 U21201 ( .A1(n18029), .A2(n18028), .B1(n18119), .B2(n18027), .ZN(
        n18030) );
  AOI211_X1 U21202 ( .C1(n18032), .C2(n18357), .A(n18031), .B(n18030), .ZN(
        n18033) );
  OAI221_X1 U21203 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18035), .C1(
        n18360), .C2(n18034), .A(n18033), .ZN(P3_U2821) );
  OAI21_X1 U21204 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18037), .A(
        n18036), .ZN(n18377) );
  NOR2_X1 U21205 ( .A1(n18407), .A2(n19032), .ZN(n18368) );
  OAI211_X1 U21206 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18038), .B(n18866), .ZN(n18040)
         );
  AOI21_X1 U21207 ( .B1(n18089), .B2(n18039), .A(n18122), .ZN(n18061) );
  OAI22_X1 U21208 ( .A1(n18041), .A2(n18040), .B1(n21294), .B2(n18061), .ZN(
        n18042) );
  AOI211_X1 U21209 ( .C1(n18043), .C2(n18129), .A(n18368), .B(n18042), .ZN(
        n18049) );
  OAI21_X1 U21210 ( .B1(n9788), .B2(n9881), .A(n18044), .ZN(n18372) );
  OAI221_X1 U21211 ( .B1(n18047), .B2(n18372), .C1(n18046), .C2(n9881), .A(
        n18045), .ZN(n18048) );
  OAI211_X1 U21212 ( .C1(n18140), .C2(n18377), .A(n18049), .B(n18048), .ZN(
        P3_U2822) );
  OAI21_X1 U21213 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18051), .A(
        n18050), .ZN(n18381) );
  OAI22_X1 U21214 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18052), .B1(
        n18139), .B2(n18381), .ZN(n18059) );
  OAI21_X1 U21215 ( .B1(n18055), .B2(n18054), .A(n18053), .ZN(n18056) );
  XOR2_X1 U21216 ( .A(n18056), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18387) );
  OAI22_X1 U21217 ( .A1(n18119), .A2(n18057), .B1(n18140), .B2(n18387), .ZN(
        n18058) );
  AOI211_X1 U21218 ( .C1(n18451), .C2(P3_REIP_REG_7__SCAN_IN), .A(n18059), .B(
        n18058), .ZN(n18060) );
  OAI21_X1 U21219 ( .B1(n18062), .B2(n18061), .A(n18060), .ZN(P3_U2823) );
  OAI21_X1 U21220 ( .B1(n18065), .B2(n18064), .A(n18063), .ZN(n18396) );
  AOI22_X1 U21221 ( .A1(n18446), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18067), 
        .B2(n18066), .ZN(n18074) );
  NOR2_X1 U21222 ( .A1(n18068), .A2(n18067), .ZN(n18084) );
  OAI21_X1 U21223 ( .B1(n18070), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18069), .ZN(n18391) );
  OAI22_X1 U21224 ( .A1(n18119), .A2(n18071), .B1(n18140), .B2(n18391), .ZN(
        n18072) );
  AOI21_X1 U21225 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18084), .A(
        n18072), .ZN(n18073) );
  OAI211_X1 U21226 ( .C1(n18139), .C2(n18396), .A(n18074), .B(n18073), .ZN(
        P3_U2824) );
  OAI21_X1 U21227 ( .B1(n18077), .B2(n18076), .A(n18075), .ZN(n18402) );
  OAI21_X1 U21228 ( .B1(n18080), .B2(n18079), .A(n18078), .ZN(n18081) );
  XOR2_X1 U21229 ( .A(n18081), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18397) );
  OAI22_X1 U21230 ( .A1(n18407), .A2(n19025), .B1(n18139), .B2(n18397), .ZN(
        n18082) );
  AOI21_X1 U21231 ( .B1(n18083), .B2(n18129), .A(n18082), .ZN(n18087) );
  OAI221_X1 U21232 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18085), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18136), .A(n18084), .ZN(n18086) );
  OAI211_X1 U21233 ( .C1(n18140), .C2(n18402), .A(n18087), .B(n18086), .ZN(
        P3_U2825) );
  AOI21_X1 U21234 ( .B1(n18089), .B2(n18088), .A(n18122), .ZN(n18108) );
  OAI21_X1 U21235 ( .B1(n18092), .B2(n18091), .A(n18090), .ZN(n18406) );
  OAI22_X1 U21236 ( .A1(n18139), .A2(n18406), .B1(n18798), .B2(n18093), .ZN(
        n18098) );
  OAI21_X1 U21237 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18095), .A(
        n18094), .ZN(n18413) );
  OAI22_X1 U21238 ( .A1(n18119), .A2(n18096), .B1(n18140), .B2(n18413), .ZN(
        n18097) );
  AOI211_X1 U21239 ( .C1(n18451), .C2(P3_REIP_REG_4__SCAN_IN), .A(n18098), .B(
        n18097), .ZN(n18099) );
  OAI21_X1 U21240 ( .B1(n18108), .B2(n18100), .A(n18099), .ZN(P3_U2826) );
  OAI21_X1 U21241 ( .B1(n18103), .B2(n18102), .A(n18101), .ZN(n18416) );
  AOI21_X1 U21242 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18136), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18107) );
  OAI21_X1 U21243 ( .B1(n18106), .B2(n18105), .A(n18104), .ZN(n18417) );
  OAI22_X1 U21244 ( .A1(n18108), .A2(n18107), .B1(n18139), .B2(n18417), .ZN(
        n18109) );
  AOI21_X1 U21245 ( .B1(n18110), .B2(n18129), .A(n18109), .ZN(n18111) );
  NAND2_X1 U21246 ( .A1(n18451), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18420) );
  OAI211_X1 U21247 ( .C1(n18140), .C2(n18416), .A(n18111), .B(n18420), .ZN(
        P3_U2827) );
  OAI21_X1 U21248 ( .B1(n18114), .B2(n18113), .A(n18112), .ZN(n18432) );
  INV_X1 U21249 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18121) );
  OAI21_X1 U21250 ( .B1(n18117), .B2(n18116), .A(n18115), .ZN(n18430) );
  OAI22_X1 U21251 ( .A1(n18119), .A2(n18118), .B1(n18140), .B2(n18430), .ZN(
        n18120) );
  AOI221_X1 U21252 ( .B1(n18122), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18866), .C2(n18121), .A(n18120), .ZN(n18123) );
  NAND2_X1 U21253 ( .A1(n18451), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18435) );
  OAI211_X1 U21254 ( .C1(n18139), .C2(n18432), .A(n18123), .B(n18435), .ZN(
        P3_U2828) );
  OAI21_X1 U21255 ( .B1(n18125), .B2(n18133), .A(n18124), .ZN(n18450) );
  NAND2_X1 U21256 ( .A1(n19118), .A2(n18134), .ZN(n18126) );
  XNOR2_X1 U21257 ( .A(n18126), .B(n18125), .ZN(n18445) );
  AOI22_X1 U21258 ( .A1(n18446), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18127), 
        .B2(n18445), .ZN(n18132) );
  AOI22_X1 U21259 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18128), .ZN(n18131) );
  OAI211_X1 U21260 ( .C1(n18139), .C2(n18450), .A(n18132), .B(n18131), .ZN(
        P3_U2829) );
  AOI21_X1 U21261 ( .B1(n18134), .B2(n19118), .A(n18133), .ZN(n18453) );
  INV_X1 U21262 ( .A(n18453), .ZN(n18455) );
  NAND3_X1 U21263 ( .A1(n19100), .A2(n18136), .A3(n18135), .ZN(n18137) );
  AOI22_X1 U21264 ( .A1(n18451), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18137), .ZN(n18138) );
  OAI221_X1 U21265 ( .B1(n18453), .B2(n18140), .C1(n18455), .C2(n18139), .A(
        n18138), .ZN(P3_U2830) );
  NOR2_X1 U21266 ( .A1(n18141), .A2(n18196), .ZN(n18152) );
  OAI22_X1 U21267 ( .A1(n18929), .A2(n18142), .B1(n18952), .B2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18143) );
  AOI211_X1 U21268 ( .C1(n18974), .C2(n18145), .A(n18144), .B(n18143), .ZN(
        n18149) );
  OAI21_X1 U21269 ( .B1(n18211), .B2(n18950), .A(n18146), .ZN(n18205) );
  NAND3_X1 U21270 ( .A1(n18147), .A2(n18203), .A3(n18205), .ZN(n18185) );
  OAI21_X1 U21271 ( .B1(n18148), .B2(n18185), .A(n10005), .ZN(n18169) );
  AOI22_X1 U21272 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18388), .B1(
        n18439), .B2(n18153), .ZN(n18155) );
  NAND2_X1 U21273 ( .A1(n18451), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18154) );
  OAI211_X1 U21274 ( .C1(n18156), .C2(n18302), .A(n18155), .B(n18154), .ZN(
        P3_U2835) );
  INV_X1 U21275 ( .A(n18196), .ZN(n18158) );
  AOI22_X1 U21276 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18159), .B1(
        n18158), .B2(n18157), .ZN(n18163) );
  AOI22_X1 U21277 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18388), .B1(
        n18373), .B2(n18160), .ZN(n18162) );
  OAI211_X1 U21278 ( .C1(n18163), .C2(n18457), .A(n18162), .B(n18161), .ZN(
        P3_U2836) );
  NOR2_X1 U21279 ( .A1(n18407), .A2(n19065), .ZN(n18172) );
  INV_X1 U21280 ( .A(n18202), .ZN(n18245) );
  AOI211_X1 U21281 ( .C1(n18947), .C2(n18165), .A(n18245), .B(n18164), .ZN(
        n18170) );
  AOI21_X1 U21282 ( .B1(n18167), .B2(n18166), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18168) );
  AOI211_X1 U21283 ( .C1(n18170), .C2(n18169), .A(n18168), .B(n18457), .ZN(
        n18171) );
  AOI211_X1 U21284 ( .C1(n18388), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18172), .B(n18171), .ZN(n18176) );
  AOI22_X1 U21285 ( .A1(n18373), .A2(n18174), .B1(n18456), .B2(n18173), .ZN(
        n18175) );
  OAI211_X1 U21286 ( .C1(n18178), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        P3_U2837) );
  NOR2_X1 U21287 ( .A1(n18179), .A2(n18457), .ZN(n18235) );
  INV_X1 U21288 ( .A(n18235), .ZN(n18181) );
  OAI22_X1 U21289 ( .A1(n18302), .A2(n18182), .B1(n18181), .B2(n18180), .ZN(
        n18183) );
  INV_X1 U21290 ( .A(n18183), .ZN(n18194) );
  INV_X1 U21291 ( .A(n18184), .ZN(n18188) );
  AOI22_X1 U21292 ( .A1(n18331), .A2(n18186), .B1(n10005), .B2(n18185), .ZN(
        n18187) );
  OAI211_X1 U21293 ( .C1(n18188), .C2(n19131), .A(n18187), .B(n18440), .ZN(
        n18191) );
  AOI211_X1 U21294 ( .C1(n18947), .C2(n18189), .A(n18245), .B(n18191), .ZN(
        n18190) );
  AOI21_X1 U21295 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18190), .A(
        n18446), .ZN(n18198) );
  OAI211_X1 U21296 ( .C1(n18367), .C2(n18191), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18198), .ZN(n18192) );
  NAND3_X1 U21297 ( .A1(n18194), .A2(n18193), .A3(n18192), .ZN(P3_U2838) );
  OAI21_X1 U21298 ( .B1(n18388), .B2(n18196), .A(n18195), .ZN(n18197) );
  AOI22_X1 U21299 ( .A1(n18373), .A2(n18199), .B1(n18198), .B2(n18197), .ZN(
        n18200) );
  OAI21_X1 U21300 ( .B1(n18407), .B2(n19062), .A(n18200), .ZN(P3_U2839) );
  OAI21_X1 U21301 ( .B1(n18244), .B2(n18229), .A(n18458), .ZN(n18201) );
  OAI211_X1 U21302 ( .C1(n18218), .C2(n18923), .A(n18202), .B(n18201), .ZN(
        n18226) );
  NAND2_X1 U21303 ( .A1(n19131), .A2(n18306), .ZN(n18246) );
  INV_X1 U21304 ( .A(n18246), .ZN(n18338) );
  OAI22_X1 U21305 ( .A1(n18220), .A2(n18340), .B1(n18203), .B2(n18338), .ZN(
        n18204) );
  NOR2_X1 U21306 ( .A1(n18226), .A2(n18204), .ZN(n18219) );
  OAI211_X1 U21307 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n18340), .A(
        n18219), .B(n18205), .ZN(n18208) );
  OAI22_X1 U21308 ( .A1(n18207), .A2(n19131), .B1(n18206), .B2(n18306), .ZN(
        n18227) );
  OAI22_X1 U21309 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18209), .B1(
        n18208), .B2(n18227), .ZN(n18215) );
  OAI22_X1 U21310 ( .A1(n18211), .A2(n18440), .B1(n18302), .B2(n18210), .ZN(
        n18212) );
  INV_X1 U21311 ( .A(n18212), .ZN(n18214) );
  OAI211_X1 U21312 ( .C1(n18457), .C2(n18215), .A(n18214), .B(n18213), .ZN(
        P3_U2840) );
  NAND2_X1 U21313 ( .A1(n18218), .A2(n18235), .ZN(n18243) );
  AOI21_X1 U21314 ( .B1(n18373), .B2(n18217), .A(n18216), .ZN(n18223) );
  AOI21_X1 U21315 ( .B1(n18266), .B2(n18218), .A(n18929), .ZN(n18228) );
  NOR2_X1 U21316 ( .A1(n18457), .A2(n18227), .ZN(n18268) );
  OAI211_X1 U21317 ( .C1(n18929), .C2(n18220), .A(n18219), .B(n18268), .ZN(
        n18221) );
  OAI211_X1 U21318 ( .C1(n18228), .C2(n18221), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18407), .ZN(n18222) );
  OAI211_X1 U21319 ( .C1(n18243), .C2(n18224), .A(n18223), .B(n18222), .ZN(
        P3_U2841) );
  INV_X1 U21320 ( .A(n18225), .ZN(n18238) );
  OR4_X1 U21321 ( .A1(n18388), .A2(n18228), .A3(n18227), .A4(n18226), .ZN(
        n18230) );
  OAI221_X1 U21322 ( .B1(n18230), .B2(n18229), .C1(n18230), .C2(n18246), .A(
        n18407), .ZN(n18241) );
  NAND2_X1 U21323 ( .A1(n18929), .A2(n18923), .ZN(n18438) );
  NAND3_X1 U21324 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18242), .A3(n18438), 
        .ZN(n18232) );
  AOI21_X1 U21325 ( .B1(n18241), .B2(n18232), .A(n18231), .ZN(n18233) );
  AOI211_X1 U21326 ( .C1(n18236), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        n18237) );
  OAI21_X1 U21327 ( .B1(n18302), .B2(n18238), .A(n18237), .ZN(P3_U2842) );
  AOI22_X1 U21328 ( .A1(n18446), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18373), 
        .B2(n18239), .ZN(n18240) );
  OAI221_X1 U21329 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18243), 
        .C1(n18242), .C2(n18241), .A(n18240), .ZN(P3_U2843) );
  NOR2_X1 U21330 ( .A1(n18929), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18403) );
  NOR3_X1 U21331 ( .A1(n18403), .A2(n18244), .A3(n15997), .ZN(n18249) );
  AOI221_X1 U21332 ( .B1(n18947), .B2(n18247), .C1(n18246), .C2(n18247), .A(
        n18245), .ZN(n18248) );
  OAI211_X1 U21333 ( .C1(n18405), .C2(n18249), .A(n18268), .B(n18248), .ZN(
        n18261) );
  OAI221_X1 U21334 ( .B1(n18261), .B2(n10005), .C1(n18261), .C2(n18250), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18260) );
  NAND2_X1 U21335 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18252) );
  OAI22_X1 U21336 ( .A1(n18923), .A2(n18425), .B1(n18252), .B2(n18251), .ZN(
        n18253) );
  OAI21_X1 U21337 ( .B1(n18320), .B2(n18319), .A(n18439), .ZN(n18361) );
  NOR2_X1 U21338 ( .A1(n18255), .A2(n18361), .ZN(n18270) );
  AOI22_X1 U21339 ( .A1(n18373), .A2(n18257), .B1(n18256), .B2(n18270), .ZN(
        n18259) );
  OAI211_X1 U21340 ( .C1(n18451), .C2(n18260), .A(n18259), .B(n18258), .ZN(
        P3_U2844) );
  NAND2_X1 U21341 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18261), .ZN(
        n18265) );
  AOI22_X1 U21342 ( .A1(n18373), .A2(n18263), .B1(n18270), .B2(n18262), .ZN(
        n18264) );
  OAI221_X1 U21343 ( .B1(n18451), .B2(n18265), .C1(n18407), .C2(n19050), .A(
        n18264), .ZN(P3_U2845) );
  INV_X1 U21344 ( .A(n18367), .ZN(n18269) );
  AOI21_X1 U21345 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18929), .A(
        n18266), .ZN(n18267) );
  NAND2_X1 U21346 ( .A1(n18458), .A2(n18353), .ZN(n18336) );
  OAI21_X1 U21347 ( .B1(n18334), .B2(n18923), .A(n18336), .ZN(n18309) );
  AOI211_X1 U21348 ( .C1(n18276), .C2(n18346), .A(n18267), .B(n18309), .ZN(
        n18282) );
  AOI221_X1 U21349 ( .B1(n18269), .B2(n18268), .C1(n18282), .C2(n18268), .A(
        n18446), .ZN(n18271) );
  AOI22_X1 U21350 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18271), .B1(
        n18270), .B2(n15997), .ZN(n18273) );
  OAI211_X1 U21351 ( .C1(n18274), .C2(n18302), .A(n18273), .B(n18272), .ZN(
        P3_U2846) );
  NAND2_X1 U21352 ( .A1(n18456), .A2(n18275), .ZN(n18287) );
  AOI22_X1 U21353 ( .A1(n18451), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18388), .ZN(n18286) );
  INV_X1 U21354 ( .A(n18276), .ZN(n18277) );
  AOI21_X1 U21355 ( .B1(n18277), .B2(n18320), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18281) );
  NAND2_X1 U21356 ( .A1(n18331), .A2(n18278), .ZN(n18279) );
  OAI22_X1 U21357 ( .A1(n18282), .A2(n18281), .B1(n18280), .B2(n18279), .ZN(
        n18284) );
  AOI22_X1 U21358 ( .A1(n18439), .A2(n18284), .B1(n18373), .B2(n18283), .ZN(
        n18285) );
  OAI211_X1 U21359 ( .C1(n18288), .C2(n18287), .A(n18286), .B(n18285), .ZN(
        P3_U2847) );
  AOI21_X1 U21360 ( .B1(n18317), .B2(n18334), .A(n18923), .ZN(n18292) );
  AOI21_X1 U21361 ( .B1(n18317), .B2(n18316), .A(n18929), .ZN(n18312) );
  INV_X1 U21362 ( .A(n18438), .ZN(n18289) );
  OAI22_X1 U21363 ( .A1(n18952), .A2(n18293), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18289), .ZN(n18290) );
  NOR4_X1 U21364 ( .A1(n18292), .A2(n18312), .A3(n18291), .A4(n18290), .ZN(
        n18295) );
  AOI21_X1 U21365 ( .B1(n18293), .B2(n18320), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18294) );
  AOI211_X1 U21366 ( .C1(n18295), .C2(n18336), .A(n18294), .B(n18457), .ZN(
        n18296) );
  AOI211_X1 U21367 ( .C1(n18388), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18297), .B(n18296), .ZN(n18301) );
  AOI22_X1 U21368 ( .A1(n18374), .A2(n18299), .B1(n18456), .B2(n18298), .ZN(
        n18300) );
  OAI211_X1 U21369 ( .C1(n18303), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2848) );
  AOI22_X1 U21370 ( .A1(n18451), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18373), 
        .B2(n18304), .ZN(n18314) );
  INV_X1 U21371 ( .A(n18341), .ZN(n18310) );
  OAI22_X1 U21372 ( .A1(n18307), .A2(n18306), .B1(n18305), .B2(n19131), .ZN(
        n18308) );
  AOI211_X1 U21373 ( .C1(n18310), .C2(n18346), .A(n18309), .B(n18308), .ZN(
        n18323) );
  OAI211_X1 U21374 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18340), .A(
        n18439), .B(n18323), .ZN(n18311) );
  OAI211_X1 U21375 ( .C1(n18312), .C2(n18311), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18407), .ZN(n18313) );
  OAI211_X1 U21376 ( .C1(n18361), .C2(n18315), .A(n18314), .B(n18313), .ZN(
        P3_U2849) );
  NAND2_X1 U21377 ( .A1(n18317), .A2(n18316), .ZN(n18318) );
  OAI21_X1 U21378 ( .B1(n18328), .B2(n18950), .A(n18318), .ZN(n18322) );
  OAI21_X1 U21379 ( .B1(n18320), .B2(n18319), .A(n18341), .ZN(n18321) );
  AOI22_X1 U21380 ( .A1(n18323), .A2(n18322), .B1(n18328), .B2(n18321), .ZN(
        n18325) );
  AOI22_X1 U21381 ( .A1(n18439), .A2(n18325), .B1(n18373), .B2(n18324), .ZN(
        n18327) );
  OAI211_X1 U21382 ( .C1(n18440), .C2(n18328), .A(n18327), .B(n18326), .ZN(
        P3_U2850) );
  AOI22_X1 U21383 ( .A1(n18446), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18373), 
        .B2(n18329), .ZN(n18344) );
  AOI22_X1 U21384 ( .A1(n18974), .A2(n18332), .B1(n18331), .B2(n18330), .ZN(
        n18333) );
  OAI211_X1 U21385 ( .C1(n18334), .C2(n18923), .A(n18439), .B(n18333), .ZN(
        n18355) );
  AOI221_X1 U21386 ( .B1(n18360), .B2(n18950), .C1(n18335), .C2(n18950), .A(
        n18355), .ZN(n18337) );
  OAI211_X1 U21387 ( .C1(n18339), .C2(n18338), .A(n18337), .B(n18336), .ZN(
        n18347) );
  OAI22_X1 U21388 ( .A1(n18929), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18341), .B2(n18340), .ZN(n18342) );
  OAI211_X1 U21389 ( .C1(n18347), .C2(n18342), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18407), .ZN(n18343) );
  OAI211_X1 U21390 ( .C1(n18345), .C2(n18361), .A(n18344), .B(n18343), .ZN(
        P3_U2851) );
  OAI221_X1 U21391 ( .B1(n18347), .B2(n18360), .C1(n18347), .C2(n18346), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18352) );
  INV_X1 U21392 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19035) );
  INV_X1 U21393 ( .A(n18361), .ZN(n18349) );
  NOR2_X1 U21394 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18360), .ZN(
        n18348) );
  AOI22_X1 U21395 ( .A1(n18373), .A2(n18350), .B1(n18349), .B2(n18348), .ZN(
        n18351) );
  OAI221_X1 U21396 ( .B1(n18451), .B2(n18352), .C1(n18407), .C2(n19035), .A(
        n18351), .ZN(P3_U2852) );
  OAI21_X1 U21397 ( .B1(n18353), .B2(n18403), .A(n10005), .ZN(n18354) );
  INV_X1 U21398 ( .A(n18354), .ZN(n18356) );
  OAI21_X1 U21399 ( .B1(n18356), .B2(n18355), .A(n18407), .ZN(n18359) );
  AOI22_X1 U21400 ( .A1(n18446), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18373), 
        .B2(n18357), .ZN(n18358) );
  OAI221_X1 U21401 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18361), .C1(
        n18360), .C2(n18359), .A(n18358), .ZN(P3_U2853) );
  INV_X1 U21402 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18378) );
  NOR2_X1 U21403 ( .A1(n18415), .A2(n18457), .ZN(n18362) );
  NAND2_X1 U21404 ( .A1(n18363), .A2(n18362), .ZN(n18392) );
  NOR3_X1 U21405 ( .A1(n18366), .A2(n18378), .A3(n18392), .ZN(n18371) );
  INV_X1 U21406 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18370) );
  AOI221_X1 U21407 ( .B1(n18425), .B2(n18947), .C1(n18379), .C2(n18947), .A(
        n18403), .ZN(n18364) );
  OAI21_X1 U21408 ( .B1(n18405), .B2(n18365), .A(n18364), .ZN(n18389) );
  AOI211_X1 U21409 ( .C1(n18367), .C2(n18378), .A(n18366), .B(n18389), .ZN(
        n18383) );
  OAI21_X1 U21410 ( .B1(n18383), .B2(n18441), .A(n18440), .ZN(n18369) );
  AOI221_X1 U21411 ( .B1(n18371), .B2(n18370), .C1(n18369), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18368), .ZN(n18376) );
  AOI22_X1 U21412 ( .A1(n9881), .A2(n18374), .B1(n18373), .B2(n18372), .ZN(
        n18375) );
  OAI211_X1 U21413 ( .C1(n18431), .C2(n18377), .A(n18376), .B(n18375), .ZN(
        P3_U2854) );
  NOR2_X1 U21414 ( .A1(n18407), .A2(n19029), .ZN(n18385) );
  NOR3_X1 U21415 ( .A1(n18415), .A2(n18379), .A3(n18378), .ZN(n18380) );
  OAI21_X1 U21416 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18380), .A(
        n18439), .ZN(n18382) );
  INV_X1 U21417 ( .A(n18454), .ZN(n18449) );
  OAI22_X1 U21418 ( .A1(n18383), .A2(n18382), .B1(n18449), .B2(n18381), .ZN(
        n18384) );
  AOI211_X1 U21419 ( .C1(n18388), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18385), .B(n18384), .ZN(n18386) );
  OAI21_X1 U21420 ( .B1(n18431), .B2(n18387), .A(n18386), .ZN(P3_U2855) );
  AOI21_X1 U21421 ( .B1(n18389), .B2(n18439), .A(n18388), .ZN(n18390) );
  INV_X1 U21422 ( .A(n18390), .ZN(n18399) );
  OAI22_X1 U21423 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18392), .B1(
        n18391), .B2(n18431), .ZN(n18393) );
  AOI21_X1 U21424 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18399), .A(
        n18393), .ZN(n18395) );
  NAND2_X1 U21425 ( .A1(n18446), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18394) );
  OAI211_X1 U21426 ( .C1(n18449), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2856) );
  OAI22_X1 U21427 ( .A1(n18407), .A2(n19025), .B1(n18449), .B2(n18397), .ZN(
        n18398) );
  AOI21_X1 U21428 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18399), .A(
        n18398), .ZN(n18401) );
  NOR3_X1 U21429 ( .A1(n18415), .A2(n18457), .A3(n18422), .ZN(n18411) );
  NAND3_X1 U21430 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18411), .A3(
        n21212), .ZN(n18400) );
  OAI211_X1 U21431 ( .C1(n18402), .C2(n18431), .A(n18401), .B(n18400), .ZN(
        P3_U2857) );
  AOI21_X1 U21432 ( .B1(n18425), .B2(n18947), .A(n18403), .ZN(n18404) );
  OAI21_X1 U21433 ( .B1(n18405), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18404), .ZN(n18423) );
  AOI211_X1 U21434 ( .C1(n10005), .C2(n18437), .A(n18422), .B(n18423), .ZN(
        n18414) );
  OAI21_X1 U21435 ( .B1(n18414), .B2(n18441), .A(n18440), .ZN(n18409) );
  OAI22_X1 U21436 ( .A1(n18407), .A2(n19023), .B1(n18449), .B2(n18406), .ZN(
        n18408) );
  AOI221_X1 U21437 ( .B1(n18411), .B2(n18410), .C1(n18409), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18408), .ZN(n18412) );
  OAI21_X1 U21438 ( .B1(n18431), .B2(n18413), .A(n18412), .ZN(P3_U2858) );
  AOI211_X1 U21439 ( .C1(n18415), .C2(n18422), .A(n18414), .B(n18457), .ZN(
        n18419) );
  OAI22_X1 U21440 ( .A1(n18449), .A2(n18417), .B1(n18431), .B2(n18416), .ZN(
        n18418) );
  NOR2_X1 U21441 ( .A1(n18419), .A2(n18418), .ZN(n18421) );
  OAI211_X1 U21442 ( .C1(n18440), .C2(n18422), .A(n18421), .B(n18420), .ZN(
        P3_U2859) );
  NOR2_X1 U21443 ( .A1(n19118), .A2(n10078), .ZN(n18424) );
  AOI21_X1 U21444 ( .B1(n18947), .B2(n18424), .A(n18423), .ZN(n18429) );
  NAND2_X1 U21445 ( .A1(n18947), .A2(n18425), .ZN(n18428) );
  NAND4_X1 U21446 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n10005), .A3(
        n18437), .A4(n18426), .ZN(n18427) );
  OAI211_X1 U21447 ( .C1(n18429), .C2(n18437), .A(n18428), .B(n18427), .ZN(
        n18434) );
  OAI22_X1 U21448 ( .A1(n18449), .A2(n18432), .B1(n18431), .B2(n18430), .ZN(
        n18433) );
  AOI21_X1 U21449 ( .B1(n18439), .B2(n18434), .A(n18433), .ZN(n18436) );
  OAI211_X1 U21450 ( .C1(n18440), .C2(n18437), .A(n18436), .B(n18435), .ZN(
        P3_U2860) );
  NAND3_X1 U21451 ( .A1(n18439), .A2(n19118), .A3(n18438), .ZN(n18460) );
  AOI21_X1 U21452 ( .B1(n18440), .B2(n18460), .A(n10078), .ZN(n18444) );
  NOR3_X1 U21453 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18442), .A3(
        n18441), .ZN(n18443) );
  AOI211_X1 U21454 ( .C1(n18456), .C2(n18445), .A(n18444), .B(n18443), .ZN(
        n18448) );
  NAND2_X1 U21455 ( .A1(n18446), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18447) );
  OAI211_X1 U21456 ( .C1(n18450), .C2(n18449), .A(n18448), .B(n18447), .ZN(
        P3_U2861) );
  AND2_X1 U21457 ( .A1(n18451), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18452) );
  AOI221_X1 U21458 ( .B1(n18456), .B2(n18455), .C1(n18454), .C2(n18453), .A(
        n18452), .ZN(n18461) );
  OAI211_X1 U21459 ( .C1(n18458), .C2(n18457), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18407), .ZN(n18459) );
  NAND3_X1 U21460 ( .A1(n18461), .A2(n18460), .A3(n18459), .ZN(P3_U2862) );
  AOI21_X1 U21461 ( .B1(n18464), .B2(n18463), .A(n18462), .ZN(n18979) );
  INV_X1 U21462 ( .A(n18465), .ZN(n18515) );
  OAI21_X1 U21463 ( .B1(n18979), .B2(n18515), .A(n18473), .ZN(n18466) );
  OAI221_X1 U21464 ( .B1(n18956), .B2(n19148), .C1(n18956), .C2(n18473), .A(
        n18466), .ZN(P3_U2863) );
  NAND2_X1 U21465 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18626) );
  AOI21_X1 U21466 ( .B1(n18626), .B2(n18468), .A(n18467), .ZN(n18472) );
  INV_X1 U21467 ( .A(n18828), .ZN(n18652) );
  AOI22_X1 U21468 ( .A1(n18652), .A2(n18473), .B1(n18469), .B2(n18468), .ZN(
        n18471) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18472), .B1(
        n18471), .B2(n18963), .ZN(P3_U2865) );
  INV_X1 U21470 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18966) );
  NAND2_X1 U21471 ( .A1(n18963), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18699) );
  INV_X1 U21472 ( .A(n18699), .ZN(n18747) );
  NAND2_X1 U21473 ( .A1(n18966), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18650) );
  INV_X1 U21474 ( .A(n18650), .ZN(n18604) );
  NOR2_X1 U21475 ( .A1(n18747), .A2(n18604), .ZN(n18470) );
  OAI22_X1 U21476 ( .A1(n18472), .A2(n18966), .B1(n18471), .B2(n18470), .ZN(
        P3_U2866) );
  NOR2_X1 U21477 ( .A1(n18967), .A2(n18473), .ZN(P3_U2867) );
  INV_X1 U21478 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18474) );
  NOR2_X1 U21479 ( .A1(n18798), .A2(n18474), .ZN(n18862) );
  NOR2_X1 U21480 ( .A1(n18966), .A2(n18626), .ZN(n18864) );
  INV_X1 U21481 ( .A(n18864), .ZN(n18860) );
  NOR2_X2 U21482 ( .A1(n18860), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18855) );
  INV_X1 U21483 ( .A(n18855), .ZN(n18531) );
  NAND2_X1 U21484 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18800) );
  NAND2_X1 U21485 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18958), .ZN(
        n18698) );
  NOR2_X2 U21486 ( .A1(n18800), .A2(n18698), .ZN(n18912) );
  NAND2_X1 U21487 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18866), .ZN(n18870) );
  INV_X1 U21488 ( .A(n18870), .ZN(n18826) );
  NOR2_X2 U21489 ( .A1(n18516), .A2(n18475), .ZN(n18861) );
  NAND2_X1 U21490 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18864), .ZN(
        n18551) );
  INV_X1 U21491 ( .A(n18551), .ZN(n18914) );
  NAND2_X1 U21492 ( .A1(n18958), .A2(n18956), .ZN(n18959) );
  NAND2_X1 U21493 ( .A1(n18963), .A2(n18966), .ZN(n18536) );
  NOR2_X2 U21494 ( .A1(n18959), .A2(n18536), .ZN(n18577) );
  NOR2_X1 U21495 ( .A1(n18914), .A2(n18577), .ZN(n18537) );
  NOR2_X1 U21496 ( .A1(n18982), .A2(n18537), .ZN(n18509) );
  AOI22_X1 U21497 ( .A1(n18912), .A2(n18826), .B1(n18861), .B2(n18509), .ZN(
        n18481) );
  INV_X1 U21498 ( .A(n18516), .ZN(n18831) );
  NOR2_X1 U21499 ( .A1(n18855), .A2(n18912), .ZN(n18827) );
  OAI21_X1 U21500 ( .B1(n18827), .B2(n18828), .A(n18537), .ZN(n18476) );
  OAI211_X1 U21501 ( .C1(n18577), .C2(n19091), .A(n18831), .B(n18476), .ZN(
        n18512) );
  NAND2_X1 U21502 ( .A1(n18478), .A2(n18477), .ZN(n18510) );
  NOR2_X2 U21503 ( .A1(n18479), .A2(n18510), .ZN(n18867) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18867), .ZN(n18480) );
  OAI211_X1 U21505 ( .C1(n18834), .C2(n18531), .A(n18481), .B(n18480), .ZN(
        P3_U2868) );
  NOR2_X1 U21506 ( .A1(n18798), .A2(n18482), .ZN(n18835) );
  NAND2_X1 U21507 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18866), .ZN(n18838) );
  INV_X1 U21508 ( .A(n18838), .ZN(n18871) );
  NOR2_X2 U21509 ( .A1(n18516), .A2(n18483), .ZN(n18872) );
  AOI22_X1 U21510 ( .A1(n18912), .A2(n18871), .B1(n18509), .B2(n18872), .ZN(
        n18486) );
  NOR2_X2 U21511 ( .A1(n18484), .A2(n18510), .ZN(n18873) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18873), .ZN(n18485) );
  OAI211_X1 U21513 ( .C1(n18531), .C2(n18876), .A(n18486), .B(n18485), .ZN(
        P3_U2869) );
  NAND2_X1 U21514 ( .A1(n18866), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18755) );
  NOR2_X1 U21515 ( .A1(n19465), .A2(n18798), .ZN(n18752) );
  NOR2_X2 U21516 ( .A1(n18516), .A2(n18487), .ZN(n18877) );
  AOI22_X1 U21517 ( .A1(n18912), .A2(n18752), .B1(n18509), .B2(n18877), .ZN(
        n18490) );
  NOR2_X2 U21518 ( .A1(n18488), .A2(n18510), .ZN(n18879) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18879), .ZN(n18489) );
  OAI211_X1 U21520 ( .C1(n18531), .C2(n18755), .A(n18490), .B(n18489), .ZN(
        P3_U2870) );
  NOR2_X1 U21521 ( .A1(n18798), .A2(n21181), .ZN(n18808) );
  INV_X1 U21522 ( .A(n18808), .ZN(n18888) );
  NAND2_X1 U21523 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18866), .ZN(n18781) );
  INV_X1 U21524 ( .A(n18781), .ZN(n18884) );
  NOR2_X2 U21525 ( .A1(n18516), .A2(n21458), .ZN(n18883) );
  AOI22_X1 U21526 ( .A1(n18912), .A2(n18884), .B1(n18509), .B2(n18883), .ZN(
        n18493) );
  NOR2_X2 U21527 ( .A1(n18491), .A2(n18510), .ZN(n18885) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18885), .ZN(n18492) );
  OAI211_X1 U21529 ( .C1(n18531), .C2(n18888), .A(n18493), .B(n18492), .ZN(
        P3_U2871) );
  INV_X1 U21530 ( .A(n18912), .ZN(n18908) );
  NAND2_X1 U21531 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18866), .ZN(n18760) );
  NOR2_X1 U21532 ( .A1(n18798), .A2(n19478), .ZN(n18811) );
  NOR2_X2 U21533 ( .A1(n18516), .A2(n18494), .ZN(n18889) );
  AOI22_X1 U21534 ( .A1(n18855), .A2(n18811), .B1(n18509), .B2(n18889), .ZN(
        n18497) );
  NOR2_X2 U21535 ( .A1(n18495), .A2(n18510), .ZN(n18891) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18891), .ZN(n18496) );
  OAI211_X1 U21537 ( .C1(n18908), .C2(n18760), .A(n18497), .B(n18496), .ZN(
        P3_U2872) );
  INV_X1 U21538 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18498) );
  NOR2_X1 U21539 ( .A1(n18498), .A2(n18798), .ZN(n18846) );
  NAND2_X1 U21540 ( .A1(n18866), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18849) );
  INV_X1 U21541 ( .A(n18849), .ZN(n18896) );
  AND2_X1 U21542 ( .A1(n18831), .A2(BUF2_REG_5__SCAN_IN), .ZN(n18895) );
  AOI22_X1 U21543 ( .A1(n18855), .A2(n18896), .B1(n18509), .B2(n18895), .ZN(
        n18501) );
  NOR2_X2 U21544 ( .A1(n18499), .A2(n18510), .ZN(n18897) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18897), .ZN(n18500) );
  OAI211_X1 U21546 ( .C1(n18908), .C2(n18900), .A(n18501), .B(n18500), .ZN(
        P3_U2873) );
  NOR2_X1 U21547 ( .A1(n18502), .A2(n18798), .ZN(n18903) );
  INV_X1 U21548 ( .A(n18903), .ZN(n18853) );
  NAND2_X1 U21549 ( .A1(n18866), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18907) );
  INV_X1 U21550 ( .A(n18907), .ZN(n18850) );
  NOR2_X2 U21551 ( .A1(n18516), .A2(n18503), .ZN(n18901) );
  AOI22_X1 U21552 ( .A1(n18855), .A2(n18850), .B1(n18509), .B2(n18901), .ZN(
        n18506) );
  NOR2_X2 U21553 ( .A1(n18504), .A2(n18510), .ZN(n18904) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18904), .ZN(n18505) );
  OAI211_X1 U21555 ( .C1(n18908), .C2(n18853), .A(n18506), .B(n18505), .ZN(
        P3_U2874) );
  INV_X1 U21556 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18507) );
  NOR2_X1 U21557 ( .A1(n18507), .A2(n18798), .ZN(n18911) );
  INV_X1 U21558 ( .A(n18911), .ZN(n18795) );
  NAND2_X1 U21559 ( .A1(n18866), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18919) );
  INV_X1 U21560 ( .A(n18919), .ZN(n18790) );
  NOR2_X2 U21561 ( .A1(n18508), .A2(n18516), .ZN(n18910) );
  AOI22_X1 U21562 ( .A1(n18912), .A2(n18790), .B1(n18509), .B2(n18910), .ZN(
        n18514) );
  NOR2_X2 U21563 ( .A1(n18511), .A2(n18510), .ZN(n18913) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18512), .B1(
        n18577), .B2(n18913), .ZN(n18513) );
  OAI211_X1 U21565 ( .C1(n18531), .C2(n18795), .A(n18514), .B(n18513), .ZN(
        P3_U2875) );
  NAND2_X1 U21566 ( .A1(n18958), .A2(n18988), .ZN(n18799) );
  NOR2_X1 U21567 ( .A1(n18536), .A2(n18799), .ZN(n18532) );
  AOI22_X1 U21568 ( .A1(n18862), .A2(n18914), .B1(n18861), .B2(n18532), .ZN(
        n18518) );
  INV_X1 U21569 ( .A(n18536), .ZN(n18558) );
  NOR2_X1 U21570 ( .A1(n18516), .A2(n18515), .ZN(n18863) );
  NAND2_X1 U21571 ( .A1(n18958), .A2(n18863), .ZN(n18796) );
  INV_X1 U21572 ( .A(n18796), .ZN(n18603) );
  AOI22_X1 U21573 ( .A1(n18866), .A2(n18864), .B1(n18558), .B2(n18603), .ZN(
        n18533) );
  NOR2_X2 U21574 ( .A1(n18536), .A2(n18698), .ZN(n18598) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18533), .B1(
        n18867), .B2(n18598), .ZN(n18517) );
  OAI211_X1 U21576 ( .C1(n18531), .C2(n18870), .A(n18518), .B(n18517), .ZN(
        P3_U2876) );
  AOI22_X1 U21577 ( .A1(n18855), .A2(n18871), .B1(n18872), .B2(n18532), .ZN(
        n18520) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18533), .B1(
        n18873), .B2(n18598), .ZN(n18519) );
  OAI211_X1 U21579 ( .C1(n18551), .C2(n18876), .A(n18520), .B(n18519), .ZN(
        P3_U2877) );
  AOI22_X1 U21580 ( .A1(n18855), .A2(n18752), .B1(n18877), .B2(n18532), .ZN(
        n18522) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18533), .B1(
        n18879), .B2(n18598), .ZN(n18521) );
  OAI211_X1 U21582 ( .C1(n18551), .C2(n18755), .A(n18522), .B(n18521), .ZN(
        P3_U2878) );
  AOI22_X1 U21583 ( .A1(n18914), .A2(n18808), .B1(n18883), .B2(n18532), .ZN(
        n18524) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18533), .B1(
        n18885), .B2(n18598), .ZN(n18523) );
  OAI211_X1 U21585 ( .C1(n18531), .C2(n18781), .A(n18524), .B(n18523), .ZN(
        P3_U2879) );
  INV_X1 U21586 ( .A(n18811), .ZN(n18894) );
  INV_X1 U21587 ( .A(n18760), .ZN(n18890) );
  AOI22_X1 U21588 ( .A1(n18855), .A2(n18890), .B1(n18889), .B2(n18532), .ZN(
        n18526) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18533), .B1(
        n18891), .B2(n18598), .ZN(n18525) );
  OAI211_X1 U21590 ( .C1(n18551), .C2(n18894), .A(n18526), .B(n18525), .ZN(
        P3_U2880) );
  AOI22_X1 U21591 ( .A1(n18855), .A2(n18846), .B1(n18895), .B2(n18532), .ZN(
        n18528) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18533), .B1(
        n18897), .B2(n18598), .ZN(n18527) );
  OAI211_X1 U21593 ( .C1(n18551), .C2(n18849), .A(n18528), .B(n18527), .ZN(
        P3_U2881) );
  AOI22_X1 U21594 ( .A1(n18914), .A2(n18850), .B1(n18901), .B2(n18532), .ZN(
        n18530) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18533), .B1(
        n18904), .B2(n18598), .ZN(n18529) );
  OAI211_X1 U21596 ( .C1(n18531), .C2(n18853), .A(n18530), .B(n18529), .ZN(
        P3_U2882) );
  AOI22_X1 U21597 ( .A1(n18855), .A2(n18790), .B1(n18910), .B2(n18532), .ZN(
        n18535) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18533), .B1(
        n18913), .B2(n18598), .ZN(n18534) );
  OAI211_X1 U21599 ( .C1(n18551), .C2(n18795), .A(n18535), .B(n18534), .ZN(
        P3_U2883) );
  INV_X1 U21600 ( .A(n18577), .ZN(n18572) );
  NOR2_X1 U21601 ( .A1(n18958), .A2(n18536), .ZN(n18605) );
  NAND2_X1 U21602 ( .A1(n18956), .A2(n18605), .ZN(n18618) );
  NOR2_X1 U21603 ( .A1(n18598), .A2(n18621), .ZN(n18581) );
  NOR2_X1 U21604 ( .A1(n18982), .A2(n18581), .ZN(n18554) );
  AOI22_X1 U21605 ( .A1(n18914), .A2(n18826), .B1(n18861), .B2(n18554), .ZN(
        n18540) );
  OAI21_X1 U21606 ( .B1(n18537), .B2(n18828), .A(n18581), .ZN(n18538) );
  OAI211_X1 U21607 ( .C1(n18621), .C2(n19091), .A(n18831), .B(n18538), .ZN(
        n18555) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18555), .B1(
        n18867), .B2(n18621), .ZN(n18539) );
  OAI211_X1 U21609 ( .C1(n18834), .C2(n18572), .A(n18540), .B(n18539), .ZN(
        P3_U2884) );
  AOI22_X1 U21610 ( .A1(n18914), .A2(n18871), .B1(n18872), .B2(n18554), .ZN(
        n18542) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18555), .B1(
        n18873), .B2(n18621), .ZN(n18541) );
  OAI211_X1 U21612 ( .C1(n18572), .C2(n18876), .A(n18542), .B(n18541), .ZN(
        P3_U2885) );
  INV_X1 U21613 ( .A(n18752), .ZN(n18882) );
  INV_X1 U21614 ( .A(n18755), .ZN(n18878) );
  AOI22_X1 U21615 ( .A1(n18577), .A2(n18878), .B1(n18877), .B2(n18554), .ZN(
        n18544) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18555), .B1(
        n18879), .B2(n18621), .ZN(n18543) );
  OAI211_X1 U21617 ( .C1(n18551), .C2(n18882), .A(n18544), .B(n18543), .ZN(
        P3_U2886) );
  AOI22_X1 U21618 ( .A1(n18914), .A2(n18884), .B1(n18883), .B2(n18554), .ZN(
        n18546) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18555), .B1(
        n18885), .B2(n18621), .ZN(n18545) );
  OAI211_X1 U21620 ( .C1(n18572), .C2(n18888), .A(n18546), .B(n18545), .ZN(
        P3_U2887) );
  AOI22_X1 U21621 ( .A1(n18577), .A2(n18811), .B1(n18889), .B2(n18554), .ZN(
        n18548) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18555), .B1(
        n18891), .B2(n18621), .ZN(n18547) );
  OAI211_X1 U21623 ( .C1(n18551), .C2(n18760), .A(n18548), .B(n18547), .ZN(
        P3_U2888) );
  AOI22_X1 U21624 ( .A1(n18577), .A2(n18896), .B1(n18895), .B2(n18554), .ZN(
        n18550) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18555), .B1(
        n18897), .B2(n18621), .ZN(n18549) );
  OAI211_X1 U21626 ( .C1(n18551), .C2(n18900), .A(n18550), .B(n18549), .ZN(
        P3_U2889) );
  AOI22_X1 U21627 ( .A1(n18914), .A2(n18903), .B1(n18901), .B2(n18554), .ZN(
        n18553) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18555), .B1(
        n18904), .B2(n18621), .ZN(n18552) );
  OAI211_X1 U21629 ( .C1(n18572), .C2(n18907), .A(n18553), .B(n18552), .ZN(
        P3_U2890) );
  AOI22_X1 U21630 ( .A1(n18914), .A2(n18790), .B1(n18910), .B2(n18554), .ZN(
        n18557) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18555), .B1(
        n18913), .B2(n18621), .ZN(n18556) );
  OAI211_X1 U21632 ( .C1(n18572), .C2(n18795), .A(n18557), .B(n18556), .ZN(
        P3_U2891) );
  OAI211_X1 U21633 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18652), .A(
        n18558), .B(n18863), .ZN(n18573) );
  INV_X1 U21634 ( .A(n18573), .ZN(n18580) );
  AND2_X1 U21635 ( .A1(n18988), .A2(n18605), .ZN(n18576) );
  AOI22_X1 U21636 ( .A1(n18577), .A2(n18826), .B1(n18861), .B2(n18576), .ZN(
        n18560) );
  NAND2_X1 U21637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18605), .ZN(
        n18648) );
  INV_X1 U21638 ( .A(n18648), .ZN(n18633) );
  AOI22_X1 U21639 ( .A1(n18862), .A2(n18598), .B1(n18867), .B2(n18633), .ZN(
        n18559) );
  OAI211_X1 U21640 ( .C1(n18580), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        P3_U2892) );
  INV_X1 U21641 ( .A(n18598), .ZN(n18593) );
  AOI22_X1 U21642 ( .A1(n18577), .A2(n18871), .B1(n18872), .B2(n18576), .ZN(
        n18563) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18573), .B1(
        n18873), .B2(n18633), .ZN(n18562) );
  OAI211_X1 U21644 ( .C1(n18876), .C2(n18593), .A(n18563), .B(n18562), .ZN(
        P3_U2893) );
  AOI22_X1 U21645 ( .A1(n18577), .A2(n18752), .B1(n18877), .B2(n18576), .ZN(
        n18565) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18573), .B1(
        n18879), .B2(n18633), .ZN(n18564) );
  OAI211_X1 U21647 ( .C1(n18755), .C2(n18593), .A(n18565), .B(n18564), .ZN(
        P3_U2894) );
  AOI22_X1 U21648 ( .A1(n18808), .A2(n18598), .B1(n18883), .B2(n18576), .ZN(
        n18567) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18573), .B1(
        n18885), .B2(n18633), .ZN(n18566) );
  OAI211_X1 U21650 ( .C1(n18572), .C2(n18781), .A(n18567), .B(n18566), .ZN(
        P3_U2895) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18573), .B1(
        n18889), .B2(n18576), .ZN(n18569) );
  AOI22_X1 U21652 ( .A1(n18577), .A2(n18890), .B1(n18891), .B2(n18633), .ZN(
        n18568) );
  OAI211_X1 U21653 ( .C1(n18894), .C2(n18593), .A(n18569), .B(n18568), .ZN(
        P3_U2896) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18573), .B1(
        n18895), .B2(n18576), .ZN(n18571) );
  AOI22_X1 U21655 ( .A1(n18897), .A2(n18633), .B1(n18896), .B2(n18598), .ZN(
        n18570) );
  OAI211_X1 U21656 ( .C1(n18572), .C2(n18900), .A(n18571), .B(n18570), .ZN(
        P3_U2897) );
  AOI22_X1 U21657 ( .A1(n18577), .A2(n18903), .B1(n18901), .B2(n18576), .ZN(
        n18575) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18573), .B1(
        n18904), .B2(n18633), .ZN(n18574) );
  OAI211_X1 U21659 ( .C1(n18907), .C2(n18593), .A(n18575), .B(n18574), .ZN(
        P3_U2898) );
  INV_X1 U21660 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21374) );
  AOI22_X1 U21661 ( .A1(n18911), .A2(n18598), .B1(n18910), .B2(n18576), .ZN(
        n18579) );
  AOI22_X1 U21662 ( .A1(n18577), .A2(n18790), .B1(n18913), .B2(n18633), .ZN(
        n18578) );
  OAI211_X1 U21663 ( .C1(n18580), .C2(n21374), .A(n18579), .B(n18578), .ZN(
        P3_U2899) );
  NOR2_X2 U21664 ( .A1(n18959), .A2(n18650), .ZN(n18665) );
  NOR2_X1 U21665 ( .A1(n18633), .A2(n18665), .ZN(n18627) );
  NOR2_X1 U21666 ( .A1(n18982), .A2(n18627), .ZN(n18599) );
  AOI22_X1 U21667 ( .A1(n18826), .A2(n18598), .B1(n18861), .B2(n18599), .ZN(
        n18584) );
  OAI21_X1 U21668 ( .B1(n18581), .B2(n18828), .A(n18627), .ZN(n18582) );
  OAI211_X1 U21669 ( .C1(n18665), .C2(n19091), .A(n18831), .B(n18582), .ZN(
        n18600) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18600), .B1(
        n18867), .B2(n18665), .ZN(n18583) );
  OAI211_X1 U21671 ( .C1(n18834), .C2(n18618), .A(n18584), .B(n18583), .ZN(
        P3_U2900) );
  AOI22_X1 U21672 ( .A1(n18872), .A2(n18599), .B1(n18871), .B2(n18598), .ZN(
        n18586) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18600), .B1(
        n18873), .B2(n18665), .ZN(n18585) );
  OAI211_X1 U21674 ( .C1(n18876), .C2(n18618), .A(n18586), .B(n18585), .ZN(
        P3_U2901) );
  AOI22_X1 U21675 ( .A1(n18752), .A2(n18598), .B1(n18877), .B2(n18599), .ZN(
        n18588) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18600), .B1(
        n18879), .B2(n18665), .ZN(n18587) );
  OAI211_X1 U21677 ( .C1(n18755), .C2(n18618), .A(n18588), .B(n18587), .ZN(
        P3_U2902) );
  AOI22_X1 U21678 ( .A1(n18808), .A2(n18621), .B1(n18883), .B2(n18599), .ZN(
        n18590) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18600), .B1(
        n18885), .B2(n18665), .ZN(n18589) );
  OAI211_X1 U21680 ( .C1(n18781), .C2(n18593), .A(n18590), .B(n18589), .ZN(
        P3_U2903) );
  AOI22_X1 U21681 ( .A1(n18811), .A2(n18621), .B1(n18889), .B2(n18599), .ZN(
        n18592) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18600), .B1(
        n18891), .B2(n18665), .ZN(n18591) );
  OAI211_X1 U21683 ( .C1(n18760), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2904) );
  AOI22_X1 U21684 ( .A1(n18846), .A2(n18598), .B1(n18895), .B2(n18599), .ZN(
        n18595) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18600), .B1(
        n18897), .B2(n18665), .ZN(n18594) );
  OAI211_X1 U21686 ( .C1(n18849), .C2(n18618), .A(n18595), .B(n18594), .ZN(
        P3_U2905) );
  AOI22_X1 U21687 ( .A1(n18903), .A2(n18598), .B1(n18901), .B2(n18599), .ZN(
        n18597) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18600), .B1(
        n18904), .B2(n18665), .ZN(n18596) );
  OAI211_X1 U21689 ( .C1(n18907), .C2(n18618), .A(n18597), .B(n18596), .ZN(
        P3_U2906) );
  AOI22_X1 U21690 ( .A1(n18910), .A2(n18599), .B1(n18790), .B2(n18598), .ZN(
        n18602) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18600), .B1(
        n18913), .B2(n18665), .ZN(n18601) );
  OAI211_X1 U21692 ( .C1(n18795), .C2(n18618), .A(n18602), .B(n18601), .ZN(
        P3_U2907) );
  NOR2_X1 U21693 ( .A1(n18650), .A2(n18799), .ZN(n18622) );
  AOI22_X1 U21694 ( .A1(n18862), .A2(n18633), .B1(n18861), .B2(n18622), .ZN(
        n18607) );
  AOI22_X1 U21695 ( .A1(n18866), .A2(n18605), .B1(n18604), .B2(n18603), .ZN(
        n18623) );
  NOR2_X2 U21696 ( .A1(n18650), .A2(n18698), .ZN(n18690) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18623), .B1(
        n18867), .B2(n18690), .ZN(n18606) );
  OAI211_X1 U21698 ( .C1(n18870), .C2(n18618), .A(n18607), .B(n18606), .ZN(
        P3_U2908) );
  AOI22_X1 U21699 ( .A1(n18835), .A2(n18633), .B1(n18872), .B2(n18622), .ZN(
        n18609) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18623), .B1(
        n18873), .B2(n18690), .ZN(n18608) );
  OAI211_X1 U21701 ( .C1(n18838), .C2(n18618), .A(n18609), .B(n18608), .ZN(
        P3_U2909) );
  AOI22_X1 U21702 ( .A1(n18878), .A2(n18633), .B1(n18877), .B2(n18622), .ZN(
        n18611) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18623), .B1(
        n18879), .B2(n18690), .ZN(n18610) );
  OAI211_X1 U21704 ( .C1(n18882), .C2(n18618), .A(n18611), .B(n18610), .ZN(
        P3_U2910) );
  AOI22_X1 U21705 ( .A1(n18884), .A2(n18621), .B1(n18883), .B2(n18622), .ZN(
        n18613) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18623), .B1(
        n18885), .B2(n18690), .ZN(n18612) );
  OAI211_X1 U21707 ( .C1(n18888), .C2(n18648), .A(n18613), .B(n18612), .ZN(
        P3_U2911) );
  AOI22_X1 U21708 ( .A1(n18890), .A2(n18621), .B1(n18889), .B2(n18622), .ZN(
        n18615) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18623), .B1(
        n18891), .B2(n18690), .ZN(n18614) );
  OAI211_X1 U21710 ( .C1(n18894), .C2(n18648), .A(n18615), .B(n18614), .ZN(
        P3_U2912) );
  AOI22_X1 U21711 ( .A1(n18896), .A2(n18633), .B1(n18895), .B2(n18622), .ZN(
        n18617) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18623), .B1(
        n18897), .B2(n18690), .ZN(n18616) );
  OAI211_X1 U21713 ( .C1(n18900), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2913) );
  AOI22_X1 U21714 ( .A1(n18903), .A2(n18621), .B1(n18901), .B2(n18622), .ZN(
        n18620) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18623), .B1(
        n18904), .B2(n18690), .ZN(n18619) );
  OAI211_X1 U21716 ( .C1(n18907), .C2(n18648), .A(n18620), .B(n18619), .ZN(
        P3_U2914) );
  AOI22_X1 U21717 ( .A1(n18910), .A2(n18622), .B1(n18790), .B2(n18621), .ZN(
        n18625) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18623), .B1(
        n18913), .B2(n18690), .ZN(n18624) );
  OAI211_X1 U21719 ( .C1(n18795), .C2(n18648), .A(n18625), .B(n18624), .ZN(
        P3_U2915) );
  INV_X1 U21720 ( .A(n18665), .ZN(n18672) );
  NOR2_X1 U21721 ( .A1(n18626), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18697) );
  NAND2_X1 U21722 ( .A1(n18956), .A2(n18697), .ZN(n18695) );
  NOR2_X1 U21723 ( .A1(n18690), .A2(n18720), .ZN(n18673) );
  NOR2_X1 U21724 ( .A1(n18982), .A2(n18673), .ZN(n18644) );
  AOI22_X1 U21725 ( .A1(n18826), .A2(n18633), .B1(n18861), .B2(n18644), .ZN(
        n18630) );
  OAI21_X1 U21726 ( .B1(n18627), .B2(n18828), .A(n18673), .ZN(n18628) );
  OAI211_X1 U21727 ( .C1(n18720), .C2(n19091), .A(n18831), .B(n18628), .ZN(
        n18645) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18645), .B1(
        n18867), .B2(n18720), .ZN(n18629) );
  OAI211_X1 U21729 ( .C1(n18834), .C2(n18672), .A(n18630), .B(n18629), .ZN(
        P3_U2916) );
  AOI22_X1 U21730 ( .A1(n18872), .A2(n18644), .B1(n18871), .B2(n18633), .ZN(
        n18632) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18645), .B1(
        n18873), .B2(n18720), .ZN(n18631) );
  OAI211_X1 U21732 ( .C1(n18876), .C2(n18672), .A(n18632), .B(n18631), .ZN(
        P3_U2917) );
  AOI22_X1 U21733 ( .A1(n18752), .A2(n18633), .B1(n18877), .B2(n18644), .ZN(
        n18635) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18645), .B1(
        n18879), .B2(n18720), .ZN(n18634) );
  OAI211_X1 U21735 ( .C1(n18755), .C2(n18672), .A(n18635), .B(n18634), .ZN(
        P3_U2918) );
  AOI22_X1 U21736 ( .A1(n18808), .A2(n18665), .B1(n18883), .B2(n18644), .ZN(
        n18637) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18645), .B1(
        n18885), .B2(n18720), .ZN(n18636) );
  OAI211_X1 U21738 ( .C1(n18781), .C2(n18648), .A(n18637), .B(n18636), .ZN(
        P3_U2919) );
  AOI22_X1 U21739 ( .A1(n18811), .A2(n18665), .B1(n18889), .B2(n18644), .ZN(
        n18639) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18645), .B1(
        n18891), .B2(n18720), .ZN(n18638) );
  OAI211_X1 U21741 ( .C1(n18760), .C2(n18648), .A(n18639), .B(n18638), .ZN(
        P3_U2920) );
  AOI22_X1 U21742 ( .A1(n18896), .A2(n18665), .B1(n18895), .B2(n18644), .ZN(
        n18641) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18645), .B1(
        n18897), .B2(n18720), .ZN(n18640) );
  OAI211_X1 U21744 ( .C1(n18900), .C2(n18648), .A(n18641), .B(n18640), .ZN(
        P3_U2921) );
  AOI22_X1 U21745 ( .A1(n18850), .A2(n18665), .B1(n18901), .B2(n18644), .ZN(
        n18643) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18645), .B1(
        n18904), .B2(n18720), .ZN(n18642) );
  OAI211_X1 U21747 ( .C1(n18853), .C2(n18648), .A(n18643), .B(n18642), .ZN(
        P3_U2922) );
  AOI22_X1 U21748 ( .A1(n18911), .A2(n18665), .B1(n18910), .B2(n18644), .ZN(
        n18647) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18645), .B1(
        n18913), .B2(n18720), .ZN(n18646) );
  OAI211_X1 U21750 ( .C1(n18919), .C2(n18648), .A(n18647), .B(n18646), .ZN(
        P3_U2923) );
  INV_X1 U21751 ( .A(n18690), .ZN(n18689) );
  INV_X1 U21752 ( .A(n18697), .ZN(n18649) );
  NOR2_X1 U21753 ( .A1(n18982), .A2(n18649), .ZN(n18668) );
  AOI22_X1 U21754 ( .A1(n18826), .A2(n18665), .B1(n18861), .B2(n18668), .ZN(
        n18654) );
  NOR2_X2 U21755 ( .A1(n18956), .A2(n18649), .ZN(n18739) );
  INV_X1 U21756 ( .A(n18739), .ZN(n18746) );
  OAI21_X1 U21757 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18650), .A(n18746), 
        .ZN(n18651) );
  OAI211_X1 U21758 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18652), .A(
        n18831), .B(n18651), .ZN(n18669) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18669), .B1(
        n18867), .B2(n18739), .ZN(n18653) );
  OAI211_X1 U21760 ( .C1(n18834), .C2(n18689), .A(n18654), .B(n18653), .ZN(
        P3_U2924) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18669), .B1(
        n18872), .B2(n18668), .ZN(n18656) );
  AOI22_X1 U21762 ( .A1(n18835), .A2(n18690), .B1(n18873), .B2(n18739), .ZN(
        n18655) );
  OAI211_X1 U21763 ( .C1(n18838), .C2(n18672), .A(n18656), .B(n18655), .ZN(
        P3_U2925) );
  AOI22_X1 U21764 ( .A1(n18752), .A2(n18665), .B1(n18877), .B2(n18668), .ZN(
        n18658) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18669), .B1(
        n18879), .B2(n18739), .ZN(n18657) );
  OAI211_X1 U21766 ( .C1(n18755), .C2(n18689), .A(n18658), .B(n18657), .ZN(
        P3_U2926) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18669), .B1(
        n18883), .B2(n18668), .ZN(n18660) );
  AOI22_X1 U21768 ( .A1(n18808), .A2(n18690), .B1(n18885), .B2(n18739), .ZN(
        n18659) );
  OAI211_X1 U21769 ( .C1(n18781), .C2(n18672), .A(n18660), .B(n18659), .ZN(
        P3_U2927) );
  AOI22_X1 U21770 ( .A1(n18890), .A2(n18665), .B1(n18889), .B2(n18668), .ZN(
        n18662) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18669), .B1(
        n18891), .B2(n18739), .ZN(n18661) );
  OAI211_X1 U21772 ( .C1(n18894), .C2(n18689), .A(n18662), .B(n18661), .ZN(
        P3_U2928) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18669), .B1(
        n18895), .B2(n18668), .ZN(n18664) );
  AOI22_X1 U21774 ( .A1(n18846), .A2(n18665), .B1(n18897), .B2(n18739), .ZN(
        n18663) );
  OAI211_X1 U21775 ( .C1(n18849), .C2(n18689), .A(n18664), .B(n18663), .ZN(
        P3_U2929) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18669), .B1(
        n18901), .B2(n18668), .ZN(n18667) );
  AOI22_X1 U21777 ( .A1(n18903), .A2(n18665), .B1(n18904), .B2(n18739), .ZN(
        n18666) );
  OAI211_X1 U21778 ( .C1(n18907), .C2(n18689), .A(n18667), .B(n18666), .ZN(
        P3_U2930) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18669), .B1(
        n18910), .B2(n18668), .ZN(n18671) );
  AOI22_X1 U21780 ( .A1(n18911), .A2(n18690), .B1(n18913), .B2(n18739), .ZN(
        n18670) );
  OAI211_X1 U21781 ( .C1(n18919), .C2(n18672), .A(n18671), .B(n18670), .ZN(
        P3_U2931) );
  NOR2_X2 U21782 ( .A1(n18959), .A2(n18699), .ZN(n18766) );
  NOR2_X1 U21783 ( .A1(n18739), .A2(n18766), .ZN(n18725) );
  NOR2_X1 U21784 ( .A1(n18982), .A2(n18725), .ZN(n18691) );
  AOI22_X1 U21785 ( .A1(n18826), .A2(n18690), .B1(n18861), .B2(n18691), .ZN(
        n18676) );
  OAI21_X1 U21786 ( .B1(n18673), .B2(n18828), .A(n18725), .ZN(n18674) );
  OAI211_X1 U21787 ( .C1(n18766), .C2(n19091), .A(n18831), .B(n18674), .ZN(
        n18692) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18692), .B1(
        n18867), .B2(n18766), .ZN(n18675) );
  OAI211_X1 U21789 ( .C1(n18834), .C2(n18695), .A(n18676), .B(n18675), .ZN(
        P3_U2932) );
  AOI22_X1 U21790 ( .A1(n18835), .A2(n18720), .B1(n18872), .B2(n18691), .ZN(
        n18678) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18692), .B1(
        n18873), .B2(n18766), .ZN(n18677) );
  OAI211_X1 U21792 ( .C1(n18838), .C2(n18689), .A(n18678), .B(n18677), .ZN(
        P3_U2933) );
  AOI22_X1 U21793 ( .A1(n18878), .A2(n18720), .B1(n18877), .B2(n18691), .ZN(
        n18680) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18692), .B1(
        n18879), .B2(n18766), .ZN(n18679) );
  OAI211_X1 U21795 ( .C1(n18882), .C2(n18689), .A(n18680), .B(n18679), .ZN(
        P3_U2934) );
  AOI22_X1 U21796 ( .A1(n18808), .A2(n18720), .B1(n18883), .B2(n18691), .ZN(
        n18682) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18692), .B1(
        n18885), .B2(n18766), .ZN(n18681) );
  OAI211_X1 U21798 ( .C1(n18781), .C2(n18689), .A(n18682), .B(n18681), .ZN(
        P3_U2935) );
  AOI22_X1 U21799 ( .A1(n18890), .A2(n18690), .B1(n18889), .B2(n18691), .ZN(
        n18684) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18692), .B1(
        n18891), .B2(n18766), .ZN(n18683) );
  OAI211_X1 U21801 ( .C1(n18894), .C2(n18695), .A(n18684), .B(n18683), .ZN(
        P3_U2936) );
  AOI22_X1 U21802 ( .A1(n18896), .A2(n18720), .B1(n18895), .B2(n18691), .ZN(
        n18686) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18692), .B1(
        n18897), .B2(n18766), .ZN(n18685) );
  OAI211_X1 U21804 ( .C1(n18900), .C2(n18689), .A(n18686), .B(n18685), .ZN(
        P3_U2937) );
  AOI22_X1 U21805 ( .A1(n18850), .A2(n18720), .B1(n18901), .B2(n18691), .ZN(
        n18688) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18692), .B1(
        n18904), .B2(n18766), .ZN(n18687) );
  OAI211_X1 U21807 ( .C1(n18853), .C2(n18689), .A(n18688), .B(n18687), .ZN(
        P3_U2938) );
  AOI22_X1 U21808 ( .A1(n18910), .A2(n18691), .B1(n18790), .B2(n18690), .ZN(
        n18694) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18692), .B1(
        n18913), .B2(n18766), .ZN(n18693) );
  OAI211_X1 U21810 ( .C1(n18795), .C2(n18695), .A(n18694), .B(n18693), .ZN(
        P3_U2939) );
  NOR2_X1 U21811 ( .A1(n18699), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18696) );
  AOI22_X1 U21812 ( .A1(n18866), .A2(n18697), .B1(n18863), .B2(n18696), .ZN(
        n18711) );
  INV_X1 U21813 ( .A(n18711), .ZN(n18723) );
  NOR2_X1 U21814 ( .A1(n18699), .A2(n18799), .ZN(n18719) );
  AOI22_X1 U21815 ( .A1(n18826), .A2(n18720), .B1(n18861), .B2(n18719), .ZN(
        n18701) );
  NOR2_X2 U21816 ( .A1(n18699), .A2(n18698), .ZN(n18789) );
  AOI22_X1 U21817 ( .A1(n18862), .A2(n18739), .B1(n18867), .B2(n18789), .ZN(
        n18700) );
  OAI211_X1 U21818 ( .C1(n18702), .C2(n18723), .A(n18701), .B(n18700), .ZN(
        P3_U2940) );
  AOI22_X1 U21819 ( .A1(n18872), .A2(n18719), .B1(n18871), .B2(n18720), .ZN(
        n18704) );
  AOI22_X1 U21820 ( .A1(n18835), .A2(n18739), .B1(n18873), .B2(n18789), .ZN(
        n18703) );
  OAI211_X1 U21821 ( .C1(n18705), .C2(n18723), .A(n18704), .B(n18703), .ZN(
        P3_U2941) );
  AOI22_X1 U21822 ( .A1(n18752), .A2(n18720), .B1(n18877), .B2(n18719), .ZN(
        n18707) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18711), .B1(
        n18879), .B2(n18789), .ZN(n18706) );
  OAI211_X1 U21824 ( .C1(n18755), .C2(n18746), .A(n18707), .B(n18706), .ZN(
        P3_U2942) );
  AOI22_X1 U21825 ( .A1(n18808), .A2(n18739), .B1(n18883), .B2(n18719), .ZN(
        n18709) );
  AOI22_X1 U21826 ( .A1(n18885), .A2(n18789), .B1(n18884), .B2(n18720), .ZN(
        n18708) );
  OAI211_X1 U21827 ( .C1(n18710), .C2(n18723), .A(n18709), .B(n18708), .ZN(
        P3_U2943) );
  AOI22_X1 U21828 ( .A1(n18890), .A2(n18720), .B1(n18889), .B2(n18719), .ZN(
        n18713) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18711), .B1(
        n18891), .B2(n18789), .ZN(n18712) );
  OAI211_X1 U21830 ( .C1(n18894), .C2(n18746), .A(n18713), .B(n18712), .ZN(
        P3_U2944) );
  AOI22_X1 U21831 ( .A1(n18896), .A2(n18739), .B1(n18895), .B2(n18719), .ZN(
        n18715) );
  AOI22_X1 U21832 ( .A1(n18846), .A2(n18720), .B1(n18897), .B2(n18789), .ZN(
        n18714) );
  OAI211_X1 U21833 ( .C1(n18716), .C2(n18723), .A(n18715), .B(n18714), .ZN(
        P3_U2945) );
  AOI22_X1 U21834 ( .A1(n18903), .A2(n18720), .B1(n18901), .B2(n18719), .ZN(
        n18718) );
  AOI22_X1 U21835 ( .A1(n18904), .A2(n18789), .B1(n18850), .B2(n18739), .ZN(
        n18717) );
  OAI211_X1 U21836 ( .C1(n21319), .C2(n18723), .A(n18718), .B(n18717), .ZN(
        P3_U2946) );
  AOI22_X1 U21837 ( .A1(n18911), .A2(n18739), .B1(n18910), .B2(n18719), .ZN(
        n18722) );
  AOI22_X1 U21838 ( .A1(n18913), .A2(n18789), .B1(n18790), .B2(n18720), .ZN(
        n18721) );
  OAI211_X1 U21839 ( .C1(n18724), .C2(n18723), .A(n18722), .B(n18721), .ZN(
        P3_U2947) );
  INV_X1 U21840 ( .A(n18766), .ZN(n18765) );
  NAND2_X1 U21841 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18747), .ZN(
        n18797) );
  NOR2_X2 U21842 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18797), .ZN(
        n18817) );
  NOR2_X1 U21843 ( .A1(n18789), .A2(n18817), .ZN(n18771) );
  NOR2_X1 U21844 ( .A1(n18982), .A2(n18771), .ZN(n18742) );
  AOI22_X1 U21845 ( .A1(n18826), .A2(n18739), .B1(n18861), .B2(n18742), .ZN(
        n18728) );
  OAI21_X1 U21846 ( .B1(n18725), .B2(n18828), .A(n18771), .ZN(n18726) );
  OAI211_X1 U21847 ( .C1(n18817), .C2(n19091), .A(n18831), .B(n18726), .ZN(
        n18743) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18743), .B1(
        n18867), .B2(n18817), .ZN(n18727) );
  OAI211_X1 U21849 ( .C1(n18834), .C2(n18765), .A(n18728), .B(n18727), .ZN(
        P3_U2948) );
  AOI22_X1 U21850 ( .A1(n18872), .A2(n18742), .B1(n18871), .B2(n18739), .ZN(
        n18730) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18743), .B1(
        n18873), .B2(n18817), .ZN(n18729) );
  OAI211_X1 U21852 ( .C1(n18876), .C2(n18765), .A(n18730), .B(n18729), .ZN(
        P3_U2949) );
  AOI22_X1 U21853 ( .A1(n18752), .A2(n18739), .B1(n18877), .B2(n18742), .ZN(
        n18732) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18743), .B1(
        n18879), .B2(n18817), .ZN(n18731) );
  OAI211_X1 U21855 ( .C1(n18755), .C2(n18765), .A(n18732), .B(n18731), .ZN(
        P3_U2950) );
  AOI22_X1 U21856 ( .A1(n18884), .A2(n18739), .B1(n18883), .B2(n18742), .ZN(
        n18734) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18743), .B1(
        n18885), .B2(n18817), .ZN(n18733) );
  OAI211_X1 U21858 ( .C1(n18888), .C2(n18765), .A(n18734), .B(n18733), .ZN(
        P3_U2951) );
  AOI22_X1 U21859 ( .A1(n18811), .A2(n18766), .B1(n18889), .B2(n18742), .ZN(
        n18736) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18743), .B1(
        n18891), .B2(n18817), .ZN(n18735) );
  OAI211_X1 U21861 ( .C1(n18760), .C2(n18746), .A(n18736), .B(n18735), .ZN(
        P3_U2952) );
  AOI22_X1 U21862 ( .A1(n18896), .A2(n18766), .B1(n18895), .B2(n18742), .ZN(
        n18738) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18743), .B1(
        n18897), .B2(n18817), .ZN(n18737) );
  OAI211_X1 U21864 ( .C1(n18900), .C2(n18746), .A(n18738), .B(n18737), .ZN(
        P3_U2953) );
  AOI22_X1 U21865 ( .A1(n18903), .A2(n18739), .B1(n18901), .B2(n18742), .ZN(
        n18741) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18743), .B1(
        n18904), .B2(n18817), .ZN(n18740) );
  OAI211_X1 U21867 ( .C1(n18907), .C2(n18765), .A(n18741), .B(n18740), .ZN(
        P3_U2954) );
  AOI22_X1 U21868 ( .A1(n18911), .A2(n18766), .B1(n18910), .B2(n18742), .ZN(
        n18745) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18743), .B1(
        n18913), .B2(n18817), .ZN(n18744) );
  OAI211_X1 U21870 ( .C1(n18919), .C2(n18746), .A(n18745), .B(n18744), .ZN(
        P3_U2955) );
  NOR2_X1 U21871 ( .A1(n18982), .A2(n18797), .ZN(n18767) );
  AOI22_X1 U21872 ( .A1(n18862), .A2(n18789), .B1(n18861), .B2(n18767), .ZN(
        n18749) );
  OAI211_X1 U21873 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18866), .A(
        n18863), .B(n18747), .ZN(n18768) );
  NOR2_X2 U21874 ( .A1(n18956), .A2(n18797), .ZN(n18845) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18768), .B1(
        n18867), .B2(n18845), .ZN(n18748) );
  OAI211_X1 U21876 ( .C1(n18870), .C2(n18765), .A(n18749), .B(n18748), .ZN(
        P3_U2956) );
  INV_X1 U21877 ( .A(n18789), .ZN(n18786) );
  AOI22_X1 U21878 ( .A1(n18872), .A2(n18767), .B1(n18871), .B2(n18766), .ZN(
        n18751) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18768), .B1(
        n18873), .B2(n18845), .ZN(n18750) );
  OAI211_X1 U21880 ( .C1(n18876), .C2(n18786), .A(n18751), .B(n18750), .ZN(
        P3_U2957) );
  AOI22_X1 U21881 ( .A1(n18752), .A2(n18766), .B1(n18877), .B2(n18767), .ZN(
        n18754) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18768), .B1(
        n18879), .B2(n18845), .ZN(n18753) );
  OAI211_X1 U21883 ( .C1(n18755), .C2(n18786), .A(n18754), .B(n18753), .ZN(
        P3_U2958) );
  AOI22_X1 U21884 ( .A1(n18884), .A2(n18766), .B1(n18883), .B2(n18767), .ZN(
        n18757) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18768), .B1(
        n18885), .B2(n18845), .ZN(n18756) );
  OAI211_X1 U21886 ( .C1(n18888), .C2(n18786), .A(n18757), .B(n18756), .ZN(
        P3_U2959) );
  AOI22_X1 U21887 ( .A1(n18811), .A2(n18789), .B1(n18889), .B2(n18767), .ZN(
        n18759) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18768), .B1(
        n18891), .B2(n18845), .ZN(n18758) );
  OAI211_X1 U21889 ( .C1(n18760), .C2(n18765), .A(n18759), .B(n18758), .ZN(
        P3_U2960) );
  AOI22_X1 U21890 ( .A1(n18846), .A2(n18766), .B1(n18895), .B2(n18767), .ZN(
        n18762) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18768), .B1(
        n18897), .B2(n18845), .ZN(n18761) );
  OAI211_X1 U21892 ( .C1(n18849), .C2(n18786), .A(n18762), .B(n18761), .ZN(
        P3_U2961) );
  AOI22_X1 U21893 ( .A1(n18850), .A2(n18789), .B1(n18901), .B2(n18767), .ZN(
        n18764) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18768), .B1(
        n18904), .B2(n18845), .ZN(n18763) );
  OAI211_X1 U21895 ( .C1(n18853), .C2(n18765), .A(n18764), .B(n18763), .ZN(
        P3_U2962) );
  AOI22_X1 U21896 ( .A1(n18910), .A2(n18767), .B1(n18790), .B2(n18766), .ZN(
        n18770) );
  AOI22_X1 U21897 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18768), .B1(
        n18913), .B2(n18845), .ZN(n18769) );
  OAI211_X1 U21898 ( .C1(n18795), .C2(n18786), .A(n18770), .B(n18769), .ZN(
        P3_U2963) );
  INV_X1 U21899 ( .A(n18817), .ZN(n18825) );
  NOR2_X2 U21900 ( .A1(n18959), .A2(n18800), .ZN(n18902) );
  NOR2_X1 U21901 ( .A1(n18845), .A2(n18902), .ZN(n18829) );
  NOR2_X1 U21902 ( .A1(n18982), .A2(n18829), .ZN(n18791) );
  AOI22_X1 U21903 ( .A1(n18826), .A2(n18789), .B1(n18861), .B2(n18791), .ZN(
        n18774) );
  OAI21_X1 U21904 ( .B1(n18771), .B2(n18828), .A(n18829), .ZN(n18772) );
  OAI211_X1 U21905 ( .C1(n18902), .C2(n19091), .A(n18831), .B(n18772), .ZN(
        n18792) );
  AOI22_X1 U21906 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18792), .B1(
        n18867), .B2(n18902), .ZN(n18773) );
  OAI211_X1 U21907 ( .C1(n18834), .C2(n18825), .A(n18774), .B(n18773), .ZN(
        P3_U2964) );
  AOI22_X1 U21908 ( .A1(n18835), .A2(n18817), .B1(n18872), .B2(n18791), .ZN(
        n18776) );
  AOI22_X1 U21909 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18792), .B1(
        n18873), .B2(n18902), .ZN(n18775) );
  OAI211_X1 U21910 ( .C1(n18838), .C2(n18786), .A(n18776), .B(n18775), .ZN(
        P3_U2965) );
  AOI22_X1 U21911 ( .A1(n18878), .A2(n18817), .B1(n18877), .B2(n18791), .ZN(
        n18778) );
  AOI22_X1 U21912 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18792), .B1(
        n18879), .B2(n18902), .ZN(n18777) );
  OAI211_X1 U21913 ( .C1(n18882), .C2(n18786), .A(n18778), .B(n18777), .ZN(
        P3_U2966) );
  AOI22_X1 U21914 ( .A1(n18808), .A2(n18817), .B1(n18883), .B2(n18791), .ZN(
        n18780) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18792), .B1(
        n18885), .B2(n18902), .ZN(n18779) );
  OAI211_X1 U21916 ( .C1(n18781), .C2(n18786), .A(n18780), .B(n18779), .ZN(
        P3_U2967) );
  AOI22_X1 U21917 ( .A1(n18890), .A2(n18789), .B1(n18889), .B2(n18791), .ZN(
        n18783) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18792), .B1(
        n18891), .B2(n18902), .ZN(n18782) );
  OAI211_X1 U21919 ( .C1(n18894), .C2(n18825), .A(n18783), .B(n18782), .ZN(
        P3_U2968) );
  AOI22_X1 U21920 ( .A1(n18896), .A2(n18817), .B1(n18895), .B2(n18791), .ZN(
        n18785) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18792), .B1(
        n18897), .B2(n18902), .ZN(n18784) );
  OAI211_X1 U21922 ( .C1(n18900), .C2(n18786), .A(n18785), .B(n18784), .ZN(
        P3_U2969) );
  AOI22_X1 U21923 ( .A1(n18903), .A2(n18789), .B1(n18901), .B2(n18791), .ZN(
        n18788) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18792), .B1(
        n18904), .B2(n18902), .ZN(n18787) );
  OAI211_X1 U21925 ( .C1(n18907), .C2(n18825), .A(n18788), .B(n18787), .ZN(
        P3_U2970) );
  AOI22_X1 U21926 ( .A1(n18910), .A2(n18791), .B1(n18790), .B2(n18789), .ZN(
        n18794) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18792), .B1(
        n18913), .B2(n18902), .ZN(n18793) );
  OAI211_X1 U21928 ( .C1(n18795), .C2(n18825), .A(n18794), .B(n18793), .ZN(
        P3_U2971) );
  OAI22_X1 U21929 ( .A1(n18798), .A2(n18797), .B1(n18800), .B2(n18796), .ZN(
        n18820) );
  NOR2_X1 U21930 ( .A1(n18800), .A2(n18799), .ZN(n18865) );
  AOI22_X1 U21931 ( .A1(n18862), .A2(n18845), .B1(n18861), .B2(n18865), .ZN(
        n18802) );
  AOI22_X1 U21932 ( .A1(n18912), .A2(n18867), .B1(n18826), .B2(n18817), .ZN(
        n18801) );
  OAI211_X1 U21933 ( .C1(n18803), .C2(n18820), .A(n18802), .B(n18801), .ZN(
        P3_U2972) );
  AOI22_X1 U21934 ( .A1(n18872), .A2(n18865), .B1(n18871), .B2(n18817), .ZN(
        n18805) );
  AOI22_X1 U21935 ( .A1(n18912), .A2(n18873), .B1(n18835), .B2(n18845), .ZN(
        n18804) );
  OAI211_X1 U21936 ( .C1(n21197), .C2(n18820), .A(n18805), .B(n18804), .ZN(
        P3_U2973) );
  AOI22_X1 U21937 ( .A1(n18878), .A2(n18845), .B1(n18877), .B2(n18865), .ZN(
        n18807) );
  INV_X1 U21938 ( .A(n18820), .ZN(n18822) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18822), .B1(
        n18912), .B2(n18879), .ZN(n18806) );
  OAI211_X1 U21940 ( .C1(n18882), .C2(n18825), .A(n18807), .B(n18806), .ZN(
        P3_U2974) );
  AOI22_X1 U21941 ( .A1(n18808), .A2(n18845), .B1(n18883), .B2(n18865), .ZN(
        n18810) );
  AOI22_X1 U21942 ( .A1(n18912), .A2(n18885), .B1(n18884), .B2(n18817), .ZN(
        n18809) );
  OAI211_X1 U21943 ( .C1(n21166), .C2(n18820), .A(n18810), .B(n18809), .ZN(
        P3_U2975) );
  AOI22_X1 U21944 ( .A1(n18890), .A2(n18817), .B1(n18889), .B2(n18865), .ZN(
        n18813) );
  AOI22_X1 U21945 ( .A1(n18912), .A2(n18891), .B1(n18811), .B2(n18845), .ZN(
        n18812) );
  OAI211_X1 U21946 ( .C1(n18814), .C2(n18820), .A(n18813), .B(n18812), .ZN(
        P3_U2976) );
  INV_X1 U21947 ( .A(n18845), .ZN(n18859) );
  AOI22_X1 U21948 ( .A1(n18846), .A2(n18817), .B1(n18895), .B2(n18865), .ZN(
        n18816) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18822), .B1(
        n18912), .B2(n18897), .ZN(n18815) );
  OAI211_X1 U21950 ( .C1(n18849), .C2(n18859), .A(n18816), .B(n18815), .ZN(
        P3_U2977) );
  AOI22_X1 U21951 ( .A1(n18850), .A2(n18845), .B1(n18901), .B2(n18865), .ZN(
        n18819) );
  AOI22_X1 U21952 ( .A1(n18912), .A2(n18904), .B1(n18903), .B2(n18817), .ZN(
        n18818) );
  OAI211_X1 U21953 ( .C1(n18821), .C2(n18820), .A(n18819), .B(n18818), .ZN(
        P3_U2978) );
  AOI22_X1 U21954 ( .A1(n18911), .A2(n18845), .B1(n18910), .B2(n18865), .ZN(
        n18824) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18822), .B1(
        n18912), .B2(n18913), .ZN(n18823) );
  OAI211_X1 U21956 ( .C1(n18919), .C2(n18825), .A(n18824), .B(n18823), .ZN(
        P3_U2979) );
  INV_X1 U21957 ( .A(n18902), .ZN(n18918) );
  NOR2_X1 U21958 ( .A1(n18982), .A2(n18827), .ZN(n18854) );
  AOI22_X1 U21959 ( .A1(n18826), .A2(n18845), .B1(n18861), .B2(n18854), .ZN(
        n18833) );
  OAI21_X1 U21960 ( .B1(n18829), .B2(n18828), .A(n18827), .ZN(n18830) );
  OAI211_X1 U21961 ( .C1(n18855), .C2(n19091), .A(n18831), .B(n18830), .ZN(
        n18856) );
  AOI22_X1 U21962 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18867), .ZN(n18832) );
  OAI211_X1 U21963 ( .C1(n18834), .C2(n18918), .A(n18833), .B(n18832), .ZN(
        P3_U2980) );
  AOI22_X1 U21964 ( .A1(n18835), .A2(n18902), .B1(n18872), .B2(n18854), .ZN(
        n18837) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18873), .ZN(n18836) );
  OAI211_X1 U21966 ( .C1(n18838), .C2(n18859), .A(n18837), .B(n18836), .ZN(
        P3_U2981) );
  AOI22_X1 U21967 ( .A1(n18878), .A2(n18902), .B1(n18877), .B2(n18854), .ZN(
        n18840) );
  AOI22_X1 U21968 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18879), .ZN(n18839) );
  OAI211_X1 U21969 ( .C1(n18882), .C2(n18859), .A(n18840), .B(n18839), .ZN(
        P3_U2982) );
  AOI22_X1 U21970 ( .A1(n18884), .A2(n18845), .B1(n18883), .B2(n18854), .ZN(
        n18842) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18885), .ZN(n18841) );
  OAI211_X1 U21972 ( .C1(n18888), .C2(n18918), .A(n18842), .B(n18841), .ZN(
        P3_U2983) );
  AOI22_X1 U21973 ( .A1(n18890), .A2(n18845), .B1(n18889), .B2(n18854), .ZN(
        n18844) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18891), .ZN(n18843) );
  OAI211_X1 U21975 ( .C1(n18894), .C2(n18918), .A(n18844), .B(n18843), .ZN(
        P3_U2984) );
  AOI22_X1 U21976 ( .A1(n18846), .A2(n18845), .B1(n18895), .B2(n18854), .ZN(
        n18848) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18897), .ZN(n18847) );
  OAI211_X1 U21978 ( .C1(n18849), .C2(n18918), .A(n18848), .B(n18847), .ZN(
        P3_U2985) );
  AOI22_X1 U21979 ( .A1(n18850), .A2(n18902), .B1(n18901), .B2(n18854), .ZN(
        n18852) );
  AOI22_X1 U21980 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18904), .ZN(n18851) );
  OAI211_X1 U21981 ( .C1(n18853), .C2(n18859), .A(n18852), .B(n18851), .ZN(
        P3_U2986) );
  AOI22_X1 U21982 ( .A1(n18911), .A2(n18902), .B1(n18910), .B2(n18854), .ZN(
        n18858) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18856), .B1(
        n18855), .B2(n18913), .ZN(n18857) );
  OAI211_X1 U21984 ( .C1(n18919), .C2(n18859), .A(n18858), .B(n18857), .ZN(
        P3_U2987) );
  NOR2_X1 U21985 ( .A1(n18982), .A2(n18860), .ZN(n18909) );
  AOI22_X1 U21986 ( .A1(n18862), .A2(n18912), .B1(n18861), .B2(n18909), .ZN(
        n18869) );
  AOI22_X1 U21987 ( .A1(n18866), .A2(n18865), .B1(n18864), .B2(n18863), .ZN(
        n18915) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18867), .ZN(n18868) );
  OAI211_X1 U21989 ( .C1(n18870), .C2(n18918), .A(n18869), .B(n18868), .ZN(
        P3_U2988) );
  AOI22_X1 U21990 ( .A1(n18872), .A2(n18909), .B1(n18871), .B2(n18902), .ZN(
        n18875) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18873), .ZN(n18874) );
  OAI211_X1 U21992 ( .C1(n18908), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        P3_U2989) );
  AOI22_X1 U21993 ( .A1(n18912), .A2(n18878), .B1(n18877), .B2(n18909), .ZN(
        n18881) );
  AOI22_X1 U21994 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18879), .ZN(n18880) );
  OAI211_X1 U21995 ( .C1(n18882), .C2(n18918), .A(n18881), .B(n18880), .ZN(
        P3_U2990) );
  AOI22_X1 U21996 ( .A1(n18884), .A2(n18902), .B1(n18883), .B2(n18909), .ZN(
        n18887) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18885), .ZN(n18886) );
  OAI211_X1 U21998 ( .C1(n18908), .C2(n18888), .A(n18887), .B(n18886), .ZN(
        P3_U2991) );
  AOI22_X1 U21999 ( .A1(n18890), .A2(n18902), .B1(n18889), .B2(n18909), .ZN(
        n18893) );
  AOI22_X1 U22000 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18891), .ZN(n18892) );
  OAI211_X1 U22001 ( .C1(n18908), .C2(n18894), .A(n18893), .B(n18892), .ZN(
        P3_U2992) );
  AOI22_X1 U22002 ( .A1(n18912), .A2(n18896), .B1(n18895), .B2(n18909), .ZN(
        n18899) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18897), .ZN(n18898) );
  OAI211_X1 U22004 ( .C1(n18900), .C2(n18918), .A(n18899), .B(n18898), .ZN(
        P3_U2993) );
  AOI22_X1 U22005 ( .A1(n18903), .A2(n18902), .B1(n18901), .B2(n18909), .ZN(
        n18906) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18904), .ZN(n18905) );
  OAI211_X1 U22007 ( .C1(n18908), .C2(n18907), .A(n18906), .B(n18905), .ZN(
        P3_U2994) );
  AOI22_X1 U22008 ( .A1(n18912), .A2(n18911), .B1(n18910), .B2(n18909), .ZN(
        n18917) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18913), .ZN(n18916) );
  OAI211_X1 U22010 ( .C1(n18919), .C2(n18918), .A(n18917), .B(n18916), .ZN(
        P3_U2995) );
  AOI21_X1 U22011 ( .B1(n18922), .B2(n18921), .A(n18920), .ZN(n19133) );
  NOR2_X1 U22012 ( .A1(n19132), .A2(n18923), .ZN(n19135) );
  AOI221_X1 U22013 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18924), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18924), .A(n19135), .ZN(n18925) );
  OAI211_X1 U22014 ( .C1(n18926), .C2(n18948), .A(n19133), .B(n18925), .ZN(
        n18972) );
  NOR2_X1 U22015 ( .A1(n18928), .A2(n18927), .ZN(n18937) );
  OAI21_X1 U22016 ( .B1(n18929), .B2(n19121), .A(n18937), .ZN(n18943) );
  AOI22_X1 U22017 ( .A1(n18947), .A2(n18930), .B1(n18944), .B2(n18943), .ZN(
        n18931) );
  NOR2_X1 U22018 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18931), .ZN(
        n19093) );
  AOI21_X1 U22019 ( .B1(n18934), .B2(n18933), .A(n18932), .ZN(n18941) );
  INV_X1 U22020 ( .A(n18935), .ZN(n18936) );
  OAI22_X1 U22021 ( .A1(n18937), .A2(n18944), .B1(n18941), .B2(n18936), .ZN(
        n18938) );
  AOI21_X1 U22022 ( .B1(n18939), .B2(n19108), .A(n18938), .ZN(n19094) );
  NAND2_X1 U22023 ( .A1(n18948), .A2(n19094), .ZN(n18940) );
  AOI22_X1 U22024 ( .A1(n18948), .A2(n19093), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18940), .ZN(n18970) );
  NOR3_X1 U22025 ( .A1(n18942), .A2(n18941), .A3(n19108), .ZN(n18946) );
  INV_X1 U22026 ( .A(n18943), .ZN(n18953) );
  AOI211_X1 U22027 ( .C1(n19114), .C2(n19108), .A(n18944), .B(n18953), .ZN(
        n18945) );
  AOI211_X1 U22028 ( .C1(n18947), .C2(n19101), .A(n18946), .B(n18945), .ZN(
        n19104) );
  AOI22_X1 U22029 ( .A1(n18961), .A2(n19108), .B1(n19104), .B2(n18948), .ZN(
        n18965) );
  INV_X1 U22030 ( .A(n18949), .ZN(n18951) );
  NOR2_X1 U22031 ( .A1(n18951), .A2(n18950), .ZN(n18955) );
  AOI22_X1 U22032 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18952), .B1(
        n18955), .B2(n19121), .ZN(n19116) );
  OAI22_X1 U22033 ( .A1(n18955), .A2(n18954), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18953), .ZN(n19112) );
  OR3_X1 U22034 ( .A1(n19116), .A2(n18958), .A3(n18956), .ZN(n18957) );
  AOI22_X1 U22035 ( .A1(n19116), .A2(n18958), .B1(n19112), .B2(n18957), .ZN(
        n18960) );
  OAI21_X1 U22036 ( .B1(n18961), .B2(n18960), .A(n18959), .ZN(n18964) );
  AND2_X1 U22037 ( .A1(n18965), .A2(n18964), .ZN(n18962) );
  OAI221_X1 U22038 ( .B1(n18965), .B2(n18964), .C1(n18963), .C2(n18962), .A(
        n18967), .ZN(n18969) );
  AOI21_X1 U22039 ( .B1(n18967), .B2(n18966), .A(n18965), .ZN(n18968) );
  AOI222_X1 U22040 ( .A1(n18970), .A2(n18969), .B1(n18970), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18969), .C2(n18968), .ZN(
        n18971) );
  NOR4_X1 U22041 ( .A1(n18974), .A2(n18973), .A3(n18972), .A4(n18971), .ZN(
        n18986) );
  AOI22_X1 U22042 ( .A1(n19143), .A2(n19152), .B1(n19115), .B2(n18975), .ZN(
        n18976) );
  INV_X1 U22043 ( .A(n18976), .ZN(n18981) );
  OAI211_X1 U22044 ( .C1(n18978), .C2(n18977), .A(n19149), .B(n18986), .ZN(
        n19090) );
  OAI21_X1 U22045 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19151), .A(n19090), 
        .ZN(n18987) );
  NOR2_X1 U22046 ( .A1(n18979), .A2(n18987), .ZN(n18980) );
  MUX2_X1 U22047 ( .A(n18981), .B(n18980), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18984) );
  NAND2_X1 U22048 ( .A1(n18990), .A2(n18982), .ZN(n18983) );
  OAI211_X1 U22049 ( .C1(n18986), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        P3_U2996) );
  NAND2_X1 U22050 ( .A1(n19143), .A2(n19152), .ZN(n18992) );
  NAND4_X1 U22051 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19143), .A4(n19142), .ZN(n18994) );
  INV_X1 U22052 ( .A(n18987), .ZN(n18989) );
  NAND3_X1 U22053 ( .A1(n18990), .A2(n18989), .A3(n18988), .ZN(n18991) );
  NAND4_X1 U22054 ( .A1(n18993), .A2(n18992), .A3(n18994), .A4(n18991), .ZN(
        P3_U2997) );
  AND4_X1 U22055 ( .A1(n19145), .A2(n18995), .A3(n18994), .A4(n19089), .ZN(
        P3_U2998) );
  AND2_X1 U22056 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18996), .ZN(
        P3_U2999) );
  AND2_X1 U22057 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18996), .ZN(
        P3_U3000) );
  AND2_X1 U22058 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18997), .ZN(
        P3_U3001) );
  AND2_X1 U22059 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18996), .ZN(
        P3_U3002) );
  AND2_X1 U22060 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18997), .ZN(
        P3_U3003) );
  AND2_X1 U22061 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18996), .ZN(
        P3_U3004) );
  AND2_X1 U22062 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18997), .ZN(
        P3_U3005) );
  AND2_X1 U22063 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18996), .ZN(
        P3_U3006) );
  AND2_X1 U22064 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18997), .ZN(
        P3_U3007) );
  AND2_X1 U22065 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18997), .ZN(
        P3_U3008) );
  AND2_X1 U22066 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18997), .ZN(
        P3_U3009) );
  AND2_X1 U22067 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18997), .ZN(
        P3_U3010) );
  AND2_X1 U22068 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18997), .ZN(
        P3_U3011) );
  AND2_X1 U22069 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18997), .ZN(
        P3_U3012) );
  AND2_X1 U22070 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18996), .ZN(
        P3_U3013) );
  AND2_X1 U22071 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18996), .ZN(
        P3_U3014) );
  AND2_X1 U22072 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18996), .ZN(
        P3_U3015) );
  AND2_X1 U22073 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18996), .ZN(
        P3_U3016) );
  AND2_X1 U22074 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18996), .ZN(
        P3_U3017) );
  AND2_X1 U22075 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18996), .ZN(
        P3_U3018) );
  AND2_X1 U22076 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18996), .ZN(
        P3_U3019) );
  AND2_X1 U22077 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18996), .ZN(
        P3_U3020) );
  AND2_X1 U22078 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18997), .ZN(P3_U3021) );
  AND2_X1 U22079 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18997), .ZN(P3_U3022) );
  AND2_X1 U22080 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18997), .ZN(P3_U3023) );
  AND2_X1 U22081 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18997), .ZN(P3_U3024) );
  AND2_X1 U22082 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18997), .ZN(P3_U3025) );
  AND2_X1 U22083 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18997), .ZN(P3_U3026) );
  AND2_X1 U22084 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18997), .ZN(P3_U3027) );
  AND2_X1 U22085 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18997), .ZN(P3_U3028) );
  NAND2_X1 U22086 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n19003) );
  NAND2_X1 U22087 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n19008) );
  AND3_X1 U22088 ( .A1(n19003), .A2(n19008), .A3(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19000) );
  NOR2_X1 U22089 ( .A1(n19151), .A2(n18998), .ZN(n19009) );
  OAI21_X1 U22090 ( .B1(n19009), .B2(n19014), .A(n19016), .ZN(n18999) );
  NAND3_X1 U22091 ( .A1(NA), .A2(n19014), .A3(n18998), .ZN(n19007) );
  OAI211_X1 U22092 ( .C1(n19083), .C2(n19000), .A(n18999), .B(n19007), .ZN(
        P3_U3029) );
  OAI21_X1 U22093 ( .B1(n19001), .B2(n21050), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19002) );
  OAI21_X1 U22094 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n19003), .A(n19002), 
        .ZN(n19004) );
  AOI22_X1 U22095 ( .A1(n19143), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19004), .ZN(n19006) );
  NAND2_X1 U22096 ( .A1(n19006), .A2(n19005), .ZN(P3_U3030) );
  AOI21_X1 U22097 ( .B1(n19014), .B2(n19007), .A(n19009), .ZN(n19015) );
  INV_X1 U22098 ( .A(n19008), .ZN(n19012) );
  INV_X1 U22099 ( .A(n19009), .ZN(n19010) );
  OAI22_X1 U22100 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19010), .ZN(n19011) );
  OAI22_X1 U22101 ( .A1(n19012), .A2(n19011), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19013) );
  OAI22_X1 U22102 ( .A1(n19015), .A2(n19016), .B1(n19014), .B2(n19013), .ZN(
        P3_U3031) );
  OAI222_X1 U22103 ( .A1(n19018), .A2(n19076), .B1(n19017), .B2(n19083), .C1(
        n19019), .C2(n19073), .ZN(P3_U3032) );
  INV_X1 U22104 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19021) );
  OAI222_X1 U22105 ( .A1(n19073), .A2(n19021), .B1(n19020), .B2(n19083), .C1(
        n19019), .C2(n19076), .ZN(P3_U3033) );
  OAI222_X1 U22106 ( .A1(n19073), .A2(n19023), .B1(n19022), .B2(n19083), .C1(
        n19021), .C2(n19076), .ZN(P3_U3034) );
  OAI222_X1 U22107 ( .A1(n19073), .A2(n19025), .B1(n19024), .B2(n19083), .C1(
        n19023), .C2(n19076), .ZN(P3_U3035) );
  OAI222_X1 U22108 ( .A1(n19073), .A2(n19027), .B1(n19026), .B2(n19083), .C1(
        n19025), .C2(n19076), .ZN(P3_U3036) );
  OAI222_X1 U22109 ( .A1(n19073), .A2(n19029), .B1(n19028), .B2(n19083), .C1(
        n19027), .C2(n19076), .ZN(P3_U3037) );
  OAI222_X1 U22110 ( .A1(n19073), .A2(n19032), .B1(n19030), .B2(n19083), .C1(
        n19029), .C2(n19076), .ZN(P3_U3038) );
  OAI222_X1 U22111 ( .A1(n19032), .A2(n19076), .B1(n19031), .B2(n19083), .C1(
        n19033), .C2(n19073), .ZN(P3_U3039) );
  OAI222_X1 U22112 ( .A1(n19073), .A2(n19035), .B1(n19034), .B2(n19083), .C1(
        n19033), .C2(n19076), .ZN(P3_U3040) );
  OAI222_X1 U22113 ( .A1(n19073), .A2(n19037), .B1(n19036), .B2(n19083), .C1(
        n19035), .C2(n19076), .ZN(P3_U3041) );
  INV_X1 U22114 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19039) );
  OAI222_X1 U22115 ( .A1(n19073), .A2(n19039), .B1(n19038), .B2(n19083), .C1(
        n19037), .C2(n19076), .ZN(P3_U3042) );
  OAI222_X1 U22116 ( .A1(n19073), .A2(n19041), .B1(n19040), .B2(n19083), .C1(
        n19039), .C2(n19076), .ZN(P3_U3043) );
  OAI222_X1 U22117 ( .A1(n19073), .A2(n19044), .B1(n19042), .B2(n19083), .C1(
        n19041), .C2(n19076), .ZN(P3_U3044) );
  OAI222_X1 U22118 ( .A1(n19044), .A2(n19076), .B1(n19043), .B2(n19083), .C1(
        n19045), .C2(n19073), .ZN(P3_U3045) );
  INV_X1 U22119 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19047) );
  OAI222_X1 U22120 ( .A1(n19073), .A2(n19047), .B1(n19046), .B2(n19083), .C1(
        n19045), .C2(n19076), .ZN(P3_U3046) );
  OAI222_X1 U22121 ( .A1(n19073), .A2(n19050), .B1(n19048), .B2(n19083), .C1(
        n19047), .C2(n19076), .ZN(P3_U3047) );
  OAI222_X1 U22122 ( .A1(n19050), .A2(n19076), .B1(n19049), .B2(n19083), .C1(
        n19051), .C2(n19073), .ZN(P3_U3048) );
  INV_X1 U22123 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19053) );
  OAI222_X1 U22124 ( .A1(n19073), .A2(n19053), .B1(n19052), .B2(n19083), .C1(
        n19051), .C2(n19076), .ZN(P3_U3049) );
  OAI222_X1 U22125 ( .A1(n19073), .A2(n19056), .B1(n19054), .B2(n19083), .C1(
        n19053), .C2(n19076), .ZN(P3_U3050) );
  OAI222_X1 U22126 ( .A1(n19056), .A2(n19076), .B1(n19055), .B2(n19083), .C1(
        n19057), .C2(n19073), .ZN(P3_U3051) );
  OAI222_X1 U22127 ( .A1(n19073), .A2(n19059), .B1(n19058), .B2(n19083), .C1(
        n19057), .C2(n19076), .ZN(P3_U3052) );
  OAI222_X1 U22128 ( .A1(n19073), .A2(n19062), .B1(n19060), .B2(n19083), .C1(
        n19059), .C2(n19076), .ZN(P3_U3053) );
  OAI222_X1 U22129 ( .A1(n19062), .A2(n19076), .B1(n19061), .B2(n19083), .C1(
        n19063), .C2(n19073), .ZN(P3_U3054) );
  OAI222_X1 U22130 ( .A1(n19073), .A2(n19065), .B1(n19064), .B2(n19083), .C1(
        n19063), .C2(n19076), .ZN(P3_U3055) );
  OAI222_X1 U22131 ( .A1(n19073), .A2(n19067), .B1(n19066), .B2(n19083), .C1(
        n19065), .C2(n19076), .ZN(P3_U3056) );
  OAI222_X1 U22132 ( .A1(n19073), .A2(n19070), .B1(n19068), .B2(n19083), .C1(
        n19067), .C2(n19076), .ZN(P3_U3057) );
  OAI222_X1 U22133 ( .A1(n19076), .A2(n19070), .B1(n19069), .B2(n19083), .C1(
        n19071), .C2(n19073), .ZN(P3_U3058) );
  OAI222_X1 U22134 ( .A1(n19073), .A2(n19074), .B1(n19072), .B2(n19083), .C1(
        n19071), .C2(n19076), .ZN(P3_U3059) );
  OAI222_X1 U22135 ( .A1(n19073), .A2(n19077), .B1(n19075), .B2(n19083), .C1(
        n19074), .C2(n19076), .ZN(P3_U3060) );
  OAI222_X1 U22136 ( .A1(n19073), .A2(n19079), .B1(n19078), .B2(n19083), .C1(
        n19077), .C2(n19076), .ZN(P3_U3061) );
  OAI22_X1 U22137 ( .A1(n19155), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19083), .ZN(n19080) );
  INV_X1 U22138 ( .A(n19080), .ZN(P3_U3274) );
  OAI22_X1 U22139 ( .A1(n19155), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19083), .ZN(n19081) );
  INV_X1 U22140 ( .A(n19081), .ZN(P3_U3275) );
  OAI22_X1 U22141 ( .A1(n19155), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19083), .ZN(n19082) );
  INV_X1 U22142 ( .A(n19082), .ZN(P3_U3276) );
  OAI22_X1 U22143 ( .A1(n19155), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19083), .ZN(n19084) );
  INV_X1 U22144 ( .A(n19084), .ZN(P3_U3277) );
  OAI21_X1 U22145 ( .B1(n19088), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19086), 
        .ZN(n19085) );
  INV_X1 U22146 ( .A(n19085), .ZN(P3_U3280) );
  OAI21_X1 U22147 ( .B1(n19088), .B2(n19087), .A(n19086), .ZN(P3_U3281) );
  OAI221_X1 U22148 ( .B1(n19091), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19091), 
        .C2(n19090), .A(n19089), .ZN(P3_U3282) );
  AOI22_X1 U22149 ( .A1(n19117), .A2(n19093), .B1(n19115), .B2(n19092), .ZN(
        n19098) );
  OAI21_X1 U22150 ( .B1(n19103), .B2(n19094), .A(n19119), .ZN(n19095) );
  INV_X1 U22151 ( .A(n19095), .ZN(n19097) );
  OAI22_X1 U22152 ( .A1(n19122), .A2(n19098), .B1(n19097), .B2(n19096), .ZN(
        P3_U3285) );
  OAI22_X1 U22153 ( .A1(n10078), .A2(n19099), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19110) );
  INV_X1 U22154 ( .A(n19110), .ZN(n19106) );
  NOR2_X1 U22155 ( .A1(n19100), .A2(n19118), .ZN(n19109) );
  OAI22_X1 U22156 ( .A1(n19104), .A2(n19103), .B1(n19102), .B2(n19101), .ZN(
        n19105) );
  AOI21_X1 U22157 ( .B1(n19106), .B2(n19109), .A(n19105), .ZN(n19107) );
  AOI22_X1 U22158 ( .A1(n19122), .A2(n19108), .B1(n19107), .B2(n19119), .ZN(
        P3_U3288) );
  AOI222_X1 U22159 ( .A1(n19112), .A2(n19117), .B1(n19115), .B2(n19111), .C1(
        n19110), .C2(n19109), .ZN(n19113) );
  AOI22_X1 U22160 ( .A1(n19122), .A2(n19114), .B1(n19113), .B2(n19119), .ZN(
        P3_U3289) );
  AOI222_X1 U22161 ( .A1(n19118), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19117), 
        .B2(n19116), .C1(n19121), .C2(n19115), .ZN(n19120) );
  AOI22_X1 U22162 ( .A1(n19122), .A2(n19121), .B1(n19120), .B2(n19119), .ZN(
        P3_U3290) );
  AOI211_X1 U22163 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19123) );
  AOI21_X1 U22164 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19123), .ZN(n19125) );
  INV_X1 U22165 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U22166 ( .A1(n19129), .A2(n19125), .B1(n19124), .B2(n19126), .ZN(
        P3_U3292) );
  NOR2_X1 U22167 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19128) );
  INV_X1 U22168 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19127) );
  AOI22_X1 U22169 ( .A1(n19129), .A2(n19128), .B1(n19127), .B2(n19126), .ZN(
        P3_U3293) );
  INV_X1 U22170 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19130) );
  AOI22_X1 U22171 ( .A1(n19083), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19130), 
        .B2(n19155), .ZN(P3_U3294) );
  INV_X1 U22172 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n19139) );
  OAI22_X1 U22173 ( .A1(n19134), .A2(n19133), .B1(n19132), .B2(n19131), .ZN(
        n19136) );
  OAI21_X1 U22174 ( .B1(n19136), .B2(n19135), .A(n19138), .ZN(n19137) );
  OAI21_X1 U22175 ( .B1(n19139), .B2(n19138), .A(n19137), .ZN(P3_U3295) );
  OAI21_X1 U22176 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19141), .A(n19140), 
        .ZN(n19144) );
  AOI211_X1 U22177 ( .C1(n19157), .C2(n19144), .A(n19143), .B(n19142), .ZN(
        n19147) );
  OAI21_X1 U22178 ( .B1(n19147), .B2(n19146), .A(n19145), .ZN(n19154) );
  NOR2_X1 U22179 ( .A1(n19149), .A2(n19148), .ZN(n19150) );
  AOI211_X1 U22180 ( .C1(n19152), .C2(n19151), .A(n19150), .B(n19162), .ZN(
        n19153) );
  MUX2_X1 U22181 ( .A(n19154), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19153), 
        .Z(P3_U3296) );
  MUX2_X1 U22182 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19155), .Z(P3_U3297) );
  OAI21_X1 U22183 ( .B1(n19159), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19158), 
        .ZN(n19156) );
  OAI21_X1 U22184 ( .B1(n19158), .B2(n19157), .A(n19156), .ZN(P3_U3298) );
  NOR2_X1 U22185 ( .A1(n19159), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19161)
         );
  OAI21_X1 U22186 ( .B1(n19162), .B2(n19161), .A(n19160), .ZN(P3_U3299) );
  INV_X1 U22187 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19167) );
  NAND2_X1 U22188 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20045), .ZN(n20035) );
  NAND2_X1 U22189 ( .A1(n19167), .A2(n19163), .ZN(n20032) );
  OAI21_X1 U22190 ( .B1(n19167), .B2(n20035), .A(n20032), .ZN(n20100) );
  AOI21_X1 U22191 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20100), .ZN(n19164) );
  INV_X1 U22192 ( .A(n19164), .ZN(P2_U2815) );
  INV_X1 U22193 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19168) );
  OAI22_X1 U22194 ( .A1(n19166), .A2(n19168), .B1(n21322), .B2(n19165), .ZN(
        P2_U2816) );
  NAND2_X1 U22195 ( .A1(n19167), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20168) );
  INV_X2 U22196 ( .A(n20168), .ZN(n20092) );
  AOI22_X1 U22197 ( .A1(n20092), .A2(n19168), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20168), .ZN(n19169) );
  OAI21_X1 U22198 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20032), .A(n19169), 
        .ZN(P2_U2817) );
  OAI21_X1 U22199 ( .B1(n20038), .B2(BS16), .A(n20100), .ZN(n20098) );
  OAI21_X1 U22200 ( .B1(n20100), .B2(n20153), .A(n20098), .ZN(P2_U2818) );
  NOR4_X1 U22201 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19173) );
  NOR4_X1 U22202 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19172) );
  NOR4_X1 U22203 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19171) );
  NOR4_X1 U22204 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19170) );
  NAND4_X1 U22205 ( .A1(n19173), .A2(n19172), .A3(n19171), .A4(n19170), .ZN(
        n19179) );
  NOR4_X1 U22206 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19177) );
  AOI211_X1 U22207 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_5__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19176) );
  NOR4_X1 U22208 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19175) );
  NOR4_X1 U22209 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19174) );
  NAND4_X1 U22210 ( .A1(n19177), .A2(n19176), .A3(n19175), .A4(n19174), .ZN(
        n19178) );
  NOR2_X1 U22211 ( .A1(n19179), .A2(n19178), .ZN(n19189) );
  INV_X1 U22212 ( .A(n19189), .ZN(n19181) );
  NOR2_X1 U22213 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19181), .ZN(n19183) );
  INV_X1 U22214 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19180) );
  AOI22_X1 U22215 ( .A1(n19183), .A2(n19342), .B1(n19181), .B2(n19180), .ZN(
        P2_U2820) );
  NOR2_X1 U22216 ( .A1(n19189), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19182)
         );
  OR4_X1 U22217 ( .A1(n19181), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19187) );
  OAI21_X1 U22218 ( .B1(n19183), .B2(n19182), .A(n19187), .ZN(P2_U2821) );
  INV_X1 U22219 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20099) );
  NAND2_X1 U22220 ( .A1(n19183), .A2(n20099), .ZN(n19186) );
  OAI21_X1 U22221 ( .B1(n20046), .B2(n19342), .A(n19189), .ZN(n19184) );
  OAI21_X1 U22222 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19189), .A(n19184), 
        .ZN(n19185) );
  OAI221_X1 U22223 ( .B1(n19186), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19186), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19185), .ZN(P2_U2822) );
  INV_X1 U22224 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19188) );
  OAI211_X1 U22225 ( .C1(n19189), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        P2_U2823) );
  NAND2_X1 U22226 ( .A1(n19327), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n19190) );
  OAI211_X1 U22227 ( .C1(n19282), .C2(n19191), .A(n19190), .B(n15303), .ZN(
        n19192) );
  AOI21_X1 U22228 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19344), .A(n19192), .ZN(
        n19193) );
  OAI21_X1 U22229 ( .B1(n19194), .B2(n19346), .A(n19193), .ZN(n19199) );
  AOI211_X1 U22230 ( .C1(n19197), .C2(n19196), .A(n20024), .B(n19195), .ZN(
        n19198) );
  AOI211_X1 U22231 ( .C1(n19339), .C2(n19200), .A(n19199), .B(n19198), .ZN(
        n19201) );
  OAI21_X1 U22232 ( .B1(n19202), .B2(n19335), .A(n19201), .ZN(P2_U2836) );
  OAI22_X1 U22233 ( .A1(n20073), .A2(n19341), .B1(n19203), .B2(n19282), .ZN(
        n19204) );
  AOI211_X1 U22234 ( .C1(n19209), .C2(n19241), .A(n19326), .B(n19204), .ZN(
        n19205) );
  OAI21_X1 U22235 ( .B1(n19206), .B2(n19306), .A(n19205), .ZN(n19207) );
  AOI21_X1 U22236 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19344), .A(n19207), .ZN(
        n19214) );
  NAND2_X1 U22237 ( .A1(n19209), .A2(n19208), .ZN(n19211) );
  AOI22_X1 U22238 ( .A1(n19212), .A2(n19211), .B1(n12566), .B2(n19210), .ZN(
        n19213) );
  OAI211_X1 U22239 ( .C1(n19215), .C2(n19335), .A(n19214), .B(n19213), .ZN(
        P2_U2838) );
  NOR2_X1 U22240 ( .A1(n19312), .A2(n19216), .ZN(n19218) );
  XOR2_X1 U22241 ( .A(n19218), .B(n19217), .Z(n19226) );
  OAI22_X1 U22242 ( .A1(n19219), .A2(n19306), .B1(n19324), .B2(n19355), .ZN(
        n19220) );
  INV_X1 U22243 ( .A(n19220), .ZN(n19221) );
  OAI211_X1 U22244 ( .C1(n15513), .C2(n19341), .A(n19221), .B(n15303), .ZN(
        n19222) );
  AOI21_X1 U22245 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19349), .A(
        n19222), .ZN(n19225) );
  OAI22_X1 U22246 ( .A1(n19359), .A2(n19346), .B1(n19335), .B2(n19399), .ZN(
        n19223) );
  INV_X1 U22247 ( .A(n19223), .ZN(n19224) );
  OAI211_X1 U22248 ( .C1(n20024), .C2(n19226), .A(n19225), .B(n19224), .ZN(
        P2_U2839) );
  NAND2_X1 U22249 ( .A1(n9751), .A2(n19227), .ZN(n19229) );
  XNOR2_X1 U22250 ( .A(n19229), .B(n19228), .ZN(n19237) );
  AOI22_X1 U22251 ( .A1(n19230), .A2(n19339), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19344), .ZN(n19231) );
  OAI211_X1 U22252 ( .C1(n15279), .C2(n19341), .A(n19231), .B(n15303), .ZN(
        n19235) );
  OAI22_X1 U22253 ( .A1(n19233), .A2(n19346), .B1(n19335), .B2(n19232), .ZN(
        n19234) );
  AOI211_X1 U22254 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19349), .A(
        n19235), .B(n19234), .ZN(n19236) );
  OAI21_X1 U22255 ( .B1(n19237), .B2(n20024), .A(n19236), .ZN(P2_U2840) );
  AOI22_X1 U22256 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19349), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19327), .ZN(n19238) );
  OAI211_X1 U22257 ( .C1(n19239), .C2(n19306), .A(n19238), .B(n15303), .ZN(
        n19240) );
  AOI21_X1 U22258 ( .B1(n9874), .B2(n19241), .A(n19240), .ZN(n19249) );
  NAND2_X1 U22259 ( .A1(n9874), .A2(n19242), .ZN(n19246) );
  OAI22_X1 U22260 ( .A1(n19244), .A2(n19335), .B1(n19346), .B2(n19243), .ZN(
        n19245) );
  AOI21_X1 U22261 ( .B1(n19247), .B2(n19246), .A(n19245), .ZN(n19248) );
  OAI211_X1 U22262 ( .C1(n19324), .C2(n12051), .A(n19249), .B(n19248), .ZN(
        P2_U2842) );
  AOI22_X1 U22263 ( .A1(n19344), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19349), .ZN(n19250) );
  OAI21_X1 U22264 ( .B1(n19251), .B2(n19306), .A(n19250), .ZN(n19252) );
  AOI211_X1 U22265 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19327), .A(n19326), 
        .B(n19252), .ZN(n19259) );
  NOR2_X1 U22266 ( .A1(n19312), .A2(n19253), .ZN(n19255) );
  XNOR2_X1 U22267 ( .A(n19255), .B(n19254), .ZN(n19257) );
  INV_X1 U22268 ( .A(n19371), .ZN(n19256) );
  AOI22_X1 U22269 ( .A1(n19257), .A2(n19336), .B1(n12566), .B2(n19256), .ZN(
        n19258) );
  OAI211_X1 U22270 ( .C1(n19411), .C2(n19335), .A(n19259), .B(n19258), .ZN(
        P2_U2843) );
  OAI22_X1 U22271 ( .A1(n19260), .A2(n19306), .B1(n19324), .B2(n13669), .ZN(
        n19261) );
  INV_X1 U22272 ( .A(n19261), .ZN(n19262) );
  OAI21_X1 U22273 ( .B1(n19263), .B2(n19282), .A(n19262), .ZN(n19264) );
  AOI211_X1 U22274 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19327), .A(n19326), 
        .B(n19264), .ZN(n19271) );
  NAND2_X1 U22275 ( .A1(n9751), .A2(n19265), .ZN(n19267) );
  XNOR2_X1 U22276 ( .A(n19267), .B(n19266), .ZN(n19269) );
  AOI22_X1 U22277 ( .A1(n19269), .A2(n19336), .B1(n12566), .B2(n19268), .ZN(
        n19270) );
  OAI211_X1 U22278 ( .C1(n19272), .C2(n19335), .A(n19271), .B(n19270), .ZN(
        P2_U2844) );
  OAI22_X1 U22279 ( .A1(n19273), .A2(n19306), .B1(n19324), .B2(n10247), .ZN(
        n19274) );
  AOI211_X1 U22280 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19327), .A(n19326), 
        .B(n19274), .ZN(n19281) );
  NOR2_X1 U22281 ( .A1(n19312), .A2(n19275), .ZN(n19276) );
  XNOR2_X1 U22282 ( .A(n19277), .B(n19276), .ZN(n19279) );
  OAI22_X1 U22283 ( .A1(n19414), .A2(n19335), .B1(n19346), .B2(n19378), .ZN(
        n19278) );
  AOI21_X1 U22284 ( .B1(n19279), .B2(n19336), .A(n19278), .ZN(n19280) );
  OAI211_X1 U22285 ( .C1(n10304), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        P2_U2845) );
  NAND2_X1 U22286 ( .A1(n9751), .A2(n19283), .ZN(n19285) );
  XOR2_X1 U22287 ( .A(n19285), .B(n19284), .Z(n19293) );
  AOI22_X1 U22288 ( .A1(n19286), .A2(n19339), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19344), .ZN(n19287) );
  OAI211_X1 U22289 ( .C1(n20061), .C2(n19341), .A(n19287), .B(n15303), .ZN(
        n19291) );
  OAI22_X1 U22290 ( .A1(n19289), .A2(n19335), .B1(n19346), .B2(n19288), .ZN(
        n19290) );
  AOI211_X1 U22291 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19349), .A(
        n19291), .B(n19290), .ZN(n19292) );
  OAI21_X1 U22292 ( .B1(n19293), .B2(n20024), .A(n19292), .ZN(P2_U2846) );
  NAND2_X1 U22293 ( .A1(n9751), .A2(n19294), .ZN(n19296) );
  XOR2_X1 U22294 ( .A(n19296), .B(n19295), .Z(n19304) );
  AOI22_X1 U22295 ( .A1(n19297), .A2(n19339), .B1(n19344), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n19298) );
  OAI211_X1 U22296 ( .C1(n20057), .C2(n19341), .A(n19298), .B(n15303), .ZN(
        n19302) );
  OAI22_X1 U22297 ( .A1(n19300), .A2(n19335), .B1(n19346), .B2(n19299), .ZN(
        n19301) );
  AOI211_X1 U22298 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19349), .A(
        n19302), .B(n19301), .ZN(n19303) );
  OAI21_X1 U22299 ( .B1(n19304), .B2(n20024), .A(n19303), .ZN(P2_U2848) );
  INV_X1 U22300 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20055) );
  OAI21_X1 U22301 ( .B1(n20055), .B2(n19341), .A(n19305), .ZN(n19310) );
  OAI22_X1 U22302 ( .A1(n19324), .A2(n19308), .B1(n19307), .B2(n19306), .ZN(
        n19309) );
  AOI211_X1 U22303 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19349), .A(
        n19310), .B(n19309), .ZN(n19318) );
  NOR2_X1 U22304 ( .A1(n19312), .A2(n19311), .ZN(n19314) );
  XNOR2_X1 U22305 ( .A(n19314), .B(n19313), .ZN(n19316) );
  AOI22_X1 U22306 ( .A1(n19316), .A2(n19336), .B1(n12566), .B2(n19315), .ZN(
        n19317) );
  OAI211_X1 U22307 ( .C1(n19335), .C2(n19319), .A(n19318), .B(n19317), .ZN(
        P2_U2849) );
  INV_X1 U22308 ( .A(n19320), .ZN(n19321) );
  AOI22_X1 U22309 ( .A1(n19321), .A2(n19339), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19349), .ZN(n19322) );
  OAI21_X1 U22310 ( .B1(n19324), .B2(n19323), .A(n19322), .ZN(n19325) );
  AOI211_X1 U22311 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19327), .A(n19326), .B(
        n19325), .ZN(n19334) );
  NAND2_X1 U22312 ( .A1(n9751), .A2(n19328), .ZN(n19329) );
  XNOR2_X1 U22313 ( .A(n19330), .B(n19329), .ZN(n19332) );
  AOI22_X1 U22314 ( .A1(n19332), .A2(n19336), .B1(n12566), .B2(n19331), .ZN(
        n19333) );
  OAI211_X1 U22315 ( .C1(n19335), .C2(n19427), .A(n19334), .B(n19333), .ZN(
        P2_U2850) );
  AOI22_X1 U22316 ( .A1(n19339), .A2(n19338), .B1(n19337), .B2(n10422), .ZN(
        n19340) );
  OAI21_X1 U22317 ( .B1(n19342), .B2(n19341), .A(n19340), .ZN(n19343) );
  AOI21_X1 U22318 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19344), .A(n19343), .ZN(
        n19345) );
  OAI21_X1 U22319 ( .B1(n9816), .B2(n19346), .A(n19345), .ZN(n19347) );
  AOI21_X1 U22320 ( .B1(n19501), .B2(n19348), .A(n19347), .ZN(n19351) );
  NAND2_X1 U22321 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19349), .ZN(
        n19350) );
  OAI211_X1 U22322 ( .C1(n19352), .C2(n16419), .A(n19351), .B(n19350), .ZN(
        P2_U2855) );
  NOR2_X1 U22323 ( .A1(n13742), .A2(n19353), .ZN(n19354) );
  OR2_X1 U22324 ( .A1(n15002), .A2(n19354), .ZN(n19401) );
  OAI22_X1 U22325 ( .A1(n19401), .A2(n19380), .B1(n19356), .B2(n19355), .ZN(
        n19357) );
  INV_X1 U22326 ( .A(n19357), .ZN(n19358) );
  OAI21_X1 U22327 ( .B1(n19385), .B2(n19359), .A(n19358), .ZN(P2_U2871) );
  AOI21_X1 U22328 ( .B1(n19366), .B2(n19361), .A(n19360), .ZN(n19362) );
  NOR3_X1 U22329 ( .A1(n19362), .A2(n9845), .A3(n19380), .ZN(n19363) );
  AOI21_X1 U22330 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19385), .A(n19363), .ZN(
        n19364) );
  OAI21_X1 U22331 ( .B1(n19365), .B2(n19385), .A(n19364), .ZN(P2_U2873) );
  AOI211_X1 U22332 ( .C1(n19368), .C2(n19367), .A(n19380), .B(n19366), .ZN(
        n19369) );
  AOI21_X1 U22333 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19385), .A(n19369), .ZN(
        n19370) );
  OAI21_X1 U22334 ( .B1(n19371), .B2(n19385), .A(n19370), .ZN(P2_U2875) );
  NOR2_X1 U22335 ( .A1(n19372), .A2(n19380), .ZN(n19376) );
  OAI21_X1 U22336 ( .B1(n13521), .B2(n19374), .A(n19373), .ZN(n19375) );
  AOI22_X1 U22337 ( .A1(n19376), .A2(n19375), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19385), .ZN(n19377) );
  OAI21_X1 U22338 ( .B1(n19378), .B2(n19385), .A(n19377), .ZN(P2_U2877) );
  INV_X1 U22339 ( .A(n19379), .ZN(n19381) );
  AOI21_X1 U22340 ( .B1(n9943), .B2(n19381), .A(n19380), .ZN(n19382) );
  AOI22_X1 U22341 ( .A1(n19382), .A2(n13521), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19385), .ZN(n19383) );
  OAI21_X1 U22342 ( .B1(n19384), .B2(n19385), .A(n19383), .ZN(P2_U2879) );
  INV_X1 U22343 ( .A(n19423), .ZN(n19387) );
  AOI22_X1 U22344 ( .A1(n19387), .A2(n19386), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19385), .ZN(n19388) );
  OAI21_X1 U22345 ( .B1(n19385), .B2(n19389), .A(n19388), .ZN(P2_U2883) );
  INV_X1 U22346 ( .A(n19390), .ZN(n19391) );
  AOI22_X1 U22347 ( .A1(n19397), .A2(BUF1_REG_31__SCAN_IN), .B1(n19392), .B2(
        n19391), .ZN(n19394) );
  AOI22_X1 U22348 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19419), .B1(n19398), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19393) );
  NAND2_X1 U22349 ( .A1(n19394), .A2(n19393), .ZN(P2_U2888) );
  INV_X1 U22350 ( .A(n19461), .ZN(n19395) );
  AOI22_X1 U22351 ( .A1(n19396), .A2(n19395), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19419), .ZN(n19405) );
  AOI22_X1 U22352 ( .A1(n19398), .A2(BUF2_REG_16__SCAN_IN), .B1(n19397), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19404) );
  OAI22_X1 U22353 ( .A1(n19401), .A2(n19422), .B1(n19400), .B2(n19399), .ZN(
        n19402) );
  INV_X1 U22354 ( .A(n19402), .ZN(n19403) );
  NAND3_X1 U22355 ( .A1(n19405), .A2(n19404), .A3(n19403), .ZN(P2_U2903) );
  AOI22_X1 U22356 ( .A1(n19421), .A2(n19406), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19419), .ZN(n19407) );
  OAI21_X1 U22357 ( .B1(n19428), .B2(n19408), .A(n19407), .ZN(P2_U2905) );
  AOI22_X1 U22358 ( .A1(n19421), .A2(n19409), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19419), .ZN(n19410) );
  OAI21_X1 U22359 ( .B1(n19428), .B2(n19411), .A(n19410), .ZN(P2_U2907) );
  AOI22_X1 U22360 ( .A1(n19421), .A2(n19412), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19419), .ZN(n19413) );
  OAI21_X1 U22361 ( .B1(n19428), .B2(n19414), .A(n19413), .ZN(P2_U2909) );
  AOI22_X1 U22362 ( .A1(n19421), .A2(n19415), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19419), .ZN(n19416) );
  OAI21_X1 U22363 ( .B1(n19428), .B2(n19417), .A(n19416), .ZN(P2_U2911) );
  INV_X1 U22364 ( .A(n19418), .ZN(n19420) );
  AOI22_X1 U22365 ( .A1(n19421), .A2(n19420), .B1(n19419), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n19426) );
  OR3_X1 U22366 ( .A1(n19424), .A2(n19423), .A3(n19422), .ZN(n19425) );
  OAI211_X1 U22367 ( .C1(n19428), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        P2_U2914) );
  AND2_X1 U22368 ( .A1(n19458), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22369 ( .A1(n13158), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19430) );
  OAI21_X1 U22370 ( .B1(n13041), .B2(n19460), .A(n19430), .ZN(P2_U2936) );
  AOI22_X1 U22371 ( .A1(n13158), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19431) );
  OAI21_X1 U22372 ( .B1(n19432), .B2(n19460), .A(n19431), .ZN(P2_U2937) );
  AOI22_X1 U22373 ( .A1(n13158), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19433) );
  OAI21_X1 U22374 ( .B1(n19434), .B2(n19460), .A(n19433), .ZN(P2_U2938) );
  AOI22_X1 U22375 ( .A1(n13158), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19435) );
  OAI21_X1 U22376 ( .B1(n19436), .B2(n19460), .A(n19435), .ZN(P2_U2939) );
  AOI22_X1 U22377 ( .A1(n13158), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19437) );
  OAI21_X1 U22378 ( .B1(n19438), .B2(n19460), .A(n19437), .ZN(P2_U2940) );
  AOI22_X1 U22379 ( .A1(n13158), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19439) );
  OAI21_X1 U22380 ( .B1(n19440), .B2(n19460), .A(n19439), .ZN(P2_U2941) );
  AOI22_X1 U22381 ( .A1(n13158), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19441) );
  OAI21_X1 U22382 ( .B1(n19442), .B2(n19460), .A(n19441), .ZN(P2_U2942) );
  AOI22_X1 U22383 ( .A1(n13158), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19443) );
  OAI21_X1 U22384 ( .B1(n19444), .B2(n19460), .A(n19443), .ZN(P2_U2943) );
  AOI22_X1 U22385 ( .A1(n13158), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22386 ( .B1(n19446), .B2(n19460), .A(n19445), .ZN(P2_U2944) );
  AOI22_X1 U22387 ( .A1(n13158), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19447) );
  OAI21_X1 U22388 ( .B1(n19448), .B2(n19460), .A(n19447), .ZN(P2_U2945) );
  INV_X1 U22389 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19450) );
  AOI22_X1 U22390 ( .A1(n13158), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19449) );
  OAI21_X1 U22391 ( .B1(n19450), .B2(n19460), .A(n19449), .ZN(P2_U2946) );
  AOI22_X1 U22392 ( .A1(n13158), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19451) );
  OAI21_X1 U22393 ( .B1(n13678), .B2(n19460), .A(n19451), .ZN(P2_U2947) );
  INV_X1 U22394 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19453) );
  AOI22_X1 U22395 ( .A1(n13158), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19452) );
  OAI21_X1 U22396 ( .B1(n19453), .B2(n19460), .A(n19452), .ZN(P2_U2948) );
  INV_X1 U22397 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19455) );
  AOI22_X1 U22398 ( .A1(n13158), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19454) );
  OAI21_X1 U22399 ( .B1(n19455), .B2(n19460), .A(n19454), .ZN(P2_U2949) );
  INV_X1 U22400 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19457) );
  AOI22_X1 U22401 ( .A1(n13158), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19456) );
  OAI21_X1 U22402 ( .B1(n19457), .B2(n19460), .A(n19456), .ZN(P2_U2950) );
  AOI22_X1 U22403 ( .A1(n13158), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19458), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19459) );
  OAI21_X1 U22404 ( .B1(n13043), .B2(n19460), .A(n19459), .ZN(P2_U2951) );
  AOI22_X1 U22405 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19494), .ZN(n19886) );
  INV_X1 U22406 ( .A(n19886), .ZN(n19962) );
  NOR2_X2 U22407 ( .A1(n19490), .A2(n9813), .ZN(n19960) );
  AOI22_X1 U22408 ( .A1(n19962), .A2(n20015), .B1(n19491), .B2(n19960), .ZN(
        n19463) );
  NOR2_X2 U22409 ( .A1(n19461), .A2(n19917), .ZN(n19961) );
  AOI22_X1 U22410 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19494), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19493), .ZN(n19820) );
  AOI22_X1 U22411 ( .A1(n19961), .A2(n19495), .B1(n19524), .B2(n19963), .ZN(
        n19462) );
  OAI211_X1 U22412 ( .C1(n19499), .C2(n19464), .A(n19463), .B(n19462), .ZN(
        P2_U3048) );
  OAI22_X2 U22413 ( .A1(n19466), .A2(n19488), .B1(n19465), .B2(n19487), .ZN(
        n19976) );
  AOI22_X1 U22414 ( .A1(n19976), .A2(n20015), .B1(n19491), .B2(n19974), .ZN(
        n19471) );
  AOI22_X2 U22415 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19494), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19493), .ZN(n19892) );
  INV_X1 U22416 ( .A(n19892), .ZN(n19975) );
  AOI22_X1 U22417 ( .A1(n19469), .A2(n19495), .B1(n19524), .B2(n19975), .ZN(
        n19470) );
  OAI211_X1 U22418 ( .C1(n19499), .C2(n19472), .A(n19471), .B(n19470), .ZN(
        P2_U3050) );
  AOI22_X1 U22419 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19494), .ZN(n19795) );
  INV_X1 U22420 ( .A(n19795), .ZN(n19982) );
  NOR2_X2 U22421 ( .A1(n19490), .A2(n11623), .ZN(n19980) );
  AOI22_X1 U22422 ( .A1(n19982), .A2(n20015), .B1(n19491), .B2(n19980), .ZN(
        n19475) );
  NOR2_X2 U22423 ( .A1(n19473), .A2(n19917), .ZN(n19981) );
  AOI22_X1 U22424 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19494), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19493), .ZN(n19895) );
  AOI22_X1 U22425 ( .A1(n19981), .A2(n19495), .B1(n19524), .B2(n19983), .ZN(
        n19474) );
  OAI211_X1 U22426 ( .C1(n19499), .C2(n12661), .A(n19475), .B(n19474), .ZN(
        P2_U3051) );
  AOI22_X2 U22427 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19494), .ZN(n19898) );
  INV_X1 U22428 ( .A(n19898), .ZN(n19989) );
  AOI22_X1 U22429 ( .A1(n19989), .A2(n20015), .B1(n19491), .B2(n19987), .ZN(
        n19480) );
  NOR2_X2 U22430 ( .A1(n19477), .A2(n19917), .ZN(n19988) );
  OAI22_X2 U22431 ( .A1(n21160), .A2(n19488), .B1(n19478), .B2(n19487), .ZN(
        n19990) );
  AOI22_X1 U22432 ( .A1(n19988), .A2(n19495), .B1(n19524), .B2(n19990), .ZN(
        n19479) );
  OAI211_X1 U22433 ( .C1(n19499), .C2(n19481), .A(n19480), .B(n19479), .ZN(
        P2_U3052) );
  AOI22_X1 U22434 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19493), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19494), .ZN(n19905) );
  NOR2_X2 U22435 ( .A1(n19490), .A2(n11548), .ZN(n20001) );
  AOI22_X1 U22436 ( .A1(n20004), .A2(n20015), .B1(n19491), .B2(n20001), .ZN(
        n19486) );
  NOR2_X2 U22437 ( .A1(n19482), .A2(n19917), .ZN(n20002) );
  AOI22_X1 U22438 ( .A1(n20002), .A2(n19495), .B1(n19524), .B2(n20003), .ZN(
        n19485) );
  OAI211_X1 U22439 ( .C1(n19499), .C2(n21331), .A(n19486), .B(n19485), .ZN(
        P2_U3054) );
  NOR2_X2 U22440 ( .A1(n19490), .A2(n10266), .ZN(n20008) );
  AOI22_X1 U22441 ( .A1(n20012), .A2(n20015), .B1(n19491), .B2(n20008), .ZN(
        n19497) );
  NOR2_X2 U22442 ( .A1(n19492), .A2(n19917), .ZN(n20010) );
  AOI22_X1 U22443 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19494), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19493), .ZN(n19911) );
  AOI22_X1 U22444 ( .A1(n20010), .A2(n19495), .B1(n19524), .B2(n20014), .ZN(
        n19496) );
  OAI211_X1 U22445 ( .C1(n19499), .C2(n19498), .A(n19497), .B(n19496), .ZN(
        P2_U3055) );
  NAND2_X1 U22446 ( .A1(n19563), .A2(n11863), .ZN(n19505) );
  INV_X1 U22447 ( .A(n20102), .ZN(n19958) );
  NOR2_X1 U22448 ( .A1(n21258), .A2(n19505), .ZN(n19527) );
  OAI21_X1 U22449 ( .B1(n19502), .B2(n19527), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19503) );
  OAI21_X1 U22450 ( .B1(n19505), .B2(n19958), .A(n19503), .ZN(n19528) );
  AOI22_X1 U22451 ( .A1(n19528), .A2(n19961), .B1(n19960), .B2(n19527), .ZN(
        n19511) );
  NAND2_X1 U22452 ( .A1(n19504), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19693) );
  OAI21_X1 U22453 ( .B1(n19693), .B2(n19750), .A(n19505), .ZN(n19509) );
  INV_X1 U22454 ( .A(n19527), .ZN(n19506) );
  OAI211_X1 U22455 ( .C1(n19507), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19506), 
        .B(n19958), .ZN(n19508) );
  NAND3_X1 U22456 ( .A1(n19509), .A2(n19952), .A3(n19508), .ZN(n19529) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n19962), .ZN(n19510) );
  OAI211_X1 U22458 ( .C1(n19820), .C2(n19562), .A(n19511), .B(n19510), .ZN(
        P2_U3056) );
  AOI22_X1 U22459 ( .A1(n19528), .A2(n19968), .B1(n19967), .B2(n19527), .ZN(
        n19514) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n19969), .ZN(n19513) );
  OAI211_X1 U22461 ( .C1(n19823), .C2(n19562), .A(n19514), .B(n19513), .ZN(
        P2_U3057) );
  AOI22_X1 U22462 ( .A1(n19528), .A2(n19469), .B1(n19974), .B2(n19527), .ZN(
        n19516) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n19976), .ZN(n19515) );
  OAI211_X1 U22464 ( .C1(n19892), .C2(n19562), .A(n19516), .B(n19515), .ZN(
        P2_U3058) );
  AOI22_X1 U22465 ( .A1(n19528), .A2(n19981), .B1(n19980), .B2(n19527), .ZN(
        n19518) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n19982), .ZN(n19517) );
  OAI211_X1 U22467 ( .C1(n19895), .C2(n19562), .A(n19518), .B(n19517), .ZN(
        P2_U3059) );
  AOI22_X1 U22468 ( .A1(n19528), .A2(n19988), .B1(n19987), .B2(n19527), .ZN(
        n19520) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19529), .B1(
        n19554), .B2(n19990), .ZN(n19519) );
  OAI211_X1 U22470 ( .C1(n19898), .C2(n19532), .A(n19520), .B(n19519), .ZN(
        P2_U3060) );
  AOI22_X1 U22471 ( .A1(n19528), .A2(n19995), .B1(n19994), .B2(n19527), .ZN(
        n19523) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n19997), .ZN(n19522) );
  OAI211_X1 U22473 ( .C1(n19864), .C2(n19562), .A(n19523), .B(n19522), .ZN(
        P2_U3061) );
  AOI22_X1 U22474 ( .A1(n19528), .A2(n20002), .B1(n20001), .B2(n19527), .ZN(
        n19526) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19529), .B1(
        n19524), .B2(n20004), .ZN(n19525) );
  OAI211_X1 U22476 ( .C1(n19835), .C2(n19562), .A(n19526), .B(n19525), .ZN(
        P2_U3062) );
  AOI22_X1 U22477 ( .A1(n19528), .A2(n20010), .B1(n20008), .B2(n19527), .ZN(
        n19531) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19529), .B1(
        n19554), .B2(n20014), .ZN(n19530) );
  OAI211_X1 U22479 ( .C1(n19842), .C2(n19532), .A(n19531), .B(n19530), .ZN(
        P2_U3063) );
  INV_X1 U22480 ( .A(n19536), .ZN(n19533) );
  NOR3_X2 U22481 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11863), .A3(
        n19565), .ZN(n19557) );
  OAI21_X1 U22482 ( .B1(n19533), .B2(n19557), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19535) );
  INV_X1 U22483 ( .A(n19781), .ZN(n19534) );
  NAND2_X1 U22484 ( .A1(n19563), .A2(n19534), .ZN(n19538) );
  NAND2_X1 U22485 ( .A1(n19535), .A2(n19538), .ZN(n19558) );
  AOI22_X1 U22486 ( .A1(n19558), .A2(n19961), .B1(n19960), .B2(n19557), .ZN(
        n19543) );
  AOI21_X1 U22487 ( .B1(n19536), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19541) );
  INV_X1 U22488 ( .A(n20103), .ZN(n19537) );
  OAI21_X1 U22489 ( .B1(n19589), .B2(n19554), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19539) );
  NAND3_X1 U22490 ( .A1(n19539), .A2(n20102), .A3(n19538), .ZN(n19540) );
  OAI211_X1 U22491 ( .C1(n19557), .C2(n19541), .A(n19540), .B(n19952), .ZN(
        n19559) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19559), .B1(
        n19589), .B2(n19963), .ZN(n19542) );
  OAI211_X1 U22493 ( .C1(n19886), .C2(n19562), .A(n19543), .B(n19542), .ZN(
        P2_U3064) );
  AOI22_X1 U22494 ( .A1(n19558), .A2(n19968), .B1(n19967), .B2(n19557), .ZN(
        n19545) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19559), .B1(
        n19589), .B2(n19970), .ZN(n19544) );
  OAI211_X1 U22496 ( .C1(n19889), .C2(n19562), .A(n19545), .B(n19544), .ZN(
        P2_U3065) );
  AOI22_X1 U22497 ( .A1(n19558), .A2(n19469), .B1(n19974), .B2(n19557), .ZN(
        n19547) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19559), .B1(
        n19554), .B2(n19976), .ZN(n19546) );
  OAI211_X1 U22499 ( .C1(n19892), .C2(n19597), .A(n19547), .B(n19546), .ZN(
        P2_U3066) );
  AOI22_X1 U22500 ( .A1(n19558), .A2(n19981), .B1(n19980), .B2(n19557), .ZN(
        n19549) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19559), .B1(
        n19589), .B2(n19983), .ZN(n19548) );
  OAI211_X1 U22502 ( .C1(n19795), .C2(n19562), .A(n19549), .B(n19548), .ZN(
        P2_U3067) );
  AOI22_X1 U22503 ( .A1(n19558), .A2(n19988), .B1(n19987), .B2(n19557), .ZN(
        n19551) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19559), .B1(
        n19589), .B2(n19990), .ZN(n19550) );
  OAI211_X1 U22505 ( .C1(n19898), .C2(n19562), .A(n19551), .B(n19550), .ZN(
        P2_U3068) );
  AOI22_X1 U22506 ( .A1(n19558), .A2(n19995), .B1(n19994), .B2(n19557), .ZN(
        n19553) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19559), .B1(
        n19554), .B2(n19997), .ZN(n19552) );
  OAI211_X1 U22508 ( .C1(n19864), .C2(n19597), .A(n19553), .B(n19552), .ZN(
        P2_U3069) );
  AOI22_X1 U22509 ( .A1(n19558), .A2(n20002), .B1(n20001), .B2(n19557), .ZN(
        n19556) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19559), .B1(
        n19554), .B2(n20004), .ZN(n19555) );
  OAI211_X1 U22511 ( .C1(n19835), .C2(n19597), .A(n19556), .B(n19555), .ZN(
        P2_U3070) );
  AOI22_X1 U22512 ( .A1(n19558), .A2(n20010), .B1(n20008), .B2(n19557), .ZN(
        n19561) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19559), .B1(
        n19589), .B2(n20014), .ZN(n19560) );
  OAI211_X1 U22514 ( .C1(n19842), .C2(n19562), .A(n19561), .B(n19560), .ZN(
        P2_U3071) );
  OAI21_X1 U22515 ( .B1(n19693), .B2(n20103), .A(n20102), .ZN(n19573) );
  NAND2_X1 U22516 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19563), .ZN(
        n19572) );
  INV_X1 U22517 ( .A(n19572), .ZN(n19564) );
  OR2_X1 U22518 ( .A1(n19573), .A2(n19564), .ZN(n19569) );
  OAI21_X1 U22519 ( .B1(n19570), .B2(n20132), .A(n20110), .ZN(n19567) );
  NOR2_X1 U22520 ( .A1(n19565), .A2(n19809), .ZN(n19592) );
  INV_X1 U22521 ( .A(n19592), .ZN(n19566) );
  AOI21_X1 U22522 ( .B1(n19567), .B2(n19566), .A(n19917), .ZN(n19568) );
  INV_X1 U22523 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19576) );
  AOI22_X1 U22524 ( .A1(n19963), .A2(n19621), .B1(n19592), .B2(n19960), .ZN(
        n19575) );
  OAI21_X1 U22525 ( .B1(n19570), .B2(n19592), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19571) );
  OAI21_X1 U22526 ( .B1(n19573), .B2(n19572), .A(n19571), .ZN(n19593) );
  AOI22_X1 U22527 ( .A1(n19961), .A2(n19593), .B1(n19589), .B2(n19962), .ZN(
        n19574) );
  OAI211_X1 U22528 ( .C1(n19582), .C2(n19576), .A(n19575), .B(n19574), .ZN(
        P2_U3072) );
  AOI22_X1 U22529 ( .A1(n19969), .A2(n19589), .B1(n19967), .B2(n19592), .ZN(
        n19578) );
  AOI22_X1 U22530 ( .A1(n19968), .A2(n19593), .B1(n19621), .B2(n19970), .ZN(
        n19577) );
  OAI211_X1 U22531 ( .C1(n19582), .C2(n11732), .A(n19578), .B(n19577), .ZN(
        P2_U3073) );
  INV_X1 U22532 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19581) );
  AOI22_X1 U22533 ( .A1(n19976), .A2(n19589), .B1(n19592), .B2(n19974), .ZN(
        n19580) );
  AOI22_X1 U22534 ( .A1(n19469), .A2(n19593), .B1(n19621), .B2(n19975), .ZN(
        n19579) );
  OAI211_X1 U22535 ( .C1(n19582), .C2(n19581), .A(n19580), .B(n19579), .ZN(
        P2_U3074) );
  AOI22_X1 U22536 ( .A1(n19983), .A2(n19621), .B1(n19592), .B2(n19980), .ZN(
        n19584) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19594), .B1(
        n19981), .B2(n19593), .ZN(n19583) );
  OAI211_X1 U22538 ( .C1(n19795), .C2(n19597), .A(n19584), .B(n19583), .ZN(
        P2_U3075) );
  AOI22_X1 U22539 ( .A1(n19990), .A2(n19621), .B1(n19592), .B2(n19987), .ZN(
        n19586) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19594), .B1(
        n19988), .B2(n19593), .ZN(n19585) );
  OAI211_X1 U22541 ( .C1(n19898), .C2(n19597), .A(n19586), .B(n19585), .ZN(
        P2_U3076) );
  AOI22_X1 U22542 ( .A1(n19996), .A2(n19621), .B1(n19994), .B2(n19592), .ZN(
        n19588) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19594), .B1(
        n19995), .B2(n19593), .ZN(n19587) );
  OAI211_X1 U22544 ( .C1(n19901), .C2(n19597), .A(n19588), .B(n19587), .ZN(
        P2_U3077) );
  AOI22_X1 U22545 ( .A1(n20004), .A2(n19589), .B1(n19592), .B2(n20001), .ZN(
        n19591) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19594), .B1(
        n20002), .B2(n19593), .ZN(n19590) );
  OAI211_X1 U22547 ( .C1(n19835), .C2(n19629), .A(n19591), .B(n19590), .ZN(
        P2_U3078) );
  AOI22_X1 U22548 ( .A1(n20014), .A2(n19621), .B1(n19592), .B2(n20008), .ZN(
        n19596) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19594), .B1(
        n20010), .B2(n19593), .ZN(n19595) );
  OAI211_X1 U22550 ( .C1(n19842), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3079) );
  INV_X1 U22551 ( .A(n19598), .ZN(n19663) );
  NAND2_X1 U22552 ( .A1(n19663), .A2(n19599), .ZN(n19849) );
  NOR2_X1 U22553 ( .A1(n19849), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19608) );
  INV_X1 U22554 ( .A(n19608), .ZN(n19601) );
  NAND2_X1 U22555 ( .A1(n20114), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19689) );
  NOR2_X1 U22556 ( .A1(n19719), .A2(n19689), .ZN(n19624) );
  OAI21_X1 U22557 ( .B1(n19603), .B2(n19624), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19600) );
  OAI21_X1 U22558 ( .B1(n19958), .B2(n19601), .A(n19600), .ZN(n19625) );
  AOI22_X1 U22559 ( .A1(n19625), .A2(n19961), .B1(n19960), .B2(n19624), .ZN(
        n19610) );
  INV_X1 U22560 ( .A(n19882), .ZN(n19602) );
  AOI21_X1 U22561 ( .B1(n19629), .B2(n19658), .A(n20153), .ZN(n19607) );
  OAI21_X1 U22562 ( .B1(n19603), .B2(n20132), .A(n20110), .ZN(n19605) );
  INV_X1 U22563 ( .A(n19624), .ZN(n19604) );
  NAND2_X1 U22564 ( .A1(n19605), .A2(n19604), .ZN(n19606) );
  OAI211_X1 U22565 ( .C1(n19608), .C2(n19607), .A(n19606), .B(n19952), .ZN(
        n19626) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19963), .ZN(n19609) );
  OAI211_X1 U22567 ( .C1(n19886), .C2(n19629), .A(n19610), .B(n19609), .ZN(
        P2_U3080) );
  AOI22_X1 U22568 ( .A1(n19625), .A2(n19968), .B1(n19967), .B2(n19624), .ZN(
        n19612) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19970), .ZN(n19611) );
  OAI211_X1 U22570 ( .C1(n19889), .C2(n19629), .A(n19612), .B(n19611), .ZN(
        P2_U3081) );
  AOI22_X1 U22571 ( .A1(n19625), .A2(n19469), .B1(n19974), .B2(n19624), .ZN(
        n19614) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19626), .B1(
        n19621), .B2(n19976), .ZN(n19613) );
  OAI211_X1 U22573 ( .C1(n19892), .C2(n19658), .A(n19614), .B(n19613), .ZN(
        P2_U3082) );
  AOI22_X1 U22574 ( .A1(n19625), .A2(n19981), .B1(n19980), .B2(n19624), .ZN(
        n19616) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19983), .ZN(n19615) );
  OAI211_X1 U22576 ( .C1(n19795), .C2(n19629), .A(n19616), .B(n19615), .ZN(
        P2_U3083) );
  AOI22_X1 U22577 ( .A1(n19625), .A2(n19988), .B1(n19987), .B2(n19624), .ZN(
        n19618) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19990), .ZN(n19617) );
  OAI211_X1 U22579 ( .C1(n19898), .C2(n19629), .A(n19618), .B(n19617), .ZN(
        P2_U3084) );
  AOI22_X1 U22580 ( .A1(n19625), .A2(n19995), .B1(n19994), .B2(n19624), .ZN(
        n19620) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n19996), .ZN(n19619) );
  OAI211_X1 U22582 ( .C1(n19901), .C2(n19629), .A(n19620), .B(n19619), .ZN(
        P2_U3085) );
  AOI22_X1 U22583 ( .A1(n19625), .A2(n20002), .B1(n20001), .B2(n19624), .ZN(
        n19623) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19626), .B1(
        n19621), .B2(n20004), .ZN(n19622) );
  OAI211_X1 U22585 ( .C1(n19835), .C2(n19658), .A(n19623), .B(n19622), .ZN(
        P2_U3086) );
  AOI22_X1 U22586 ( .A1(n19625), .A2(n20010), .B1(n20008), .B2(n19624), .ZN(
        n19628) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19626), .B1(
        n19650), .B2(n20014), .ZN(n19627) );
  OAI211_X1 U22588 ( .C1(n19842), .C2(n19629), .A(n19628), .B(n19627), .ZN(
        P2_U3087) );
  NOR2_X1 U22589 ( .A1(n19689), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19633) );
  INV_X1 U22590 ( .A(n19633), .ZN(n19636) );
  NOR2_X1 U22591 ( .A1(n21258), .A2(n19636), .ZN(n19653) );
  AOI22_X1 U22592 ( .A1(n19963), .A2(n19680), .B1(n19960), .B2(n19653), .ZN(
        n19639) );
  OAI21_X1 U22593 ( .B1(n19693), .B2(n19882), .A(n20102), .ZN(n19637) );
  OAI21_X1 U22594 ( .B1(n19634), .B2(n20132), .A(n20110), .ZN(n19631) );
  INV_X1 U22595 ( .A(n19653), .ZN(n19630) );
  AOI21_X1 U22596 ( .B1(n19631), .B2(n19630), .A(n19917), .ZN(n19632) );
  OAI21_X1 U22597 ( .B1(n19637), .B2(n19633), .A(n19632), .ZN(n19655) );
  OAI21_X1 U22598 ( .B1(n19634), .B2(n19653), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19635) );
  OAI21_X1 U22599 ( .B1(n19637), .B2(n19636), .A(n19635), .ZN(n19654) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19655), .B1(
        n19961), .B2(n19654), .ZN(n19638) );
  OAI211_X1 U22601 ( .C1(n19886), .C2(n19658), .A(n19639), .B(n19638), .ZN(
        P2_U3088) );
  AOI22_X1 U22602 ( .A1(n19970), .A2(n19680), .B1(n19967), .B2(n19653), .ZN(
        n19641) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19655), .B1(
        n19968), .B2(n19654), .ZN(n19640) );
  OAI211_X1 U22604 ( .C1(n19889), .C2(n19658), .A(n19641), .B(n19640), .ZN(
        P2_U3089) );
  AOI22_X1 U22605 ( .A1(n19976), .A2(n19650), .B1(n19653), .B2(n19974), .ZN(
        n19643) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19655), .B1(
        n19469), .B2(n19654), .ZN(n19642) );
  OAI211_X1 U22607 ( .C1(n19892), .C2(n19688), .A(n19643), .B(n19642), .ZN(
        P2_U3090) );
  AOI22_X1 U22608 ( .A1(n19983), .A2(n19680), .B1(n19653), .B2(n19980), .ZN(
        n19645) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19655), .B1(
        n19981), .B2(n19654), .ZN(n19644) );
  OAI211_X1 U22610 ( .C1(n19795), .C2(n19658), .A(n19645), .B(n19644), .ZN(
        P2_U3091) );
  AOI22_X1 U22611 ( .A1(n19990), .A2(n19680), .B1(n19653), .B2(n19987), .ZN(
        n19647) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19655), .B1(
        n19988), .B2(n19654), .ZN(n19646) );
  OAI211_X1 U22613 ( .C1(n19898), .C2(n19658), .A(n19647), .B(n19646), .ZN(
        P2_U3092) );
  AOI22_X1 U22614 ( .A1(n19997), .A2(n19650), .B1(n19994), .B2(n19653), .ZN(
        n19649) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19655), .B1(
        n19995), .B2(n19654), .ZN(n19648) );
  OAI211_X1 U22616 ( .C1(n19864), .C2(n19688), .A(n19649), .B(n19648), .ZN(
        P2_U3093) );
  AOI22_X1 U22617 ( .A1(n20004), .A2(n19650), .B1(n19653), .B2(n20001), .ZN(
        n19652) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19655), .B1(
        n20002), .B2(n19654), .ZN(n19651) );
  OAI211_X1 U22619 ( .C1(n19835), .C2(n19688), .A(n19652), .B(n19651), .ZN(
        P2_U3094) );
  AOI22_X1 U22620 ( .A1(n20014), .A2(n19680), .B1(n19653), .B2(n20008), .ZN(
        n19657) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19655), .B1(
        n20010), .B2(n19654), .ZN(n19656) );
  OAI211_X1 U22622 ( .C1(n19842), .C2(n19658), .A(n19657), .B(n19656), .ZN(
        P2_U3095) );
  INV_X1 U22623 ( .A(n11936), .ZN(n19659) );
  NOR3_X2 U22624 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19948), .ZN(n19683) );
  OAI21_X1 U22625 ( .B1(n19659), .B2(n19683), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19660) );
  OAI21_X1 U22626 ( .B1(n19689), .B2(n19781), .A(n19660), .ZN(n19684) );
  AOI22_X1 U22627 ( .A1(n19684), .A2(n19961), .B1(n19960), .B2(n19683), .ZN(
        n19669) );
  AOI21_X1 U22628 ( .B1(n19688), .B2(n19718), .A(n20153), .ZN(n19667) );
  NOR2_X1 U22629 ( .A1(n19663), .A2(n19689), .ZN(n19666) );
  INV_X1 U22630 ( .A(n19683), .ZN(n19664) );
  OAI211_X1 U22631 ( .C1(n11936), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19664), 
        .B(n19958), .ZN(n19665) );
  OAI211_X1 U22632 ( .C1(n19667), .C2(n19666), .A(n19665), .B(n19952), .ZN(
        n19685) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n19963), .ZN(n19668) );
  OAI211_X1 U22634 ( .C1(n19886), .C2(n19688), .A(n19669), .B(n19668), .ZN(
        P2_U3096) );
  AOI22_X1 U22635 ( .A1(n19684), .A2(n19968), .B1(n19967), .B2(n19683), .ZN(
        n19671) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n19970), .ZN(n19670) );
  OAI211_X1 U22637 ( .C1(n19889), .C2(n19688), .A(n19671), .B(n19670), .ZN(
        P2_U3097) );
  AOI22_X1 U22638 ( .A1(n19684), .A2(n19469), .B1(n19974), .B2(n19683), .ZN(
        n19673) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19685), .B1(
        n19680), .B2(n19976), .ZN(n19672) );
  OAI211_X1 U22640 ( .C1(n19892), .C2(n19718), .A(n19673), .B(n19672), .ZN(
        P2_U3098) );
  AOI22_X1 U22641 ( .A1(n19684), .A2(n19981), .B1(n19980), .B2(n19683), .ZN(
        n19675) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n19983), .ZN(n19674) );
  OAI211_X1 U22643 ( .C1(n19795), .C2(n19688), .A(n19675), .B(n19674), .ZN(
        P2_U3099) );
  AOI22_X1 U22644 ( .A1(n19684), .A2(n19988), .B1(n19987), .B2(n19683), .ZN(
        n19677) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n19990), .ZN(n19676) );
  OAI211_X1 U22646 ( .C1(n19898), .C2(n19688), .A(n19677), .B(n19676), .ZN(
        P2_U3100) );
  AOI22_X1 U22647 ( .A1(n19684), .A2(n19995), .B1(n19994), .B2(n19683), .ZN(
        n19679) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n19996), .ZN(n19678) );
  OAI211_X1 U22649 ( .C1(n19901), .C2(n19688), .A(n19679), .B(n19678), .ZN(
        P2_U3101) );
  AOI22_X1 U22650 ( .A1(n19684), .A2(n20002), .B1(n20001), .B2(n19683), .ZN(
        n19682) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19685), .B1(
        n19680), .B2(n20004), .ZN(n19681) );
  OAI211_X1 U22652 ( .C1(n19835), .C2(n19718), .A(n19682), .B(n19681), .ZN(
        P2_U3102) );
  AOI22_X1 U22653 ( .A1(n19684), .A2(n20010), .B1(n20008), .B2(n19683), .ZN(
        n19687) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19685), .B1(
        n19711), .B2(n20014), .ZN(n19686) );
  OAI211_X1 U22655 ( .C1(n19842), .C2(n19688), .A(n19687), .B(n19686), .ZN(
        P2_U3103) );
  NOR2_X1 U22656 ( .A1(n19809), .A2(n19689), .ZN(n19726) );
  NOR2_X1 U22657 ( .A1(n19726), .A2(n20132), .ZN(n19690) );
  NAND2_X1 U22658 ( .A1(n11941), .A2(n19690), .ZN(n19694) );
  NOR2_X1 U22659 ( .A1(n19948), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19697) );
  INV_X1 U22660 ( .A(n19697), .ZN(n19691) );
  OAI21_X1 U22661 ( .B1(n19691), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20132), 
        .ZN(n19692) );
  AND2_X1 U22662 ( .A1(n19694), .A2(n19692), .ZN(n19714) );
  AOI22_X1 U22663 ( .A1(n19714), .A2(n19961), .B1(n19726), .B2(n19960), .ZN(
        n19700) );
  NOR2_X1 U22664 ( .A1(n19693), .A2(n19949), .ZN(n20101) );
  OAI211_X1 U22665 ( .C1(n19726), .C2(n20110), .A(n19694), .B(n19952), .ZN(
        n19695) );
  INV_X1 U22666 ( .A(n19695), .ZN(n19696) );
  OAI21_X1 U22667 ( .B1(n19697), .B2(n20101), .A(n19696), .ZN(n19715) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19715), .B1(
        n19741), .B2(n19963), .ZN(n19699) );
  OAI211_X1 U22669 ( .C1(n19886), .C2(n19718), .A(n19700), .B(n19699), .ZN(
        P2_U3104) );
  AOI22_X1 U22670 ( .A1(n19714), .A2(n19968), .B1(n19967), .B2(n19726), .ZN(
        n19702) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19715), .B1(
        n19711), .B2(n19969), .ZN(n19701) );
  OAI211_X1 U22672 ( .C1(n19823), .C2(n19749), .A(n19702), .B(n19701), .ZN(
        P2_U3105) );
  AOI22_X1 U22673 ( .A1(n19714), .A2(n19469), .B1(n19726), .B2(n19974), .ZN(
        n19704) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19715), .B1(
        n19711), .B2(n19976), .ZN(n19703) );
  OAI211_X1 U22675 ( .C1(n19892), .C2(n19749), .A(n19704), .B(n19703), .ZN(
        P2_U3106) );
  AOI22_X1 U22676 ( .A1(n19714), .A2(n19981), .B1(n19726), .B2(n19980), .ZN(
        n19706) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19715), .B1(
        n19711), .B2(n19982), .ZN(n19705) );
  OAI211_X1 U22678 ( .C1(n19895), .C2(n19749), .A(n19706), .B(n19705), .ZN(
        P2_U3107) );
  AOI22_X1 U22679 ( .A1(n19714), .A2(n19988), .B1(n19726), .B2(n19987), .ZN(
        n19708) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19715), .B1(
        n19741), .B2(n19990), .ZN(n19707) );
  OAI211_X1 U22681 ( .C1(n19898), .C2(n19718), .A(n19708), .B(n19707), .ZN(
        P2_U3108) );
  AOI22_X1 U22682 ( .A1(n19714), .A2(n19995), .B1(n19994), .B2(n19726), .ZN(
        n19710) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19715), .B1(
        n19711), .B2(n19997), .ZN(n19709) );
  OAI211_X1 U22684 ( .C1(n19864), .C2(n19749), .A(n19710), .B(n19709), .ZN(
        P2_U3109) );
  AOI22_X1 U22685 ( .A1(n19714), .A2(n20002), .B1(n19726), .B2(n20001), .ZN(
        n19713) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19715), .B1(
        n19711), .B2(n20004), .ZN(n19712) );
  OAI211_X1 U22687 ( .C1(n19835), .C2(n19749), .A(n19713), .B(n19712), .ZN(
        P2_U3110) );
  AOI22_X1 U22688 ( .A1(n19714), .A2(n20010), .B1(n19726), .B2(n20008), .ZN(
        n19717) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19715), .B1(
        n19741), .B2(n20014), .ZN(n19716) );
  OAI211_X1 U22690 ( .C1(n19842), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3111) );
  NAND2_X1 U22691 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20121), .ZN(
        n19812) );
  NOR2_X1 U22692 ( .A1(n19719), .A2(n19812), .ZN(n19744) );
  AOI22_X1 U22693 ( .A1(n19963), .A2(n19774), .B1(n19960), .B2(n19744), .ZN(
        n19730) );
  AOI21_X1 U22694 ( .B1(n19749), .B2(n19773), .A(n20153), .ZN(n19720) );
  NOR2_X1 U22695 ( .A1(n19720), .A2(n19958), .ZN(n19725) );
  INV_X1 U22696 ( .A(n19726), .ZN(n19723) );
  AOI21_X1 U22697 ( .B1(n10121), .B2(n20110), .A(n20102), .ZN(n19722) );
  AOI21_X1 U22698 ( .B1(n19725), .B2(n19723), .A(n19722), .ZN(n19724) );
  OAI21_X1 U22699 ( .B1(n19744), .B2(n19724), .A(n19952), .ZN(n19746) );
  OAI21_X1 U22700 ( .B1(n19726), .B2(n19744), .A(n19725), .ZN(n19728) );
  OAI21_X1 U22701 ( .B1(n10121), .B2(n19744), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19727) );
  NAND2_X1 U22702 ( .A1(n19728), .A2(n19727), .ZN(n19745) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19746), .B1(
        n19961), .B2(n19745), .ZN(n19729) );
  OAI211_X1 U22704 ( .C1(n19886), .C2(n19749), .A(n19730), .B(n19729), .ZN(
        P2_U3112) );
  AOI22_X1 U22705 ( .A1(n19970), .A2(n19774), .B1(n19967), .B2(n19744), .ZN(
        n19732) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19968), .ZN(n19731) );
  OAI211_X1 U22707 ( .C1(n19889), .C2(n19749), .A(n19732), .B(n19731), .ZN(
        P2_U3113) );
  AOI22_X1 U22708 ( .A1(n19976), .A2(n19741), .B1(n19974), .B2(n19744), .ZN(
        n19734) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19469), .ZN(n19733) );
  OAI211_X1 U22710 ( .C1(n19892), .C2(n19773), .A(n19734), .B(n19733), .ZN(
        P2_U3114) );
  AOI22_X1 U22711 ( .A1(n19983), .A2(n19774), .B1(n19980), .B2(n19744), .ZN(
        n19736) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19981), .ZN(n19735) );
  OAI211_X1 U22713 ( .C1(n19795), .C2(n19749), .A(n19736), .B(n19735), .ZN(
        P2_U3115) );
  AOI22_X1 U22714 ( .A1(n19990), .A2(n19774), .B1(n19987), .B2(n19744), .ZN(
        n19738) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19988), .ZN(n19737) );
  OAI211_X1 U22716 ( .C1(n19898), .C2(n19749), .A(n19738), .B(n19737), .ZN(
        P2_U3116) );
  AOI22_X1 U22717 ( .A1(n19997), .A2(n19741), .B1(n19994), .B2(n19744), .ZN(
        n19740) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19995), .ZN(n19739) );
  OAI211_X1 U22719 ( .C1(n19864), .C2(n19773), .A(n19740), .B(n19739), .ZN(
        P2_U3117) );
  AOI22_X1 U22720 ( .A1(n20004), .A2(n19741), .B1(n19744), .B2(n20001), .ZN(
        n19743) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20002), .ZN(n19742) );
  OAI211_X1 U22722 ( .C1(n19835), .C2(n19773), .A(n19743), .B(n19742), .ZN(
        P2_U3118) );
  AOI22_X1 U22723 ( .A1(n20014), .A2(n19774), .B1(n20008), .B2(n19744), .ZN(
        n19748) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20010), .ZN(n19747) );
  OAI211_X1 U22725 ( .C1(n19842), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P2_U3119) );
  NOR3_X2 U22726 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21258), .A3(
        n19812), .ZN(n19782) );
  AOI22_X1 U22727 ( .A1(n19962), .A2(n19774), .B1(n19960), .B2(n19782), .ZN(
        n19760) );
  NAND2_X1 U22728 ( .A1(n20106), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19950) );
  OAI21_X1 U22729 ( .B1(n19950), .B2(n19750), .A(n20102), .ZN(n19758) );
  NOR2_X1 U22730 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19812), .ZN(
        n19753) );
  INV_X1 U22731 ( .A(n19782), .ZN(n19751) );
  OAI211_X1 U22732 ( .C1(n19754), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19751), 
        .B(n19958), .ZN(n19752) );
  OAI211_X1 U22733 ( .C1(n19758), .C2(n19753), .A(n19952), .B(n19752), .ZN(
        n19776) );
  INV_X1 U22734 ( .A(n19753), .ZN(n19757) );
  INV_X1 U22735 ( .A(n19754), .ZN(n19755) );
  OAI21_X1 U22736 ( .B1(n19755), .B2(n19782), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19756) );
  OAI21_X1 U22737 ( .B1(n19758), .B2(n19757), .A(n19756), .ZN(n19775) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19776), .B1(
        n19961), .B2(n19775), .ZN(n19759) );
  OAI211_X1 U22739 ( .C1(n19820), .C2(n19808), .A(n19760), .B(n19759), .ZN(
        P2_U3120) );
  AOI22_X1 U22740 ( .A1(n19969), .A2(n19774), .B1(n19967), .B2(n19782), .ZN(
        n19762) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19776), .B1(
        n19968), .B2(n19775), .ZN(n19761) );
  OAI211_X1 U22742 ( .C1(n19823), .C2(n19808), .A(n19762), .B(n19761), .ZN(
        P2_U3121) );
  AOI22_X1 U22743 ( .A1(n19976), .A2(n19774), .B1(n19974), .B2(n19782), .ZN(
        n19764) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19776), .B1(
        n19469), .B2(n19775), .ZN(n19763) );
  OAI211_X1 U22745 ( .C1(n19892), .C2(n19808), .A(n19764), .B(n19763), .ZN(
        P2_U3122) );
  AOI22_X1 U22746 ( .A1(n19982), .A2(n19774), .B1(n19980), .B2(n19782), .ZN(
        n19766) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19776), .B1(
        n19981), .B2(n19775), .ZN(n19765) );
  OAI211_X1 U22748 ( .C1(n19895), .C2(n19808), .A(n19766), .B(n19765), .ZN(
        P2_U3123) );
  AOI22_X1 U22749 ( .A1(n19990), .A2(n19800), .B1(n19987), .B2(n19782), .ZN(
        n19768) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19776), .B1(
        n19988), .B2(n19775), .ZN(n19767) );
  OAI211_X1 U22751 ( .C1(n19898), .C2(n19773), .A(n19768), .B(n19767), .ZN(
        P2_U3124) );
  AOI22_X1 U22752 ( .A1(n19996), .A2(n19800), .B1(n19994), .B2(n19782), .ZN(
        n19770) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19776), .B1(
        n19995), .B2(n19775), .ZN(n19769) );
  OAI211_X1 U22754 ( .C1(n19901), .C2(n19773), .A(n19770), .B(n19769), .ZN(
        P2_U3125) );
  AOI22_X1 U22755 ( .A1(n20003), .A2(n19800), .B1(n20001), .B2(n19782), .ZN(
        n19772) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19776), .B1(
        n20002), .B2(n19775), .ZN(n19771) );
  OAI211_X1 U22757 ( .C1(n19905), .C2(n19773), .A(n19772), .B(n19771), .ZN(
        P2_U3126) );
  AOI22_X1 U22758 ( .A1(n20012), .A2(n19774), .B1(n20008), .B2(n19782), .ZN(
        n19778) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19776), .B1(
        n20010), .B2(n19775), .ZN(n19777) );
  OAI211_X1 U22760 ( .C1(n19911), .C2(n19808), .A(n19778), .B(n19777), .ZN(
        P2_U3127) );
  INV_X1 U22761 ( .A(n19783), .ZN(n19779) );
  NOR3_X2 U22762 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11863), .A3(
        n19812), .ZN(n19803) );
  OAI21_X1 U22763 ( .B1(n19779), .B2(n19803), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19780) );
  OAI21_X1 U22764 ( .B1(n19812), .B2(n19781), .A(n19780), .ZN(n19804) );
  AOI22_X1 U22765 ( .A1(n19804), .A2(n19961), .B1(n19960), .B2(n19803), .ZN(
        n19788) );
  AOI221_X1 U22766 ( .B1(n19800), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19832), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19782), .ZN(n19784) );
  MUX2_X1 U22767 ( .A(n19784), .B(n19783), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19785) );
  NOR2_X1 U22768 ( .A1(n19785), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19786) );
  OAI21_X1 U22769 ( .B1(n19786), .B2(n19803), .A(n19952), .ZN(n19805) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19805), .B1(
        n19832), .B2(n19963), .ZN(n19787) );
  OAI211_X1 U22771 ( .C1(n19886), .C2(n19808), .A(n19788), .B(n19787), .ZN(
        P2_U3128) );
  AOI22_X1 U22772 ( .A1(n19804), .A2(n19968), .B1(n19967), .B2(n19803), .ZN(
        n19790) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19805), .B1(
        n19832), .B2(n19970), .ZN(n19789) );
  OAI211_X1 U22774 ( .C1(n19889), .C2(n19808), .A(n19790), .B(n19789), .ZN(
        P2_U3129) );
  INV_X1 U22775 ( .A(n19832), .ZN(n19841) );
  AOI22_X1 U22776 ( .A1(n19804), .A2(n19469), .B1(n19974), .B2(n19803), .ZN(
        n19792) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19805), .B1(
        n19800), .B2(n19976), .ZN(n19791) );
  OAI211_X1 U22778 ( .C1(n19892), .C2(n19841), .A(n19792), .B(n19791), .ZN(
        P2_U3130) );
  AOI22_X1 U22779 ( .A1(n19804), .A2(n19981), .B1(n19980), .B2(n19803), .ZN(
        n19794) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19805), .B1(
        n19832), .B2(n19983), .ZN(n19793) );
  OAI211_X1 U22781 ( .C1(n19795), .C2(n19808), .A(n19794), .B(n19793), .ZN(
        P2_U3131) );
  AOI22_X1 U22782 ( .A1(n19804), .A2(n19988), .B1(n19987), .B2(n19803), .ZN(
        n19797) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19805), .B1(
        n19832), .B2(n19990), .ZN(n19796) );
  OAI211_X1 U22784 ( .C1(n19898), .C2(n19808), .A(n19797), .B(n19796), .ZN(
        P2_U3132) );
  AOI22_X1 U22785 ( .A1(n19804), .A2(n19995), .B1(n19994), .B2(n19803), .ZN(
        n19799) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19805), .B1(
        n19800), .B2(n19997), .ZN(n19798) );
  OAI211_X1 U22787 ( .C1(n19864), .C2(n19841), .A(n19799), .B(n19798), .ZN(
        P2_U3133) );
  AOI22_X1 U22788 ( .A1(n19804), .A2(n20002), .B1(n20001), .B2(n19803), .ZN(
        n19802) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19805), .B1(
        n19800), .B2(n20004), .ZN(n19801) );
  OAI211_X1 U22790 ( .C1(n19835), .C2(n19841), .A(n19802), .B(n19801), .ZN(
        P2_U3134) );
  AOI22_X1 U22791 ( .A1(n19804), .A2(n20010), .B1(n20008), .B2(n19803), .ZN(
        n19807) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19805), .B1(
        n19832), .B2(n20014), .ZN(n19806) );
  OAI211_X1 U22793 ( .C1(n19842), .C2(n19808), .A(n19807), .B(n19806), .ZN(
        P2_U3135) );
  INV_X1 U22794 ( .A(n19870), .ZN(n19867) );
  NOR2_X1 U22795 ( .A1(n19809), .A2(n19812), .ZN(n19836) );
  NOR2_X1 U22796 ( .A1(n19836), .A2(n20132), .ZN(n19810) );
  NAND2_X1 U22797 ( .A1(n19811), .A2(n19810), .ZN(n19815) );
  OR2_X1 U22798 ( .A1(n11863), .A2(n19812), .ZN(n19814) );
  OAI21_X1 U22799 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19814), .A(n20132), 
        .ZN(n19813) );
  AOI22_X1 U22800 ( .A1(n19837), .A2(n19961), .B1(n19960), .B2(n19836), .ZN(
        n19819) );
  OAI21_X1 U22801 ( .B1(n19950), .B2(n20103), .A(n19814), .ZN(n19816) );
  AND2_X1 U22802 ( .A1(n19816), .A2(n19815), .ZN(n19817) );
  OAI211_X1 U22803 ( .C1(n19836), .C2(n20110), .A(n19952), .B(n19817), .ZN(
        n19838) );
  AOI22_X1 U22804 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19838), .B1(
        n19832), .B2(n19962), .ZN(n19818) );
  OAI211_X1 U22805 ( .C1(n19820), .C2(n19867), .A(n19819), .B(n19818), .ZN(
        P2_U3136) );
  AOI22_X1 U22806 ( .A1(n19837), .A2(n19968), .B1(n19967), .B2(n19836), .ZN(
        n19822) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19838), .B1(
        n19832), .B2(n19969), .ZN(n19821) );
  OAI211_X1 U22808 ( .C1(n19823), .C2(n19867), .A(n19822), .B(n19821), .ZN(
        P2_U3137) );
  AOI22_X1 U22809 ( .A1(n19837), .A2(n19469), .B1(n19974), .B2(n19836), .ZN(
        n19825) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19838), .B1(
        n19832), .B2(n19976), .ZN(n19824) );
  OAI211_X1 U22811 ( .C1(n19892), .C2(n19867), .A(n19825), .B(n19824), .ZN(
        P2_U3138) );
  AOI22_X1 U22812 ( .A1(n19837), .A2(n19981), .B1(n19980), .B2(n19836), .ZN(
        n19827) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19838), .B1(
        n19832), .B2(n19982), .ZN(n19826) );
  OAI211_X1 U22814 ( .C1(n19895), .C2(n19867), .A(n19827), .B(n19826), .ZN(
        P2_U3139) );
  AOI22_X1 U22815 ( .A1(n19837), .A2(n19988), .B1(n19987), .B2(n19836), .ZN(
        n19829) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19838), .B1(
        n19870), .B2(n19990), .ZN(n19828) );
  OAI211_X1 U22817 ( .C1(n19898), .C2(n19841), .A(n19829), .B(n19828), .ZN(
        P2_U3140) );
  AOI22_X1 U22818 ( .A1(n19837), .A2(n19995), .B1(n19994), .B2(n19836), .ZN(
        n19831) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19838), .B1(
        n19870), .B2(n19996), .ZN(n19830) );
  OAI211_X1 U22820 ( .C1(n19901), .C2(n19841), .A(n19831), .B(n19830), .ZN(
        P2_U3141) );
  AOI22_X1 U22821 ( .A1(n19837), .A2(n20002), .B1(n20001), .B2(n19836), .ZN(
        n19834) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19838), .B1(
        n19832), .B2(n20004), .ZN(n19833) );
  OAI211_X1 U22823 ( .C1(n19835), .C2(n19867), .A(n19834), .B(n19833), .ZN(
        P2_U3142) );
  AOI22_X1 U22824 ( .A1(n19837), .A2(n20010), .B1(n20008), .B2(n19836), .ZN(
        n19840) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19838), .B1(
        n19870), .B2(n20014), .ZN(n19839) );
  OAI211_X1 U22826 ( .C1(n19842), .C2(n19841), .A(n19840), .B(n19839), .ZN(
        P2_U3143) );
  INV_X1 U22827 ( .A(n19843), .ZN(n19846) );
  INV_X1 U22828 ( .A(n19847), .ZN(n19844) );
  NAND3_X1 U22829 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n11863), .ZN(n19878) );
  NOR2_X1 U22830 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19878), .ZN(
        n19868) );
  OAI21_X1 U22831 ( .B1(n19844), .B2(n19868), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19845) );
  OAI21_X1 U22832 ( .B1(n19846), .B2(n19849), .A(n19845), .ZN(n19869) );
  AOI22_X1 U22833 ( .A1(n19869), .A2(n19961), .B1(n19960), .B2(n19868), .ZN(
        n19853) );
  AOI21_X1 U22834 ( .B1(n19847), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19851) );
  OAI21_X1 U22835 ( .B1(n19907), .B2(n19870), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19848) );
  OAI21_X1 U22836 ( .B1(n19849), .B2(n20114), .A(n19848), .ZN(n19850) );
  OAI211_X1 U22837 ( .C1(n19868), .C2(n19851), .A(n19850), .B(n19952), .ZN(
        n19871) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19871), .B1(
        n19907), .B2(n19963), .ZN(n19852) );
  OAI211_X1 U22839 ( .C1(n19886), .C2(n19867), .A(n19853), .B(n19852), .ZN(
        P2_U3144) );
  AOI22_X1 U22840 ( .A1(n19869), .A2(n19968), .B1(n19967), .B2(n19868), .ZN(
        n19855) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19871), .B1(
        n19907), .B2(n19970), .ZN(n19854) );
  OAI211_X1 U22842 ( .C1(n19889), .C2(n19867), .A(n19855), .B(n19854), .ZN(
        P2_U3145) );
  AOI22_X1 U22843 ( .A1(n19869), .A2(n19469), .B1(n19974), .B2(n19868), .ZN(
        n19857) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19871), .B1(
        n19870), .B2(n19976), .ZN(n19856) );
  OAI211_X1 U22845 ( .C1(n19892), .C2(n19904), .A(n19857), .B(n19856), .ZN(
        P2_U3146) );
  AOI22_X1 U22846 ( .A1(n19869), .A2(n19981), .B1(n19980), .B2(n19868), .ZN(
        n19859) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19871), .B1(
        n19870), .B2(n19982), .ZN(n19858) );
  OAI211_X1 U22848 ( .C1(n19895), .C2(n19904), .A(n19859), .B(n19858), .ZN(
        P2_U3147) );
  AOI22_X1 U22849 ( .A1(n19869), .A2(n19988), .B1(n19987), .B2(n19868), .ZN(
        n19861) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19871), .B1(
        n19907), .B2(n19990), .ZN(n19860) );
  OAI211_X1 U22851 ( .C1(n19898), .C2(n19867), .A(n19861), .B(n19860), .ZN(
        P2_U3148) );
  AOI22_X1 U22852 ( .A1(n19869), .A2(n19995), .B1(n19994), .B2(n19868), .ZN(
        n19863) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19871), .B1(
        n19870), .B2(n19997), .ZN(n19862) );
  OAI211_X1 U22854 ( .C1(n19864), .C2(n19904), .A(n19863), .B(n19862), .ZN(
        P2_U3149) );
  AOI22_X1 U22855 ( .A1(n19869), .A2(n20002), .B1(n20001), .B2(n19868), .ZN(
        n19866) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19871), .B1(
        n19907), .B2(n20003), .ZN(n19865) );
  OAI211_X1 U22857 ( .C1(n19905), .C2(n19867), .A(n19866), .B(n19865), .ZN(
        P2_U3150) );
  AOI22_X1 U22858 ( .A1(n19869), .A2(n20010), .B1(n20008), .B2(n19868), .ZN(
        n19873) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19871), .B1(
        n19870), .B2(n20012), .ZN(n19872) );
  OAI211_X1 U22860 ( .C1(n19911), .C2(n19904), .A(n19873), .B(n19872), .ZN(
        P2_U3151) );
  NOR2_X1 U22861 ( .A1(n21258), .A2(n19878), .ZN(n19915) );
  INV_X1 U22862 ( .A(n19915), .ZN(n19874) );
  AND2_X1 U22863 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19874), .ZN(n19875) );
  NAND2_X1 U22864 ( .A1(n19876), .A2(n19875), .ZN(n19879) );
  OAI21_X1 U22865 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19878), .A(n20132), 
        .ZN(n19877) );
  AND2_X1 U22866 ( .A1(n19879), .A2(n19877), .ZN(n19906) );
  AOI22_X1 U22867 ( .A1(n19906), .A2(n19961), .B1(n19960), .B2(n19915), .ZN(
        n19885) );
  OAI21_X1 U22868 ( .B1(n19950), .B2(n19882), .A(n19878), .ZN(n19880) );
  AND2_X1 U22869 ( .A1(n19880), .A2(n19879), .ZN(n19881) );
  OAI211_X1 U22870 ( .C1(n19915), .C2(n20110), .A(n19952), .B(n19881), .ZN(
        n19908) );
  AOI22_X1 U22871 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19908), .B1(
        n19942), .B2(n19963), .ZN(n19884) );
  OAI211_X1 U22872 ( .C1(n19886), .C2(n19904), .A(n19885), .B(n19884), .ZN(
        P2_U3152) );
  AOI22_X1 U22873 ( .A1(n19906), .A2(n19968), .B1(n19967), .B2(n19915), .ZN(
        n19888) );
  AOI22_X1 U22874 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19908), .B1(
        n19942), .B2(n19970), .ZN(n19887) );
  OAI211_X1 U22875 ( .C1(n19889), .C2(n19904), .A(n19888), .B(n19887), .ZN(
        P2_U3153) );
  AOI22_X1 U22876 ( .A1(n19906), .A2(n19469), .B1(n19974), .B2(n19915), .ZN(
        n19891) );
  AOI22_X1 U22877 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n19976), .ZN(n19890) );
  OAI211_X1 U22878 ( .C1(n19892), .C2(n19913), .A(n19891), .B(n19890), .ZN(
        P2_U3154) );
  AOI22_X1 U22879 ( .A1(n19906), .A2(n19981), .B1(n19980), .B2(n19915), .ZN(
        n19894) );
  AOI22_X1 U22880 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n19982), .ZN(n19893) );
  OAI211_X1 U22881 ( .C1(n19895), .C2(n19913), .A(n19894), .B(n19893), .ZN(
        P2_U3155) );
  AOI22_X1 U22882 ( .A1(n19906), .A2(n19988), .B1(n19987), .B2(n19915), .ZN(
        n19897) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19908), .B1(
        n19942), .B2(n19990), .ZN(n19896) );
  OAI211_X1 U22884 ( .C1(n19898), .C2(n19904), .A(n19897), .B(n19896), .ZN(
        P2_U3156) );
  AOI22_X1 U22885 ( .A1(n19906), .A2(n19995), .B1(n19994), .B2(n19915), .ZN(
        n19900) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19908), .B1(
        n19942), .B2(n19996), .ZN(n19899) );
  OAI211_X1 U22887 ( .C1(n19901), .C2(n19904), .A(n19900), .B(n19899), .ZN(
        P2_U3157) );
  AOI22_X1 U22888 ( .A1(n19906), .A2(n20002), .B1(n20001), .B2(n19915), .ZN(
        n19903) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19908), .B1(
        n19942), .B2(n20003), .ZN(n19902) );
  OAI211_X1 U22890 ( .C1(n19905), .C2(n19904), .A(n19903), .B(n19902), .ZN(
        P2_U3158) );
  AOI22_X1 U22891 ( .A1(n19906), .A2(n20010), .B1(n20008), .B2(n19915), .ZN(
        n19910) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n20012), .ZN(n19909) );
  OAI211_X1 U22893 ( .C1(n19911), .C2(n19913), .A(n19910), .B(n19909), .ZN(
        P2_U3159) );
  AOI21_X1 U22894 ( .B1(n19919), .B2(n19913), .A(n20153), .ZN(n19914) );
  NOR2_X1 U22895 ( .A1(n19914), .A2(n19958), .ZN(n19920) );
  NOR3_X2 U22896 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20114), .A3(
        n19948), .ZN(n19941) );
  NOR2_X1 U22897 ( .A1(n19941), .A2(n19915), .ZN(n19923) );
  INV_X1 U22898 ( .A(n19916), .ZN(n19921) );
  AOI211_X1 U22899 ( .C1(n19921), .C2(n20110), .A(n19941), .B(n20102), .ZN(
        n19918) );
  INV_X1 U22900 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21446) );
  AOI22_X1 U22901 ( .A1(n19963), .A2(n20013), .B1(n19960), .B2(n19941), .ZN(
        n19926) );
  INV_X1 U22902 ( .A(n19920), .ZN(n19924) );
  OAI21_X1 U22903 ( .B1(n19921), .B2(n19941), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19922) );
  AOI22_X1 U22904 ( .A1(n19961), .A2(n19943), .B1(n19942), .B2(n19962), .ZN(
        n19925) );
  OAI211_X1 U22905 ( .C1(n19947), .C2(n21446), .A(n19926), .B(n19925), .ZN(
        P2_U3160) );
  AOI22_X1 U22906 ( .A1(n19969), .A2(n19942), .B1(n19967), .B2(n19941), .ZN(
        n19928) );
  AOI22_X1 U22907 ( .A1(n19968), .A2(n19943), .B1(n20013), .B2(n19970), .ZN(
        n19927) );
  OAI211_X1 U22908 ( .C1(n19947), .C2(n11718), .A(n19928), .B(n19927), .ZN(
        P2_U3161) );
  INV_X1 U22909 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U22910 ( .A1(n19975), .A2(n20013), .B1(n19974), .B2(n19941), .ZN(
        n19930) );
  AOI22_X1 U22911 ( .A1(n19469), .A2(n19943), .B1(n19942), .B2(n19976), .ZN(
        n19929) );
  OAI211_X1 U22912 ( .C1(n19947), .C2(n19931), .A(n19930), .B(n19929), .ZN(
        P2_U3162) );
  AOI22_X1 U22913 ( .A1(n19983), .A2(n20013), .B1(n19980), .B2(n19941), .ZN(
        n19933) );
  AOI22_X1 U22914 ( .A1(n19981), .A2(n19943), .B1(n19942), .B2(n19982), .ZN(
        n19932) );
  OAI211_X1 U22915 ( .C1(n19947), .C2(n11810), .A(n19933), .B(n19932), .ZN(
        P2_U3163) );
  INV_X1 U22916 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19936) );
  AOI22_X1 U22917 ( .A1(n19989), .A2(n19942), .B1(n19987), .B2(n19941), .ZN(
        n19935) );
  AOI22_X1 U22918 ( .A1(n19988), .A2(n19943), .B1(n20013), .B2(n19990), .ZN(
        n19934) );
  OAI211_X1 U22919 ( .C1(n19947), .C2(n19936), .A(n19935), .B(n19934), .ZN(
        P2_U3164) );
  AOI22_X1 U22920 ( .A1(n19997), .A2(n19942), .B1(n19994), .B2(n19941), .ZN(
        n19938) );
  AOI22_X1 U22921 ( .A1(n19995), .A2(n19943), .B1(n20013), .B2(n19996), .ZN(
        n19937) );
  OAI211_X1 U22922 ( .C1(n19947), .C2(n11932), .A(n19938), .B(n19937), .ZN(
        P2_U3165) );
  AOI22_X1 U22923 ( .A1(n20004), .A2(n19942), .B1(n20001), .B2(n19941), .ZN(
        n19940) );
  AOI22_X1 U22924 ( .A1(n20002), .A2(n19943), .B1(n20013), .B2(n20003), .ZN(
        n19939) );
  OAI211_X1 U22925 ( .C1(n19947), .C2(n11983), .A(n19940), .B(n19939), .ZN(
        P2_U3166) );
  INV_X1 U22926 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19946) );
  AOI22_X1 U22927 ( .A1(n20012), .A2(n19942), .B1(n20008), .B2(n19941), .ZN(
        n19945) );
  AOI22_X1 U22928 ( .A1(n20010), .A2(n19943), .B1(n20013), .B2(n20014), .ZN(
        n19944) );
  OAI211_X1 U22929 ( .C1(n19947), .C2(n19946), .A(n19945), .B(n19944), .ZN(
        P2_U3167) );
  OR2_X1 U22930 ( .A1(n20114), .A2(n19948), .ZN(n19959) );
  OAI21_X1 U22931 ( .B1(n19950), .B2(n19949), .A(n19959), .ZN(n19953) );
  OAI211_X1 U22932 ( .C1(n19954), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19955), 
        .B(n19958), .ZN(n19951) );
  AND3_X1 U22933 ( .A1(n19953), .A2(n19952), .A3(n19951), .ZN(n20019) );
  INV_X1 U22934 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19966) );
  INV_X1 U22935 ( .A(n19954), .ZN(n19956) );
  INV_X1 U22936 ( .A(n19955), .ZN(n20009) );
  OAI21_X1 U22937 ( .B1(n19956), .B2(n20009), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19957) );
  OAI21_X1 U22938 ( .B1(n19959), .B2(n19958), .A(n19957), .ZN(n20011) );
  AOI22_X1 U22939 ( .A1(n20011), .A2(n19961), .B1(n20009), .B2(n19960), .ZN(
        n19965) );
  AOI22_X1 U22940 ( .A1(n20015), .A2(n19963), .B1(n20013), .B2(n19962), .ZN(
        n19964) );
  OAI211_X1 U22941 ( .C1(n20019), .C2(n19966), .A(n19965), .B(n19964), .ZN(
        P2_U3168) );
  AOI22_X1 U22942 ( .A1(n20011), .A2(n19968), .B1(n20009), .B2(n19967), .ZN(
        n19972) );
  AOI22_X1 U22943 ( .A1(n20015), .A2(n19970), .B1(n20013), .B2(n19969), .ZN(
        n19971) );
  OAI211_X1 U22944 ( .C1(n20019), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P2_U3169) );
  INV_X1 U22945 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U22946 ( .A1(n20011), .A2(n19469), .B1(n20009), .B2(n19974), .ZN(
        n19978) );
  AOI22_X1 U22947 ( .A1(n20013), .A2(n19976), .B1(n20015), .B2(n19975), .ZN(
        n19977) );
  OAI211_X1 U22948 ( .C1(n20019), .C2(n19979), .A(n19978), .B(n19977), .ZN(
        P2_U3170) );
  INV_X1 U22949 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U22950 ( .A1(n20011), .A2(n19981), .B1(n20009), .B2(n19980), .ZN(
        n19985) );
  AOI22_X1 U22951 ( .A1(n20015), .A2(n19983), .B1(n20013), .B2(n19982), .ZN(
        n19984) );
  OAI211_X1 U22952 ( .C1(n20019), .C2(n19986), .A(n19985), .B(n19984), .ZN(
        P2_U3171) );
  INV_X1 U22953 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U22954 ( .A1(n20011), .A2(n19988), .B1(n20009), .B2(n19987), .ZN(
        n19992) );
  AOI22_X1 U22955 ( .A1(n20015), .A2(n19990), .B1(n20013), .B2(n19989), .ZN(
        n19991) );
  OAI211_X1 U22956 ( .C1(n20019), .C2(n19993), .A(n19992), .B(n19991), .ZN(
        P2_U3172) );
  INV_X1 U22957 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20000) );
  AOI22_X1 U22958 ( .A1(n20011), .A2(n19995), .B1(n20009), .B2(n19994), .ZN(
        n19999) );
  AOI22_X1 U22959 ( .A1(n20013), .A2(n19997), .B1(n20015), .B2(n19996), .ZN(
        n19998) );
  OAI211_X1 U22960 ( .C1(n20019), .C2(n20000), .A(n19999), .B(n19998), .ZN(
        P2_U3173) );
  AOI22_X1 U22961 ( .A1(n20011), .A2(n20002), .B1(n20009), .B2(n20001), .ZN(
        n20006) );
  AOI22_X1 U22962 ( .A1(n20013), .A2(n20004), .B1(n20015), .B2(n20003), .ZN(
        n20005) );
  OAI211_X1 U22963 ( .C1(n20019), .C2(n20007), .A(n20006), .B(n20005), .ZN(
        P2_U3174) );
  INV_X1 U22964 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U22965 ( .A1(n20011), .A2(n20010), .B1(n20009), .B2(n20008), .ZN(
        n20017) );
  AOI22_X1 U22966 ( .A1(n20015), .A2(n20014), .B1(n20013), .B2(n20012), .ZN(
        n20016) );
  OAI211_X1 U22967 ( .C1(n20019), .C2(n20018), .A(n20017), .B(n20016), .ZN(
        P2_U3175) );
  AOI21_X1 U22968 ( .B1(n20021), .B2(n20020), .A(n20165), .ZN(n20026) );
  OAI211_X1 U22969 ( .C1(n20022), .C2(n20025), .A(n20150), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20023) );
  OAI211_X1 U22970 ( .C1(n20026), .C2(n20025), .A(n20024), .B(n20023), .ZN(
        P2_U3177) );
  AND2_X1 U22971 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20027), .ZN(
        P2_U3179) );
  AND2_X1 U22972 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20027), .ZN(
        P2_U3180) );
  AND2_X1 U22973 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20027), .ZN(
        P2_U3181) );
  AND2_X1 U22974 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20027), .ZN(
        P2_U3182) );
  AND2_X1 U22975 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20027), .ZN(
        P2_U3183) );
  AND2_X1 U22976 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20027), .ZN(
        P2_U3184) );
  AND2_X1 U22977 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20027), .ZN(
        P2_U3185) );
  AND2_X1 U22978 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20027), .ZN(
        P2_U3186) );
  AND2_X1 U22979 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20027), .ZN(
        P2_U3187) );
  AND2_X1 U22980 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20027), .ZN(
        P2_U3188) );
  AND2_X1 U22981 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20027), .ZN(
        P2_U3189) );
  AND2_X1 U22982 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20027), .ZN(
        P2_U3190) );
  AND2_X1 U22983 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20027), .ZN(
        P2_U3191) );
  AND2_X1 U22984 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20027), .ZN(
        P2_U3192) );
  AND2_X1 U22985 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20027), .ZN(
        P2_U3193) );
  AND2_X1 U22986 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20027), .ZN(
        P2_U3194) );
  AND2_X1 U22987 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20027), .ZN(
        P2_U3195) );
  AND2_X1 U22988 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20027), .ZN(
        P2_U3196) );
  AND2_X1 U22989 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20027), .ZN(
        P2_U3197) );
  AND2_X1 U22990 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20027), .ZN(
        P2_U3198) );
  AND2_X1 U22991 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20027), .ZN(
        P2_U3199) );
  AND2_X1 U22992 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20027), .ZN(
        P2_U3200) );
  AND2_X1 U22993 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20027), .ZN(P2_U3201) );
  AND2_X1 U22994 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20027), .ZN(P2_U3202) );
  AND2_X1 U22995 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20027), .ZN(P2_U3203) );
  AND2_X1 U22996 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20027), .ZN(P2_U3204) );
  AND2_X1 U22997 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20027), .ZN(P2_U3205) );
  AND2_X1 U22998 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20027), .ZN(P2_U3206) );
  AND2_X1 U22999 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20027), .ZN(P2_U3207) );
  AND2_X1 U23000 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20027), .ZN(P2_U3208) );
  NAND2_X1 U23001 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20150), .ZN(n20039) );
  NAND3_X1 U23002 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20039), .ZN(n20029) );
  AOI211_X1 U23003 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21050), .A(
        n20038), .B(n20092), .ZN(n20028) );
  INV_X1 U23004 ( .A(NA), .ZN(n21034) );
  NOR2_X1 U23005 ( .A1(n21034), .A2(n20032), .ZN(n20044) );
  AOI211_X1 U23006 ( .C1(n20045), .C2(n20029), .A(n20028), .B(n20044), .ZN(
        n20030) );
  INV_X1 U23007 ( .A(n20030), .ZN(P2_U3209) );
  INV_X1 U23008 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20031) );
  AOI21_X1 U23009 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21050), .A(n20045), 
        .ZN(n20036) );
  NOR2_X1 U23010 ( .A1(n20031), .A2(n20036), .ZN(n20033) );
  AOI21_X1 U23011 ( .B1(n20033), .B2(n20032), .A(n20151), .ZN(n20034) );
  OAI211_X1 U23012 ( .C1(n21050), .C2(n20035), .A(n20034), .B(n20039), .ZN(
        P2_U3210) );
  AOI21_X1 U23013 ( .B1(n20150), .B2(n20037), .A(n20036), .ZN(n20043) );
  INV_X1 U23014 ( .A(n20038), .ZN(n20040) );
  OAI22_X1 U23015 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20040), .B1(NA), 
        .B2(n20039), .ZN(n20041) );
  OAI211_X1 U23016 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20041), .ZN(n20042) );
  OAI21_X1 U23017 ( .B1(n20044), .B2(n20043), .A(n20042), .ZN(P2_U3211) );
  OAI222_X1 U23018 ( .A1(n20094), .A2(n20048), .B1(n20047), .B2(n20092), .C1(
        n20046), .C2(n20091), .ZN(P2_U3212) );
  OAI222_X1 U23019 ( .A1(n20094), .A2(n13639), .B1(n20049), .B2(n20092), .C1(
        n20048), .C2(n20091), .ZN(P2_U3213) );
  OAI222_X1 U23020 ( .A1(n20094), .A2(n20051), .B1(n20050), .B2(n20092), .C1(
        n13639), .C2(n20091), .ZN(P2_U3214) );
  INV_X1 U23021 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20053) );
  OAI222_X1 U23022 ( .A1(n20094), .A2(n20053), .B1(n20052), .B2(n20092), .C1(
        n20051), .C2(n20091), .ZN(P2_U3215) );
  OAI222_X1 U23023 ( .A1(n20094), .A2(n20055), .B1(n20054), .B2(n20092), .C1(
        n20053), .C2(n20091), .ZN(P2_U3216) );
  OAI222_X1 U23024 ( .A1(n20094), .A2(n20057), .B1(n20056), .B2(n20092), .C1(
        n20055), .C2(n20091), .ZN(P2_U3217) );
  OAI222_X1 U23025 ( .A1(n20094), .A2(n20059), .B1(n20058), .B2(n20092), .C1(
        n20057), .C2(n20091), .ZN(P2_U3218) );
  OAI222_X1 U23026 ( .A1(n20094), .A2(n20061), .B1(n20060), .B2(n20092), .C1(
        n20059), .C2(n20091), .ZN(P2_U3219) );
  OAI222_X1 U23027 ( .A1(n20094), .A2(n20063), .B1(n20062), .B2(n20092), .C1(
        n20061), .C2(n20091), .ZN(P2_U3220) );
  OAI222_X1 U23028 ( .A1(n20094), .A2(n15313), .B1(n20064), .B2(n20092), .C1(
        n20063), .C2(n20091), .ZN(P2_U3221) );
  OAI222_X1 U23029 ( .A1(n20094), .A2(n20066), .B1(n20065), .B2(n20092), .C1(
        n15313), .C2(n20091), .ZN(P2_U3222) );
  OAI222_X1 U23030 ( .A1(n20094), .A2(n15288), .B1(n20067), .B2(n20092), .C1(
        n20066), .C2(n20091), .ZN(P2_U3223) );
  INV_X1 U23031 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20069) );
  OAI222_X1 U23032 ( .A1(n20094), .A2(n20069), .B1(n20068), .B2(n20092), .C1(
        n15288), .C2(n20091), .ZN(P2_U3224) );
  OAI222_X1 U23033 ( .A1(n20094), .A2(n15279), .B1(n20070), .B2(n20092), .C1(
        n20069), .C2(n20091), .ZN(P2_U3225) );
  OAI222_X1 U23034 ( .A1(n20094), .A2(n15513), .B1(n20071), .B2(n20092), .C1(
        n15279), .C2(n20091), .ZN(P2_U3226) );
  OAI222_X1 U23035 ( .A1(n20094), .A2(n20073), .B1(n20072), .B2(n20092), .C1(
        n15513), .C2(n20091), .ZN(P2_U3227) );
  OAI222_X1 U23036 ( .A1(n20094), .A2(n20075), .B1(n20074), .B2(n20092), .C1(
        n20073), .C2(n20091), .ZN(P2_U3228) );
  OAI222_X1 U23037 ( .A1(n20094), .A2(n21162), .B1(n20076), .B2(n20092), .C1(
        n20075), .C2(n20091), .ZN(P2_U3229) );
  OAI222_X1 U23038 ( .A1(n20094), .A2(n15225), .B1(n20077), .B2(n20092), .C1(
        n21162), .C2(n20091), .ZN(P2_U3230) );
  OAI222_X1 U23039 ( .A1(n20094), .A2(n12223), .B1(n20078), .B2(n20092), .C1(
        n15225), .C2(n20091), .ZN(P2_U3231) );
  OAI222_X1 U23040 ( .A1(n20094), .A2(n12523), .B1(n20079), .B2(n20092), .C1(
        n12223), .C2(n20091), .ZN(P2_U3232) );
  OAI222_X1 U23041 ( .A1(n20094), .A2(n12232), .B1(n20080), .B2(n20092), .C1(
        n12523), .C2(n20091), .ZN(P2_U3233) );
  OAI222_X1 U23042 ( .A1(n20094), .A2(n20082), .B1(n20081), .B2(n20092), .C1(
        n12232), .C2(n20091), .ZN(P2_U3234) );
  INV_X1 U23043 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21317) );
  OAI222_X1 U23044 ( .A1(n20094), .A2(n21317), .B1(n20083), .B2(n20092), .C1(
        n20082), .C2(n20091), .ZN(P2_U3235) );
  OAI222_X1 U23045 ( .A1(n20094), .A2(n16453), .B1(n20084), .B2(n20092), .C1(
        n21317), .C2(n20091), .ZN(P2_U3236) );
  OAI222_X1 U23046 ( .A1(n20094), .A2(n20087), .B1(n20085), .B2(n20092), .C1(
        n16453), .C2(n20091), .ZN(P2_U3237) );
  INV_X1 U23047 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n21150) );
  OAI222_X1 U23048 ( .A1(n20091), .A2(n20087), .B1(n20086), .B2(n20092), .C1(
        n21150), .C2(n20094), .ZN(P2_U3238) );
  OAI222_X1 U23049 ( .A1(n20094), .A2(n20089), .B1(n20088), .B2(n20092), .C1(
        n21150), .C2(n20091), .ZN(P2_U3239) );
  OAI222_X1 U23050 ( .A1(n20094), .A2(n15138), .B1(n20090), .B2(n20092), .C1(
        n20089), .C2(n20091), .ZN(P2_U3240) );
  OAI222_X1 U23051 ( .A1(n20094), .A2(n20093), .B1(n21261), .B2(n20092), .C1(
        n15138), .C2(n20091), .ZN(P2_U3241) );
  OAI22_X1 U23052 ( .A1(n20168), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20092), .ZN(n20095) );
  INV_X1 U23053 ( .A(n20095), .ZN(P2_U3585) );
  MUX2_X1 U23054 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20168), .Z(P2_U3586) );
  MUX2_X1 U23055 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .B(P2_BE_N_REG_1__SCAN_IN), .S(n20168), .Z(P2_U3587) );
  OAI22_X1 U23056 ( .A1(n20168), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20092), .ZN(n20096) );
  INV_X1 U23057 ( .A(n20096), .ZN(P2_U3588) );
  OAI21_X1 U23058 ( .B1(n20100), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20098), 
        .ZN(n20097) );
  INV_X1 U23059 ( .A(n20097), .ZN(P2_U3591) );
  OAI21_X1 U23060 ( .B1(n20100), .B2(n20099), .A(n20098), .ZN(P2_U3592) );
  INV_X1 U23061 ( .A(n20137), .ZN(n20136) );
  NAND2_X1 U23062 ( .A1(n20101), .A2(n20102), .ZN(n20109) );
  NAND2_X1 U23063 ( .A1(n20102), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20126) );
  OR2_X1 U23064 ( .A1(n20103), .A2(n20126), .ZN(n20115) );
  NAND3_X1 U23065 ( .A1(n20127), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20104), 
        .ZN(n20105) );
  NAND2_X1 U23066 ( .A1(n20105), .A2(n20122), .ZN(n20116) );
  NAND2_X1 U23067 ( .A1(n20115), .A2(n20116), .ZN(n20107) );
  NAND2_X1 U23068 ( .A1(n20107), .A2(n20106), .ZN(n20108) );
  OAI211_X1 U23069 ( .C1(n20111), .C2(n20110), .A(n20109), .B(n20108), .ZN(
        n20112) );
  INV_X1 U23070 ( .A(n20112), .ZN(n20113) );
  AOI22_X1 U23071 ( .A1(n20136), .A2(n20114), .B1(n20113), .B2(n20137), .ZN(
        P2_U3602) );
  OAI21_X1 U23072 ( .B1(n20117), .B2(n20116), .A(n20115), .ZN(n20118) );
  AOI21_X1 U23073 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20119), .A(n20118), 
        .ZN(n20120) );
  AOI22_X1 U23074 ( .A1(n20136), .A2(n20121), .B1(n20120), .B2(n20137), .ZN(
        P2_U3603) );
  INV_X1 U23075 ( .A(n20122), .ZN(n20164) );
  OR3_X1 U23076 ( .A1(n20124), .A2(n20164), .A3(n20123), .ZN(n20125) );
  OAI21_X1 U23077 ( .B1(n20127), .B2(n20126), .A(n20125), .ZN(n20128) );
  AOI21_X1 U23078 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20129), .A(n20128), 
        .ZN(n20130) );
  AOI22_X1 U23079 ( .A1(n20136), .A2(n11863), .B1(n20130), .B2(n20137), .ZN(
        P2_U3604) );
  OAI22_X1 U23080 ( .A1(n20133), .A2(n20164), .B1(n20132), .B2(n20131), .ZN(
        n20134) );
  AOI21_X1 U23081 ( .B1(n21258), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20134), 
        .ZN(n20135) );
  OAI22_X1 U23082 ( .A1(n21258), .A2(n20137), .B1(n20136), .B2(n20135), .ZN(
        P2_U3605) );
  INV_X1 U23083 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20138) );
  AOI22_X1 U23084 ( .A1(n20092), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20138), 
        .B2(n20168), .ZN(P2_U3608) );
  INV_X1 U23085 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20148) );
  AOI22_X1 U23086 ( .A1(n20142), .A2(n20141), .B1(n20140), .B2(n20139), .ZN(
        n20144) );
  NOR2_X1 U23087 ( .A1(n20144), .A2(n20143), .ZN(n20146) );
  OAI21_X1 U23088 ( .B1(n20146), .B2(n20145), .A(n20149), .ZN(n20147) );
  OAI21_X1 U23089 ( .B1(n20149), .B2(n20148), .A(n20147), .ZN(P2_U3609) );
  NOR2_X1 U23090 ( .A1(n20150), .A2(n20132), .ZN(n20160) );
  INV_X1 U23091 ( .A(n20151), .ZN(n20154) );
  OAI21_X1 U23092 ( .B1(n20154), .B2(n20153), .A(n20152), .ZN(n20157) );
  NAND3_X1 U23093 ( .A1(n9812), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20154), 
        .ZN(n20156) );
  MUX2_X1 U23094 ( .A(n20157), .B(n20156), .S(n20155), .Z(n20158) );
  OAI21_X1 U23095 ( .B1(n20160), .B2(n20159), .A(n20158), .ZN(n20167) );
  NAND4_X1 U23096 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .A3(n21322), .A4(n20161), .ZN(n20163) );
  OAI211_X1 U23097 ( .C1(n20165), .C2(n20164), .A(n20163), .B(n20162), .ZN(
        n20166) );
  MUX2_X1 U23098 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n20167), .S(n20166), 
        .Z(P2_U3610) );
  OAI22_X1 U23099 ( .A1(n20168), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20092), .ZN(n20169) );
  INV_X1 U23100 ( .A(n20169), .ZN(P2_U3611) );
  AOI21_X1 U23101 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21051), .A(n21043), 
        .ZN(n21042) );
  INV_X1 U23102 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20170) );
  AOI21_X1 U23103 ( .B1(n21042), .B2(n20170), .A(n21116), .ZN(P1_U2802) );
  NAND2_X1 U23104 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21102), .ZN(n20174) );
  OAI21_X1 U23105 ( .B1(n20172), .B2(n20171), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20173) );
  OAI21_X1 U23106 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20174), .A(n20173), 
        .ZN(P1_U2803) );
  INV_X1 U23107 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n21352) );
  NAND2_X1 U23108 ( .A1(n21051), .A2(n21043), .ZN(n21038) );
  INV_X1 U23109 ( .A(n21038), .ZN(n20176) );
  NOR2_X1 U23110 ( .A1(n21116), .A2(n20176), .ZN(n20175) );
  AOI22_X1 U23111 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n21116), .B1(n21352), 
        .B2(n20175), .ZN(P1_U2804) );
  NOR2_X1 U23112 ( .A1(n21116), .A2(n21042), .ZN(n21099) );
  OAI21_X1 U23113 ( .B1(BS16), .B2(n20176), .A(n21099), .ZN(n21097) );
  OAI21_X1 U23114 ( .B1(n21099), .B2(n20894), .A(n21097), .ZN(P1_U2805) );
  AOI21_X1 U23115 ( .B1(n20177), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20369), .ZN(
        n20178) );
  INV_X1 U23116 ( .A(n20178), .ZN(P1_U2806) );
  NOR4_X1 U23117 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_18__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20182) );
  NOR4_X1 U23118 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20181) );
  NOR4_X1 U23119 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20180) );
  NOR4_X1 U23120 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_22__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_24__SCAN_IN), .ZN(n20179) );
  NAND4_X1 U23121 ( .A1(n20182), .A2(n20181), .A3(n20180), .A4(n20179), .ZN(
        n20188) );
  NOR4_X1 U23122 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20186) );
  AOI211_X1 U23123 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_8__SCAN_IN), .B(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20185) );
  NOR4_X1 U23124 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20184) );
  NOR4_X1 U23125 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20183) );
  NAND4_X1 U23126 ( .A1(n20186), .A2(n20185), .A3(n20184), .A4(n20183), .ZN(
        n20187) );
  NOR2_X1 U23127 ( .A1(n20188), .A2(n20187), .ZN(n21114) );
  INV_X1 U23128 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20190) );
  NOR3_X1 U23129 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20191) );
  OAI21_X1 U23130 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20191), .A(n21114), .ZN(
        n20189) );
  OAI21_X1 U23131 ( .B1(n21114), .B2(n20190), .A(n20189), .ZN(P1_U2807) );
  INV_X1 U23132 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21098) );
  AOI21_X1 U23133 ( .B1(n21107), .B2(n21098), .A(n20191), .ZN(n20193) );
  INV_X1 U23134 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20192) );
  INV_X1 U23135 ( .A(n21114), .ZN(n21109) );
  AOI22_X1 U23136 ( .A1(n21114), .A2(n20193), .B1(n20192), .B2(n21109), .ZN(
        P1_U2808) );
  AOI22_X1 U23137 ( .A1(n20261), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n20257), .B2(
        n20194), .ZN(n20203) );
  AOI22_X1 U23138 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20271), .B1(
        n20260), .B2(n20286), .ZN(n20202) );
  INV_X1 U23139 ( .A(n20195), .ZN(n20199) );
  OAI21_X1 U23140 ( .B1(n20273), .B2(n20197), .A(n20196), .ZN(n20198) );
  AOI22_X1 U23141 ( .A1(n20200), .A2(n20210), .B1(n20199), .B2(n20198), .ZN(
        n20201) );
  NAND4_X1 U23142 ( .A1(n20203), .A2(n20202), .A3(n20201), .A4(n20243), .ZN(
        P1_U2831) );
  OAI21_X1 U23143 ( .B1(n20270), .B2(n20205), .A(n20224), .ZN(n20217) );
  INV_X1 U23144 ( .A(n20204), .ZN(n20293) );
  NOR3_X1 U23145 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20273), .A3(n20205), .ZN(
        n20209) );
  AOI22_X1 U23146 ( .A1(n20261), .A2(P1_EBX_REG_7__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20271), .ZN(n20206) );
  OAI211_X1 U23147 ( .C1(n20285), .C2(n20207), .A(n20206), .B(n20243), .ZN(
        n20208) );
  AOI211_X1 U23148 ( .C1(n20293), .C2(n20260), .A(n20209), .B(n20208), .ZN(
        n20212) );
  NAND2_X1 U23149 ( .A1(n20294), .A2(n20210), .ZN(n20211) );
  OAI211_X1 U23150 ( .C1(n20217), .C2(n21242), .A(n20212), .B(n20211), .ZN(
        P1_U2833) );
  AOI22_X1 U23151 ( .A1(n20213), .A2(n20260), .B1(n20261), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20223) );
  NAND3_X1 U23152 ( .A1(n20236), .A2(n20214), .A3(n21058), .ZN(n20215) );
  OAI211_X1 U23153 ( .C1(n20285), .C2(n20216), .A(n20243), .B(n20215), .ZN(
        n20221) );
  OAI22_X1 U23154 ( .A1(n20219), .A2(n20218), .B1(n21058), .B2(n20217), .ZN(
        n20220) );
  AOI211_X1 U23155 ( .C1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20271), .A(
        n20221), .B(n20220), .ZN(n20222) );
  NAND2_X1 U23156 ( .A1(n20223), .A2(n20222), .ZN(P1_U2834) );
  OAI21_X1 U23157 ( .B1(n20270), .B2(n20235), .A(n20224), .ZN(n20245) );
  AOI22_X1 U23158 ( .A1(n20261), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n20297), .B2(
        n20260), .ZN(n20233) );
  INV_X1 U23159 ( .A(n20235), .ZN(n20225) );
  NAND2_X1 U23160 ( .A1(n20225), .A2(n20234), .ZN(n20230) );
  NAND2_X1 U23161 ( .A1(n20257), .A2(n20226), .ZN(n20228) );
  NAND2_X1 U23162 ( .A1(n20271), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20227) );
  AND3_X1 U23163 ( .A1(n20228), .A2(n20227), .A3(n20243), .ZN(n20229) );
  OAI21_X1 U23164 ( .B1(n20273), .B2(n20230), .A(n20229), .ZN(n20231) );
  AOI21_X1 U23165 ( .B1(n20300), .B2(n20281), .A(n20231), .ZN(n20232) );
  OAI211_X1 U23166 ( .C1(n20245), .C2(n20234), .A(n20233), .B(n20232), .ZN(
        P1_U2835) );
  NAND3_X1 U23167 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20255) );
  NAND2_X1 U23168 ( .A1(n20236), .A2(n20235), .ZN(n20254) );
  INV_X1 U23169 ( .A(n20237), .ZN(n20238) );
  AOI22_X1 U23170 ( .A1(n20261), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20260), .B2(
        n20238), .ZN(n20253) );
  OAI22_X1 U23171 ( .A1(n20242), .A2(n20241), .B1(n20240), .B2(n20239), .ZN(
        n20251) );
  OAI21_X1 U23172 ( .B1(n20285), .B2(n20244), .A(n20243), .ZN(n20250) );
  OAI22_X1 U23173 ( .A1(n20248), .A2(n20247), .B1(n20246), .B2(n20245), .ZN(
        n20249) );
  NOR3_X1 U23174 ( .A1(n20251), .A2(n20250), .A3(n20249), .ZN(n20252) );
  OAI211_X1 U23175 ( .C1(n20255), .C2(n20254), .A(n20253), .B(n20252), .ZN(
        P1_U2836) );
  INV_X1 U23176 ( .A(n20256), .ZN(n20258) );
  AOI222_X1 U23177 ( .A1(n20680), .A2(n20275), .B1(n20258), .B2(n20257), .C1(
        n20271), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20269) );
  AOI22_X1 U23178 ( .A1(n20261), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20260), .B2(
        n20259), .ZN(n20268) );
  AOI22_X1 U23179 ( .A1(n20263), .A2(n20281), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20262), .ZN(n20267) );
  NAND2_X1 U23180 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20264) );
  OAI211_X1 U23181 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20265), .B(n20264), .ZN(n20266) );
  NAND4_X1 U23182 ( .A1(n20269), .A2(n20268), .A3(n20267), .A4(n20266), .ZN(
        P1_U2837) );
  AOI22_X1 U23183 ( .A1(n20271), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20270), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20272) );
  OAI21_X1 U23184 ( .B1(n20273), .B2(P1_REIP_REG_1__SCAN_IN), .A(n20272), .ZN(
        n20274) );
  AOI21_X1 U23185 ( .B1(n20896), .B2(n20275), .A(n20274), .ZN(n20284) );
  OAI22_X1 U23186 ( .A1(n20279), .A2(n20278), .B1(n20277), .B2(n20276), .ZN(
        n20280) );
  AOI21_X1 U23187 ( .B1(n20282), .B2(n20281), .A(n20280), .ZN(n20283) );
  OAI211_X1 U23188 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20285), .A(
        n20284), .B(n20283), .ZN(P1_U2839) );
  INV_X1 U23189 ( .A(n20286), .ZN(n20287) );
  OAI22_X1 U23190 ( .A1(n20289), .A2(n14452), .B1(n20288), .B2(n20287), .ZN(
        n20290) );
  INV_X1 U23191 ( .A(n20290), .ZN(n20291) );
  OAI21_X1 U23192 ( .B1(n20302), .B2(n20292), .A(n20291), .ZN(P1_U2863) );
  AOI22_X1 U23193 ( .A1(n20294), .A2(n20299), .B1(n20298), .B2(n20293), .ZN(
        n20295) );
  OAI21_X1 U23194 ( .B1(n20302), .B2(n20296), .A(n20295), .ZN(P1_U2865) );
  AOI22_X1 U23195 ( .A1(n20300), .A2(n20299), .B1(n20298), .B2(n20297), .ZN(
        n20301) );
  OAI21_X1 U23196 ( .B1(n20302), .B2(n21135), .A(n20301), .ZN(P1_U2867) );
  AOI22_X1 U23197 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20306), .B1(n20331), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20303) );
  OAI21_X1 U23198 ( .B1(n20305), .B2(n20304), .A(n20303), .ZN(P1_U2921) );
  AOI22_X1 U23199 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20307) );
  OAI21_X1 U23200 ( .B1(n14547), .B2(n20334), .A(n20307), .ZN(P1_U2922) );
  INV_X1 U23201 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20309) );
  AOI22_X1 U23202 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20308) );
  OAI21_X1 U23203 ( .B1(n20309), .B2(n20334), .A(n20308), .ZN(P1_U2923) );
  INV_X1 U23204 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20311) );
  AOI22_X1 U23205 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20310) );
  OAI21_X1 U23206 ( .B1(n20311), .B2(n20334), .A(n20310), .ZN(P1_U2924) );
  INV_X1 U23207 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20313) );
  AOI22_X1 U23208 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20312) );
  OAI21_X1 U23209 ( .B1(n20313), .B2(n20334), .A(n20312), .ZN(P1_U2925) );
  INV_X1 U23210 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20315) );
  AOI22_X1 U23211 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20314) );
  OAI21_X1 U23212 ( .B1(n20315), .B2(n20334), .A(n20314), .ZN(P1_U2926) );
  AOI22_X1 U23213 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20316) );
  OAI21_X1 U23214 ( .B1(n13938), .B2(n20334), .A(n20316), .ZN(P1_U2927) );
  INV_X1 U23215 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20318) );
  AOI22_X1 U23216 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20317) );
  OAI21_X1 U23217 ( .B1(n20318), .B2(n20334), .A(n20317), .ZN(P1_U2928) );
  AOI22_X1 U23218 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20319) );
  OAI21_X1 U23219 ( .B1(n20320), .B2(n20334), .A(n20319), .ZN(P1_U2929) );
  AOI22_X1 U23220 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20321) );
  OAI21_X1 U23221 ( .B1(n20322), .B2(n20334), .A(n20321), .ZN(P1_U2930) );
  AOI22_X1 U23222 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20323) );
  OAI21_X1 U23223 ( .B1(n13753), .B2(n20334), .A(n20323), .ZN(P1_U2931) );
  AOI22_X1 U23224 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20324) );
  OAI21_X1 U23225 ( .B1(n21336), .B2(n20334), .A(n20324), .ZN(P1_U2932) );
  AOI22_X1 U23226 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20325) );
  OAI21_X1 U23227 ( .B1(n20326), .B2(n20334), .A(n20325), .ZN(P1_U2933) );
  AOI22_X1 U23228 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20327) );
  OAI21_X1 U23229 ( .B1(n20328), .B2(n20334), .A(n20327), .ZN(P1_U2934) );
  AOI22_X1 U23230 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20329) );
  OAI21_X1 U23231 ( .B1(n20330), .B2(n20334), .A(n20329), .ZN(P1_U2935) );
  AOI22_X1 U23232 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20332), .B1(n20331), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20333) );
  OAI21_X1 U23233 ( .B1(n20335), .B2(n20334), .A(n20333), .ZN(P1_U2936) );
  AOI22_X1 U23234 ( .A1(n20363), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20360), .ZN(n20337) );
  NAND2_X1 U23235 ( .A1(n20348), .A2(n20336), .ZN(n20350) );
  NAND2_X1 U23236 ( .A1(n20337), .A2(n20350), .ZN(P1_U2945) );
  AOI22_X1 U23237 ( .A1(n20363), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20360), .ZN(n20339) );
  NAND2_X1 U23238 ( .A1(n20348), .A2(n20338), .ZN(n20354) );
  NAND2_X1 U23239 ( .A1(n20339), .A2(n20354), .ZN(P1_U2947) );
  AOI22_X1 U23240 ( .A1(n20363), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20360), .ZN(n20341) );
  NAND2_X1 U23241 ( .A1(n20348), .A2(n20340), .ZN(n20356) );
  NAND2_X1 U23242 ( .A1(n20341), .A2(n20356), .ZN(P1_U2948) );
  AOI22_X1 U23243 ( .A1(n20363), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20360), .ZN(n20343) );
  NAND2_X1 U23244 ( .A1(n20348), .A2(n20342), .ZN(n20358) );
  NAND2_X1 U23245 ( .A1(n20343), .A2(n20358), .ZN(P1_U2949) );
  AOI22_X1 U23246 ( .A1(n20363), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20360), .ZN(n20345) );
  NAND2_X1 U23247 ( .A1(n20348), .A2(n20344), .ZN(n20361) );
  NAND2_X1 U23248 ( .A1(n20345), .A2(n20361), .ZN(P1_U2950) );
  AOI22_X1 U23249 ( .A1(n20363), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20360), .ZN(n20349) );
  INV_X1 U23250 ( .A(n20346), .ZN(n20347) );
  NAND2_X1 U23251 ( .A1(n20348), .A2(n20347), .ZN(n20364) );
  NAND2_X1 U23252 ( .A1(n20349), .A2(n20364), .ZN(P1_U2951) );
  AOI22_X1 U23253 ( .A1(n20363), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20360), .ZN(n20351) );
  NAND2_X1 U23254 ( .A1(n20351), .A2(n20350), .ZN(P1_U2960) );
  AOI22_X1 U23255 ( .A1(n20363), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20360), .ZN(n20353) );
  NAND2_X1 U23256 ( .A1(n20353), .A2(n20352), .ZN(P1_U2961) );
  AOI22_X1 U23257 ( .A1(n20363), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20360), .ZN(n20355) );
  NAND2_X1 U23258 ( .A1(n20355), .A2(n20354), .ZN(P1_U2962) );
  AOI22_X1 U23259 ( .A1(n20363), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20360), .ZN(n20357) );
  NAND2_X1 U23260 ( .A1(n20357), .A2(n20356), .ZN(P1_U2963) );
  AOI22_X1 U23261 ( .A1(n20363), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20360), .ZN(n20359) );
  NAND2_X1 U23262 ( .A1(n20359), .A2(n20358), .ZN(P1_U2964) );
  AOI22_X1 U23263 ( .A1(n20363), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20360), .ZN(n20362) );
  NAND2_X1 U23264 ( .A1(n20362), .A2(n20361), .ZN(P1_U2965) );
  AOI22_X1 U23265 ( .A1(n20363), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20360), .ZN(n20365) );
  NAND2_X1 U23266 ( .A1(n20365), .A2(n20364), .ZN(P1_U2966) );
  OR2_X1 U23267 ( .A1(n20367), .A2(n20366), .ZN(n20368) );
  AOI22_X1 U23268 ( .A1(n20370), .A2(n20369), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20368), .ZN(n20372) );
  OAI211_X1 U23269 ( .C1(n20374), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P1_U2999) );
  NOR2_X1 U23270 ( .A1(n20376), .A2(n20375), .ZN(P1_U3032) );
  NAND2_X1 U23271 ( .A1(n20378), .A2(n20377), .ZN(n20403) );
  NAND2_X1 U23272 ( .A1(n20379), .A2(n20378), .ZN(n20402) );
  INV_X1 U23273 ( .A(n20402), .ZN(n20422) );
  AOI22_X1 U23274 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20423), .B1(DATAI_16_), 
        .B2(n20422), .ZN(n20906) );
  NAND2_X1 U23275 ( .A1(n13604), .A2(n20382), .ZN(n20796) );
  INV_X1 U23276 ( .A(n20796), .ZN(n20636) );
  AOI22_X1 U23277 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20423), .B1(DATAI_24_), 
        .B2(n20422), .ZN(n20972) );
  INV_X1 U23278 ( .A(n20972), .ZN(n20903) );
  NAND2_X1 U23279 ( .A1(n20425), .A2(n9755), .ZN(n20964) );
  INV_X1 U23280 ( .A(n20964), .ZN(n20892) );
  NAND2_X1 U23281 ( .A1(n10574), .A2(n20679), .ZN(n20500) );
  OR2_X1 U23282 ( .A1(n20833), .A2(n20500), .ZN(n20388) );
  INV_X1 U23283 ( .A(n20388), .ZN(n20426) );
  AOI22_X1 U23284 ( .A1(n21021), .A2(n20903), .B1(n20892), .B2(n20426), .ZN(
        n20397) );
  INV_X1 U23285 ( .A(n20747), .ZN(n20384) );
  OR2_X1 U23286 ( .A1(n20681), .A2(n20384), .ZN(n20393) );
  INV_X1 U23287 ( .A(n20393), .ZN(n20536) );
  NAND2_X1 U23288 ( .A1(n20392), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20889) );
  INV_X1 U23289 ( .A(n21021), .ZN(n20385) );
  NAND3_X1 U23290 ( .A1(n20385), .A2(n20826), .A3(n20442), .ZN(n20386) );
  NAND2_X1 U23291 ( .A1(n20826), .A2(n20894), .ZN(n20828) );
  NAND2_X1 U23292 ( .A1(n20386), .A2(n20828), .ZN(n20391) );
  OR2_X1 U23293 ( .A1(n20680), .A2(n20387), .ZN(n20499) );
  OR2_X1 U23294 ( .A1(n20499), .A2(n20896), .ZN(n20394) );
  AOI22_X1 U23295 ( .A1(n20391), .A2(n20394), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20388), .ZN(n20389) );
  NAND2_X1 U23296 ( .A1(n20390), .A2(n20427), .ZN(n20963) );
  INV_X1 U23297 ( .A(n20963), .ZN(n20891) );
  INV_X1 U23298 ( .A(n20391), .ZN(n20395) );
  OR2_X1 U23299 ( .A1(n20392), .A2(n21030), .ZN(n20543) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20430), .B1(
        n20891), .B2(n20429), .ZN(n20396) );
  OAI211_X1 U23301 ( .C1(n20906), .C2(n20442), .A(n20397), .B(n20396), .ZN(
        P1_U3033) );
  AOI22_X1 U23302 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20423), .B1(DATAI_17_), 
        .B2(n20422), .ZN(n20912) );
  AOI22_X1 U23303 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20423), .B1(DATAI_25_), 
        .B2(n20422), .ZN(n20979) );
  INV_X1 U23304 ( .A(n20979), .ZN(n20909) );
  NAND2_X1 U23305 ( .A1(n20425), .A2(n20398), .ZN(n20974) );
  INV_X1 U23306 ( .A(n20974), .ZN(n20908) );
  AOI22_X1 U23307 ( .A1(n21021), .A2(n20909), .B1(n20908), .B2(n20426), .ZN(
        n20401) );
  NAND2_X1 U23308 ( .A1(n20399), .A2(n20427), .ZN(n20973) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20430), .B1(
        n20907), .B2(n20429), .ZN(n20400) );
  OAI211_X1 U23310 ( .C1(n20912), .C2(n20442), .A(n20401), .B(n20400), .ZN(
        P1_U3034) );
  OAI22_X1 U23311 ( .A1(n20404), .A2(n20403), .B1(n14529), .B2(n20402), .ZN(
        n20983) );
  INV_X1 U23312 ( .A(n20983), .ZN(n20918) );
  AOI22_X1 U23313 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20423), .B1(DATAI_26_), 
        .B2(n20422), .ZN(n20986) );
  INV_X1 U23314 ( .A(n20986), .ZN(n20915) );
  NAND2_X1 U23315 ( .A1(n20425), .A2(n10063), .ZN(n20981) );
  INV_X1 U23316 ( .A(n20981), .ZN(n20914) );
  AOI22_X1 U23317 ( .A1(n21021), .A2(n20915), .B1(n20914), .B2(n20426), .ZN(
        n20407) );
  NAND2_X1 U23318 ( .A1(n20405), .A2(n20427), .ZN(n20980) );
  INV_X1 U23319 ( .A(n20980), .ZN(n20913) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20430), .B1(
        n20913), .B2(n20429), .ZN(n20406) );
  OAI211_X1 U23321 ( .C1(n20918), .C2(n20442), .A(n20407), .B(n20406), .ZN(
        P1_U3035) );
  AOI22_X1 U23322 ( .A1(DATAI_19_), .A2(n20422), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20423), .ZN(n20924) );
  AOI22_X1 U23323 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20423), .B1(DATAI_27_), 
        .B2(n20422), .ZN(n20993) );
  INV_X1 U23324 ( .A(n20993), .ZN(n20921) );
  NAND2_X1 U23325 ( .A1(n20425), .A2(n20408), .ZN(n20988) );
  INV_X1 U23326 ( .A(n20988), .ZN(n20920) );
  AOI22_X1 U23327 ( .A1(n21021), .A2(n20921), .B1(n20920), .B2(n20426), .ZN(
        n20411) );
  NAND2_X1 U23328 ( .A1(n20409), .A2(n20427), .ZN(n20987) );
  INV_X1 U23329 ( .A(n20987), .ZN(n20919) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20430), .B1(
        n20919), .B2(n20429), .ZN(n20410) );
  OAI211_X1 U23331 ( .C1(n20924), .C2(n20442), .A(n20411), .B(n20410), .ZN(
        P1_U3036) );
  AOI22_X1 U23332 ( .A1(DATAI_20_), .A2(n20422), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20423), .ZN(n20930) );
  AOI22_X1 U23333 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20423), .B1(DATAI_28_), 
        .B2(n20422), .ZN(n21000) );
  INV_X1 U23334 ( .A(n21000), .ZN(n20927) );
  NAND2_X1 U23335 ( .A1(n20425), .A2(n9779), .ZN(n20995) );
  INV_X1 U23336 ( .A(n20995), .ZN(n20926) );
  AOI22_X1 U23337 ( .A1(n21021), .A2(n20927), .B1(n20926), .B2(n20426), .ZN(
        n20415) );
  NAND2_X1 U23338 ( .A1(n20413), .A2(n20427), .ZN(n20994) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20430), .B1(
        n20925), .B2(n20429), .ZN(n20414) );
  OAI211_X1 U23340 ( .C1(n20930), .C2(n20442), .A(n20415), .B(n20414), .ZN(
        P1_U3037) );
  AOI22_X1 U23341 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20423), .B1(DATAI_21_), 
        .B2(n20422), .ZN(n20936) );
  AOI22_X1 U23342 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20423), .B1(DATAI_29_), 
        .B2(n20422), .ZN(n21007) );
  INV_X1 U23343 ( .A(n21007), .ZN(n20933) );
  NAND2_X1 U23344 ( .A1(n20425), .A2(n10552), .ZN(n21002) );
  INV_X1 U23345 ( .A(n21002), .ZN(n20932) );
  AOI22_X1 U23346 ( .A1(n21021), .A2(n20933), .B1(n20932), .B2(n20426), .ZN(
        n20418) );
  NAND2_X1 U23347 ( .A1(n20416), .A2(n20427), .ZN(n21001) );
  INV_X1 U23348 ( .A(n21001), .ZN(n20931) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20430), .B1(
        n20931), .B2(n20429), .ZN(n20417) );
  OAI211_X1 U23350 ( .C1(n20936), .C2(n20442), .A(n20418), .B(n20417), .ZN(
        P1_U3038) );
  AOI22_X1 U23351 ( .A1(DATAI_22_), .A2(n20422), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20423), .ZN(n20942) );
  AOI22_X1 U23352 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20423), .B1(DATAI_30_), 
        .B2(n20422), .ZN(n21014) );
  INV_X1 U23353 ( .A(n21014), .ZN(n20939) );
  NAND2_X1 U23354 ( .A1(n20425), .A2(n10623), .ZN(n21009) );
  INV_X1 U23355 ( .A(n21009), .ZN(n20938) );
  AOI22_X1 U23356 ( .A1(n21021), .A2(n20939), .B1(n20938), .B2(n20426), .ZN(
        n20421) );
  NAND2_X1 U23357 ( .A1(n20419), .A2(n20427), .ZN(n21008) );
  INV_X1 U23358 ( .A(n21008), .ZN(n20937) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20430), .B1(
        n20937), .B2(n20429), .ZN(n20420) );
  OAI211_X1 U23360 ( .C1(n20942), .C2(n20442), .A(n20421), .B(n20420), .ZN(
        P1_U3039) );
  AOI22_X1 U23361 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20423), .B1(DATAI_23_), 
        .B2(n20422), .ZN(n20952) );
  AOI22_X1 U23362 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20423), .B1(DATAI_31_), 
        .B2(n20422), .ZN(n21026) );
  INV_X1 U23363 ( .A(n21026), .ZN(n20947) );
  NAND2_X1 U23364 ( .A1(n20425), .A2(n20424), .ZN(n21018) );
  INV_X1 U23365 ( .A(n21018), .ZN(n20946) );
  AOI22_X1 U23366 ( .A1(n21021), .A2(n20947), .B1(n20946), .B2(n20426), .ZN(
        n20432) );
  NAND2_X1 U23367 ( .A1(n20428), .A2(n20427), .ZN(n21016) );
  INV_X1 U23368 ( .A(n21016), .ZN(n20944) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20430), .B1(
        n20944), .B2(n20429), .ZN(n20431) );
  OAI211_X1 U23370 ( .C1(n20952), .C2(n20442), .A(n20432), .B(n20431), .ZN(
        P1_U3040) );
  NOR2_X1 U23371 ( .A1(n20500), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20437) );
  INV_X1 U23372 ( .A(n20437), .ZN(n20434) );
  NOR2_X1 U23373 ( .A1(n21321), .A2(n20434), .ZN(n20454) );
  INV_X1 U23374 ( .A(n20499), .ZN(n20433) );
  INV_X1 U23375 ( .A(n20861), .ZN(n20718) );
  AOI21_X1 U23376 ( .B1(n20433), .B2(n20718), .A(n20454), .ZN(n20435) );
  OAI22_X1 U23377 ( .A1(n20435), .A2(n20958), .B1(n20434), .B2(n21030), .ZN(
        n20453) );
  AOI22_X1 U23378 ( .A1(n20892), .A2(n20454), .B1(n20891), .B2(n20453), .ZN(
        n20439) );
  INV_X1 U23379 ( .A(n20494), .ZN(n20504) );
  OAI21_X1 U23380 ( .B1(n20504), .B2(n20894), .A(n20435), .ZN(n20436) );
  OAI221_X1 U23381 ( .B1(n20826), .B2(n20437), .C1(n20958), .C2(n20436), .A(
        n20966), .ZN(n20456) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20903), .ZN(n20438) );
  OAI211_X1 U23383 ( .C1(n20906), .C2(n20487), .A(n20439), .B(n20438), .ZN(
        P1_U3041) );
  AOI22_X1 U23384 ( .A1(n20908), .A2(n20454), .B1(n20907), .B2(n20453), .ZN(
        n20441) );
  INV_X1 U23385 ( .A(n20487), .ZN(n20460) );
  INV_X1 U23386 ( .A(n20912), .ZN(n20976) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20456), .B1(
        n20460), .B2(n20976), .ZN(n20440) );
  OAI211_X1 U23388 ( .C1(n20979), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P1_U3042) );
  AOI22_X1 U23389 ( .A1(n20914), .A2(n20454), .B1(n20913), .B2(n20453), .ZN(
        n20444) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20915), .ZN(n20443) );
  OAI211_X1 U23391 ( .C1(n20918), .C2(n20487), .A(n20444), .B(n20443), .ZN(
        P1_U3043) );
  AOI22_X1 U23392 ( .A1(n20920), .A2(n20454), .B1(n20919), .B2(n20453), .ZN(
        n20446) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20921), .ZN(n20445) );
  OAI211_X1 U23394 ( .C1(n20924), .C2(n20487), .A(n20446), .B(n20445), .ZN(
        P1_U3044) );
  AOI22_X1 U23395 ( .A1(n20926), .A2(n20454), .B1(n20925), .B2(n20453), .ZN(
        n20448) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20927), .ZN(n20447) );
  OAI211_X1 U23397 ( .C1(n20930), .C2(n20487), .A(n20448), .B(n20447), .ZN(
        P1_U3045) );
  AOI22_X1 U23398 ( .A1(n20932), .A2(n20454), .B1(n20931), .B2(n20453), .ZN(
        n20450) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20933), .ZN(n20449) );
  OAI211_X1 U23400 ( .C1(n20936), .C2(n20487), .A(n20450), .B(n20449), .ZN(
        P1_U3046) );
  AOI22_X1 U23401 ( .A1(n20938), .A2(n20454), .B1(n20937), .B2(n20453), .ZN(
        n20452) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20939), .ZN(n20451) );
  OAI211_X1 U23403 ( .C1(n20942), .C2(n20487), .A(n20452), .B(n20451), .ZN(
        P1_U3047) );
  AOI22_X1 U23404 ( .A1(n20946), .A2(n20454), .B1(n20944), .B2(n20453), .ZN(
        n20458) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20947), .ZN(n20457) );
  OAI211_X1 U23406 ( .C1(n20952), .C2(n20487), .A(n20458), .B(n20457), .ZN(
        P1_U3048) );
  NAND2_X1 U23407 ( .A1(n13604), .A2(n20381), .ZN(n20745) );
  OR3_X1 U23408 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20957), .A3(
        n20500), .ZN(n20486) );
  OAI22_X1 U23409 ( .A1(n20487), .A2(n20972), .B1(n20964), .B2(n20486), .ZN(
        n20459) );
  INV_X1 U23410 ( .A(n20459), .ZN(n20467) );
  OAI21_X1 U23411 ( .B1(n20522), .B2(n20460), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20461) );
  NAND2_X1 U23412 ( .A1(n20461), .A2(n20826), .ZN(n20465) );
  INV_X1 U23413 ( .A(n20465), .ZN(n20462) );
  OR2_X1 U23414 ( .A1(n20499), .A2(n14186), .ZN(n20464) );
  AOI22_X1 U23415 ( .A1(n20462), .A2(n20464), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20486), .ZN(n20463) );
  OR2_X1 U23416 ( .A1(n20747), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20606) );
  NAND2_X1 U23417 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20606), .ZN(n20603) );
  NAND3_X1 U23418 ( .A1(n20755), .A2(n20463), .A3(n20603), .ZN(n20490) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20490), .B1(
        n20891), .B2(n20489), .ZN(n20466) );
  OAI211_X1 U23420 ( .C1(n20906), .C2(n20529), .A(n20467), .B(n20466), .ZN(
        P1_U3049) );
  OAI22_X1 U23421 ( .A1(n20487), .A2(n20979), .B1(n20486), .B2(n20974), .ZN(
        n20468) );
  INV_X1 U23422 ( .A(n20468), .ZN(n20470) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20490), .B1(
        n20907), .B2(n20489), .ZN(n20469) );
  OAI211_X1 U23424 ( .C1(n20912), .C2(n20529), .A(n20470), .B(n20469), .ZN(
        P1_U3050) );
  OAI22_X1 U23425 ( .A1(n20529), .A2(n20918), .B1(n20486), .B2(n20981), .ZN(
        n20471) );
  INV_X1 U23426 ( .A(n20471), .ZN(n20473) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20490), .B1(
        n20913), .B2(n20489), .ZN(n20472) );
  OAI211_X1 U23428 ( .C1(n20986), .C2(n20487), .A(n20473), .B(n20472), .ZN(
        P1_U3051) );
  OAI22_X1 U23429 ( .A1(n20529), .A2(n20924), .B1(n20486), .B2(n20988), .ZN(
        n20474) );
  INV_X1 U23430 ( .A(n20474), .ZN(n20476) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20490), .B1(
        n20919), .B2(n20489), .ZN(n20475) );
  OAI211_X1 U23432 ( .C1(n20993), .C2(n20487), .A(n20476), .B(n20475), .ZN(
        P1_U3052) );
  OAI22_X1 U23433 ( .A1(n20487), .A2(n21000), .B1(n20486), .B2(n20995), .ZN(
        n20477) );
  INV_X1 U23434 ( .A(n20477), .ZN(n20479) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20490), .B1(
        n20925), .B2(n20489), .ZN(n20478) );
  OAI211_X1 U23436 ( .C1(n20930), .C2(n20529), .A(n20479), .B(n20478), .ZN(
        P1_U3053) );
  OAI22_X1 U23437 ( .A1(n20529), .A2(n20936), .B1(n20486), .B2(n21002), .ZN(
        n20480) );
  INV_X1 U23438 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20490), .B1(
        n20931), .B2(n20489), .ZN(n20481) );
  OAI211_X1 U23440 ( .C1(n21007), .C2(n20487), .A(n20482), .B(n20481), .ZN(
        P1_U3054) );
  OAI22_X1 U23441 ( .A1(n20487), .A2(n21014), .B1(n20486), .B2(n21009), .ZN(
        n20483) );
  INV_X1 U23442 ( .A(n20483), .ZN(n20485) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20490), .B1(
        n20937), .B2(n20489), .ZN(n20484) );
  OAI211_X1 U23444 ( .C1(n20942), .C2(n20529), .A(n20485), .B(n20484), .ZN(
        P1_U3055) );
  OAI22_X1 U23445 ( .A1(n20487), .A2(n21026), .B1(n20486), .B2(n21018), .ZN(
        n20488) );
  INV_X1 U23446 ( .A(n20488), .ZN(n20492) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20490), .B1(
        n20944), .B2(n20489), .ZN(n20491) );
  OAI211_X1 U23448 ( .C1(n20952), .C2(n20529), .A(n20492), .B(n20491), .ZN(
        P1_U3056) );
  NOR2_X1 U23449 ( .A1(n20957), .A2(n20500), .ZN(n20508) );
  AOI21_X1 U23450 ( .B1(n20494), .B2(n20493), .A(n20958), .ZN(n20506) );
  INV_X1 U23451 ( .A(n20495), .ZN(n20497) );
  AND2_X1 U23452 ( .A1(n20497), .A2(n20496), .ZN(n20961) );
  INV_X1 U23453 ( .A(n20961), .ZN(n20498) );
  OR2_X1 U23454 ( .A1(n20499), .A2(n20498), .ZN(n20502) );
  INV_X1 U23455 ( .A(n20500), .ZN(n20501) );
  NAND2_X1 U23456 ( .A1(n20954), .A2(n20501), .ZN(n20528) );
  AND2_X1 U23457 ( .A1(n20502), .A2(n20528), .ZN(n20505) );
  INV_X1 U23458 ( .A(n20505), .ZN(n20503) );
  INV_X1 U23459 ( .A(n20906), .ZN(n20969) );
  INV_X1 U23460 ( .A(n20528), .ZN(n20521) );
  AOI22_X1 U23461 ( .A1(n20570), .A2(n20969), .B1(n20892), .B2(n20521), .ZN(
        n20510) );
  NAND2_X1 U23462 ( .A1(n20506), .A2(n20505), .ZN(n20507) );
  OAI211_X1 U23463 ( .C1(n20826), .C2(n20508), .A(n20966), .B(n20507), .ZN(
        n20531) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20531), .B1(
        n20522), .B2(n20903), .ZN(n20509) );
  OAI211_X1 U23465 ( .C1(n20534), .C2(n20963), .A(n20510), .B(n20509), .ZN(
        P1_U3057) );
  AOI22_X1 U23466 ( .A1(n20570), .A2(n20976), .B1(n20908), .B2(n20521), .ZN(
        n20512) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20531), .B1(
        n20522), .B2(n20909), .ZN(n20511) );
  OAI211_X1 U23468 ( .C1(n20534), .C2(n20973), .A(n20512), .B(n20511), .ZN(
        P1_U3058) );
  AOI22_X1 U23469 ( .A1(n20570), .A2(n20983), .B1(n20521), .B2(n20914), .ZN(
        n20514) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20531), .B1(
        n20522), .B2(n20915), .ZN(n20513) );
  OAI211_X1 U23471 ( .C1(n20534), .C2(n20980), .A(n20514), .B(n20513), .ZN(
        P1_U3059) );
  OAI22_X1 U23472 ( .A1(n20529), .A2(n20993), .B1(n20528), .B2(n20988), .ZN(
        n20515) );
  INV_X1 U23473 ( .A(n20515), .ZN(n20517) );
  INV_X1 U23474 ( .A(n20924), .ZN(n20990) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20531), .B1(
        n20570), .B2(n20990), .ZN(n20516) );
  OAI211_X1 U23476 ( .C1(n20534), .C2(n20987), .A(n20517), .B(n20516), .ZN(
        P1_U3060) );
  OAI22_X1 U23477 ( .A1(n20529), .A2(n21000), .B1(n20995), .B2(n20528), .ZN(
        n20518) );
  INV_X1 U23478 ( .A(n20518), .ZN(n20520) );
  INV_X1 U23479 ( .A(n20930), .ZN(n20997) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20531), .B1(
        n20570), .B2(n20997), .ZN(n20519) );
  OAI211_X1 U23481 ( .C1(n20534), .C2(n20994), .A(n20520), .B(n20519), .ZN(
        P1_U3061) );
  INV_X1 U23482 ( .A(n20936), .ZN(n21004) );
  AOI22_X1 U23483 ( .A1(n20570), .A2(n21004), .B1(n20521), .B2(n20932), .ZN(
        n20524) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20531), .B1(
        n20522), .B2(n20933), .ZN(n20523) );
  OAI211_X1 U23485 ( .C1(n20534), .C2(n21001), .A(n20524), .B(n20523), .ZN(
        P1_U3062) );
  OAI22_X1 U23486 ( .A1(n20529), .A2(n21014), .B1(n21009), .B2(n20528), .ZN(
        n20525) );
  INV_X1 U23487 ( .A(n20525), .ZN(n20527) );
  INV_X1 U23488 ( .A(n20942), .ZN(n21011) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20531), .B1(
        n20570), .B2(n21011), .ZN(n20526) );
  OAI211_X1 U23490 ( .C1(n20534), .C2(n21008), .A(n20527), .B(n20526), .ZN(
        P1_U3063) );
  OAI22_X1 U23491 ( .A1(n20529), .A2(n21026), .B1(n21018), .B2(n20528), .ZN(
        n20530) );
  INV_X1 U23492 ( .A(n20530), .ZN(n20533) );
  INV_X1 U23493 ( .A(n20952), .ZN(n21020) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20531), .B1(
        n20570), .B2(n21020), .ZN(n20532) );
  OAI211_X1 U23495 ( .C1(n20534), .C2(n21016), .A(n20533), .B(n20532), .ZN(
        P1_U3064) );
  OR2_X1 U23496 ( .A1(n20833), .A2(n20600), .ZN(n20568) );
  NOR2_X1 U23497 ( .A1(n20831), .A2(n20535), .ZN(n20639) );
  NAND3_X1 U23498 ( .A1(n20639), .A2(n20826), .A3(n14186), .ZN(n20538) );
  INV_X1 U23499 ( .A(n20889), .ZN(n20832) );
  NAND2_X1 U23500 ( .A1(n20536), .A2(n20832), .ZN(n20537) );
  AND2_X1 U23501 ( .A1(n20538), .A2(n20537), .ZN(n20567) );
  OAI22_X1 U23502 ( .A1(n20964), .A2(n20568), .B1(n20963), .B2(n20567), .ZN(
        n20539) );
  INV_X1 U23503 ( .A(n20539), .ZN(n20548) );
  INV_X1 U23504 ( .A(n20568), .ZN(n20546) );
  INV_X1 U23505 ( .A(n20639), .ZN(n20542) );
  INV_X1 U23506 ( .A(n20599), .ZN(n20540) );
  OAI21_X1 U23507 ( .B1(n20570), .B2(n20540), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20541) );
  OAI21_X1 U23508 ( .B1(n20896), .B2(n20542), .A(n20541), .ZN(n20545) );
  INV_X1 U23509 ( .A(n20543), .ZN(n20748) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20903), .ZN(n20547) );
  OAI211_X1 U23511 ( .C1(n20906), .C2(n20599), .A(n20548), .B(n20547), .ZN(
        P1_U3065) );
  OAI22_X1 U23512 ( .A1(n20974), .A2(n20568), .B1(n20973), .B2(n20567), .ZN(
        n20549) );
  INV_X1 U23513 ( .A(n20549), .ZN(n20551) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20909), .ZN(n20550) );
  OAI211_X1 U23515 ( .C1(n20912), .C2(n20599), .A(n20551), .B(n20550), .ZN(
        P1_U3066) );
  OAI22_X1 U23516 ( .A1(n20981), .A2(n20568), .B1(n20980), .B2(n20567), .ZN(
        n20552) );
  INV_X1 U23517 ( .A(n20552), .ZN(n20554) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20915), .ZN(n20553) );
  OAI211_X1 U23519 ( .C1(n20918), .C2(n20599), .A(n20554), .B(n20553), .ZN(
        P1_U3067) );
  OAI22_X1 U23520 ( .A1(n20988), .A2(n20568), .B1(n20987), .B2(n20567), .ZN(
        n20555) );
  INV_X1 U23521 ( .A(n20555), .ZN(n20557) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20921), .ZN(n20556) );
  OAI211_X1 U23523 ( .C1(n20924), .C2(n20599), .A(n20557), .B(n20556), .ZN(
        P1_U3068) );
  OAI22_X1 U23524 ( .A1(n20995), .A2(n20568), .B1(n20994), .B2(n20567), .ZN(
        n20558) );
  INV_X1 U23525 ( .A(n20558), .ZN(n20560) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20927), .ZN(n20559) );
  OAI211_X1 U23527 ( .C1(n20930), .C2(n20599), .A(n20560), .B(n20559), .ZN(
        P1_U3069) );
  OAI22_X1 U23528 ( .A1(n21002), .A2(n20568), .B1(n21001), .B2(n20567), .ZN(
        n20561) );
  INV_X1 U23529 ( .A(n20561), .ZN(n20563) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20933), .ZN(n20562) );
  OAI211_X1 U23531 ( .C1(n20936), .C2(n20599), .A(n20563), .B(n20562), .ZN(
        P1_U3070) );
  OAI22_X1 U23532 ( .A1(n21009), .A2(n20568), .B1(n21008), .B2(n20567), .ZN(
        n20564) );
  INV_X1 U23533 ( .A(n20564), .ZN(n20566) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20939), .ZN(n20565) );
  OAI211_X1 U23535 ( .C1(n20942), .C2(n20599), .A(n20566), .B(n20565), .ZN(
        P1_U3071) );
  OAI22_X1 U23536 ( .A1(n21018), .A2(n20568), .B1(n21016), .B2(n20567), .ZN(
        n20569) );
  INV_X1 U23537 ( .A(n20569), .ZN(n20573) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20947), .ZN(n20572) );
  OAI211_X1 U23539 ( .C1(n20952), .C2(n20599), .A(n20573), .B(n20572), .ZN(
        P1_U3072) );
  NOR2_X1 U23540 ( .A1(n20600), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20578) );
  INV_X1 U23541 ( .A(n20578), .ZN(n20574) );
  NOR2_X1 U23542 ( .A1(n21321), .A2(n20574), .ZN(n20594) );
  AOI21_X1 U23543 ( .B1(n20639), .B2(n20718), .A(n20594), .ZN(n20575) );
  OAI22_X1 U23544 ( .A1(n20575), .A2(n20958), .B1(n20574), .B2(n21030), .ZN(
        n20593) );
  AOI22_X1 U23545 ( .A1(n20892), .A2(n20594), .B1(n20891), .B2(n20593), .ZN(
        n20580) );
  INV_X1 U23546 ( .A(n20637), .ZN(n20576) );
  OAI21_X1 U23547 ( .B1(n20576), .B2(n20894), .A(n20575), .ZN(n20577) );
  OAI221_X1 U23548 ( .B1(n20826), .B2(n20578), .C1(n20958), .C2(n20577), .A(
        n20966), .ZN(n20596) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n20969), .ZN(n20579) );
  OAI211_X1 U23550 ( .C1(n20972), .C2(n20599), .A(n20580), .B(n20579), .ZN(
        P1_U3073) );
  AOI22_X1 U23551 ( .A1(n20908), .A2(n20594), .B1(n20907), .B2(n20593), .ZN(
        n20582) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n20976), .ZN(n20581) );
  OAI211_X1 U23553 ( .C1(n20979), .C2(n20599), .A(n20582), .B(n20581), .ZN(
        P1_U3074) );
  AOI22_X1 U23554 ( .A1(n20914), .A2(n20594), .B1(n20913), .B2(n20593), .ZN(
        n20584) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n20983), .ZN(n20583) );
  OAI211_X1 U23556 ( .C1(n20986), .C2(n20599), .A(n20584), .B(n20583), .ZN(
        P1_U3075) );
  AOI22_X1 U23557 ( .A1(n20920), .A2(n20594), .B1(n20919), .B2(n20593), .ZN(
        n20586) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n20990), .ZN(n20585) );
  OAI211_X1 U23559 ( .C1(n20993), .C2(n20599), .A(n20586), .B(n20585), .ZN(
        P1_U3076) );
  AOI22_X1 U23560 ( .A1(n20926), .A2(n20594), .B1(n20925), .B2(n20593), .ZN(
        n20588) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n20997), .ZN(n20587) );
  OAI211_X1 U23562 ( .C1(n21000), .C2(n20599), .A(n20588), .B(n20587), .ZN(
        P1_U3077) );
  AOI22_X1 U23563 ( .A1(n20932), .A2(n20594), .B1(n20931), .B2(n20593), .ZN(
        n20590) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n21004), .ZN(n20589) );
  OAI211_X1 U23565 ( .C1(n21007), .C2(n20599), .A(n20590), .B(n20589), .ZN(
        P1_U3078) );
  AOI22_X1 U23566 ( .A1(n20938), .A2(n20594), .B1(n20937), .B2(n20593), .ZN(
        n20592) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n21011), .ZN(n20591) );
  OAI211_X1 U23568 ( .C1(n21014), .C2(n20599), .A(n20592), .B(n20591), .ZN(
        P1_U3079) );
  AOI22_X1 U23569 ( .A1(n20946), .A2(n20594), .B1(n20944), .B2(n20593), .ZN(
        n20598) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20596), .B1(
        n20595), .B2(n21020), .ZN(n20597) );
  OAI211_X1 U23571 ( .C1(n21026), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P1_U3080) );
  NOR2_X1 U23572 ( .A1(n20957), .A2(n20600), .ZN(n20648) );
  NAND2_X1 U23573 ( .A1(n21321), .A2(n20648), .ZN(n20629) );
  OAI22_X1 U23574 ( .A1(n20630), .A2(n20972), .B1(n20964), .B2(n20629), .ZN(
        n20601) );
  INV_X1 U23575 ( .A(n20601), .ZN(n20610) );
  NAND2_X1 U23576 ( .A1(n20666), .A2(n20630), .ZN(n20602) );
  AOI21_X1 U23577 ( .B1(n20602), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20958), 
        .ZN(n20605) );
  NAND2_X1 U23578 ( .A1(n20639), .A2(n20896), .ZN(n20607) );
  AOI22_X1 U23579 ( .A1(n20605), .A2(n20607), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20629), .ZN(n20604) );
  NAND3_X1 U23580 ( .A1(n20900), .A2(n20604), .A3(n20603), .ZN(n20633) );
  INV_X1 U23581 ( .A(n20605), .ZN(n20608) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20633), .B1(
        n20891), .B2(n20632), .ZN(n20609) );
  OAI211_X1 U23583 ( .C1(n20906), .C2(n20666), .A(n20610), .B(n20609), .ZN(
        P1_U3081) );
  OAI22_X1 U23584 ( .A1(n20666), .A2(n20912), .B1(n20974), .B2(n20629), .ZN(
        n20611) );
  INV_X1 U23585 ( .A(n20611), .ZN(n20613) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20633), .B1(
        n20907), .B2(n20632), .ZN(n20612) );
  OAI211_X1 U23587 ( .C1(n20979), .C2(n20630), .A(n20613), .B(n20612), .ZN(
        P1_U3082) );
  OAI22_X1 U23588 ( .A1(n20666), .A2(n20918), .B1(n20981), .B2(n20629), .ZN(
        n20614) );
  INV_X1 U23589 ( .A(n20614), .ZN(n20616) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20633), .B1(
        n20913), .B2(n20632), .ZN(n20615) );
  OAI211_X1 U23591 ( .C1(n20986), .C2(n20630), .A(n20616), .B(n20615), .ZN(
        P1_U3083) );
  OAI22_X1 U23592 ( .A1(n20630), .A2(n20993), .B1(n20988), .B2(n20629), .ZN(
        n20617) );
  INV_X1 U23593 ( .A(n20617), .ZN(n20619) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20633), .B1(
        n20919), .B2(n20632), .ZN(n20618) );
  OAI211_X1 U23595 ( .C1(n20924), .C2(n20666), .A(n20619), .B(n20618), .ZN(
        P1_U3084) );
  OAI22_X1 U23596 ( .A1(n20630), .A2(n21000), .B1(n20995), .B2(n20629), .ZN(
        n20620) );
  INV_X1 U23597 ( .A(n20620), .ZN(n20622) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20633), .B1(
        n20925), .B2(n20632), .ZN(n20621) );
  OAI211_X1 U23599 ( .C1(n20930), .C2(n20666), .A(n20622), .B(n20621), .ZN(
        P1_U3085) );
  OAI22_X1 U23600 ( .A1(n20630), .A2(n21007), .B1(n21002), .B2(n20629), .ZN(
        n20623) );
  INV_X1 U23601 ( .A(n20623), .ZN(n20625) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20633), .B1(
        n20931), .B2(n20632), .ZN(n20624) );
  OAI211_X1 U23603 ( .C1(n20936), .C2(n20666), .A(n20625), .B(n20624), .ZN(
        P1_U3086) );
  OAI22_X1 U23604 ( .A1(n20630), .A2(n21014), .B1(n21009), .B2(n20629), .ZN(
        n20626) );
  INV_X1 U23605 ( .A(n20626), .ZN(n20628) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20633), .B1(
        n20937), .B2(n20632), .ZN(n20627) );
  OAI211_X1 U23607 ( .C1(n20942), .C2(n20666), .A(n20628), .B(n20627), .ZN(
        P1_U3087) );
  OAI22_X1 U23608 ( .A1(n20630), .A2(n21026), .B1(n21018), .B2(n20629), .ZN(
        n20631) );
  INV_X1 U23609 ( .A(n20631), .ZN(n20635) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20633), .B1(
        n20944), .B2(n20632), .ZN(n20634) );
  OAI211_X1 U23611 ( .C1(n20952), .C2(n20666), .A(n20635), .B(n20634), .ZN(
        P1_U3088) );
  NAND2_X1 U23612 ( .A1(n20637), .A2(n20636), .ZN(n20677) );
  INV_X1 U23613 ( .A(n20671), .ZN(n20638) );
  AOI21_X1 U23614 ( .B1(n20639), .B2(n20961), .A(n20638), .ZN(n20645) );
  OR2_X1 U23615 ( .A1(n20645), .A2(n20958), .ZN(n20641) );
  NAND2_X1 U23616 ( .A1(n20648), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20640) );
  OAI22_X1 U23617 ( .A1(n20964), .A2(n20671), .B1(n20963), .B2(n20670), .ZN(
        n20642) );
  INV_X1 U23618 ( .A(n20642), .ZN(n20650) );
  INV_X1 U23619 ( .A(n20888), .ZN(n20643) );
  NOR3_X1 U23620 ( .A1(n20643), .A2(n20958), .A3(n20793), .ZN(n20967) );
  OAI21_X1 U23621 ( .B1(n13603), .B2(n20793), .A(n20826), .ZN(n20644) );
  INV_X1 U23622 ( .A(n20644), .ZN(n20646) );
  OAI21_X1 U23623 ( .B1(n20967), .B2(n20646), .A(n20645), .ZN(n20647) );
  OAI211_X1 U23624 ( .C1(n20826), .C2(n20648), .A(n20966), .B(n20647), .ZN(
        n20674) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20903), .ZN(n20649) );
  OAI211_X1 U23626 ( .C1(n20906), .C2(n20677), .A(n20650), .B(n20649), .ZN(
        P1_U3089) );
  OAI22_X1 U23627 ( .A1(n20974), .A2(n20671), .B1(n20973), .B2(n20670), .ZN(
        n20651) );
  INV_X1 U23628 ( .A(n20651), .ZN(n20653) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20909), .ZN(n20652) );
  OAI211_X1 U23630 ( .C1(n20912), .C2(n20677), .A(n20653), .B(n20652), .ZN(
        P1_U3090) );
  OAI22_X1 U23631 ( .A1(n20981), .A2(n20671), .B1(n20980), .B2(n20670), .ZN(
        n20654) );
  INV_X1 U23632 ( .A(n20654), .ZN(n20656) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20674), .B1(
        n20713), .B2(n20983), .ZN(n20655) );
  OAI211_X1 U23634 ( .C1(n20986), .C2(n20666), .A(n20656), .B(n20655), .ZN(
        P1_U3091) );
  OAI22_X1 U23635 ( .A1(n20988), .A2(n20671), .B1(n20987), .B2(n20670), .ZN(
        n20657) );
  INV_X1 U23636 ( .A(n20657), .ZN(n20659) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20921), .ZN(n20658) );
  OAI211_X1 U23638 ( .C1(n20924), .C2(n20677), .A(n20659), .B(n20658), .ZN(
        P1_U3092) );
  OAI22_X1 U23639 ( .A1(n20995), .A2(n20671), .B1(n20994), .B2(n20670), .ZN(
        n20660) );
  INV_X1 U23640 ( .A(n20660), .ZN(n20662) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20927), .ZN(n20661) );
  OAI211_X1 U23642 ( .C1(n20930), .C2(n20677), .A(n20662), .B(n20661), .ZN(
        P1_U3093) );
  OAI22_X1 U23643 ( .A1(n21002), .A2(n20671), .B1(n21001), .B2(n20670), .ZN(
        n20663) );
  INV_X1 U23644 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20674), .B1(
        n20713), .B2(n21004), .ZN(n20664) );
  OAI211_X1 U23646 ( .C1(n21007), .C2(n20666), .A(n20665), .B(n20664), .ZN(
        P1_U3094) );
  OAI22_X1 U23647 ( .A1(n21009), .A2(n20671), .B1(n21008), .B2(n20670), .ZN(
        n20667) );
  INV_X1 U23648 ( .A(n20667), .ZN(n20669) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20939), .ZN(n20668) );
  OAI211_X1 U23650 ( .C1(n20942), .C2(n20677), .A(n20669), .B(n20668), .ZN(
        P1_U3095) );
  OAI22_X1 U23651 ( .A1(n21018), .A2(n20671), .B1(n21016), .B2(n20670), .ZN(
        n20672) );
  INV_X1 U23652 ( .A(n20672), .ZN(n20676) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20947), .ZN(n20675) );
  OAI211_X1 U23654 ( .C1(n20952), .C2(n20677), .A(n20676), .B(n20675), .ZN(
        P1_U3096) );
  INV_X1 U23655 ( .A(n20797), .ZN(n20678) );
  NAND2_X1 U23656 ( .A1(n20679), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20785) );
  OR2_X1 U23657 ( .A1(n20833), .A2(n20785), .ZN(n20711) );
  AND2_X1 U23658 ( .A1(n20680), .A2(n20831), .ZN(n20787) );
  INV_X1 U23659 ( .A(n20711), .ZN(n20689) );
  AOI21_X1 U23660 ( .B1(n20787), .B2(n14186), .A(n20689), .ZN(n20686) );
  OR2_X1 U23661 ( .A1(n20686), .A2(n20958), .ZN(n20683) );
  AND2_X1 U23662 ( .A1(n20681), .A2(n20747), .ZN(n20835) );
  NAND2_X1 U23663 ( .A1(n20748), .A2(n20835), .ZN(n20682) );
  OAI22_X1 U23664 ( .A1(n20964), .A2(n20711), .B1(n20963), .B2(n20710), .ZN(
        n20684) );
  INV_X1 U23665 ( .A(n20684), .ZN(n20691) );
  INV_X1 U23666 ( .A(n20744), .ZN(n20685) );
  OAI21_X1 U23667 ( .B1(n20685), .B2(n20713), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20687) );
  NAND2_X1 U23668 ( .A1(n20687), .A2(n20686), .ZN(n20688) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20903), .ZN(n20690) );
  OAI211_X1 U23670 ( .C1(n20906), .C2(n20744), .A(n20691), .B(n20690), .ZN(
        P1_U3097) );
  OAI22_X1 U23671 ( .A1(n20974), .A2(n20711), .B1(n20710), .B2(n20973), .ZN(
        n20692) );
  INV_X1 U23672 ( .A(n20692), .ZN(n20694) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20909), .ZN(n20693) );
  OAI211_X1 U23674 ( .C1(n20912), .C2(n20744), .A(n20694), .B(n20693), .ZN(
        P1_U3098) );
  OAI22_X1 U23675 ( .A1(n20981), .A2(n20711), .B1(n20710), .B2(n20980), .ZN(
        n20695) );
  INV_X1 U23676 ( .A(n20695), .ZN(n20697) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20915), .ZN(n20696) );
  OAI211_X1 U23678 ( .C1(n20918), .C2(n20744), .A(n20697), .B(n20696), .ZN(
        P1_U3099) );
  OAI22_X1 U23679 ( .A1(n20988), .A2(n20711), .B1(n20710), .B2(n20987), .ZN(
        n20698) );
  INV_X1 U23680 ( .A(n20698), .ZN(n20700) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20921), .ZN(n20699) );
  OAI211_X1 U23682 ( .C1(n20924), .C2(n20744), .A(n20700), .B(n20699), .ZN(
        P1_U3100) );
  OAI22_X1 U23683 ( .A1(n20995), .A2(n20711), .B1(n20710), .B2(n20994), .ZN(
        n20701) );
  INV_X1 U23684 ( .A(n20701), .ZN(n20703) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20927), .ZN(n20702) );
  OAI211_X1 U23686 ( .C1(n20930), .C2(n20744), .A(n20703), .B(n20702), .ZN(
        P1_U3101) );
  OAI22_X1 U23687 ( .A1(n21002), .A2(n20711), .B1(n20710), .B2(n21001), .ZN(
        n20704) );
  INV_X1 U23688 ( .A(n20704), .ZN(n20706) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20933), .ZN(n20705) );
  OAI211_X1 U23690 ( .C1(n20936), .C2(n20744), .A(n20706), .B(n20705), .ZN(
        P1_U3102) );
  OAI22_X1 U23691 ( .A1(n21009), .A2(n20711), .B1(n20710), .B2(n21008), .ZN(
        n20707) );
  INV_X1 U23692 ( .A(n20707), .ZN(n20709) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20939), .ZN(n20708) );
  OAI211_X1 U23694 ( .C1(n20942), .C2(n20744), .A(n20709), .B(n20708), .ZN(
        P1_U3103) );
  OAI22_X1 U23695 ( .A1(n21018), .A2(n20711), .B1(n20710), .B2(n21016), .ZN(
        n20712) );
  INV_X1 U23696 ( .A(n20712), .ZN(n20716) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20714), .B1(
        n20713), .B2(n20947), .ZN(n20715) );
  OAI211_X1 U23698 ( .C1(n20952), .C2(n20744), .A(n20716), .B(n20715), .ZN(
        P1_U3104) );
  NOR2_X1 U23699 ( .A1(n20785), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20723) );
  INV_X1 U23700 ( .A(n20723), .ZN(n20717) );
  NOR2_X1 U23701 ( .A1(n21321), .A2(n20717), .ZN(n20740) );
  AOI21_X1 U23702 ( .B1(n20787), .B2(n20718), .A(n20740), .ZN(n20721) );
  OR2_X1 U23703 ( .A1(n20721), .A2(n20958), .ZN(n20720) );
  NAND2_X1 U23704 ( .A1(n20723), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20719) );
  NAND2_X1 U23705 ( .A1(n20720), .A2(n20719), .ZN(n20739) );
  AOI22_X1 U23706 ( .A1(n20892), .A2(n20740), .B1(n20891), .B2(n20739), .ZN(
        n20726) );
  OAI21_X1 U23707 ( .B1(n20797), .B2(n20894), .A(n20721), .ZN(n20722) );
  OAI221_X1 U23708 ( .B1(n20826), .B2(n20723), .C1(n20958), .C2(n20722), .A(
        n20966), .ZN(n20741) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n20969), .ZN(n20725) );
  OAI211_X1 U23710 ( .C1(n20972), .C2(n20744), .A(n20726), .B(n20725), .ZN(
        P1_U3105) );
  AOI22_X1 U23711 ( .A1(n20908), .A2(n20740), .B1(n20907), .B2(n20739), .ZN(
        n20728) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n20976), .ZN(n20727) );
  OAI211_X1 U23713 ( .C1(n20979), .C2(n20744), .A(n20728), .B(n20727), .ZN(
        P1_U3106) );
  AOI22_X1 U23714 ( .A1(n20914), .A2(n20740), .B1(n20913), .B2(n20739), .ZN(
        n20730) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n20983), .ZN(n20729) );
  OAI211_X1 U23716 ( .C1(n20986), .C2(n20744), .A(n20730), .B(n20729), .ZN(
        P1_U3107) );
  AOI22_X1 U23717 ( .A1(n20920), .A2(n20740), .B1(n20919), .B2(n20739), .ZN(
        n20732) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n20990), .ZN(n20731) );
  OAI211_X1 U23719 ( .C1(n20993), .C2(n20744), .A(n20732), .B(n20731), .ZN(
        P1_U3108) );
  AOI22_X1 U23720 ( .A1(n20926), .A2(n20740), .B1(n20925), .B2(n20739), .ZN(
        n20734) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n20997), .ZN(n20733) );
  OAI211_X1 U23722 ( .C1(n21000), .C2(n20744), .A(n20734), .B(n20733), .ZN(
        P1_U3109) );
  AOI22_X1 U23723 ( .A1(n20932), .A2(n20740), .B1(n20931), .B2(n20739), .ZN(
        n20736) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n21004), .ZN(n20735) );
  OAI211_X1 U23725 ( .C1(n21007), .C2(n20744), .A(n20736), .B(n20735), .ZN(
        P1_U3110) );
  AOI22_X1 U23726 ( .A1(n20938), .A2(n20740), .B1(n20937), .B2(n20739), .ZN(
        n20738) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n21011), .ZN(n20737) );
  OAI211_X1 U23728 ( .C1(n21014), .C2(n20744), .A(n20738), .B(n20737), .ZN(
        P1_U3111) );
  AOI22_X1 U23729 ( .A1(n20946), .A2(n20740), .B1(n20944), .B2(n20739), .ZN(
        n20743) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20741), .B1(
        n20780), .B2(n21020), .ZN(n20742) );
  OAI211_X1 U23731 ( .C1(n21026), .C2(n20744), .A(n20743), .B(n20742), .ZN(
        P1_U3112) );
  NAND3_X1 U23732 ( .A1(n20824), .A2(n20773), .A3(n20826), .ZN(n20746) );
  NAND2_X1 U23733 ( .A1(n20746), .A2(n20828), .ZN(n20753) );
  AND2_X1 U23734 ( .A1(n20787), .A2(n20896), .ZN(n20751) );
  OR2_X1 U23735 ( .A1(n20747), .A2(n10574), .ZN(n20890) );
  INV_X1 U23736 ( .A(n20890), .ZN(n20749) );
  NOR2_X1 U23737 ( .A1(n20957), .A2(n20785), .ZN(n20794) );
  NAND2_X1 U23738 ( .A1(n21321), .A2(n20794), .ZN(n20778) );
  OAI22_X1 U23739 ( .A1(n20824), .A2(n20906), .B1(n20964), .B2(n20778), .ZN(
        n20750) );
  INV_X1 U23740 ( .A(n20750), .ZN(n20757) );
  INV_X1 U23741 ( .A(n20751), .ZN(n20752) );
  AOI22_X1 U23742 ( .A1(n20753), .A2(n20752), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20778), .ZN(n20754) );
  NAND2_X1 U23743 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20890), .ZN(n20899) );
  NAND3_X1 U23744 ( .A1(n20755), .A2(n20754), .A3(n20899), .ZN(n20781) );
  AOI22_X1 U23745 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20903), .ZN(n20756) );
  OAI211_X1 U23746 ( .C1(n20784), .C2(n20963), .A(n20757), .B(n20756), .ZN(
        P1_U3113) );
  OAI22_X1 U23747 ( .A1(n20824), .A2(n20912), .B1(n20974), .B2(n20778), .ZN(
        n20758) );
  INV_X1 U23748 ( .A(n20758), .ZN(n20760) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20909), .ZN(n20759) );
  OAI211_X1 U23750 ( .C1(n20784), .C2(n20973), .A(n20760), .B(n20759), .ZN(
        P1_U3114) );
  OAI22_X1 U23751 ( .A1(n20824), .A2(n20918), .B1(n20981), .B2(n20778), .ZN(
        n20761) );
  INV_X1 U23752 ( .A(n20761), .ZN(n20763) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20915), .ZN(n20762) );
  OAI211_X1 U23754 ( .C1(n20784), .C2(n20980), .A(n20763), .B(n20762), .ZN(
        P1_U3115) );
  OAI22_X1 U23755 ( .A1(n20773), .A2(n20993), .B1(n20988), .B2(n20778), .ZN(
        n20764) );
  INV_X1 U23756 ( .A(n20764), .ZN(n20766) );
  INV_X1 U23757 ( .A(n20824), .ZN(n20775) );
  AOI22_X1 U23758 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20781), .B1(
        n20775), .B2(n20990), .ZN(n20765) );
  OAI211_X1 U23759 ( .C1(n20784), .C2(n20987), .A(n20766), .B(n20765), .ZN(
        P1_U3116) );
  OAI22_X1 U23760 ( .A1(n20824), .A2(n20930), .B1(n20995), .B2(n20778), .ZN(
        n20767) );
  INV_X1 U23761 ( .A(n20767), .ZN(n20769) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20927), .ZN(n20768) );
  OAI211_X1 U23763 ( .C1(n20784), .C2(n20994), .A(n20769), .B(n20768), .ZN(
        P1_U3117) );
  OAI22_X1 U23764 ( .A1(n20824), .A2(n20936), .B1(n21002), .B2(n20778), .ZN(
        n20770) );
  INV_X1 U23765 ( .A(n20770), .ZN(n20772) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20933), .ZN(n20771) );
  OAI211_X1 U23767 ( .C1(n20784), .C2(n21001), .A(n20772), .B(n20771), .ZN(
        P1_U3118) );
  OAI22_X1 U23768 ( .A1(n20773), .A2(n21014), .B1(n21009), .B2(n20778), .ZN(
        n20774) );
  INV_X1 U23769 ( .A(n20774), .ZN(n20777) );
  AOI22_X1 U23770 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20781), .B1(
        n20775), .B2(n21011), .ZN(n20776) );
  OAI211_X1 U23771 ( .C1(n20784), .C2(n21008), .A(n20777), .B(n20776), .ZN(
        P1_U3119) );
  OAI22_X1 U23772 ( .A1(n20824), .A2(n20952), .B1(n21018), .B2(n20778), .ZN(
        n20779) );
  INV_X1 U23773 ( .A(n20779), .ZN(n20783) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20781), .B1(
        n20780), .B2(n20947), .ZN(n20782) );
  OAI211_X1 U23775 ( .C1(n20784), .C2(n21016), .A(n20783), .B(n20782), .ZN(
        P1_U3120) );
  INV_X1 U23776 ( .A(n20785), .ZN(n20786) );
  NAND2_X1 U23777 ( .A1(n20954), .A2(n20786), .ZN(n20819) );
  NAND2_X1 U23778 ( .A1(n20787), .A2(n20961), .ZN(n20788) );
  NAND2_X1 U23779 ( .A1(n20788), .A2(n20819), .ZN(n20789) );
  NAND2_X1 U23780 ( .A1(n20789), .A2(n20826), .ZN(n20791) );
  NAND2_X1 U23781 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20794), .ZN(n20790) );
  OAI22_X1 U23782 ( .A1(n20964), .A2(n20819), .B1(n20963), .B2(n20818), .ZN(
        n20792) );
  INV_X1 U23783 ( .A(n20792), .ZN(n20799) );
  NOR3_X1 U23784 ( .A1(n20797), .A2(n20958), .A3(n20793), .ZN(n20795) );
  OAI21_X1 U23785 ( .B1(n20795), .B2(n20794), .A(n20966), .ZN(n20821) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n20969), .ZN(n20798) );
  OAI211_X1 U23787 ( .C1(n20972), .C2(n20824), .A(n20799), .B(n20798), .ZN(
        P1_U3121) );
  OAI22_X1 U23788 ( .A1(n20974), .A2(n20819), .B1(n20973), .B2(n20818), .ZN(
        n20800) );
  INV_X1 U23789 ( .A(n20800), .ZN(n20802) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n20976), .ZN(n20801) );
  OAI211_X1 U23791 ( .C1(n20979), .C2(n20824), .A(n20802), .B(n20801), .ZN(
        P1_U3122) );
  OAI22_X1 U23792 ( .A1(n20981), .A2(n20819), .B1(n20980), .B2(n20818), .ZN(
        n20803) );
  INV_X1 U23793 ( .A(n20803), .ZN(n20805) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n20983), .ZN(n20804) );
  OAI211_X1 U23795 ( .C1(n20986), .C2(n20824), .A(n20805), .B(n20804), .ZN(
        P1_U3123) );
  OAI22_X1 U23796 ( .A1(n20988), .A2(n20819), .B1(n20987), .B2(n20818), .ZN(
        n20806) );
  INV_X1 U23797 ( .A(n20806), .ZN(n20808) );
  AOI22_X1 U23798 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n20990), .ZN(n20807) );
  OAI211_X1 U23799 ( .C1(n20993), .C2(n20824), .A(n20808), .B(n20807), .ZN(
        P1_U3124) );
  OAI22_X1 U23800 ( .A1(n20995), .A2(n20819), .B1(n20994), .B2(n20818), .ZN(
        n20809) );
  INV_X1 U23801 ( .A(n20809), .ZN(n20811) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n20997), .ZN(n20810) );
  OAI211_X1 U23803 ( .C1(n21000), .C2(n20824), .A(n20811), .B(n20810), .ZN(
        P1_U3125) );
  OAI22_X1 U23804 ( .A1(n21002), .A2(n20819), .B1(n21001), .B2(n20818), .ZN(
        n20812) );
  INV_X1 U23805 ( .A(n20812), .ZN(n20814) );
  AOI22_X1 U23806 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n21004), .ZN(n20813) );
  OAI211_X1 U23807 ( .C1(n21007), .C2(n20824), .A(n20814), .B(n20813), .ZN(
        P1_U3126) );
  OAI22_X1 U23808 ( .A1(n21009), .A2(n20819), .B1(n21008), .B2(n20818), .ZN(
        n20815) );
  INV_X1 U23809 ( .A(n20815), .ZN(n20817) );
  AOI22_X1 U23810 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n21011), .ZN(n20816) );
  OAI211_X1 U23811 ( .C1(n21014), .C2(n20824), .A(n20817), .B(n20816), .ZN(
        P1_U3127) );
  OAI22_X1 U23812 ( .A1(n21018), .A2(n20819), .B1(n21016), .B2(n20818), .ZN(
        n20820) );
  INV_X1 U23813 ( .A(n20820), .ZN(n20823) );
  AOI22_X1 U23814 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20821), .B1(
        n20855), .B2(n21020), .ZN(n20822) );
  OAI211_X1 U23815 ( .C1(n21026), .C2(n20824), .A(n20823), .B(n20822), .ZN(
        P1_U3128) );
  INV_X1 U23816 ( .A(n20883), .ZN(n20827) );
  NAND3_X1 U23817 ( .A1(n20827), .A2(n20826), .A3(n20825), .ZN(n20829) );
  NAND2_X1 U23818 ( .A1(n20829), .A2(n20828), .ZN(n20838) );
  OR2_X1 U23819 ( .A1(n20831), .A2(n20830), .ZN(n20893) );
  NOR2_X1 U23820 ( .A1(n20893), .A2(n20896), .ZN(n20834) );
  NAND2_X1 U23821 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U23822 ( .A1(n20883), .A2(n20969), .B1(n20892), .B2(n10410), .ZN(
        n20842) );
  INV_X1 U23823 ( .A(n20834), .ZN(n20837) );
  INV_X1 U23824 ( .A(n20835), .ZN(n20836) );
  AOI22_X1 U23825 ( .A1(n20838), .A2(n20837), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20836), .ZN(n20839) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20903), .ZN(n20841) );
  OAI211_X1 U23827 ( .C1(n20859), .C2(n20963), .A(n20842), .B(n20841), .ZN(
        P1_U3129) );
  AOI22_X1 U23828 ( .A1(n20883), .A2(n20976), .B1(n20908), .B2(n10410), .ZN(
        n20844) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20909), .ZN(n20843) );
  OAI211_X1 U23830 ( .C1(n20859), .C2(n20973), .A(n20844), .B(n20843), .ZN(
        P1_U3130) );
  AOI22_X1 U23831 ( .A1(n20883), .A2(n20983), .B1(n20914), .B2(n10410), .ZN(
        n20846) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20915), .ZN(n20845) );
  OAI211_X1 U23833 ( .C1(n20859), .C2(n20980), .A(n20846), .B(n20845), .ZN(
        P1_U3131) );
  AOI22_X1 U23834 ( .A1(n20883), .A2(n20990), .B1(n20920), .B2(n10410), .ZN(
        n20848) );
  AOI22_X1 U23835 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20921), .ZN(n20847) );
  OAI211_X1 U23836 ( .C1(n20859), .C2(n20987), .A(n20848), .B(n20847), .ZN(
        P1_U3132) );
  AOI22_X1 U23837 ( .A1(n20883), .A2(n20997), .B1(n20926), .B2(n10410), .ZN(
        n20850) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20927), .ZN(n20849) );
  OAI211_X1 U23839 ( .C1(n20859), .C2(n20994), .A(n20850), .B(n20849), .ZN(
        P1_U3133) );
  AOI22_X1 U23840 ( .A1(n20883), .A2(n21004), .B1(n20932), .B2(n10410), .ZN(
        n20852) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20933), .ZN(n20851) );
  OAI211_X1 U23842 ( .C1(n20859), .C2(n21001), .A(n20852), .B(n20851), .ZN(
        P1_U3134) );
  AOI22_X1 U23843 ( .A1(n20883), .A2(n21011), .B1(n20938), .B2(n10410), .ZN(
        n20854) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20939), .ZN(n20853) );
  OAI211_X1 U23845 ( .C1(n20859), .C2(n21008), .A(n20854), .B(n20853), .ZN(
        P1_U3135) );
  AOI22_X1 U23846 ( .A1(n20883), .A2(n21020), .B1(n20946), .B2(n10410), .ZN(
        n20858) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20856), .B1(
        n20855), .B2(n20947), .ZN(n20857) );
  OAI211_X1 U23848 ( .C1(n20859), .C2(n21016), .A(n20858), .B(n20857), .ZN(
        P1_U3136) );
  NOR3_X2 U23849 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21321), .A3(
        n20956), .ZN(n20882) );
  INV_X1 U23850 ( .A(n20882), .ZN(n20863) );
  NOR2_X1 U23851 ( .A1(n20956), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20865) );
  INV_X1 U23852 ( .A(n20865), .ZN(n20862) );
  OR2_X1 U23853 ( .A1(n20893), .A2(n20958), .ZN(n20955) );
  OAI222_X1 U23854 ( .A1(n20863), .A2(n20958), .B1(n21030), .B2(n20862), .C1(
        n20861), .C2(n20955), .ZN(n20881) );
  AOI22_X1 U23855 ( .A1(n20892), .A2(n20882), .B1(n20891), .B2(n20881), .ZN(
        n20868) );
  NOR3_X1 U23856 ( .A1(n20864), .A2(n20958), .A3(n20894), .ZN(n20866) );
  OAI21_X1 U23857 ( .B1(n20866), .B2(n20865), .A(n20966), .ZN(n20884) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20903), .ZN(n20867) );
  OAI211_X1 U23859 ( .C1(n20906), .C2(n20902), .A(n20868), .B(n20867), .ZN(
        P1_U3137) );
  AOI22_X1 U23860 ( .A1(n20908), .A2(n20882), .B1(n20907), .B2(n20881), .ZN(
        n20870) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20909), .ZN(n20869) );
  OAI211_X1 U23862 ( .C1(n20912), .C2(n20902), .A(n20870), .B(n20869), .ZN(
        P1_U3138) );
  AOI22_X1 U23863 ( .A1(n20914), .A2(n20882), .B1(n20913), .B2(n20881), .ZN(
        n20872) );
  AOI22_X1 U23864 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20915), .ZN(n20871) );
  OAI211_X1 U23865 ( .C1(n20918), .C2(n20902), .A(n20872), .B(n20871), .ZN(
        P1_U3139) );
  AOI22_X1 U23866 ( .A1(n20920), .A2(n20882), .B1(n20919), .B2(n20881), .ZN(
        n20874) );
  AOI22_X1 U23867 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20921), .ZN(n20873) );
  OAI211_X1 U23868 ( .C1(n20924), .C2(n20902), .A(n20874), .B(n20873), .ZN(
        P1_U3140) );
  AOI22_X1 U23869 ( .A1(n20926), .A2(n20882), .B1(n20925), .B2(n20881), .ZN(
        n20876) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20927), .ZN(n20875) );
  OAI211_X1 U23871 ( .C1(n20930), .C2(n20902), .A(n20876), .B(n20875), .ZN(
        P1_U3141) );
  AOI22_X1 U23872 ( .A1(n20932), .A2(n20882), .B1(n20931), .B2(n20881), .ZN(
        n20878) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20933), .ZN(n20877) );
  OAI211_X1 U23874 ( .C1(n20936), .C2(n20902), .A(n20878), .B(n20877), .ZN(
        P1_U3142) );
  AOI22_X1 U23875 ( .A1(n20938), .A2(n20882), .B1(n20937), .B2(n20881), .ZN(
        n20880) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20939), .ZN(n20879) );
  OAI211_X1 U23877 ( .C1(n20942), .C2(n20902), .A(n20880), .B(n20879), .ZN(
        P1_U3143) );
  AOI22_X1 U23878 ( .A1(n20946), .A2(n20882), .B1(n20944), .B2(n20881), .ZN(
        n20886) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20884), .B1(
        n20883), .B2(n20947), .ZN(n20885) );
  OAI211_X1 U23880 ( .C1(n20952), .C2(n20902), .A(n20886), .B(n20885), .ZN(
        P1_U3144) );
  NOR3_X2 U23881 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20957), .A3(
        n20956), .ZN(n20945) );
  OAI22_X1 U23882 ( .A1(n20955), .A2(n14186), .B1(n20890), .B2(n20889), .ZN(
        n20943) );
  AOI22_X1 U23883 ( .A1(n20892), .A2(n20945), .B1(n20891), .B2(n20943), .ZN(
        n20905) );
  INV_X1 U23884 ( .A(n20893), .ZN(n20897) );
  AOI21_X1 U23885 ( .B1(n20902), .B2(n21025), .A(n20894), .ZN(n20895) );
  AOI21_X1 U23886 ( .B1(n20897), .B2(n20896), .A(n20895), .ZN(n20898) );
  NOR2_X1 U23887 ( .A1(n20898), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20903), .ZN(n20904) );
  OAI211_X1 U23889 ( .C1(n20906), .C2(n21025), .A(n20905), .B(n20904), .ZN(
        P1_U3145) );
  AOI22_X1 U23890 ( .A1(n20908), .A2(n20945), .B1(n20907), .B2(n20943), .ZN(
        n20911) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20909), .ZN(n20910) );
  OAI211_X1 U23892 ( .C1(n20912), .C2(n21025), .A(n20911), .B(n20910), .ZN(
        P1_U3146) );
  AOI22_X1 U23893 ( .A1(n20914), .A2(n20945), .B1(n20913), .B2(n20943), .ZN(
        n20917) );
  AOI22_X1 U23894 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20915), .ZN(n20916) );
  OAI211_X1 U23895 ( .C1(n20918), .C2(n21025), .A(n20917), .B(n20916), .ZN(
        P1_U3147) );
  AOI22_X1 U23896 ( .A1(n20920), .A2(n20945), .B1(n20919), .B2(n20943), .ZN(
        n20923) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20921), .ZN(n20922) );
  OAI211_X1 U23898 ( .C1(n20924), .C2(n21025), .A(n20923), .B(n20922), .ZN(
        P1_U3148) );
  AOI22_X1 U23899 ( .A1(n20926), .A2(n20945), .B1(n20925), .B2(n20943), .ZN(
        n20929) );
  AOI22_X1 U23900 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20927), .ZN(n20928) );
  OAI211_X1 U23901 ( .C1(n20930), .C2(n21025), .A(n20929), .B(n20928), .ZN(
        P1_U3149) );
  AOI22_X1 U23902 ( .A1(n20932), .A2(n20945), .B1(n20931), .B2(n20943), .ZN(
        n20935) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20933), .ZN(n20934) );
  OAI211_X1 U23904 ( .C1(n20936), .C2(n21025), .A(n20935), .B(n20934), .ZN(
        P1_U3150) );
  AOI22_X1 U23905 ( .A1(n20938), .A2(n20945), .B1(n20937), .B2(n20943), .ZN(
        n20941) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20939), .ZN(n20940) );
  OAI211_X1 U23907 ( .C1(n20942), .C2(n21025), .A(n20941), .B(n20940), .ZN(
        P1_U3151) );
  AOI22_X1 U23908 ( .A1(n20946), .A2(n20945), .B1(n20944), .B2(n20943), .ZN(
        n20951) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20949), .B1(
        n20948), .B2(n20947), .ZN(n20950) );
  OAI211_X1 U23910 ( .C1(n20952), .C2(n21025), .A(n20951), .B(n20950), .ZN(
        P1_U3152) );
  INV_X1 U23911 ( .A(n20956), .ZN(n20953) );
  NAND2_X1 U23912 ( .A1(n20954), .A2(n20953), .ZN(n21017) );
  INV_X1 U23913 ( .A(n20955), .ZN(n20962) );
  NOR2_X1 U23914 ( .A1(n20957), .A2(n20956), .ZN(n20968) );
  INV_X1 U23915 ( .A(n20968), .ZN(n20959) );
  OAI22_X1 U23916 ( .A1(n20959), .A2(n21030), .B1(n20958), .B2(n21017), .ZN(
        n20960) );
  AOI21_X1 U23917 ( .B1(n20962), .B2(n20961), .A(n20960), .ZN(n21015) );
  OAI22_X1 U23918 ( .A1(n20964), .A2(n21017), .B1(n20963), .B2(n21015), .ZN(
        n20965) );
  INV_X1 U23919 ( .A(n20965), .ZN(n20971) );
  OAI21_X1 U23920 ( .B1(n20968), .B2(n20967), .A(n20966), .ZN(n21022) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n20969), .ZN(n20970) );
  OAI211_X1 U23922 ( .C1(n20972), .C2(n21025), .A(n20971), .B(n20970), .ZN(
        P1_U3153) );
  OAI22_X1 U23923 ( .A1(n20974), .A2(n21017), .B1(n20973), .B2(n21015), .ZN(
        n20975) );
  INV_X1 U23924 ( .A(n20975), .ZN(n20978) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n20976), .ZN(n20977) );
  OAI211_X1 U23926 ( .C1(n20979), .C2(n21025), .A(n20978), .B(n20977), .ZN(
        P1_U3154) );
  OAI22_X1 U23927 ( .A1(n20981), .A2(n21017), .B1(n20980), .B2(n21015), .ZN(
        n20982) );
  INV_X1 U23928 ( .A(n20982), .ZN(n20985) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n20983), .ZN(n20984) );
  OAI211_X1 U23930 ( .C1(n20986), .C2(n21025), .A(n20985), .B(n20984), .ZN(
        P1_U3155) );
  OAI22_X1 U23931 ( .A1(n20988), .A2(n21017), .B1(n20987), .B2(n21015), .ZN(
        n20989) );
  INV_X1 U23932 ( .A(n20989), .ZN(n20992) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n20990), .ZN(n20991) );
  OAI211_X1 U23934 ( .C1(n20993), .C2(n21025), .A(n20992), .B(n20991), .ZN(
        P1_U3156) );
  OAI22_X1 U23935 ( .A1(n20995), .A2(n21017), .B1(n20994), .B2(n21015), .ZN(
        n20996) );
  INV_X1 U23936 ( .A(n20996), .ZN(n20999) );
  AOI22_X1 U23937 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n20997), .ZN(n20998) );
  OAI211_X1 U23938 ( .C1(n21000), .C2(n21025), .A(n20999), .B(n20998), .ZN(
        P1_U3157) );
  OAI22_X1 U23939 ( .A1(n21002), .A2(n21017), .B1(n21001), .B2(n21015), .ZN(
        n21003) );
  INV_X1 U23940 ( .A(n21003), .ZN(n21006) );
  AOI22_X1 U23941 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n21004), .ZN(n21005) );
  OAI211_X1 U23942 ( .C1(n21007), .C2(n21025), .A(n21006), .B(n21005), .ZN(
        P1_U3158) );
  OAI22_X1 U23943 ( .A1(n21009), .A2(n21017), .B1(n21008), .B2(n21015), .ZN(
        n21010) );
  INV_X1 U23944 ( .A(n21010), .ZN(n21013) );
  AOI22_X1 U23945 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n21011), .ZN(n21012) );
  OAI211_X1 U23946 ( .C1(n21014), .C2(n21025), .A(n21013), .B(n21012), .ZN(
        P1_U3159) );
  OAI22_X1 U23947 ( .A1(n21018), .A2(n21017), .B1(n21016), .B2(n21015), .ZN(
        n21019) );
  INV_X1 U23948 ( .A(n21019), .ZN(n21024) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21022), .B1(
        n21021), .B2(n21020), .ZN(n21023) );
  OAI211_X1 U23950 ( .C1(n21026), .C2(n21025), .A(n21024), .B(n21023), .ZN(
        P1_U3160) );
  NOR2_X1 U23951 ( .A1(n21027), .A2(n21324), .ZN(n21031) );
  INV_X1 U23952 ( .A(n21028), .ZN(n21029) );
  OAI21_X1 U23953 ( .B1(n21031), .B2(n21030), .A(n21029), .ZN(P1_U3163) );
  AND2_X1 U23954 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P1_U3164) );
  AND2_X1 U23955 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21032), .ZN(
        P1_U3165) );
  AND2_X1 U23956 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(
        P1_U3166) );
  AND2_X1 U23957 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21032), .ZN(
        P1_U3167) );
  AND2_X1 U23958 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21032), .ZN(
        P1_U3168) );
  AND2_X1 U23959 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21032), .ZN(
        P1_U3169) );
  AND2_X1 U23960 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_25__SCAN_IN), .ZN(
        P1_U3170) );
  AND2_X1 U23961 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21032), .ZN(
        P1_U3171) );
  AND2_X1 U23962 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21032), .ZN(
        P1_U3172) );
  AND2_X1 U23963 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21032), .ZN(
        P1_U3173) );
  AND2_X1 U23964 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21032), .ZN(
        P1_U3174) );
  AND2_X1 U23965 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21032), .ZN(
        P1_U3175) );
  AND2_X1 U23966 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21032), .ZN(
        P1_U3176) );
  AND2_X1 U23967 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21032), .ZN(
        P1_U3177) );
  AND2_X1 U23968 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21032), .ZN(
        P1_U3178) );
  AND2_X1 U23969 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21032), .ZN(
        P1_U3179) );
  AND2_X1 U23970 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21032), .ZN(
        P1_U3180) );
  AND2_X1 U23971 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21032), .ZN(
        P1_U3181) );
  AND2_X1 U23972 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21032), .ZN(
        P1_U3182) );
  AND2_X1 U23973 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21032), .ZN(
        P1_U3183) );
  AND2_X1 U23974 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P1_U3184) );
  AND2_X1 U23975 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P1_U3185) );
  AND2_X1 U23976 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21032), .ZN(P1_U3186) );
  AND2_X1 U23977 ( .A1(n21032), .A2(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(P1_U3187) );
  AND2_X1 U23978 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21032), .ZN(P1_U3188) );
  AND2_X1 U23979 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21032), .ZN(P1_U3189) );
  AND2_X1 U23980 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21032), .ZN(P1_U3190) );
  AND2_X1 U23981 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21032), .ZN(P1_U3191) );
  AND2_X1 U23982 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21032), .ZN(P1_U3192) );
  AND2_X1 U23983 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21032), .ZN(P1_U3193) );
  NAND2_X1 U23984 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21051), .ZN(n21039) );
  NAND2_X1 U23985 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n21033) );
  OAI211_X1 U23986 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21034), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n21033), .ZN(n21035) );
  INV_X2 U23987 ( .A(n21116), .ZN(n21128) );
  OAI21_X1 U23988 ( .B1(n21036), .B2(n21035), .A(n21128), .ZN(n21037) );
  OAI211_X1 U23989 ( .C1(n21119), .C2(n21039), .A(n21038), .B(n21037), .ZN(
        P1_U3194) );
  NOR3_X1 U23990 ( .A1(NA), .A2(n21043), .A3(n21119), .ZN(n21041) );
  INV_X1 U23991 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21040) );
  OAI22_X1 U23992 ( .A1(n21042), .A2(n21041), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21040), .ZN(n21049) );
  NOR2_X1 U23993 ( .A1(NA), .A2(n21043), .ZN(n21047) );
  INV_X1 U23994 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21045) );
  OAI221_X1 U23995 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(NA), .C1(
        P1_STATE_REG_0__SCAN_IN), .C2(n21045), .A(n21044), .ZN(n21046) );
  OAI221_X1 U23996 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(P1_STATE_REG_2__SCAN_IN), .C2(
        n21047), .A(n21046), .ZN(n21048) );
  OAI21_X1 U23997 ( .B1(n21050), .B2(n21049), .A(n21048), .ZN(P1_U3196) );
  NOR2_X1 U23998 ( .A1(n21128), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21086) );
  INV_X1 U23999 ( .A(n21086), .ZN(n21076) );
  OR2_X1 U24000 ( .A1(n21051), .A2(n21128), .ZN(n21073) );
  INV_X1 U24001 ( .A(n21073), .ZN(n21090) );
  AOI222_X1 U24002 ( .A1(n21089), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21090), .ZN(n21052) );
  INV_X1 U24003 ( .A(n21052), .ZN(P1_U3197) );
  AOI22_X1 U24004 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21128), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21086), .ZN(n21053) );
  OAI21_X1 U24005 ( .B1(n21054), .B2(n21073), .A(n21053), .ZN(P1_U3198) );
  AOI222_X1 U24006 ( .A1(n21090), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21086), .ZN(n21055) );
  INV_X1 U24007 ( .A(n21055), .ZN(P1_U3199) );
  AOI222_X1 U24008 ( .A1(n21090), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n21086), .ZN(n21056) );
  INV_X1 U24009 ( .A(n21056), .ZN(P1_U3200) );
  AOI222_X1 U24010 ( .A1(n21090), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21086), .ZN(n21057) );
  INV_X1 U24011 ( .A(n21057), .ZN(P1_U3201) );
  INV_X1 U24012 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21287) );
  OAI222_X1 U24013 ( .A1(n21073), .A2(n21058), .B1(n21287), .B2(n21116), .C1(
        n21242), .C2(n21076), .ZN(P1_U3202) );
  AOI222_X1 U24014 ( .A1(n21090), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21089), .ZN(n21059) );
  INV_X1 U24015 ( .A(n21059), .ZN(P1_U3203) );
  AOI222_X1 U24016 ( .A1(n21090), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n21089), .ZN(n21060) );
  INV_X1 U24017 ( .A(n21060), .ZN(P1_U3204) );
  AOI222_X1 U24018 ( .A1(n21090), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21089), .ZN(n21061) );
  INV_X1 U24019 ( .A(n21061), .ZN(P1_U3205) );
  AOI222_X1 U24020 ( .A1(n21090), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n21089), .ZN(n21062) );
  INV_X1 U24021 ( .A(n21062), .ZN(P1_U3206) );
  AOI222_X1 U24022 ( .A1(n21090), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21089), .ZN(n21063) );
  INV_X1 U24023 ( .A(n21063), .ZN(P1_U3207) );
  INV_X1 U24024 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21277) );
  OAI222_X1 U24025 ( .A1(n21073), .A2(n21065), .B1(n21277), .B2(n21116), .C1(
        n21064), .C2(n21076), .ZN(P1_U3208) );
  AOI222_X1 U24026 ( .A1(n21090), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21089), .ZN(n21066) );
  INV_X1 U24027 ( .A(n21066), .ZN(P1_U3209) );
  AOI222_X1 U24028 ( .A1(n21089), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21090), .ZN(n21067) );
  INV_X1 U24029 ( .A(n21067), .ZN(P1_U3210) );
  AOI222_X1 U24030 ( .A1(n21090), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21089), .ZN(n21068) );
  INV_X1 U24031 ( .A(n21068), .ZN(P1_U3211) );
  AOI22_X1 U24032 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21128), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21086), .ZN(n21069) );
  OAI21_X1 U24033 ( .B1(n21070), .B2(n21073), .A(n21069), .ZN(P1_U3212) );
  AOI22_X1 U24034 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21128), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21090), .ZN(n21071) );
  OAI21_X1 U24035 ( .B1(n21074), .B2(n21076), .A(n21071), .ZN(P1_U3213) );
  AOI22_X1 U24036 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21128), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21089), .ZN(n21072) );
  OAI21_X1 U24037 ( .B1(n21074), .B2(n21073), .A(n21072), .ZN(P1_U3214) );
  AOI22_X1 U24038 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21128), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21090), .ZN(n21075) );
  OAI21_X1 U24039 ( .B1(n21077), .B2(n21076), .A(n21075), .ZN(P1_U3215) );
  AOI222_X1 U24040 ( .A1(n21090), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21089), .ZN(n21078) );
  INV_X1 U24041 ( .A(n21078), .ZN(P1_U3216) );
  AOI222_X1 U24042 ( .A1(n21090), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21089), .ZN(n21079) );
  INV_X1 U24043 ( .A(n21079), .ZN(P1_U3217) );
  AOI222_X1 U24044 ( .A1(n21090), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21089), .ZN(n21080) );
  INV_X1 U24045 ( .A(n21080), .ZN(P1_U3218) );
  AOI222_X1 U24046 ( .A1(n21090), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n21086), .ZN(n21081) );
  INV_X1 U24047 ( .A(n21081), .ZN(P1_U3219) );
  AOI222_X1 U24048 ( .A1(n21090), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21089), .ZN(n21082) );
  INV_X1 U24049 ( .A(n21082), .ZN(P1_U3220) );
  AOI222_X1 U24050 ( .A1(n21090), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21086), .ZN(n21083) );
  INV_X1 U24051 ( .A(n21083), .ZN(P1_U3221) );
  AOI222_X1 U24052 ( .A1(n21090), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21086), .ZN(n21084) );
  INV_X1 U24053 ( .A(n21084), .ZN(P1_U3222) );
  AOI222_X1 U24054 ( .A1(n21090), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21086), .ZN(n21085) );
  INV_X1 U24055 ( .A(n21085), .ZN(P1_U3223) );
  AOI222_X1 U24056 ( .A1(n21090), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21086), .ZN(n21087) );
  INV_X1 U24057 ( .A(n21087), .ZN(P1_U3224) );
  AOI222_X1 U24058 ( .A1(n21089), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21090), .ZN(n21088) );
  INV_X1 U24059 ( .A(n21088), .ZN(P1_U3225) );
  AOI222_X1 U24060 ( .A1(n21090), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21128), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21089), .ZN(n21091) );
  INV_X1 U24061 ( .A(n21091), .ZN(P1_U3226) );
  OAI22_X1 U24062 ( .A1(n21128), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21116), .ZN(n21092) );
  INV_X1 U24063 ( .A(n21092), .ZN(P1_U3458) );
  OAI22_X1 U24064 ( .A1(n21128), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21116), .ZN(n21093) );
  INV_X1 U24065 ( .A(n21093), .ZN(P1_U3459) );
  OAI22_X1 U24066 ( .A1(n21128), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21116), .ZN(n21094) );
  INV_X1 U24067 ( .A(n21094), .ZN(P1_U3460) );
  OAI22_X1 U24068 ( .A1(n21128), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21116), .ZN(n21095) );
  INV_X1 U24069 ( .A(n21095), .ZN(P1_U3461) );
  OAI21_X1 U24070 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21099), .A(n21097), 
        .ZN(n21096) );
  INV_X1 U24071 ( .A(n21096), .ZN(P1_U3464) );
  OAI21_X1 U24072 ( .B1(n21099), .B2(n21098), .A(n21097), .ZN(P1_U3465) );
  AOI22_X1 U24073 ( .A1(n21103), .A2(n21102), .B1(n21101), .B2(n21100), .ZN(
        n21104) );
  INV_X1 U24074 ( .A(n21104), .ZN(n21106) );
  MUX2_X1 U24075 ( .A(n21106), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21105), .Z(P1_U3469) );
  AOI21_X1 U24076 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21108) );
  AOI22_X1 U24077 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21108), .B2(n21107), .ZN(n21111) );
  INV_X1 U24078 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21110) );
  AOI22_X1 U24079 ( .A1(n21114), .A2(n21111), .B1(n21110), .B2(n21109), .ZN(
        P1_U3481) );
  INV_X1 U24080 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21113) );
  OAI21_X1 U24081 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21114), .ZN(n21112) );
  OAI21_X1 U24082 ( .B1(n21114), .B2(n21113), .A(n21112), .ZN(P1_U3482) );
  AOI22_X1 U24083 ( .A1(n21116), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21115), 
        .B2(n21128), .ZN(P1_U3483) );
  AOI211_X1 U24084 ( .C1(n20332), .C2(n21119), .A(n21118), .B(n21117), .ZN(
        n21127) );
  INV_X1 U24085 ( .A(n21120), .ZN(n21121) );
  NAND3_X1 U24086 ( .A1(n21122), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21121), 
        .ZN(n21124) );
  AOI21_X1 U24087 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21124), .A(n21123), 
        .ZN(n21126) );
  NAND2_X1 U24088 ( .A1(n21127), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21125) );
  OAI21_X1 U24089 ( .B1(n21127), .B2(n21126), .A(n21125), .ZN(P1_U3485) );
  MUX2_X1 U24090 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21128), .Z(P1_U3486) );
  INV_X1 U24091 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n21130) );
  AOI22_X1 U24092 ( .A1(n21131), .A2(keyinput79), .B1(keyinput66), .B2(n21130), 
        .ZN(n21129) );
  OAI221_X1 U24093 ( .B1(n21131), .B2(keyinput79), .C1(n21130), .C2(keyinput66), .A(n21129), .ZN(n21143) );
  INV_X1 U24094 ( .A(keyinput123), .ZN(n21133) );
  AOI22_X1 U24095 ( .A1(n13691), .A2(keyinput45), .B1(P3_LWORD_REG_2__SCAN_IN), 
        .B2(n21133), .ZN(n21132) );
  OAI221_X1 U24096 ( .B1(n13691), .B2(keyinput45), .C1(n21133), .C2(
        P3_LWORD_REG_2__SCAN_IN), .A(n21132), .ZN(n21142) );
  INV_X1 U24097 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n21136) );
  AOI22_X1 U24098 ( .A1(n21136), .A2(keyinput70), .B1(n21135), .B2(keyinput28), 
        .ZN(n21134) );
  OAI221_X1 U24099 ( .B1(n21136), .B2(keyinput70), .C1(n21135), .C2(keyinput28), .A(n21134), .ZN(n21141) );
  NOR4_X1 U24100 ( .A1(n21143), .A2(n21142), .A3(n21141), .A4(n21140), .ZN(
        n21191) );
  AOI22_X1 U24101 ( .A1(n11795), .A2(keyinput17), .B1(keyinput87), .B2(n21145), 
        .ZN(n21144) );
  OAI221_X1 U24102 ( .B1(n11795), .B2(keyinput17), .C1(n21145), .C2(keyinput87), .A(n21144), .ZN(n21157) );
  AOI22_X1 U24103 ( .A1(n21147), .A2(keyinput5), .B1(n12319), .B2(keyinput0), 
        .ZN(n21146) );
  OAI221_X1 U24104 ( .B1(n21147), .B2(keyinput5), .C1(n12319), .C2(keyinput0), 
        .A(n21146), .ZN(n21156) );
  AOI22_X1 U24105 ( .A1(n21150), .A2(keyinput48), .B1(n21149), .B2(keyinput114), .ZN(n21148) );
  OAI221_X1 U24106 ( .B1(n21150), .B2(keyinput48), .C1(n21149), .C2(
        keyinput114), .A(n21148), .ZN(n21155) );
  INV_X1 U24107 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21151) );
  XOR2_X1 U24108 ( .A(n21151), .B(keyinput1), .Z(n21153) );
  XNOR2_X1 U24109 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B(keyinput29), .ZN(
        n21152) );
  NAND2_X1 U24110 ( .A1(n21153), .A2(n21152), .ZN(n21154) );
  NOR4_X1 U24111 ( .A1(n21157), .A2(n21156), .A3(n21155), .A4(n21154), .ZN(
        n21190) );
  INV_X1 U24112 ( .A(keyinput71), .ZN(n21159) );
  AOI22_X1 U24113 ( .A1(n21160), .A2(keyinput24), .B1(P3_LWORD_REG_12__SCAN_IN), .B2(n21159), .ZN(n21158) );
  OAI221_X1 U24114 ( .B1(n21160), .B2(keyinput24), .C1(n21159), .C2(
        P3_LWORD_REG_12__SCAN_IN), .A(n21158), .ZN(n21172) );
  AOI22_X1 U24115 ( .A1(n21163), .A2(keyinput32), .B1(n21162), .B2(keyinput20), 
        .ZN(n21161) );
  OAI221_X1 U24116 ( .B1(n21163), .B2(keyinput32), .C1(n21162), .C2(keyinput20), .A(n21161), .ZN(n21171) );
  INV_X1 U24117 ( .A(keyinput25), .ZN(n21165) );
  AOI22_X1 U24118 ( .A1(n21166), .A2(keyinput104), .B1(
        P1_DATAWIDTH_REG_11__SCAN_IN), .B2(n21165), .ZN(n21164) );
  OAI221_X1 U24119 ( .B1(n21166), .B2(keyinput104), .C1(n21165), .C2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A(n21164), .ZN(n21170) );
  INV_X1 U24120 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21168) );
  AOI22_X1 U24121 ( .A1(n11852), .A2(keyinput31), .B1(keyinput44), .B2(n21168), 
        .ZN(n21167) );
  OAI221_X1 U24122 ( .B1(n11852), .B2(keyinput31), .C1(n21168), .C2(keyinput44), .A(n21167), .ZN(n21169) );
  NOR4_X1 U24123 ( .A1(n21172), .A2(n21171), .A3(n21170), .A4(n21169), .ZN(
        n21189) );
  INV_X1 U24124 ( .A(keyinput84), .ZN(n21174) );
  AOI22_X1 U24125 ( .A1(n21175), .A2(keyinput127), .B1(P2_W_R_N_REG_SCAN_IN), 
        .B2(n21174), .ZN(n21173) );
  OAI221_X1 U24126 ( .B1(n21175), .B2(keyinput127), .C1(n21174), .C2(
        P2_W_R_N_REG_SCAN_IN), .A(n21173), .ZN(n21187) );
  INV_X1 U24127 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21178) );
  INV_X1 U24128 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n21177) );
  AOI22_X1 U24129 ( .A1(n21178), .A2(keyinput22), .B1(n21177), .B2(keyinput69), 
        .ZN(n21176) );
  OAI221_X1 U24130 ( .B1(n21178), .B2(keyinput22), .C1(n21177), .C2(keyinput69), .A(n21176), .ZN(n21186) );
  INV_X1 U24131 ( .A(keyinput8), .ZN(n21180) );
  AOI22_X1 U24132 ( .A1(n21181), .A2(keyinput101), .B1(P3_DATAO_REG_6__SCAN_IN), .B2(n21180), .ZN(n21179) );
  OAI221_X1 U24133 ( .B1(n21181), .B2(keyinput101), .C1(n21180), .C2(
        P3_DATAO_REG_6__SCAN_IN), .A(n21179), .ZN(n21185) );
  INV_X1 U24134 ( .A(DATAI_7_), .ZN(n21183) );
  AOI22_X1 U24135 ( .A1(n21183), .A2(keyinput67), .B1(n11922), .B2(keyinput109), .ZN(n21182) );
  OAI221_X1 U24136 ( .B1(n21183), .B2(keyinput67), .C1(n11922), .C2(
        keyinput109), .A(n21182), .ZN(n21184) );
  NOR4_X1 U24137 ( .A1(n21187), .A2(n21186), .A3(n21185), .A4(n21184), .ZN(
        n21188) );
  NAND4_X1 U24138 ( .A1(n21191), .A2(n21190), .A3(n21189), .A4(n21188), .ZN(
        n21454) );
  INV_X1 U24139 ( .A(keyinput74), .ZN(n21193) );
  AOI22_X1 U24140 ( .A1(n21194), .A2(keyinput98), .B1(
        P1_DATAWIDTH_REG_25__SCAN_IN), .B2(n21193), .ZN(n21192) );
  OAI221_X1 U24141 ( .B1(n21194), .B2(keyinput98), .C1(n21193), .C2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A(n21192), .ZN(n21206) );
  INV_X1 U24142 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n21196) );
  AOI22_X1 U24143 ( .A1(n21197), .A2(keyinput47), .B1(keyinput15), .B2(n21196), 
        .ZN(n21195) );
  OAI221_X1 U24144 ( .B1(n21197), .B2(keyinput47), .C1(n21196), .C2(keyinput15), .A(n21195), .ZN(n21205) );
  INV_X1 U24145 ( .A(keyinput62), .ZN(n21402) );
  AOI22_X1 U24146 ( .A1(n21199), .A2(keyinput94), .B1(
        P1_DATAWIDTH_REG_29__SCAN_IN), .B2(n21402), .ZN(n21198) );
  OAI221_X1 U24147 ( .B1(n21199), .B2(keyinput94), .C1(n21402), .C2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A(n21198), .ZN(n21204) );
  INV_X1 U24148 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21202) );
  AOI22_X1 U24149 ( .A1(n21202), .A2(keyinput111), .B1(n21201), .B2(keyinput65), .ZN(n21200) );
  OAI221_X1 U24150 ( .B1(n21202), .B2(keyinput111), .C1(n21201), .C2(
        keyinput65), .A(n21200), .ZN(n21203) );
  NOR4_X1 U24151 ( .A1(n21206), .A2(n21205), .A3(n21204), .A4(n21203), .ZN(
        n21256) );
  INV_X1 U24152 ( .A(keyinput7), .ZN(n21208) );
  AOI22_X1 U24153 ( .A1(n21209), .A2(keyinput56), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n21208), .ZN(n21207) );
  OAI221_X1 U24154 ( .B1(n21209), .B2(keyinput56), .C1(n21208), .C2(
        P3_ADDRESS_REG_10__SCAN_IN), .A(n21207), .ZN(n21221) );
  INV_X1 U24155 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21211) );
  AOI22_X1 U24156 ( .A1(n21212), .A2(keyinput14), .B1(n21211), .B2(keyinput121), .ZN(n21210) );
  OAI221_X1 U24157 ( .B1(n21212), .B2(keyinput14), .C1(n21211), .C2(
        keyinput121), .A(n21210), .ZN(n21220) );
  AOI22_X1 U24158 ( .A1(n21215), .A2(keyinput19), .B1(n21214), .B2(keyinput96), 
        .ZN(n21213) );
  OAI221_X1 U24159 ( .B1(n21215), .B2(keyinput19), .C1(n21214), .C2(keyinput96), .A(n21213), .ZN(n21219) );
  INV_X1 U24160 ( .A(keyinput10), .ZN(n21217) );
  AOI22_X1 U24161 ( .A1(n13406), .A2(keyinput119), .B1(P3_DATAO_REG_8__SCAN_IN), .B2(n21217), .ZN(n21216) );
  OAI221_X1 U24162 ( .B1(n13406), .B2(keyinput119), .C1(n21217), .C2(
        P3_DATAO_REG_8__SCAN_IN), .A(n21216), .ZN(n21218) );
  NOR4_X1 U24163 ( .A1(n21221), .A2(n21220), .A3(n21219), .A4(n21218), .ZN(
        n21255) );
  AOI22_X1 U24164 ( .A1(n21224), .A2(keyinput42), .B1(keyinput63), .B2(n21223), 
        .ZN(n21222) );
  OAI221_X1 U24165 ( .B1(n21224), .B2(keyinput42), .C1(n21223), .C2(keyinput63), .A(n21222), .ZN(n21236) );
  INV_X1 U24166 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21227) );
  AOI22_X1 U24167 ( .A1(n21227), .A2(keyinput58), .B1(keyinput61), .B2(n21226), 
        .ZN(n21225) );
  OAI221_X1 U24168 ( .B1(n21227), .B2(keyinput58), .C1(n21226), .C2(keyinput61), .A(n21225), .ZN(n21235) );
  AOI22_X1 U24169 ( .A1(n21230), .A2(keyinput59), .B1(n21229), .B2(keyinput105), .ZN(n21228) );
  OAI221_X1 U24170 ( .B1(n21230), .B2(keyinput59), .C1(n21229), .C2(
        keyinput105), .A(n21228), .ZN(n21234) );
  AOI22_X1 U24171 ( .A1(n21232), .A2(keyinput92), .B1(keyinput9), .B2(n11469), 
        .ZN(n21231) );
  OAI221_X1 U24172 ( .B1(n21232), .B2(keyinput92), .C1(n11469), .C2(keyinput9), 
        .A(n21231), .ZN(n21233) );
  NOR4_X1 U24173 ( .A1(n21236), .A2(n21235), .A3(n21234), .A4(n21233), .ZN(
        n21254) );
  INV_X1 U24174 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21239) );
  AOI22_X1 U24175 ( .A1(n21239), .A2(keyinput116), .B1(keyinput50), .B2(n21238), .ZN(n21237) );
  OAI221_X1 U24176 ( .B1(n21239), .B2(keyinput116), .C1(n21238), .C2(
        keyinput50), .A(n21237), .ZN(n21252) );
  INV_X1 U24177 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n21241) );
  AOI22_X1 U24178 ( .A1(n21242), .A2(keyinput54), .B1(keyinput55), .B2(n21241), 
        .ZN(n21240) );
  OAI221_X1 U24179 ( .B1(n21242), .B2(keyinput54), .C1(n21241), .C2(keyinput55), .A(n21240), .ZN(n21251) );
  INV_X1 U24180 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n21245) );
  AOI22_X1 U24181 ( .A1(n21245), .A2(keyinput91), .B1(n21244), .B2(keyinput108), .ZN(n21243) );
  OAI221_X1 U24182 ( .B1(n21245), .B2(keyinput91), .C1(n21244), .C2(
        keyinput108), .A(n21243), .ZN(n21250) );
  INV_X1 U24183 ( .A(DATAI_12_), .ZN(n21248) );
  AOI22_X1 U24184 ( .A1(n21248), .A2(keyinput102), .B1(keyinput112), .B2(
        n21247), .ZN(n21246) );
  OAI221_X1 U24185 ( .B1(n21248), .B2(keyinput102), .C1(n21247), .C2(
        keyinput112), .A(n21246), .ZN(n21249) );
  NOR4_X1 U24186 ( .A1(n21252), .A2(n21251), .A3(n21250), .A4(n21249), .ZN(
        n21253) );
  NAND4_X1 U24187 ( .A1(n21256), .A2(n21255), .A3(n21254), .A4(n21253), .ZN(
        n21453) );
  AOI22_X1 U24188 ( .A1(n21259), .A2(keyinput23), .B1(n21258), .B2(keyinput40), 
        .ZN(n21257) );
  OAI221_X1 U24189 ( .B1(n21259), .B2(keyinput23), .C1(n21258), .C2(keyinput40), .A(n21257), .ZN(n21264) );
  XNOR2_X1 U24190 ( .A(n21260), .B(keyinput36), .ZN(n21263) );
  XNOR2_X1 U24191 ( .A(n21261), .B(keyinput38), .ZN(n21262) );
  OR3_X1 U24192 ( .A1(n21264), .A2(n21263), .A3(n21262), .ZN(n21272) );
  AOI22_X1 U24193 ( .A1(n21266), .A2(keyinput103), .B1(n13339), .B2(keyinput88), .ZN(n21265) );
  OAI221_X1 U24194 ( .B1(n21266), .B2(keyinput103), .C1(n13339), .C2(
        keyinput88), .A(n21265), .ZN(n21271) );
  INV_X1 U24195 ( .A(keyinput39), .ZN(n21268) );
  AOI22_X1 U24196 ( .A1(n21269), .A2(keyinput120), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n21268), .ZN(n21267) );
  OAI221_X1 U24197 ( .B1(n21269), .B2(keyinput120), .C1(n21268), .C2(
        P3_ADDRESS_REG_4__SCAN_IN), .A(n21267), .ZN(n21270) );
  NOR3_X1 U24198 ( .A1(n21272), .A2(n21271), .A3(n21270), .ZN(n21451) );
  AOI22_X1 U24199 ( .A1(n10161), .A2(keyinput89), .B1(n21274), .B2(keyinput11), 
        .ZN(n21273) );
  OAI221_X1 U24200 ( .B1(n10161), .B2(keyinput89), .C1(n21274), .C2(keyinput11), .A(n21273), .ZN(n21285) );
  INV_X1 U24201 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n21276) );
  AOI22_X1 U24202 ( .A1(n21277), .A2(keyinput117), .B1(n21276), .B2(keyinput86), .ZN(n21275) );
  OAI221_X1 U24203 ( .B1(n21277), .B2(keyinput117), .C1(n21276), .C2(
        keyinput86), .A(n21275), .ZN(n21284) );
  AOI22_X1 U24204 ( .A1(n21279), .A2(keyinput100), .B1(keyinput99), .B2(n14529), .ZN(n21278) );
  OAI221_X1 U24205 ( .B1(n21279), .B2(keyinput100), .C1(n14529), .C2(
        keyinput99), .A(n21278), .ZN(n21283) );
  INV_X1 U24206 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n21281) );
  AOI22_X1 U24207 ( .A1(n13046), .A2(keyinput64), .B1(n21281), .B2(keyinput125), .ZN(n21280) );
  OAI221_X1 U24208 ( .B1(n13046), .B2(keyinput64), .C1(n21281), .C2(
        keyinput125), .A(n21280), .ZN(n21282) );
  NOR4_X1 U24209 ( .A1(n21285), .A2(n21284), .A3(n21283), .A4(n21282), .ZN(
        n21450) );
  AOI22_X1 U24210 ( .A1(n21287), .A2(keyinput77), .B1(n10919), .B2(keyinput73), 
        .ZN(n21286) );
  OAI221_X1 U24211 ( .B1(n21287), .B2(keyinput77), .C1(n10919), .C2(keyinput73), .A(n21286), .ZN(n21298) );
  AOI22_X1 U24212 ( .A1(n11976), .A2(keyinput53), .B1(keyinput13), .B2(n21289), 
        .ZN(n21288) );
  OAI221_X1 U24213 ( .B1(n11976), .B2(keyinput53), .C1(n21289), .C2(keyinput13), .A(n21288), .ZN(n21297) );
  INV_X1 U24214 ( .A(DATAI_29_), .ZN(n21291) );
  AOI22_X1 U24215 ( .A1(n11800), .A2(keyinput80), .B1(keyinput51), .B2(n21291), 
        .ZN(n21290) );
  OAI221_X1 U24216 ( .B1(n11800), .B2(keyinput80), .C1(n21291), .C2(keyinput51), .A(n21290), .ZN(n21296) );
  INV_X1 U24217 ( .A(keyinput76), .ZN(n21293) );
  AOI22_X1 U24218 ( .A1(n21294), .A2(keyinput93), .B1(P3_LWORD_REG_7__SCAN_IN), 
        .B2(n21293), .ZN(n21292) );
  OAI221_X1 U24219 ( .B1(n21294), .B2(keyinput93), .C1(n21293), .C2(
        P3_LWORD_REG_7__SCAN_IN), .A(n21292), .ZN(n21295) );
  NOR4_X1 U24220 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21346) );
  INV_X1 U24221 ( .A(keyinput46), .ZN(n21301) );
  INV_X1 U24222 ( .A(keyinput118), .ZN(n21300) );
  AOI22_X1 U24223 ( .A1(n21301), .A2(P3_DATAWIDTH_REG_2__SCAN_IN), .B1(
        P1_DATAWIDTH_REG_10__SCAN_IN), .B2(n21300), .ZN(n21299) );
  OAI221_X1 U24224 ( .B1(n21301), .B2(P3_DATAWIDTH_REG_2__SCAN_IN), .C1(n21300), .C2(P1_DATAWIDTH_REG_10__SCAN_IN), .A(n21299), .ZN(n21314) );
  AOI22_X1 U24225 ( .A1(n21304), .A2(keyinput106), .B1(n21303), .B2(keyinput83), .ZN(n21302) );
  OAI221_X1 U24226 ( .B1(n21304), .B2(keyinput106), .C1(n21303), .C2(
        keyinput83), .A(n21302), .ZN(n21313) );
  INV_X1 U24227 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n21307) );
  INV_X1 U24228 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n21306) );
  AOI22_X1 U24229 ( .A1(n21307), .A2(keyinput107), .B1(keyinput81), .B2(n21306), .ZN(n21305) );
  OAI221_X1 U24230 ( .B1(n21307), .B2(keyinput107), .C1(n21306), .C2(
        keyinput81), .A(n21305), .ZN(n21312) );
  INV_X1 U24231 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21310) );
  INV_X1 U24232 ( .A(keyinput16), .ZN(n21309) );
  AOI22_X1 U24233 ( .A1(n21310), .A2(keyinput60), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n21309), .ZN(n21308) );
  OAI221_X1 U24234 ( .B1(n21310), .B2(keyinput60), .C1(n21309), .C2(
        P3_ADDRESS_REG_26__SCAN_IN), .A(n21308), .ZN(n21311) );
  NOR4_X1 U24235 ( .A1(n21314), .A2(n21313), .A3(n21312), .A4(n21311), .ZN(
        n21345) );
  AOI22_X1 U24236 ( .A1(n21317), .A2(keyinput12), .B1(keyinput3), .B2(n21316), 
        .ZN(n21315) );
  OAI221_X1 U24237 ( .B1(n21317), .B2(keyinput12), .C1(n21316), .C2(keyinput3), 
        .A(n21315), .ZN(n21329) );
  AOI22_X1 U24238 ( .A1(n21319), .A2(keyinput90), .B1(n14427), .B2(keyinput27), 
        .ZN(n21318) );
  OAI221_X1 U24239 ( .B1(n21319), .B2(keyinput90), .C1(n14427), .C2(keyinput27), .A(n21318), .ZN(n21328) );
  AOI22_X1 U24240 ( .A1(n21322), .A2(keyinput122), .B1(keyinput85), .B2(n21321), .ZN(n21320) );
  OAI221_X1 U24241 ( .B1(n21322), .B2(keyinput122), .C1(n21321), .C2(
        keyinput85), .A(n21320), .ZN(n21327) );
  AOI22_X1 U24242 ( .A1(n21325), .A2(keyinput57), .B1(n21324), .B2(keyinput113), .ZN(n21323) );
  OAI221_X1 U24243 ( .B1(n21325), .B2(keyinput57), .C1(n21324), .C2(
        keyinput113), .A(n21323), .ZN(n21326) );
  NOR4_X1 U24244 ( .A1(n21329), .A2(n21328), .A3(n21327), .A4(n21326), .ZN(
        n21344) );
  AOI22_X1 U24245 ( .A1(n21331), .A2(keyinput4), .B1(keyinput21), .B2(n11259), 
        .ZN(n21330) );
  OAI221_X1 U24246 ( .B1(n21331), .B2(keyinput4), .C1(n11259), .C2(keyinput21), 
        .A(n21330), .ZN(n21342) );
  INV_X1 U24247 ( .A(keyinput26), .ZN(n21415) );
  AOI22_X1 U24248 ( .A1(n21333), .A2(keyinput30), .B1(
        P1_DATAWIDTH_REG_31__SCAN_IN), .B2(n21415), .ZN(n21332) );
  OAI221_X1 U24249 ( .B1(n21333), .B2(keyinput30), .C1(n21415), .C2(
        P1_DATAWIDTH_REG_31__SCAN_IN), .A(n21332), .ZN(n21341) );
  AOI22_X1 U24250 ( .A1(n11789), .A2(keyinput52), .B1(keyinput95), .B2(n21338), 
        .ZN(n21337) );
  OAI221_X1 U24251 ( .B1(n11789), .B2(keyinput52), .C1(n21338), .C2(keyinput95), .A(n21337), .ZN(n21339) );
  NOR4_X1 U24252 ( .A1(n21342), .A2(n21341), .A3(n21340), .A4(n21339), .ZN(
        n21343) );
  NAND4_X1 U24253 ( .A1(n21346), .A2(n21345), .A3(n21344), .A4(n21343), .ZN(
        n21380) );
  INV_X1 U24254 ( .A(keyinput34), .ZN(n21351) );
  INV_X1 U24255 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21349) );
  AOI22_X1 U24256 ( .A1(n21349), .A2(keyinput75), .B1(keyinput97), .B2(n21348), 
        .ZN(n21347) );
  OAI221_X1 U24257 ( .B1(n21349), .B2(keyinput75), .C1(n21348), .C2(keyinput97), .A(n21347), .ZN(n21350) );
  AOI221_X1 U24258 ( .B1(keyinput34), .B2(n21352), .C1(n21351), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21350), .ZN(n21370) );
  INV_X1 U24259 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n21354) );
  AOI22_X1 U24260 ( .A1(n21355), .A2(keyinput2), .B1(n21354), .B2(keyinput37), 
        .ZN(n21353) );
  OAI221_X1 U24261 ( .B1(n21355), .B2(keyinput2), .C1(n21354), .C2(keyinput37), 
        .A(n21353), .ZN(n21368) );
  INV_X1 U24262 ( .A(keyinput33), .ZN(n21357) );
  AOI22_X1 U24263 ( .A1(n21358), .A2(keyinput115), .B1(
        P1_DATAWIDTH_REG_8__SCAN_IN), .B2(n21357), .ZN(n21356) );
  OAI221_X1 U24264 ( .B1(n21358), .B2(keyinput115), .C1(n21357), .C2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A(n21356), .ZN(n21367) );
  AOI22_X1 U24265 ( .A1(n21361), .A2(keyinput110), .B1(n21360), .B2(keyinput72), .ZN(n21359) );
  OAI221_X1 U24266 ( .B1(n21361), .B2(keyinput110), .C1(n21360), .C2(
        keyinput72), .A(n21359), .ZN(n21366) );
  INV_X1 U24267 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21363) );
  AOI22_X1 U24268 ( .A1(n21364), .A2(keyinput82), .B1(n21363), .B2(keyinput41), 
        .ZN(n21362) );
  OAI221_X1 U24269 ( .B1(n21364), .B2(keyinput82), .C1(n21363), .C2(keyinput41), .A(n21362), .ZN(n21365) );
  NOR4_X1 U24270 ( .A1(n21368), .A2(n21367), .A3(n21366), .A4(n21365), .ZN(
        n21369) );
  OAI211_X1 U24271 ( .C1(keyinput126), .C2(n21446), .A(n21370), .B(n21369), 
        .ZN(n21379) );
  INV_X1 U24272 ( .A(keyinput43), .ZN(n21372) );
  AOI22_X1 U24273 ( .A1(n11981), .A2(keyinput6), .B1(
        P2_DATAWIDTH_REG_5__SCAN_IN), .B2(n21372), .ZN(n21371) );
  OAI221_X1 U24274 ( .B1(n11981), .B2(keyinput6), .C1(n21372), .C2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A(n21371), .ZN(n21373) );
  INV_X1 U24275 ( .A(n21373), .ZN(n21377) );
  XOR2_X1 U24276 ( .A(keyinput18), .B(n21374), .Z(n21376) );
  XNOR2_X1 U24277 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B(keyinput35), .ZN(
        n21375) );
  NAND3_X1 U24278 ( .A1(n21377), .A2(n21376), .A3(n21375), .ZN(n21378) );
  NOR3_X1 U24279 ( .A1(n21380), .A2(n21379), .A3(n21378), .ZN(n21449) );
  NAND4_X1 U24280 ( .A1(keyinput34), .A2(keyinput18), .A3(keyinput35), .A4(
        keyinput43), .ZN(n21381) );
  NOR2_X1 U24281 ( .A1(keyinput102), .A2(n21381), .ZN(n21393) );
  NAND2_X1 U24282 ( .A1(keyinput36), .A2(keyinput120), .ZN(n21382) );
  NOR3_X1 U24283 ( .A1(keyinput40), .A2(keyinput23), .A3(n21382), .ZN(n21383)
         );
  NAND3_X1 U24284 ( .A1(keyinput88), .A2(keyinput39), .A3(n21383), .ZN(n21391)
         );
  NAND2_X1 U24285 ( .A1(keyinput41), .A2(keyinput2), .ZN(n21384) );
  NOR3_X1 U24286 ( .A1(keyinput115), .A2(keyinput110), .A3(n21384), .ZN(n21389) );
  NOR4_X1 U24287 ( .A1(keyinput6), .A2(keyinput33), .A3(keyinput37), .A4(
        keyinput82), .ZN(n21388) );
  AND4_X1 U24288 ( .A1(keyinput86), .A2(keyinput89), .A3(keyinput11), .A4(
        keyinput64), .ZN(n21387) );
  INV_X1 U24289 ( .A(keyinput72), .ZN(n21385) );
  NOR4_X1 U24290 ( .A1(keyinput125), .A2(keyinput117), .A3(keyinput100), .A4(
        n21385), .ZN(n21386) );
  NAND4_X1 U24291 ( .A1(n21389), .A2(n21388), .A3(n21387), .A4(n21386), .ZN(
        n21390) );
  NOR4_X1 U24292 ( .A1(keyinput99), .A2(keyinput103), .A3(n21391), .A4(n21390), 
        .ZN(n21392) );
  NAND4_X1 U24293 ( .A1(keyinput75), .A2(keyinput97), .A3(n21393), .A4(n21392), 
        .ZN(n21445) );
  NAND2_X1 U24294 ( .A1(keyinput92), .A2(keyinput61), .ZN(n21394) );
  NOR3_X1 U24295 ( .A1(keyinput105), .A2(keyinput59), .A3(n21394), .ZN(n21401)
         );
  NAND2_X1 U24296 ( .A1(keyinput58), .A2(keyinput42), .ZN(n21395) );
  NOR3_X1 U24297 ( .A1(keyinput10), .A2(keyinput63), .A3(n21395), .ZN(n21400)
         );
  NAND2_X1 U24298 ( .A1(keyinput108), .A2(keyinput91), .ZN(n21396) );
  NOR3_X1 U24299 ( .A1(keyinput55), .A2(keyinput112), .A3(n21396), .ZN(n21399)
         );
  INV_X1 U24300 ( .A(keyinput116), .ZN(n21397) );
  NOR4_X1 U24301 ( .A1(keyinput9), .A2(keyinput50), .A3(keyinput54), .A4(
        n21397), .ZN(n21398) );
  NAND4_X1 U24302 ( .A1(n21401), .A2(n21400), .A3(n21399), .A4(n21398), .ZN(
        n21444) );
  NOR4_X1 U24303 ( .A1(keyinput15), .A2(keyinput94), .A3(keyinput111), .A4(
        n21402), .ZN(n21409) );
  NAND2_X1 U24304 ( .A1(keyinput98), .A2(keyinput109), .ZN(n21403) );
  NOR3_X1 U24305 ( .A1(keyinput74), .A2(keyinput47), .A3(n21403), .ZN(n21408)
         );
  NAND2_X1 U24306 ( .A1(keyinput96), .A2(keyinput121), .ZN(n21404) );
  NOR3_X1 U24307 ( .A1(keyinput19), .A2(keyinput119), .A3(n21404), .ZN(n21407)
         );
  NAND2_X1 U24308 ( .A1(keyinput14), .A2(keyinput56), .ZN(n21405) );
  NOR3_X1 U24309 ( .A1(keyinput65), .A2(keyinput7), .A3(n21405), .ZN(n21406)
         );
  NAND4_X1 U24310 ( .A1(n21409), .A2(n21408), .A3(n21407), .A4(n21406), .ZN(
        n21443) );
  NAND2_X1 U24311 ( .A1(keyinput80), .A2(keyinput73), .ZN(n21410) );
  NOR3_X1 U24312 ( .A1(keyinput93), .A2(keyinput76), .A3(n21410), .ZN(n21441)
         );
  INV_X1 U24313 ( .A(keyinput81), .ZN(n21411) );
  NOR4_X1 U24314 ( .A1(keyinput13), .A2(keyinput53), .A3(keyinput77), .A4(
        n21411), .ZN(n21440) );
  INV_X1 U24315 ( .A(keyinput60), .ZN(n21412) );
  NAND4_X1 U24316 ( .A1(keyinput118), .A2(keyinput16), .A3(keyinput107), .A4(
        n21412), .ZN(n21422) );
  NOR2_X1 U24317 ( .A1(keyinput38), .A2(keyinput83), .ZN(n21413) );
  NAND3_X1 U24318 ( .A1(keyinput106), .A2(keyinput46), .A3(n21413), .ZN(n21421) );
  NAND2_X1 U24319 ( .A1(keyinput68), .A2(keyinput21), .ZN(n21414) );
  NOR3_X1 U24320 ( .A1(keyinput95), .A2(keyinput52), .A3(n21414), .ZN(n21419)
         );
  NOR4_X1 U24321 ( .A1(keyinput51), .A2(keyinput30), .A3(keyinput4), .A4(
        n21415), .ZN(n21418) );
  NOR4_X1 U24322 ( .A1(keyinput27), .A2(keyinput12), .A3(keyinput3), .A4(
        keyinput57), .ZN(n21417) );
  AND4_X1 U24323 ( .A1(keyinput78), .A2(keyinput90), .A3(keyinput113), .A4(
        keyinput122), .ZN(n21416) );
  NAND4_X1 U24324 ( .A1(n21419), .A2(n21418), .A3(n21417), .A4(n21416), .ZN(
        n21420) );
  NOR3_X1 U24325 ( .A1(n21422), .A2(n21421), .A3(n21420), .ZN(n21439) );
  INV_X1 U24326 ( .A(keyinput104), .ZN(n21423) );
  NOR4_X1 U24327 ( .A1(keyinput20), .A2(keyinput25), .A3(keyinput31), .A4(
        n21423), .ZN(n21424) );
  NAND3_X1 U24328 ( .A1(keyinput24), .A2(keyinput32), .A3(n21424), .ZN(n21437)
         );
  NOR4_X1 U24329 ( .A1(keyinput29), .A2(keyinput48), .A3(keyinput114), .A4(
        keyinput5), .ZN(n21435) );
  NAND2_X1 U24330 ( .A1(keyinput0), .A2(keyinput124), .ZN(n21425) );
  NOR3_X1 U24331 ( .A1(keyinput1), .A2(keyinput17), .A3(n21425), .ZN(n21434)
         );
  NAND4_X1 U24332 ( .A1(keyinput45), .A2(keyinput70), .A3(keyinput28), .A4(
        keyinput49), .ZN(n21432) );
  NOR2_X1 U24333 ( .A1(keyinput85), .A2(keyinput66), .ZN(n21426) );
  NAND3_X1 U24334 ( .A1(keyinput79), .A2(keyinput123), .A3(n21426), .ZN(n21431) );
  NOR2_X1 U24335 ( .A1(keyinput101), .A2(keyinput67), .ZN(n21427) );
  NAND3_X1 U24336 ( .A1(keyinput69), .A2(keyinput8), .A3(n21427), .ZN(n21430)
         );
  INV_X1 U24337 ( .A(keyinput127), .ZN(n21428) );
  NAND4_X1 U24338 ( .A1(keyinput44), .A2(keyinput84), .A3(keyinput22), .A4(
        n21428), .ZN(n21429) );
  NOR4_X1 U24339 ( .A1(n21432), .A2(n21431), .A3(n21430), .A4(n21429), .ZN(
        n21433) );
  NAND3_X1 U24340 ( .A1(n21435), .A2(n21434), .A3(n21433), .ZN(n21436) );
  NOR4_X1 U24341 ( .A1(keyinput87), .A2(keyinput71), .A3(n21437), .A4(n21436), 
        .ZN(n21438) );
  NAND4_X1 U24342 ( .A1(n21441), .A2(n21440), .A3(n21439), .A4(n21438), .ZN(
        n21442) );
  NOR4_X1 U24343 ( .A1(n21445), .A2(n21444), .A3(n21443), .A4(n21442), .ZN(
        n21447) );
  OAI21_X1 U24344 ( .B1(keyinput126), .B2(n21447), .A(n21446), .ZN(n21448) );
  NAND4_X1 U24345 ( .A1(n21451), .A2(n21450), .A3(n21449), .A4(n21448), .ZN(
        n21452) );
  NOR3_X1 U24346 ( .A1(n21454), .A2(n21453), .A3(n21452), .ZN(n21461) );
  OAI22_X1 U24347 ( .A1(n21458), .A2(n21457), .B1(n21456), .B2(n21455), .ZN(
        n21459) );
  AOI21_X1 U24348 ( .B1(P3_UWORD_REG_3__SCAN_IN), .B2(n17752), .A(n21459), 
        .ZN(n21460) );
  XNOR2_X1 U24349 ( .A(n21461), .B(n21460), .ZN(P3_U2771) );
  INV_X1 U11587 ( .A(n11369), .ZN(n9786) );
  INV_X1 U11298 ( .A(n9789), .ZN(n20141) );
  INV_X2 U11524 ( .A(n15718), .ZN(n17379) );
  INV_X4 U11331 ( .A(n13976), .ZN(n17418) );
  NOR2_X1 U12971 ( .A1(n15862), .A2(n10134), .ZN(n17648) );
  AND2_X1 U14599 ( .A1(n11686), .A2(n12166), .ZN(n12165) );
  BUF_X1 U11202 ( .A(n12381), .Z(n9754) );
  CLKBUF_X2 U11193 ( .A(n11627), .Z(n9813) );
  CLKBUF_X1 U11203 ( .A(n11405), .Z(n9809) );
  CLKBUF_X1 U11218 ( .A(n11694), .Z(n9783) );
  INV_X2 U11225 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16597) );
  CLKBUF_X1 U11227 ( .A(n11627), .Z(n9811) );
  AND2_X1 U11229 ( .A1(n12351), .A2(n10298), .ZN(n12353) );
  CLKBUF_X1 U11253 ( .A(n11627), .Z(n9812) );
  CLKBUF_X1 U11269 ( .A(n10132), .Z(n9784) );
  CLKBUF_X1 U11281 ( .A(n13788), .Z(n9751) );
  NAND2_X1 U11288 ( .A1(n14973), .A2(n14972), .ZN(n14971) );
  NAND2_X1 U11289 ( .A1(n17985), .A2(n17856), .ZN(n18129) );
  CLKBUF_X1 U11311 ( .A(n12665), .Z(n9816) );
  INV_X1 U11338 ( .A(n18129), .ZN(n18119) );
  CLKBUF_X1 U11507 ( .A(n16792), .Z(n16808) );
  INV_X1 U11525 ( .A(n10466), .ZN(n11297) );
endmodule

