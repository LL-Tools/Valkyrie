

module b21_C_AntiSAT_k_256_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418;

  CLKBUF_X2 U4958 ( .A(n5298), .Z(n9045) );
  NAND2_X2 U4959 ( .A1(n6051), .A2(n6050), .ZN(n7647) );
  INV_X1 U4960 ( .A(n5734), .ZN(n5892) );
  CLKBUF_X2 U4961 ( .A(n6793), .Z(n8436) );
  NAND2_X1 U4962 ( .A1(n4588), .A2(n4586), .ZN(n6507) );
  CLKBUF_X1 U4963 ( .A(n8534), .Z(n4453) );
  OAI21_X1 U4964 ( .B1(n6806), .B2(n7261), .A(n8882), .ZN(n8534) );
  AND2_X1 U4965 ( .A1(n7051), .A2(n6514), .ZN(n5215) );
  NAND2_X1 U4966 ( .A1(n9419), .A2(n8260), .ZN(n9409) );
  INV_X2 U4967 ( .A(n8436), .ZN(n8429) );
  INV_X2 U4968 ( .A(n5848), .ZN(n5814) );
  INV_X1 U4969 ( .A(n5846), .ZN(n6600) );
  NAND2_X2 U4970 ( .A1(n5216), .A2(n6555), .ZN(n8161) );
  NAND2_X1 U4971 ( .A1(n6833), .A2(n7051), .ZN(n5374) );
  XNOR2_X1 U4972 ( .A(n5924), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5925) );
  CLKBUF_X2 U4973 ( .A(n4839), .Z(n8163) );
  XNOR2_X1 U4974 ( .A(n4561), .B(n9012), .ZN(n5927) );
  AND2_X1 U4975 ( .A1(n6047), .A2(n6355), .ZN(n4454) );
  XNOR2_X1 U4976 ( .A(n6312), .B(n4921), .ZN(n6748) );
  NAND2_X2 U4977 ( .A1(n7802), .A2(n7801), .ZN(n7916) );
  NAND2_X2 U4978 ( .A1(n7763), .A2(n7764), .ZN(n7802) );
  OR2_X2 U4979 ( .A1(n4914), .A2(n4913), .ZN(n8063) );
  INV_X2 U4980 ( .A(n8063), .ZN(n4457) );
  CLKBUF_X1 U4981 ( .A(n6748), .Z(n4455) );
  XNOR2_X2 U4982 ( .A(n5140), .B(n5139), .ZN(n8349) );
  XNOR2_X1 U4983 ( .A(n8436), .B(n4457), .ZN(n4918) );
  INV_X2 U4985 ( .A(n4460), .ZN(n4919) );
  MUX2_X1 U4986 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5136), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5138) );
  CLKBUF_X2 U4987 ( .A(n6464), .Z(n4460) );
  NAND2_X4 U4988 ( .A1(n6508), .A2(n6507), .ZN(n6902) );
  INV_X2 U4989 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI211_X1 U4990 ( .C1(n9445), .C2(n10212), .A(n8056), .B(n8055), .ZN(n8057)
         );
  AND2_X1 U4991 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  AOI21_X1 U4992 ( .B1(n8054), .B2(n9985), .A(n8053), .ZN(n9447) );
  NOR2_X1 U4993 ( .A1(n4609), .A2(n4607), .ZN(n4606) );
  OAI21_X1 U4994 ( .B1(n9321), .B2(n4827), .A(n4825), .ZN(n9272) );
  INV_X1 U4995 ( .A(n4820), .ZN(n4819) );
  NAND2_X1 U4996 ( .A1(n4828), .A2(n8329), .ZN(n4823) );
  OAI21_X1 U4997 ( .B1(n8835), .B2(n6399), .A(n6466), .ZN(n8819) );
  NAND2_X1 U4998 ( .A1(n6065), .A2(n6064), .ZN(n7734) );
  NAND2_X1 U4999 ( .A1(n6102), .A2(n6101), .ZN(n8977) );
  NAND2_X1 U5000 ( .A1(n6090), .A2(n6089), .ZN(n8984) );
  NAND2_X1 U5001 ( .A1(n6981), .A2(n6982), .ZN(n6980) );
  AOI21_X1 U5002 ( .B1(n7151), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7150), .ZN(
        n7152) );
  NAND2_X1 U5003 ( .A1(n6038), .A2(n6037), .ZN(n7630) );
  NAND2_X1 U5004 ( .A1(n4662), .A2(n8232), .ZN(n7414) );
  NAND2_X1 U5005 ( .A1(n6998), .A2(n8312), .ZN(n7447) );
  INV_X2 U5006 ( .A(n10279), .ZN(n4456) );
  AND2_X1 U5007 ( .A1(n6942), .A2(n6791), .ZN(n6797) );
  AND2_X1 U5008 ( .A1(n6330), .A2(n6335), .ZN(n6753) );
  NAND2_X1 U5009 ( .A1(n4551), .A2(n5304), .ZN(n5320) );
  INV_X2 U5010 ( .A(n5175), .ZN(n9049) );
  AND3_X1 U5011 ( .A1(n5985), .A2(n4571), .A3(n5984), .ZN(n7368) );
  NAND2_X1 U5012 ( .A1(n5254), .A2(n5253), .ZN(n5276) );
  NAND4_X1 U5013 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n6946)
         );
  INV_X1 U5014 ( .A(n6944), .ZN(n7025) );
  INV_X2 U5015 ( .A(n4465), .ZN(n5928) );
  INV_X4 U5016 ( .A(n8161), .ZN(n4841) );
  INV_X2 U5017 ( .A(n6285), .ZN(n6258) );
  CLKBUF_X2 U5018 ( .A(n6026), .Z(n4465) );
  INV_X1 U5019 ( .A(n6026), .ZN(n4464) );
  AND2_X2 U5020 ( .A1(n5926), .A2(n9020), .ZN(n6285) );
  XNOR2_X1 U5021 ( .A(n5147), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9342) );
  INV_X2 U5022 ( .A(n5216), .ZN(n4458) );
  INV_X1 U5023 ( .A(n5925), .ZN(n9020) );
  NAND2_X1 U5024 ( .A1(n5153), .A2(n9882), .ZN(n9887) );
  INV_X2 U5025 ( .A(n7950), .ZN(n4459) );
  AND2_X1 U5026 ( .A1(n6158), .A2(n6157), .ZN(n6310) );
  OR2_X1 U5027 ( .A1(n6294), .A2(n6156), .ZN(n6158) );
  INV_X1 U5028 ( .A(n5128), .ZN(n5255) );
  NAND2_X1 U5029 ( .A1(n4990), .A2(n4989), .ZN(n5128) );
  AND3_X1 U5030 ( .A1(n5089), .A2(n5247), .A3(n4499), .ZN(n5068) );
  NAND2_X1 U5031 ( .A1(n5125), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4989) );
  AND3_X1 U5032 ( .A1(n4584), .A2(n4578), .A3(n4577), .ZN(n4581) );
  AND2_X1 U5033 ( .A1(n10290), .A2(n4936), .ZN(n5956) );
  AND2_X1 U5034 ( .A1(n5922), .A2(n5028), .ZN(n5027) );
  INV_X1 U5035 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5110) );
  INV_X1 U5036 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5933) );
  INV_X1 U5037 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5595) );
  NOR2_X1 U5038 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4583) );
  NOR2_X1 U5039 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4582) );
  NOR2_X1 U5040 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4584) );
  NOR2_X1 U5041 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4578) );
  NOR2_X1 U5042 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4577) );
  NOR2_X1 U5043 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5087) );
  NOR2_X1 U5044 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5088) );
  NOR2_X1 U5045 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4585) );
  NOR2_X1 U5046 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6123) );
  INV_X1 U5047 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5105) );
  INV_X4 U5048 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5049 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U5050 ( .A1(n6902), .A2(n6556), .ZN(n4461) );
  NAND2_X1 U5051 ( .A1(n6902), .A2(n6556), .ZN(n4462) );
  NAND2_X1 U5052 ( .A1(n6902), .A2(n6556), .ZN(n5976) );
  NAND2_X1 U5053 ( .A1(n5926), .A2(n5925), .ZN(n4463) );
  AOI21_X2 U5054 ( .B1(n8843), .B2(n6148), .A(n6147), .ZN(n8835) );
  NAND2_X1 U5055 ( .A1(n5927), .A2(n9020), .ZN(n6026) );
  AOI21_X1 U5056 ( .B1(n4768), .B2(n4770), .A(n4767), .ZN(n4766) );
  INV_X1 U5057 ( .A(n5700), .ZN(n4767) );
  INV_X1 U5058 ( .A(n4772), .ZN(n4768) );
  NAND2_X1 U5059 ( .A1(n5592), .A2(n4971), .ZN(n4970) );
  NOR2_X1 U5060 ( .A1(n5620), .A2(n4972), .ZN(n4971) );
  INV_X1 U5061 ( .A(n5591), .ZN(n4972) );
  INV_X1 U5062 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5026) );
  AND2_X1 U5063 ( .A1(n5092), .A2(n4480), .ZN(n5145) );
  OAI211_X1 U5064 ( .C1(n7414), .C2(n8170), .A(n8187), .B(n4660), .ZN(n8084)
         );
  NAND2_X1 U5065 ( .A1(n4661), .A2(n8170), .ZN(n4660) );
  INV_X1 U5066 ( .A(n4662), .ZN(n4661) );
  OAI21_X1 U5067 ( .B1(n6337), .B2(n6331), .A(n4697), .ZN(n6332) );
  NAND2_X1 U5068 ( .A1(n4574), .A2(n4680), .ZN(n6359) );
  INV_X1 U5069 ( .A(n6341), .ZN(n4680) );
  NAND2_X1 U5070 ( .A1(n4575), .A2(n6342), .ZN(n4574) );
  MUX2_X1 U5071 ( .A(n8130), .B(n8129), .S(n8170), .Z(n8132) );
  NOR2_X1 U5072 ( .A1(n6433), .A2(n8728), .ZN(n6441) );
  MUX2_X1 U5073 ( .A(n6432), .B(n6431), .S(n6430), .Z(n6433) );
  NAND2_X1 U5074 ( .A1(n6743), .A2(n8063), .ZN(n6324) );
  NOR2_X1 U5075 ( .A1(n5458), .A2(n4979), .ZN(n4978) );
  INV_X1 U5076 ( .A(n5439), .ZN(n4979) );
  INV_X1 U5077 ( .A(n7915), .ZN(n4951) );
  OR2_X1 U5078 ( .A1(n8900), .A2(n8444), .ZN(n6452) );
  NAND2_X1 U5079 ( .A1(n8714), .A2(n4632), .ZN(n4631) );
  AOI21_X1 U5080 ( .B1(n5001), .B2(n4999), .A(n4506), .ZN(n4998) );
  INV_X1 U5081 ( .A(n5003), .ZN(n4999) );
  INV_X1 U5082 ( .A(n5001), .ZN(n5000) );
  OR2_X1 U5083 ( .A1(n8977), .A2(n7805), .ZN(n6377) );
  OAI21_X1 U5084 ( .B1(n7652), .B2(n5012), .A(n7810), .ZN(n5011) );
  INV_X1 U5085 ( .A(n7666), .ZN(n6747) );
  NAND2_X1 U5086 ( .A1(n7368), .A2(n7468), .ZN(n6474) );
  NAND2_X1 U5087 ( .A1(n8566), .A2(n7122), .ZN(n6473) );
  INV_X1 U5088 ( .A(n6756), .ZN(n6743) );
  NAND2_X1 U5089 ( .A1(n6463), .A2(n7666), .ZN(n6804) );
  NOR2_X1 U5090 ( .A1(n9085), .A2(n5052), .ZN(n5051) );
  INV_X1 U5091 ( .A(n5564), .ZN(n5052) );
  INV_X1 U5092 ( .A(n9887), .ZN(n4657) );
  INV_X1 U5093 ( .A(n8139), .ZN(n4832) );
  NOR2_X1 U5094 ( .A1(n4910), .A2(n8027), .ZN(n4909) );
  INV_X1 U5095 ( .A(n9288), .ZN(n4910) );
  NOR2_X1 U5096 ( .A1(n7710), .A2(n7679), .ZN(n4804) );
  INV_X1 U5097 ( .A(n7412), .ZN(n4902) );
  XNOR2_X1 U5098 ( .A(n6302), .B(n6301), .ZN(n6300) );
  OAI21_X1 U5099 ( .B1(n5807), .B2(n5806), .A(n5805), .ZN(n5834) );
  AND2_X1 U5100 ( .A1(n5835), .A2(n5811), .ZN(n5833) );
  INV_X1 U5101 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5132) );
  NOR2_X1 U5102 ( .A1(n5107), .A2(n5106), .ZN(n5108) );
  INV_X1 U5103 ( .A(SI_21_), .ZN(n5703) );
  INV_X1 U5104 ( .A(n4770), .ZN(n4769) );
  AND2_X1 U5105 ( .A1(n4968), .A2(n4773), .ZN(n4772) );
  INV_X1 U5106 ( .A(n5664), .ZN(n4773) );
  AOI21_X1 U5107 ( .B1(n4772), .B2(n5641), .A(n4771), .ZN(n4770) );
  INV_X1 U5108 ( .A(n5663), .ZN(n4771) );
  AND2_X1 U5109 ( .A1(n5702), .A2(n5669), .ZN(n5700) );
  NAND2_X1 U5110 ( .A1(n4784), .A2(n4489), .ZN(n4783) );
  NOR2_X1 U5111 ( .A1(n5540), .A2(n4789), .ZN(n4788) );
  INV_X1 U5112 ( .A(n5511), .ZN(n4789) );
  INV_X1 U5113 ( .A(n5513), .ZN(n5092) );
  AND3_X1 U5114 ( .A1(n5031), .A2(n5030), .A3(n5029), .ZN(n5089) );
  NOR2_X1 U5115 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5031) );
  NOR2_X1 U5116 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5030) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5029) );
  NAND2_X1 U5118 ( .A1(n4778), .A2(n4779), .ZN(n5416) );
  INV_X1 U5119 ( .A(n4780), .ZN(n4779) );
  OR2_X1 U5120 ( .A1(n7917), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U5121 ( .A1(n7917), .A2(n4951), .ZN(n4949) );
  NAND2_X1 U5122 ( .A1(n6174), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6183) );
  INV_X1 U5123 ( .A(n6175), .ZN(n6174) );
  NAND2_X1 U5124 ( .A1(n4920), .A2(n6747), .ZN(n6784) );
  NAND2_X1 U5125 ( .A1(n6748), .A2(n4919), .ZN(n6798) );
  INV_X1 U5126 ( .A(n5969), .ZN(n5948) );
  CLKBUF_X1 U5127 ( .A(n5969), .Z(n6287) );
  NAND2_X1 U5128 ( .A1(n5927), .A2(n5925), .ZN(n5969) );
  NAND2_X1 U5129 ( .A1(n8817), .A2(n7988), .ZN(n7990) );
  OR2_X1 U5130 ( .A1(n8951), .A2(n8836), .ZN(n7988) );
  OAI21_X1 U5131 ( .B1(n5006), .B2(n4596), .A(n4594), .ZN(n8866) );
  INV_X1 U5132 ( .A(n4595), .ZN(n4594) );
  AND2_X1 U5133 ( .A1(n6086), .A2(n7785), .ZN(n4637) );
  INV_X1 U5134 ( .A(n4641), .ZN(n4639) );
  OAI21_X1 U5135 ( .B1(n6088), .B2(n4642), .A(n6098), .ZN(n4641) );
  INV_X1 U5136 ( .A(n5976), .ZN(n6159) );
  INV_X1 U5137 ( .A(n6902), .ZN(n6584) );
  NAND2_X1 U5138 ( .A1(n6902), .A2(n6555), .ZN(n5975) );
  OR2_X1 U5139 ( .A1(n10301), .A2(n6738), .ZN(n7032) );
  INV_X1 U5140 ( .A(n5027), .ZN(n4870) );
  AND2_X1 U5141 ( .A1(n4991), .A2(n4582), .ZN(n4580) );
  AND2_X1 U5142 ( .A1(n4585), .A2(n4583), .ZN(n4579) );
  INV_X1 U5143 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4991) );
  AOI21_X1 U5144 ( .B1(n4719), .B2(n4721), .A(n5057), .ZN(n4717) );
  NAND2_X2 U5145 ( .A1(n5886), .A2(n8349), .ZN(n5216) );
  AND2_X1 U5146 ( .A1(n9438), .A2(n8173), .ZN(n8339) );
  NAND2_X1 U5147 ( .A1(n4658), .A2(n4657), .ZN(n5895) );
  AOI21_X1 U5148 ( .B1(n6654), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6650), .ZN(
        n6651) );
  OR2_X1 U5149 ( .A1(n9465), .A2(n9104), .ZN(n9271) );
  OR2_X1 U5150 ( .A1(n9465), .A2(n9306), .ZN(n4912) );
  NAND2_X1 U5151 ( .A1(n7877), .A2(n8201), .ZN(n4876) );
  INV_X1 U5152 ( .A(n9985), .ZN(n9421) );
  XNOR2_X1 U5153 ( .A(n6838), .B(n8305), .ZN(n8182) );
  NAND2_X1 U5154 ( .A1(n7944), .A2(n5120), .ZN(n6514) );
  NAND2_X1 U5155 ( .A1(n5154), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5155) );
  XNOR2_X1 U5156 ( .A(n4794), .B(n5781), .ZN(n7823) );
  OAI21_X1 U5157 ( .B1(n5745), .B2(n4964), .A(n4961), .ZN(n4794) );
  AND2_X1 U5158 ( .A1(n5764), .A2(n5749), .ZN(n5762) );
  AOI21_X1 U5159 ( .B1(n5096), .B2(P1_IR_REG_31__SCAN_IN), .A(n4709), .ZN(
        n4708) );
  NAND2_X1 U5160 ( .A1(n4710), .A2(n5097), .ZN(n4709) );
  NAND2_X1 U5161 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4710) );
  NAND2_X1 U5163 ( .A1(n8080), .A2(n8320), .ZN(n4676) );
  NAND2_X1 U5164 ( .A1(n4700), .A2(n4698), .ZN(n6337) );
  MUX2_X1 U5165 ( .A(n8095), .B(n8094), .S(n8170), .Z(n8108) );
  MUX2_X1 U5166 ( .A(n6364), .B(n6363), .S(n6432), .Z(n6365) );
  NAND2_X1 U5167 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  INV_X1 U5168 ( .A(n6366), .ZN(n4707) );
  NOR2_X1 U5169 ( .A1(n6372), .A2(n4642), .ZN(n4704) );
  INV_X1 U5170 ( .A(n6412), .ZN(n4565) );
  AOI21_X1 U5171 ( .B1(n4495), .B2(n4566), .A(n6397), .ZN(n6413) );
  NOR2_X1 U5172 ( .A1(n8845), .A2(n6392), .ZN(n4566) );
  OAI21_X1 U5173 ( .B1(n8132), .B2(n8131), .A(n8133), .ZN(n4673) );
  AOI21_X1 U5174 ( .B1(n8132), .B2(n8268), .A(n4671), .ZN(n4670) );
  INV_X1 U5175 ( .A(n6440), .ZN(n4694) );
  INV_X1 U5176 ( .A(n4689), .ZN(n4688) );
  INV_X1 U5177 ( .A(n7621), .ZN(n4926) );
  INV_X1 U5178 ( .A(n6486), .ZN(n4695) );
  NAND2_X1 U5179 ( .A1(n4696), .A2(n4690), .ZN(n4689) );
  NAND2_X1 U5180 ( .A1(n6451), .A2(n4691), .ZN(n4690) );
  NOR2_X1 U5181 ( .A1(n6450), .A2(n8369), .ZN(n4696) );
  NAND2_X1 U5182 ( .A1(n7996), .A2(n6439), .ZN(n4691) );
  OR2_X1 U5183 ( .A1(n4668), .A2(n9255), .ZN(n4667) );
  NOR2_X1 U5184 ( .A1(n9485), .A2(n9489), .ZN(n4810) );
  AND2_X1 U5185 ( .A1(n4967), .A2(n5762), .ZN(n4966) );
  NAND2_X1 U5186 ( .A1(n5744), .A2(n5743), .ZN(n4967) );
  INV_X1 U5187 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5487) );
  AND2_X1 U5188 ( .A1(n4973), .A2(n5381), .ZN(n4775) );
  NOR2_X1 U5189 ( .A1(n4977), .A2(n4974), .ZN(n4973) );
  INV_X1 U5190 ( .A(n5415), .ZN(n4974) );
  INV_X1 U5191 ( .A(n4978), .ZN(n4977) );
  INV_X1 U5192 ( .A(n5080), .ZN(n4976) );
  INV_X1 U5193 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5440) );
  OAI21_X1 U5194 ( .B1(n5380), .B2(n4781), .A(n5082), .ZN(n4780) );
  NAND2_X1 U5195 ( .A1(n4922), .A2(n7270), .ZN(n6793) );
  NAND2_X1 U5196 ( .A1(n4515), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U5197 ( .A1(n4856), .A2(n6299), .ZN(n4649) );
  OAI21_X1 U5198 ( .B1(n6454), .B2(n4646), .A(n6457), .ZN(n4645) );
  NAND2_X1 U5199 ( .A1(n4857), .A2(n6299), .ZN(n4646) );
  OR2_X1 U5200 ( .A1(n8909), .A2(n8443), .ZN(n6247) );
  NAND2_X1 U5201 ( .A1(n4633), .A2(n4475), .ZN(n8713) );
  NAND2_X1 U5202 ( .A1(n8756), .A2(n4893), .ZN(n4633) );
  AND2_X1 U5203 ( .A1(n4895), .A2(n4899), .ZN(n4893) );
  AOI21_X1 U5204 ( .B1(n5019), .B2(n5018), .A(n7994), .ZN(n5017) );
  NOR2_X1 U5205 ( .A1(n8924), .A2(n7993), .ZN(n7994) );
  NOR2_X1 U5206 ( .A1(n8924), .A2(n4750), .ZN(n4749) );
  INV_X1 U5207 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U5208 ( .A1(n5010), .A2(n7811), .ZN(n5009) );
  NOR2_X1 U5209 ( .A1(n4760), .A2(n7647), .ZN(n4759) );
  INV_X1 U5210 ( .A(n4761), .ZN(n4760) );
  NOR2_X1 U5211 ( .A1(n7630), .A2(n7479), .ZN(n4761) );
  OAI22_X1 U5212 ( .A1(n7067), .A2(n6258), .B1(n5968), .B2(n7011), .ZN(n4572)
         );
  OR3_X1 U5213 ( .A1(n7825), .A2(n7929), .A3(n7949), .ZN(n6812) );
  OAI21_X1 U5214 ( .B1(n6313), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6493) );
  AND2_X1 U5215 ( .A1(n5070), .A2(n4958), .ZN(n4957) );
  NOR2_X1 U5216 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4958) );
  INV_X1 U5217 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6122) );
  INV_X1 U5218 ( .A(n5483), .ZN(n5058) );
  NOR2_X1 U5219 ( .A1(n5043), .A2(n9101), .ZN(n5039) );
  INV_X1 U5220 ( .A(n5045), .ZN(n5043) );
  NOR2_X1 U5221 ( .A1(n5046), .A2(n9148), .ZN(n5045) );
  INV_X1 U5222 ( .A(n9076), .ZN(n5046) );
  NAND2_X1 U5223 ( .A1(n4714), .A2(n4716), .ZN(n4711) );
  NOR2_X1 U5224 ( .A1(n9193), .A2(n10128), .ZN(n9194) );
  NOR2_X1 U5225 ( .A1(n9451), .A2(n4798), .ZN(n4797) );
  INV_X1 U5226 ( .A(n4799), .ZN(n4798) );
  INV_X1 U5227 ( .A(n4912), .ZN(n4908) );
  INV_X1 U5228 ( .A(n8024), .ZN(n4862) );
  OR2_X1 U5229 ( .A1(n9485), .A2(n9324), .ZN(n8274) );
  OR2_X1 U5230 ( .A1(n9510), .A2(n10009), .ZN(n4814) );
  INV_X1 U5231 ( .A(n4874), .ZN(n4873) );
  OAI21_X1 U5232 ( .B1(n9996), .B2(n4875), .A(n8010), .ZN(n4874) );
  INV_X1 U5233 ( .A(n8009), .ZN(n4875) );
  OR2_X1 U5234 ( .A1(n10009), .A2(n9422), .ZN(n8257) );
  OR2_X1 U5235 ( .A1(n7941), .A2(n7905), .ZN(n8250) );
  NAND2_X1 U5236 ( .A1(n4804), .A2(n4803), .ZN(n4802) );
  NAND2_X1 U5237 ( .A1(n4651), .A2(n10211), .ZN(n4653) );
  INV_X1 U5238 ( .A(n6606), .ZN(n4651) );
  OR2_X1 U5239 ( .A1(n7563), .A2(n7594), .ZN(n7564) );
  INV_X1 U5240 ( .A(n6559), .ZN(n4838) );
  NAND2_X1 U5241 ( .A1(n4458), .A2(n6531), .ZN(n4836) );
  AND2_X1 U5242 ( .A1(n5066), .A2(n5065), .ZN(n5064) );
  INV_X1 U5243 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U5244 ( .A1(n6263), .A2(n6262), .ZN(n4986) );
  AND2_X1 U5245 ( .A1(n4737), .A2(n5105), .ZN(n4736) );
  INV_X1 U5246 ( .A(SI_10_), .ZN(n5417) );
  NAND2_X1 U5247 ( .A1(n5356), .A2(n5355), .ZN(n5378) );
  OR2_X1 U5248 ( .A1(n6798), .A2(n6804), .ZN(n6944) );
  INV_X1 U5249 ( .A(n6130), .ZN(n6128) );
  INV_X1 U5250 ( .A(n4949), .ZN(n4948) );
  AND2_X1 U5251 ( .A1(n7919), .A2(n4946), .ZN(n4945) );
  NAND2_X1 U5252 ( .A1(n4947), .A2(n4949), .ZN(n4946) );
  INV_X1 U5253 ( .A(n8468), .ZN(n4942) );
  OR2_X1 U5254 ( .A1(n6183), .A2(n8476), .ZN(n6192) );
  NOR2_X1 U5255 ( .A1(n6809), .A2(n10293), .ZN(n6803) );
  OR2_X1 U5256 ( .A1(n5969), .A2(n10359), .ZN(n5941) );
  AND2_X1 U5257 ( .A1(n5072), .A2(n5940), .ZN(n5943) );
  OR2_X1 U5258 ( .A1(n8719), .A2(n4739), .ZN(n8689) );
  NAND2_X1 U5259 ( .A1(n8691), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U5260 ( .A1(n6268), .A2(n6267), .ZN(n8900) );
  NOR2_X1 U5261 ( .A1(n8719), .A2(n4738), .ZN(n8690) );
  INV_X1 U5262 ( .A(n4740), .ZN(n4738) );
  AOI21_X1 U5263 ( .B1(n4895), .B2(n8758), .A(n6409), .ZN(n4894) );
  NOR2_X1 U5264 ( .A1(n8747), .A2(n4896), .ZN(n4895) );
  INV_X1 U5265 ( .A(n6424), .ZN(n4896) );
  OAI22_X1 U5266 ( .A1(n8768), .A2(n4599), .B1(n4601), .B2(n4598), .ZN(n8729)
         );
  AND2_X1 U5267 ( .A1(n5019), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5268 ( .A1(n5017), .A2(n4603), .ZN(n4599) );
  INV_X1 U5269 ( .A(n5017), .ZN(n4598) );
  NAND2_X1 U5270 ( .A1(n4898), .A2(n5018), .ZN(n4897) );
  INV_X1 U5271 ( .A(n8756), .ZN(n4898) );
  INV_X1 U5272 ( .A(n8780), .ZN(n8749) );
  INV_X1 U5273 ( .A(n4885), .ZN(n4884) );
  OAI21_X1 U5274 ( .B1(n8808), .B2(n4886), .A(n6180), .ZN(n4885) );
  NOR2_X1 U5275 ( .A1(n7991), .A2(n5004), .ZN(n5003) );
  INV_X1 U5276 ( .A(n5074), .ZN(n5004) );
  NAND2_X1 U5277 ( .A1(n5002), .A2(n5005), .ZN(n5001) );
  INV_X1 U5278 ( .A(n6400), .ZN(n4888) );
  OR2_X1 U5279 ( .A1(n7989), .A2(n8810), .ZN(n5074) );
  OR2_X1 U5280 ( .A1(n6164), .A2(n6163), .ZN(n6175) );
  AND2_X1 U5281 ( .A1(n4590), .A2(n4537), .ZN(n8817) );
  NAND2_X1 U5282 ( .A1(n8828), .A2(n7987), .ZN(n4590) );
  INV_X1 U5283 ( .A(n5009), .ZN(n4593) );
  INV_X1 U5284 ( .A(n5007), .ZN(n5006) );
  OAI21_X1 U5285 ( .B1(n5011), .B2(n4513), .A(n4479), .ZN(n5007) );
  AND2_X1 U5286 ( .A1(n4639), .A2(n7858), .ZN(n4638) );
  INV_X1 U5287 ( .A(n5011), .ZN(n5010) );
  INV_X1 U5288 ( .A(n7782), .ZN(n5014) );
  NAND2_X1 U5289 ( .A1(n7504), .A2(n4503), .ZN(n7649) );
  OR2_X1 U5290 ( .A1(n7489), .A2(n7490), .ZN(n7504) );
  AND2_X1 U5291 ( .A1(n6347), .A2(n6355), .ZN(n7490) );
  NAND2_X1 U5292 ( .A1(n6748), .A2(n6747), .ZN(n7270) );
  OR2_X1 U5293 ( .A1(n6784), .A2(n6757), .ZN(n8852) );
  OR2_X1 U5294 ( .A1(n6784), .A2(n6509), .ZN(n8850) );
  OAI211_X1 U5295 ( .C1(n7385), .C2(n4994), .A(n6936), .B(n4993), .ZN(n7124)
         );
  INV_X1 U5296 ( .A(n6930), .ZN(n4994) );
  NAND2_X1 U5297 ( .A1(n6929), .A2(n4474), .ZN(n4993) );
  NAND2_X1 U5298 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  OR2_X1 U5299 ( .A1(n7442), .A2(n8063), .ZN(n7280) );
  INV_X1 U5300 ( .A(n8852), .ZN(n8873) );
  AND2_X1 U5301 ( .A1(n6783), .A2(n6737), .ZN(n7033) );
  NAND2_X1 U5302 ( .A1(n8901), .A2(n8985), .ZN(n4608) );
  NAND2_X1 U5303 ( .A1(n8900), .A2(n9980), .ZN(n4793) );
  INV_X1 U5304 ( .A(n10348), .ZN(n9980) );
  NAND2_X1 U5305 ( .A1(n6798), .A2(n10308), .ZN(n10348) );
  OR2_X1 U5306 ( .A1(n6804), .A2(n6314), .ZN(n10350) );
  AND2_X1 U5307 ( .A1(n6733), .A2(n6732), .ZN(n10292) );
  OR2_X1 U5308 ( .A1(n5935), .A2(n6156), .ZN(n5934) );
  OR2_X1 U5309 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  INV_X1 U5310 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4956) );
  AOI21_X1 U5311 ( .B1(n4722), .B2(n4720), .A(n4497), .ZN(n4719) );
  INV_X1 U5312 ( .A(n7671), .ZN(n4720) );
  INV_X1 U5313 ( .A(n4722), .ZN(n4721) );
  NOR2_X1 U5314 ( .A1(n5779), .A2(n5780), .ZN(n5042) );
  NAND2_X1 U5315 ( .A1(n9158), .A2(n5561), .ZN(n5053) );
  INV_X1 U5316 ( .A(n4728), .ZN(n4727) );
  OAI21_X1 U5317 ( .B1(n5051), .B2(n4729), .A(n9094), .ZN(n4728) );
  NOR2_X1 U5318 ( .A1(n9023), .A2(n9026), .ZN(n5049) );
  INV_X1 U5319 ( .A(n4715), .ZN(n4714) );
  OAI21_X1 U5320 ( .B1(n5350), .B2(n4716), .A(n7588), .ZN(n4715) );
  NAND2_X1 U5321 ( .A1(n5349), .A2(n7312), .ZN(n7315) );
  NAND2_X1 U5322 ( .A1(n7315), .A2(n4471), .ZN(n7586) );
  NOR2_X1 U5323 ( .A1(n5063), .A2(n5160), .ZN(n8071) );
  AND2_X1 U5324 ( .A1(n9049), .A2(n6606), .ZN(n5063) );
  NAND2_X1 U5325 ( .A1(n4731), .A2(n4730), .ZN(n9124) );
  AOI21_X1 U5326 ( .B1(n4732), .B2(n4734), .A(n4526), .ZN(n4730) );
  AND2_X1 U5327 ( .A1(n6676), .A2(n10234), .ZN(n5884) );
  AND2_X1 U5328 ( .A1(n8343), .A2(n10200), .ZN(n7043) );
  NOR2_X1 U5329 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5133), .ZN(n5067) );
  INV_X1 U5330 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5131) );
  MUX2_X1 U5331 ( .A(n8172), .B(n8171), .S(n8170), .Z(n8176) );
  AOI21_X1 U5332 ( .B1(n4664), .B2(n8215), .A(n8169), .ZN(n8171) );
  NAND2_X1 U5333 ( .A1(n8295), .A2(n9342), .ZN(n8293) );
  OR2_X1 U5334 ( .A1(n8292), .A2(n9342), .ZN(n8294) );
  NAND2_X1 U5335 ( .A1(n4510), .A2(n4658), .ZN(n4656) );
  AND2_X1 U5336 ( .A1(n5708), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U5337 ( .A1(n8352), .A2(n8304), .ZN(n8177) );
  NOR2_X1 U5338 ( .A1(n6633), .A2(n6632), .ZN(n6631) );
  NAND2_X1 U5339 ( .A1(n6577), .A2(n4617), .ZN(n4616) );
  INV_X1 U5340 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4617) );
  INV_X1 U5341 ( .A(n4616), .ZN(n4615) );
  AND2_X1 U5342 ( .A1(n10104), .A2(n4614), .ZN(n4613) );
  OR2_X1 U5343 ( .A1(n6615), .A2(n4615), .ZN(n4614) );
  AOI21_X1 U5344 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6636), .A(n6631), .ZN(
        n6614) );
  NAND2_X1 U5345 ( .A1(n6614), .A2(n6615), .ZN(n6613) );
  NOR2_X1 U5346 ( .A1(n6651), .A2(n6652), .ZN(n6701) );
  NAND2_X1 U5347 ( .A1(n9190), .A2(n9189), .ZN(n4621) );
  NAND2_X1 U5348 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  INV_X1 U5349 ( .A(n10116), .ZN(n4620) );
  NAND2_X1 U5350 ( .A1(n5092), .A2(n4735), .ZN(n5572) );
  OR2_X1 U5351 ( .A1(n10165), .A2(n4627), .ZN(n4626) );
  AND2_X1 U5352 ( .A1(n10170), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5353 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5354 ( .A(n10180), .ZN(n4625) );
  AND2_X1 U5355 ( .A1(n8286), .A2(n8284), .ZN(n9244) );
  OR2_X1 U5356 ( .A1(n8211), .A2(n8210), .ZN(n9274) );
  INV_X1 U5357 ( .A(n8138), .ZN(n4829) );
  NAND2_X1 U5358 ( .A1(n4911), .A2(n4909), .ZN(n9281) );
  AOI21_X1 U5359 ( .B1(n9321), .B2(n8178), .A(n9318), .ZN(n9299) );
  NAND2_X1 U5360 ( .A1(n9333), .A2(n8023), .ZN(n4863) );
  NOR2_X1 U5361 ( .A1(n8179), .A2(n8221), .ZN(n4833) );
  AOI21_X1 U5362 ( .B1(n9401), .B2(n8021), .A(n4491), .ZN(n9350) );
  NAND2_X1 U5363 ( .A1(n9393), .A2(n9394), .ZN(n4834) );
  NOR2_X1 U5364 ( .A1(n9389), .A2(n9493), .ZN(n9375) );
  OR2_X1 U5365 ( .A1(n8180), .A2(n8179), .ZN(n9373) );
  AND2_X1 U5366 ( .A1(n9408), .A2(n8260), .ZN(n9418) );
  OR2_X1 U5367 ( .A1(n7872), .A2(n9169), .ZN(n9998) );
  NOR2_X1 U5368 ( .A1(n9998), .A2(n10009), .ZN(n10002) );
  NAND2_X1 U5369 ( .A1(n9997), .A2(n9996), .ZN(n9995) );
  AND2_X1 U5370 ( .A1(n8256), .A2(n8254), .ZN(n8203) );
  NAND2_X1 U5371 ( .A1(n7846), .A2(n7845), .ZN(n7877) );
  NAND2_X1 U5372 ( .A1(n4866), .A2(n4864), .ZN(n7846) );
  NOR2_X1 U5373 ( .A1(n4527), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U5374 ( .A1(n7720), .A2(n8196), .ZN(n4866) );
  NAND2_X1 U5375 ( .A1(n5443), .A2(n5442), .ZN(n7710) );
  NOR2_X1 U5376 ( .A1(n7564), .A2(n10262), .ZN(n7536) );
  AOI21_X1 U5377 ( .B1(n8193), .B2(n4467), .A(n4477), .ZN(n4900) );
  NAND2_X1 U5378 ( .A1(n4817), .A2(n8091), .ZN(n7601) );
  NOR2_X1 U5379 ( .A1(n8189), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5380 ( .A1(n7414), .A2(n8314), .ZN(n4848) );
  NAND2_X1 U5381 ( .A1(n6872), .A2(n6879), .ZN(n6994) );
  OR2_X1 U5382 ( .A1(n8177), .A2(n5886), .ZN(n9423) );
  AND2_X1 U5383 ( .A1(n7965), .A2(n10235), .ZN(n7967) );
  OR2_X1 U5384 ( .A1(n5859), .A2(n6844), .ZN(n7051) );
  NAND2_X1 U5385 ( .A1(n6841), .A2(n6840), .ZN(n9985) );
  INV_X1 U5386 ( .A(n9423), .ZN(n9988) );
  INV_X1 U5387 ( .A(n9425), .ZN(n9990) );
  INV_X1 U5388 ( .A(n9253), .ZN(n9455) );
  OR2_X1 U5389 ( .A1(n6831), .A2(n6830), .ZN(n6853) );
  NAND3_X1 U5390 ( .A1(n5112), .A2(n5152), .A3(n5064), .ZN(n5154) );
  XNOR2_X1 U5391 ( .A(n4987), .B(n6305), .ZN(n8160) );
  OAI21_X1 U5392 ( .B1(n6300), .B2(n4988), .A(n6303), .ZN(n4987) );
  XNOR2_X1 U5393 ( .A(n6300), .B(SI_30_), .ZN(n8451) );
  AND2_X1 U5394 ( .A1(n5112), .A2(n5064), .ZN(n5149) );
  INV_X1 U5395 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5396 ( .A1(n5836), .A2(n5835), .ZN(n6249) );
  AND2_X1 U5397 ( .A1(n6250), .A2(n5840), .ZN(n6248) );
  NAND2_X1 U5398 ( .A1(n5112), .A2(n5111), .ZN(n5134) );
  NAND2_X1 U5399 ( .A1(n5114), .A2(n5132), .ZN(n5116) );
  NAND2_X1 U5400 ( .A1(n4764), .A2(n4763), .ZN(n5724) );
  AOI21_X1 U5401 ( .B1(n4766), .B2(n4769), .A(n4535), .ZN(n4763) );
  XNOR2_X1 U5402 ( .A(n5879), .B(n5110), .ZN(n7744) );
  INV_X1 U5403 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5097) );
  INV_X1 U5404 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5405 ( .A1(n4765), .A2(n4770), .ZN(n5701) );
  NAND2_X1 U5406 ( .A1(n4970), .A2(n4772), .ZN(n4765) );
  NAND2_X1 U5407 ( .A1(n4774), .A2(n4968), .ZN(n5665) );
  OAI21_X1 U5408 ( .B1(n5512), .B2(n4489), .A(n4784), .ZN(n5590) );
  NAND2_X1 U5409 ( .A1(n4787), .A2(n5539), .ZN(n5567) );
  NAND2_X1 U5410 ( .A1(n5512), .A2(n4788), .ZN(n4787) );
  NOR2_X1 U5411 ( .A1(n5393), .A2(n5392), .ZN(n6654) );
  XNOR2_X1 U5412 ( .A(n5378), .B(n5379), .ZN(n6579) );
  NAND2_X1 U5413 ( .A1(n6202), .A2(n6201), .ZN(n8930) );
  NAND2_X1 U5414 ( .A1(n6182), .A2(n6181), .ZN(n8939) );
  NAND2_X1 U5415 ( .A1(n4683), .A2(n4500), .ZN(n4576) );
  NAND2_X1 U5416 ( .A1(n4468), .A2(n4684), .ZN(n4683) );
  NOR2_X1 U5417 ( .A1(n4548), .A2(n10308), .ZN(n4684) );
  NOR2_X1 U5418 ( .A1(n4468), .A2(n6489), .ZN(n4635) );
  NAND2_X1 U5419 ( .A1(n4492), .A2(n5995), .ZN(n8565) );
  NAND4_X1 U5420 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8567)
         );
  NAND2_X1 U5421 ( .A1(n5952), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5953) );
  OR2_X1 U5422 ( .A1(n5969), .A2(n6898), .ZN(n5931) );
  XNOR2_X1 U5423 ( .A(n8367), .B(n8369), .ZN(n8903) );
  NAND2_X1 U5424 ( .A1(n6139), .A2(n6138), .ZN(n8961) );
  INV_X1 U5425 ( .A(n8865), .ZN(n8760) );
  INV_X1 U5426 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9012) );
  INV_X1 U5427 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4560) );
  NOR2_X1 U5428 ( .A1(n5935), .A2(n4587), .ZN(n4586) );
  OR2_X1 U5429 ( .A1(n4869), .A2(n4589), .ZN(n4588) );
  NOR2_X1 U5430 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4587) );
  OR2_X1 U5431 ( .A1(n5219), .A2(n6558), .ZN(n4868) );
  OAI22_X1 U5432 ( .A1(n4458), .A2(n4476), .B1(n5216), .B2(n10056), .ZN(n4867)
         );
  NAND2_X1 U5433 ( .A1(n5788), .A2(n5787), .ZN(n9465) );
  XNOR2_X1 U5434 ( .A(n5144), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U5435 ( .A1(n5143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U5436 ( .A1(n5898), .A2(n5897), .ZN(n9257) );
  INV_X1 U5437 ( .A(n9151), .ZN(n9275) );
  NAND2_X1 U5438 ( .A1(n5798), .A2(n5797), .ZN(n9306) );
  OR2_X1 U5439 ( .A1(n9284), .A2(n5734), .ZN(n5798) );
  NAND4_X2 U5440 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n9187)
         );
  NAND2_X1 U5441 ( .A1(n5183), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U5442 ( .A1(n5751), .A2(n5750), .ZN(n9480) );
  OR2_X1 U5443 ( .A1(n9937), .A2(n5882), .ZN(n10221) );
  CLKBUF_X1 U5444 ( .A(n5154), .Z(n9882) );
  INV_X1 U5445 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5390) );
  OAI211_X1 U5446 ( .C1(n8085), .C2(n8170), .A(n8086), .B(n4674), .ZN(n8090)
         );
  NAND2_X1 U5447 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NOR2_X1 U5448 ( .A1(n4843), .A2(n8158), .ZN(n4675) );
  INV_X1 U5449 ( .A(n4681), .ZN(n4575) );
  AOI21_X1 U5450 ( .B1(n6333), .B2(n6334), .A(n4682), .ZN(n4681) );
  AOI21_X1 U5451 ( .B1(n6359), .B2(n4573), .A(n6346), .ZN(n6351) );
  NOR2_X1 U5452 ( .A1(n7483), .A2(n6344), .ZN(n4573) );
  OAI21_X1 U5453 ( .B1(n8108), .B2(n8107), .A(n8106), .ZN(n8114) );
  AOI21_X1 U5454 ( .B1(n4703), .B2(n4702), .A(n4498), .ZN(n6388) );
  NOR2_X1 U5455 ( .A1(n7811), .A2(n6376), .ZN(n4702) );
  OAI21_X1 U5456 ( .B1(n4705), .B2(n6365), .A(n4704), .ZN(n4703) );
  NAND2_X1 U5457 ( .A1(n4564), .A2(n4563), .ZN(n6407) );
  AND2_X1 U5458 ( .A1(n6414), .A2(n6411), .ZN(n4563) );
  OAI21_X1 U5459 ( .B1(n6413), .B2(n6398), .A(n4565), .ZN(n4564) );
  OAI21_X1 U5460 ( .B1(n4672), .B2(n4669), .A(n8145), .ZN(n8153) );
  OAI21_X1 U5461 ( .B1(n4670), .B2(n4472), .A(n4501), .ZN(n4669) );
  AOI211_X1 U5462 ( .C1(n4673), .C2(n8274), .A(n8170), .B(n9319), .ZN(n4672)
         );
  OAI21_X1 U5463 ( .B1(n6441), .B2(n4693), .A(n4688), .ZN(n4570) );
  NAND2_X1 U5464 ( .A1(n6473), .A2(n6934), .ZN(n4699) );
  NAND2_X1 U5465 ( .A1(n6946), .A2(n7276), .ZN(n6335) );
  INV_X1 U5466 ( .A(n5718), .ZN(n5033) );
  OR2_X1 U5467 ( .A1(n9444), .A2(n8033), .ZN(n8287) );
  INV_X1 U5468 ( .A(SI_19_), .ZN(n5645) );
  INV_X1 U5469 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5593) );
  INV_X1 U5470 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5594) );
  INV_X1 U5471 ( .A(SI_12_), .ZN(n5460) );
  OAI21_X1 U5472 ( .B1(n7758), .B2(n4925), .A(n4470), .ZN(n4924) );
  NAND2_X1 U5473 ( .A1(n4926), .A2(n7638), .ZN(n4925) );
  INV_X1 U5474 ( .A(n7638), .ZN(n4928) );
  INV_X1 U5475 ( .A(n4950), .ZN(n4947) );
  OR2_X1 U5476 ( .A1(n8683), .A2(n8685), .ZN(n6315) );
  NAND2_X1 U5477 ( .A1(n4567), .A2(n6457), .ZN(n6460) );
  NAND2_X1 U5478 ( .A1(n4568), .A2(n4856), .ZN(n4567) );
  NAND2_X1 U5479 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NOR2_X1 U5480 ( .A1(n4857), .A2(n6453), .ZN(n4569) );
  NAND2_X1 U5481 ( .A1(n4687), .A2(n4695), .ZN(n4686) );
  NAND2_X1 U5482 ( .A1(n6285), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5940) );
  NOR3_X1 U5483 ( .A1(n10290), .A2(n5939), .A3(n9909), .ZN(n9907) );
  NOR2_X1 U5484 ( .A1(n4741), .A2(n8900), .ZN(n4740) );
  OR2_X1 U5485 ( .A1(n8904), .A2(n8705), .ZN(n6261) );
  NAND2_X1 U5486 ( .A1(n8364), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U5487 ( .A1(n8777), .A2(n4603), .ZN(n4602) );
  NOR2_X1 U5488 ( .A1(n8930), .A2(n6200), .ZN(n4751) );
  NOR2_X1 U5489 ( .A1(n6419), .A2(n4882), .ZN(n4881) );
  INV_X1 U5490 ( .A(n4887), .ZN(n4882) );
  NOR2_X1 U5491 ( .A1(n8775), .A2(n8795), .ZN(n6418) );
  NOR2_X1 U5492 ( .A1(n8961), .A2(n8964), .ZN(n4746) );
  NOR2_X1 U5493 ( .A1(n8954), .A2(n4745), .ZN(n4744) );
  INV_X1 U5494 ( .A(n4746), .ZN(n4745) );
  OR2_X1 U5495 ( .A1(n8961), .A2(n8532), .ZN(n6393) );
  AND2_X1 U5496 ( .A1(n7860), .A2(n7650), .ZN(n4591) );
  INV_X1 U5497 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5498 ( .A1(n7125), .A2(n7132), .ZN(n6340) );
  INV_X1 U5499 ( .A(n8565), .ZN(n7125) );
  AND2_X1 U5500 ( .A1(n6340), .A2(n6338), .ZN(n6472) );
  NAND2_X1 U5501 ( .A1(n7276), .A2(n4457), .ZN(n4757) );
  AND2_X1 U5502 ( .A1(n8787), .A2(n4487), .ZN(n8733) );
  NAND2_X1 U5503 ( .A1(n8888), .A2(n8887), .ZN(n8890) );
  INV_X1 U5504 ( .A(n6781), .ZN(n7259) );
  INV_X1 U5505 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U5506 ( .A1(n6494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U5507 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  INV_X1 U5508 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6495) );
  INV_X1 U5509 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6492) );
  INV_X1 U5510 ( .A(n5588), .ZN(n4729) );
  NOR2_X1 U5511 ( .A1(n4729), .A2(n4726), .ZN(n4725) );
  INV_X1 U5512 ( .A(n5561), .ZN(n4726) );
  INV_X1 U5513 ( .A(n4733), .ZN(n4732) );
  OAI21_X1 U5514 ( .B1(n5699), .B2(n4734), .A(n5032), .ZN(n4733) );
  NOR2_X1 U5515 ( .A1(n5035), .A2(n5033), .ZN(n5032) );
  NOR2_X1 U5516 ( .A1(n9125), .A2(n5034), .ZN(n5035) );
  AND2_X1 U5517 ( .A1(n5067), .A2(n5139), .ZN(n5066) );
  NAND2_X1 U5518 ( .A1(n4665), .A2(n4663), .ZN(n8167) );
  AOI21_X1 U5519 ( .B1(n4666), .B2(n4668), .A(n4664), .ZN(n4663) );
  AND2_X1 U5520 ( .A1(n4667), .A2(n4518), .ZN(n4666) );
  INV_X1 U5521 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5324) );
  AND2_X1 U5522 ( .A1(n4619), .A2(n4618), .ZN(n9192) );
  NAND2_X1 U5523 ( .A1(n10120), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4618) );
  OAI21_X1 U5524 ( .B1(n4825), .B2(n4822), .A(n4821), .ZN(n4820) );
  INV_X1 U5525 ( .A(n8281), .ZN(n4821) );
  INV_X1 U5526 ( .A(n8329), .ZN(n4822) );
  NOR2_X1 U5527 ( .A1(n9455), .A2(n9460), .ZN(n4799) );
  NOR2_X1 U5528 ( .A1(n9480), .A2(n4809), .ZN(n4808) );
  INV_X1 U5529 ( .A(n4810), .ZN(n4809) );
  OR2_X1 U5530 ( .A1(n9471), .A2(n9325), .ZN(n8138) );
  INV_X1 U5531 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5094) );
  NOR2_X1 U5532 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4735) );
  NOR2_X1 U5533 ( .A1(n9503), .A2(n4814), .ZN(n4812) );
  INV_X1 U5534 ( .A(n9998), .ZN(n4813) );
  INV_X1 U5535 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5520) );
  INV_X1 U5536 ( .A(n7721), .ZN(n4865) );
  INV_X1 U5537 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6663) );
  INV_X1 U5538 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5396) );
  OR2_X1 U5539 ( .A1(n5397), .A2(n5396), .ZN(n5424) );
  AND2_X1 U5540 ( .A1(n8314), .A2(n8319), .ZN(n8187) );
  INV_X1 U5541 ( .A(n6875), .ZN(n4654) );
  NAND2_X1 U5542 ( .A1(n9375), .A2(n4810), .ZN(n9339) );
  INV_X1 U5543 ( .A(SI_28_), .ZN(n9735) );
  INV_X1 U5544 ( .A(SI_30_), .ZN(n4988) );
  NAND2_X1 U5545 ( .A1(n4960), .A2(n4959), .ZN(n5807) );
  AOI21_X1 U5546 ( .B1(n4484), .B2(n4964), .A(n4534), .ZN(n4959) );
  AOI21_X1 U5547 ( .B1(n4966), .B2(n4963), .A(n4962), .ZN(n4961) );
  INV_X1 U5548 ( .A(n5764), .ZN(n4962) );
  INV_X1 U5549 ( .A(n5743), .ZN(n4963) );
  INV_X1 U5550 ( .A(n4966), .ZN(n4964) );
  AOI21_X1 U5551 ( .B1(n5642), .B2(n4969), .A(n4511), .ZN(n4968) );
  INV_X1 U5552 ( .A(n5619), .ZN(n4969) );
  INV_X1 U5553 ( .A(SI_16_), .ZN(n5568) );
  INV_X1 U5554 ( .A(n5539), .ZN(n4786) );
  INV_X1 U5555 ( .A(n4785), .ZN(n4784) );
  OAI21_X1 U5556 ( .B1(n4788), .B2(n4489), .A(n5565), .ZN(n4785) );
  INV_X1 U5557 ( .A(SI_13_), .ZN(n5488) );
  AOI21_X1 U5558 ( .B1(n4976), .B2(n4978), .A(n4512), .ZN(n4975) );
  NAND2_X1 U5559 ( .A1(n4973), .A2(n4780), .ZN(n4776) );
  AND2_X1 U5560 ( .A1(n4679), .A2(n4678), .ZN(n5303) );
  NAND2_X1 U5561 ( .A1(n5128), .A2(n6570), .ZN(n4679) );
  NAND2_X1 U5562 ( .A1(n6556), .A2(n6566), .ZN(n4678) );
  INV_X1 U5563 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5124) );
  NAND2_X1 U5564 ( .A1(n5123), .A2(n8682), .ZN(n4990) );
  INV_X1 U5565 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5122) );
  INV_X1 U5566 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5121) );
  NAND2_X1 U5567 ( .A1(n8528), .A2(n8527), .ZN(n4943) );
  NAND2_X1 U5568 ( .A1(n7622), .A2(n7621), .ZN(n7639) );
  NAND2_X1 U5569 ( .A1(n6190), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6203) );
  OR2_X1 U5570 ( .A1(n6067), .A2(n6066), .ZN(n6079) );
  NOR2_X1 U5571 ( .A1(n7017), .A2(n6960), .ZN(n4932) );
  NAND2_X1 U5572 ( .A1(n6956), .A2(n7007), .ZN(n4931) );
  NAND2_X1 U5573 ( .A1(n8482), .A2(n8424), .ZN(n4952) );
  NAND2_X1 U5574 ( .A1(n4647), .A2(n4644), .ZN(n6308) );
  INV_X1 U5575 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U5576 ( .A1(n5948), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U5577 ( .A1(n6285), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5950) );
  NOR2_X1 U5578 ( .A1(n8585), .A2(n8584), .ZN(n8583) );
  NOR2_X1 U5579 ( .A1(n8598), .A2(n8597), .ZN(n8596) );
  NOR2_X1 U5580 ( .A1(n7208), .A2(n7209), .ZN(n7207) );
  NAND2_X1 U5581 ( .A1(n7296), .A2(n7297), .ZN(n7573) );
  NAND2_X1 U5582 ( .A1(n7573), .A2(n4553), .ZN(n8616) );
  NAND2_X1 U5583 ( .A1(n7577), .A2(n6106), .ZN(n4553) );
  NOR2_X1 U5584 ( .A1(n8620), .A2(n8621), .ZN(n8643) );
  NAND2_X1 U5585 ( .A1(n8673), .A2(n8674), .ZN(n4552) );
  NAND2_X1 U5586 ( .A1(n6261), .A2(n6446), .ZN(n8365) );
  OR2_X1 U5587 ( .A1(n8719), .A2(n4741), .ZN(n8375) );
  NOR2_X1 U5588 ( .A1(n8702), .A2(n8703), .ZN(n4629) );
  NAND2_X1 U5589 ( .A1(n6247), .A2(n6442), .ZN(n8702) );
  INV_X1 U5590 ( .A(n4630), .ZN(n8716) );
  OAI22_X1 U5591 ( .A1(n8729), .A2(n4899), .B1(n8554), .B2(n8921), .ZN(n8712)
         );
  NAND2_X1 U5592 ( .A1(n8787), .A2(n4749), .ZN(n8742) );
  NAND2_X1 U5593 ( .A1(n4880), .A2(n4877), .ZN(n8778) );
  NAND2_X1 U5594 ( .A1(n4879), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U5595 ( .A1(n8819), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U5596 ( .A1(n4884), .A2(n8792), .ZN(n4879) );
  NAND2_X1 U5597 ( .A1(n8787), .A2(n8775), .ZN(n8769) );
  AOI21_X1 U5598 ( .B1(n4998), .B2(n5000), .A(n4507), .ZN(n4996) );
  NAND2_X1 U5599 ( .A1(n7990), .A2(n4998), .ZN(n4995) );
  NOR2_X1 U5600 ( .A1(n8801), .A2(n8939), .ZN(n8787) );
  NAND2_X1 U5601 ( .A1(n4891), .A2(n4890), .ZN(n4889) );
  INV_X1 U5602 ( .A(n8818), .ZN(n4890) );
  INV_X1 U5603 ( .A(n8819), .ZN(n4891) );
  NAND2_X1 U5604 ( .A1(n4889), .A2(n6400), .ZN(n8809) );
  AND2_X1 U5605 ( .A1(n8888), .A2(n4743), .ZN(n8822) );
  AND2_X1 U5606 ( .A1(n4744), .A2(n7989), .ZN(n4743) );
  INV_X1 U5607 ( .A(n6141), .ZN(n6140) );
  NAND2_X1 U5608 ( .A1(n8888), .A2(n4744), .ZN(n8829) );
  NAND2_X1 U5609 ( .A1(n5023), .A2(n5022), .ZN(n8828) );
  AOI21_X1 U5610 ( .B1(n4469), .B2(n8870), .A(n4509), .ZN(n5022) );
  OR2_X1 U5611 ( .A1(n8866), .A2(n8870), .ZN(n5024) );
  AND2_X1 U5612 ( .A1(n6389), .A2(n8844), .ZN(n8870) );
  AND2_X1 U5613 ( .A1(n7851), .A2(n7853), .ZN(n8888) );
  NAND2_X1 U5614 ( .A1(n7816), .A2(n6377), .ZN(n7849) );
  NOR2_X1 U5615 ( .A1(n7812), .A2(n8977), .ZN(n7851) );
  NAND2_X1 U5616 ( .A1(n6077), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6092) );
  INV_X1 U5617 ( .A(n6079), .ZN(n6077) );
  INV_X1 U5618 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6091) );
  OR2_X1 U5619 ( .A1(n6092), .A2(n6091), .ZN(n6104) );
  OR2_X1 U5620 ( .A1(n7792), .A2(n8984), .ZN(n7812) );
  NAND2_X1 U5621 ( .A1(n7507), .A2(n6086), .ZN(n4643) );
  AND2_X1 U5622 ( .A1(n7339), .A2(n4481), .ZN(n7698) );
  NAND2_X1 U5623 ( .A1(n7649), .A2(n7648), .ZN(n7693) );
  NAND2_X1 U5624 ( .A1(n7339), .A2(n4759), .ZN(n7699) );
  INV_X1 U5625 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6040) );
  OR2_X1 U5626 ( .A1(n6041), .A2(n6040), .ZN(n6053) );
  NAND2_X1 U5627 ( .A1(n7339), .A2(n10337), .ZN(n7494) );
  AND2_X1 U5628 ( .A1(n6343), .A2(n6358), .ZN(n7129) );
  INV_X1 U5629 ( .A(n7129), .ZN(n7480) );
  AND2_X1 U5630 ( .A1(n7133), .A2(n7545), .ZN(n7339) );
  INV_X1 U5631 ( .A(n4572), .ZN(n4571) );
  NAND2_X1 U5632 ( .A1(n4756), .A2(n4753), .ZN(n7370) );
  AND3_X1 U5633 ( .A1(n7122), .A2(n10323), .A3(n4754), .ZN(n4753) );
  INV_X1 U5634 ( .A(n4757), .ZN(n4754) );
  NAND2_X1 U5635 ( .A1(n4756), .A2(n4755), .ZN(n7380) );
  NOR2_X1 U5636 ( .A1(n4757), .A2(n6953), .ZN(n4755) );
  NAND2_X1 U5637 ( .A1(n6929), .A2(n6928), .ZN(n7386) );
  NAND2_X1 U5638 ( .A1(n7283), .A2(n6744), .ZN(n6746) );
  NAND2_X1 U5639 ( .A1(n6746), .A2(n6745), .ZN(n6929) );
  NOR2_X1 U5640 ( .A1(n7442), .A2(n4757), .ZN(n7381) );
  NOR2_X1 U5641 ( .A1(n10350), .A2(n4919), .ZN(n6807) );
  NAND2_X1 U5642 ( .A1(n7285), .A2(n7284), .ZN(n7283) );
  CLKBUF_X1 U5643 ( .A(n6467), .Z(n7284) );
  NAND2_X1 U5644 ( .A1(n7260), .A2(n7259), .ZN(n7263) );
  NAND2_X1 U5645 ( .A1(n6470), .A2(n6469), .ZN(n7438) );
  NAND2_X1 U5646 ( .A1(n6225), .A2(n6224), .ZN(n8916) );
  INV_X1 U5647 ( .A(n10350), .ZN(n8985) );
  NAND2_X1 U5648 ( .A1(n6812), .A2(n10306), .ZN(n10293) );
  NAND2_X1 U5649 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4589) );
  NAND2_X1 U5650 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  NAND2_X1 U5651 ( .A1(n5921), .A2(n4954), .ZN(n6313) );
  AND2_X1 U5652 ( .A1(n4957), .A2(n6293), .ZN(n4954) );
  NAND2_X1 U5653 ( .A1(n5921), .A2(n5070), .ZN(n6136) );
  AND2_X1 U5654 ( .A1(n4582), .A2(n4583), .ZN(n5987) );
  INV_X1 U5655 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4936) );
  OR2_X1 U5656 ( .A1(n5752), .A2(n9028), .ZN(n5768) );
  NAND2_X1 U5657 ( .A1(n5628), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5652) );
  INV_X1 U5658 ( .A(n5629), .ZN(n5628) );
  AOI21_X1 U5659 ( .B1(n5045), .B2(n5042), .A(n5044), .ZN(n5041) );
  NAND2_X1 U5660 ( .A1(n9024), .A2(n5039), .ZN(n5037) );
  OAI21_X1 U5661 ( .B1(n5050), .B2(n9148), .A(n9146), .ZN(n5044) );
  NAND2_X1 U5662 ( .A1(n4712), .A2(n4505), .ZN(n7683) );
  OR2_X1 U5663 ( .A1(n9035), .A2(n9036), .ZN(n9109) );
  NAND2_X1 U5664 ( .A1(n5719), .A2(n5718), .ZN(n5036) );
  NAND2_X1 U5665 ( .A1(n9067), .A2(n9068), .ZN(n5719) );
  AND2_X1 U5666 ( .A1(n4546), .A2(n7773), .ZN(n4722) );
  NAND2_X1 U5667 ( .A1(n7670), .A2(n7671), .ZN(n4723) );
  OR2_X1 U5668 ( .A1(n5424), .A2(n6663), .ZN(n5471) );
  OR2_X1 U5669 ( .A1(n6838), .A2(n5175), .ZN(n5177) );
  OR2_X1 U5670 ( .A1(n8309), .A2(n5175), .ZN(n5078) );
  NAND2_X1 U5671 ( .A1(n5289), .A2(n5288), .ZN(n7214) );
  OR2_X1 U5672 ( .A1(n8177), .A2(n7043), .ZN(n7042) );
  OR2_X1 U5673 ( .A1(n5521), .A2(n5520), .ZN(n5551) );
  NAND2_X1 U5674 ( .A1(n8352), .A2(n10200), .ZN(n6833) );
  CLKBUF_X1 U5675 ( .A(n5216), .Z(n6640) );
  NOR2_X1 U5676 ( .A1(n10054), .A2(n10076), .ZN(n10053) );
  AOI21_X1 U5677 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n9895), .A(n9896), .ZN(
        n10088) );
  OR2_X1 U5678 ( .A1(n6681), .A2(n6682), .ZN(n4612) );
  INV_X1 U5679 ( .A(n5886), .ZN(n6842) );
  NAND2_X1 U5680 ( .A1(n4612), .A2(n4611), .ZN(n6633) );
  NAND2_X1 U5681 ( .A1(n6565), .A2(n10209), .ZN(n4611) );
  INV_X1 U5682 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5326) );
  OAI22_X1 U5683 ( .A1(n6614), .A2(n4532), .B1(n4613), .B2(n4485), .ZN(n6526)
         );
  NAND2_X1 U5684 ( .A1(n5089), .A2(n5247), .ZN(n5391) );
  NOR2_X1 U5685 ( .A1(n6701), .A2(n4542), .ZN(n6703) );
  NAND2_X1 U5686 ( .A1(n6703), .A2(n6704), .ZN(n6773) );
  AND2_X1 U5687 ( .A1(n9208), .A2(n9207), .ZN(n10134) );
  XNOR2_X1 U5688 ( .A(n9192), .B(n9210), .ZN(n10129) );
  NOR2_X1 U5689 ( .A1(n9195), .A2(n10141), .ZN(n10154) );
  XNOR2_X1 U5690 ( .A(n4622), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U5691 ( .A1(n4624), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5692 ( .A1(n10185), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4623) );
  AND2_X1 U5693 ( .A1(n9283), .A2(n4536), .ZN(n8036) );
  AND2_X1 U5694 ( .A1(n5891), .A2(n8037), .ZN(n9239) );
  NAND2_X1 U5695 ( .A1(n9283), .A2(n4797), .ZN(n9236) );
  NAND2_X1 U5696 ( .A1(n4903), .A2(n4904), .ZN(n9249) );
  INV_X1 U5697 ( .A(n4905), .ZN(n4904) );
  OAI21_X1 U5698 ( .B1(n4909), .B2(n4906), .A(n8209), .ZN(n4905) );
  AND2_X1 U5699 ( .A1(n8283), .A2(n9242), .ZN(n9255) );
  AOI21_X1 U5700 ( .B1(n4831), .B2(n4828), .A(n4826), .ZN(n4825) );
  NAND2_X1 U5701 ( .A1(n9283), .A2(n9270), .ZN(n9264) );
  NAND2_X1 U5702 ( .A1(n9375), .A2(n4806), .ZN(n9309) );
  NOR2_X1 U5703 ( .A1(n9471), .A2(n4807), .ZN(n4806) );
  INV_X1 U5704 ( .A(n4808), .ZN(n4807) );
  NOR2_X1 U5705 ( .A1(n9465), .A2(n9309), .ZN(n9283) );
  NOR2_X1 U5706 ( .A1(n4862), .A2(n4494), .ZN(n4861) );
  AND2_X1 U5707 ( .A1(n8138), .A2(n8141), .ZN(n9302) );
  NAND2_X1 U5708 ( .A1(n5730), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5752) );
  INV_X1 U5709 ( .A(n5732), .ZN(n5730) );
  AND2_X1 U5710 ( .A1(n8268), .A2(n8133), .ZN(n9363) );
  NAND2_X1 U5711 ( .A1(n9375), .A2(n9359), .ZN(n9353) );
  OR2_X1 U5712 ( .A1(n8020), .A2(n8019), .ZN(n9348) );
  NAND2_X1 U5713 ( .A1(n4813), .A2(n4811), .ZN(n9389) );
  AND2_X1 U5714 ( .A1(n4812), .A2(n4815), .ZN(n4811) );
  NOR2_X1 U5715 ( .A1(n9998), .A2(n4814), .ZN(n9426) );
  NAND2_X1 U5716 ( .A1(n4813), .A2(n4812), .ZN(n9402) );
  NAND2_X1 U5717 ( .A1(n4872), .A2(n4871), .ZN(n9401) );
  AOI21_X1 U5718 ( .B1(n4873), .B2(n4875), .A(n4528), .ZN(n4871) );
  NAND2_X1 U5719 ( .A1(n5549), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5602) );
  INV_X1 U5720 ( .A(n5551), .ZN(n5549) );
  AND2_X1 U5721 ( .A1(n4801), .A2(n7536), .ZN(n7841) );
  NOR2_X1 U5722 ( .A1(n4802), .A2(n7907), .ZN(n4801) );
  INV_X1 U5723 ( .A(n4802), .ZN(n4800) );
  NAND2_X1 U5724 ( .A1(n7536), .A2(n4804), .ZN(n7714) );
  NAND2_X1 U5725 ( .A1(n4816), .A2(n8241), .ZN(n7709) );
  NAND2_X1 U5726 ( .A1(n7600), .A2(n7599), .ZN(n7707) );
  NAND2_X1 U5727 ( .A1(n7536), .A2(n9939), .ZN(n7603) );
  AOI21_X1 U5728 ( .B1(n4846), .B2(n4844), .A(n4843), .ZN(n4842) );
  INV_X1 U5729 ( .A(n4846), .ZN(n4845) );
  AND3_X1 U5730 ( .A1(n4805), .A2(n10197), .A3(n4486), .ZN(n7428) );
  NAND2_X1 U5731 ( .A1(n7428), .A2(n7518), .ZN(n7563) );
  NAND2_X1 U5732 ( .A1(n7410), .A2(n7409), .ZN(n7427) );
  NAND2_X1 U5733 ( .A1(n7186), .A2(n4915), .ZN(n7410) );
  NOR2_X1 U5734 ( .A1(n8187), .A2(n4916), .ZN(n4915) );
  INV_X1 U5735 ( .A(n7185), .ZN(n4916) );
  NAND2_X1 U5736 ( .A1(n7447), .A2(n6999), .ZN(n4835) );
  AND2_X1 U5737 ( .A1(n8234), .A2(n8232), .ZN(n8186) );
  NAND2_X1 U5738 ( .A1(n4859), .A2(n4858), .ZN(n6997) );
  NAND2_X1 U5739 ( .A1(n6999), .A2(n6995), .ZN(n4858) );
  NAND2_X1 U5740 ( .A1(n6994), .A2(n4860), .ZN(n4859) );
  AND2_X1 U5741 ( .A1(n6995), .A2(n6993), .ZN(n4860) );
  NAND2_X1 U5742 ( .A1(n6997), .A2(n6996), .ZN(n7186) );
  NAND2_X1 U5743 ( .A1(n4805), .A2(n10241), .ZN(n7458) );
  NAND2_X1 U5744 ( .A1(n4652), .A2(n6875), .ZN(n7957) );
  NAND2_X1 U5745 ( .A1(n6874), .A2(n6873), .ZN(n4652) );
  NOR2_X1 U5746 ( .A1(n8305), .A2(n10211), .ZN(n7965) );
  INV_X1 U5747 ( .A(n4653), .ZN(n6873) );
  NAND2_X1 U5748 ( .A1(n5671), .A2(n5670), .ZN(n9493) );
  INV_X1 U5749 ( .A(n10265), .ZN(n9999) );
  NAND2_X1 U5750 ( .A1(n4841), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U5751 ( .A1(n4839), .A2(n4838), .ZN(n4837) );
  OR2_X1 U5752 ( .A1(n7044), .A2(n6844), .ZN(n10265) );
  INV_X1 U5753 ( .A(n10222), .ZN(n5877) );
  XNOR2_X1 U5754 ( .A(n6274), .B(n6266), .ZN(n9017) );
  NAND2_X1 U5755 ( .A1(n4986), .A2(n6265), .ZN(n6274) );
  XNOR2_X1 U5756 ( .A(n6263), .B(n6262), .ZN(n8449) );
  NAND2_X1 U5757 ( .A1(n4985), .A2(n5702), .ZN(n5720) );
  NAND2_X1 U5758 ( .A1(n4762), .A2(n4766), .ZN(n4985) );
  OR2_X1 U5759 ( .A1(n4970), .A2(n4769), .ZN(n4762) );
  NAND2_X1 U5760 ( .A1(n4970), .A2(n5619), .ZN(n5643) );
  NOR2_X1 U5761 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5090) );
  INV_X1 U5762 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U5763 ( .A1(n5092), .A2(n5514), .ZN(n5516) );
  AND3_X1 U5764 ( .A1(n5089), .A2(n5247), .A3(n4737), .ZN(n5109) );
  NAND2_X1 U5765 ( .A1(n4980), .A2(n5439), .ZN(n5459) );
  NAND2_X1 U5766 ( .A1(n5438), .A2(n5080), .ZN(n4980) );
  XNOR2_X1 U5767 ( .A(n5303), .B(n4677), .ZN(n5301) );
  INV_X1 U5768 ( .A(SI_5_), .ZN(n4677) );
  INV_X1 U5769 ( .A(n8558), .ZN(n7767) );
  OR2_X1 U5770 ( .A1(n8546), .A2(n8852), .ZN(n8530) );
  XNOR2_X1 U5771 ( .A(n8414), .B(n5085), .ZN(n8502) );
  NAND2_X1 U5772 ( .A1(n4943), .A2(n8391), .ZN(n8469) );
  NOR2_X1 U5773 ( .A1(n5975), .A2(n6558), .ZN(n4604) );
  NAND2_X1 U5774 ( .A1(n4944), .A2(n4949), .ZN(n7918) );
  NAND2_X1 U5775 ( .A1(n7916), .A2(n4950), .ZN(n4944) );
  NAND2_X1 U5776 ( .A1(n7823), .A2(n6171), .ZN(n6211) );
  NAND2_X1 U5777 ( .A1(n4935), .A2(n4934), .ZN(n7015) );
  OR2_X1 U5778 ( .A1(n7248), .A2(n7249), .ZN(n7250) );
  NAND2_X1 U5779 ( .A1(n7247), .A2(n7246), .ZN(n7254) );
  AOI21_X1 U5780 ( .B1(n4940), .B2(n4939), .A(n4938), .ZN(n4937) );
  INV_X1 U5781 ( .A(n8397), .ZN(n4938) );
  INV_X1 U5782 ( .A(n8527), .ZN(n4939) );
  NAND2_X1 U5783 ( .A1(n6173), .A2(n6172), .ZN(n8944) );
  NAND2_X1 U5784 ( .A1(n7639), .A2(n7638), .ZN(n7757) );
  OAI22_X1 U5785 ( .A1(n5975), .A2(n6559), .B1(n6902), .B2(n6912), .ZN(n4914)
         );
  NOR2_X1 U5786 ( .A1(n4462), .A2(n6560), .ZN(n4913) );
  XNOR2_X1 U5787 ( .A(n4918), .B(n6945), .ZN(n8059) );
  NAND2_X1 U5788 ( .A1(n4559), .A2(n4930), .ZN(n6981) );
  NAND2_X1 U5789 ( .A1(n4933), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U5790 ( .A1(n4935), .A2(n4932), .ZN(n4559) );
  INV_X1 U5791 ( .A(n6960), .ZN(n4933) );
  AND2_X1 U5792 ( .A1(n4953), .A2(n4952), .ZN(n8542) );
  INV_X1 U5793 ( .A(n8537), .ZN(n8539) );
  NAND2_X1 U5794 ( .A1(n6803), .A2(n6785), .ZN(n8537) );
  NAND2_X1 U5795 ( .A1(n6967), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8522) );
  NAND2_X1 U5796 ( .A1(n6116), .A2(n6115), .ZN(n8972) );
  OR2_X1 U5797 ( .A1(n8698), .A2(n4463), .ZN(n6246) );
  CLKBUF_X1 U5798 ( .A(n6317), .Z(n8569) );
  NOR2_X1 U5799 ( .A1(n7088), .A2(n7087), .ZN(n7086) );
  NOR2_X1 U5800 ( .A1(n7073), .A2(n7072), .ZN(n7099) );
  NOR2_X1 U5801 ( .A1(n7104), .A2(n7103), .ZN(n7150) );
  OR2_X1 U5802 ( .A1(n9913), .A2(n8682), .ZN(n4556) );
  INV_X1 U5803 ( .A(n8916), .ZN(n8725) );
  NAND2_X1 U5804 ( .A1(n8756), .A2(n4895), .ZN(n4892) );
  NAND2_X1 U5805 ( .A1(n4897), .A2(n6424), .ZN(n8748) );
  AND2_X1 U5806 ( .A1(n8759), .A2(n5019), .ZN(n8739) );
  AND2_X1 U5807 ( .A1(n4883), .A2(n4884), .ZN(n8793) );
  NAND2_X1 U5808 ( .A1(n8819), .A2(n4887), .ZN(n4883) );
  NAND2_X1 U5809 ( .A1(n4997), .A2(n5001), .ZN(n8786) );
  NAND2_X1 U5810 ( .A1(n7990), .A2(n5003), .ZN(n4997) );
  NAND2_X1 U5811 ( .A1(n7990), .A2(n5074), .ZN(n8800) );
  NAND2_X1 U5812 ( .A1(n6161), .A2(n6160), .ZN(n8951) );
  NAND2_X1 U5813 ( .A1(n7861), .A2(n7860), .ZN(n7986) );
  NAND2_X1 U5814 ( .A1(n4597), .A2(n5006), .ZN(n7861) );
  NAND2_X1 U5815 ( .A1(n4593), .A2(n5016), .ZN(n4597) );
  AND2_X1 U5816 ( .A1(n4640), .A2(n4639), .ZN(n7817) );
  NAND2_X1 U5817 ( .A1(n5008), .A2(n5010), .ZN(n7859) );
  NAND2_X1 U5818 ( .A1(n7783), .A2(n5013), .ZN(n5008) );
  NAND2_X1 U5819 ( .A1(n5015), .A2(n7782), .ZN(n7784) );
  NAND2_X1 U5820 ( .A1(n5016), .A2(n7652), .ZN(n5015) );
  NAND2_X1 U5821 ( .A1(n7504), .A2(n7503), .ZN(n7506) );
  NAND2_X1 U5822 ( .A1(n6579), .A2(n6171), .ZN(n4636) );
  INV_X1 U5823 ( .A(n8861), .ZN(n8886) );
  INV_X1 U5824 ( .A(n7132), .ZN(n10329) );
  NAND2_X1 U5825 ( .A1(n7384), .A2(n6930), .ZN(n6931) );
  AND2_X1 U5826 ( .A1(n8894), .A2(n7272), .ZN(n8865) );
  AND2_X2 U5827 ( .A1(n7033), .A2(n6740), .ZN(n10370) );
  AOI211_X1 U5828 ( .C1(n9980), .C2(n6297), .A(n9979), .B(n9978), .ZN(n9982)
         );
  NAND2_X1 U5829 ( .A1(n4610), .A2(n4606), .ZN(n8991) );
  OR2_X1 U5830 ( .A1(n8903), .A2(n8981), .ZN(n4610) );
  NAND2_X1 U5831 ( .A1(n4608), .A2(n4793), .ZN(n4607) );
  AND2_X2 U5832 ( .A1(n7260), .A2(n7035), .ZN(n10358) );
  AND2_X1 U5833 ( .A1(n6811), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10306) );
  INV_X1 U5834 ( .A(n10299), .ZN(n10303) );
  NAND2_X1 U5835 ( .A1(n4562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4561) );
  CLKBUF_X1 U5836 ( .A(n6508), .Z(n6509) );
  INV_X1 U5837 ( .A(n4869), .ZN(n6505) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7931) );
  INV_X1 U5839 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7824) );
  XNOR2_X1 U5840 ( .A(n6500), .B(n6499), .ZN(n7825) );
  INV_X1 U5841 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U5842 ( .A1(n6498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6500) );
  INV_X1 U5843 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7751) );
  INV_X1 U5844 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8068) );
  XNOR2_X1 U5845 ( .A(n6296), .B(n6295), .ZN(n7666) );
  INV_X1 U5846 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U5847 ( .A1(n6313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  INV_X1 U5848 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5849 ( .A1(n6311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6312) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8361) );
  AND2_X1 U5851 ( .A1(n5070), .A2(n4956), .ZN(n4955) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9781) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6925) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6722) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6718) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6609) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9602) );
  INV_X1 U5858 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6589) );
  INV_X1 U5859 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6580) );
  OR2_X1 U5860 ( .A1(n6514), .A2(n6515), .ZN(n6546) );
  AOI21_X1 U5861 ( .B1(n5056), .B2(n7888), .A(n4530), .ZN(n5054) );
  NAND2_X1 U5862 ( .A1(n7315), .A2(n5350), .ZN(n4713) );
  INV_X1 U5863 ( .A(n5042), .ZN(n5040) );
  NAND2_X1 U5864 ( .A1(n9024), .A2(n5048), .ZN(n5038) );
  NAND2_X1 U5865 ( .A1(n9083), .A2(n5588), .ZN(n9093) );
  NAND2_X1 U5866 ( .A1(n5047), .A2(n9024), .ZN(n9100) );
  OAI21_X1 U5867 ( .B1(n7315), .B2(n4716), .A(n4714), .ZN(n5377) );
  INV_X1 U5868 ( .A(n9138), .ZN(n9164) );
  NAND2_X1 U5869 ( .A1(n7886), .A2(n5483), .ZN(n7898) );
  NAND2_X1 U5870 ( .A1(n5036), .A2(n5742), .ZN(n9127) );
  INV_X1 U5871 ( .A(n9180), .ZN(n7776) );
  NAND2_X1 U5872 ( .A1(n4723), .A2(n4722), .ZN(n7772) );
  INV_X1 U5873 ( .A(n6713), .ZN(n5061) );
  INV_X1 U5874 ( .A(n6712), .ZN(n5062) );
  AND2_X1 U5875 ( .A1(n5907), .A2(n6842), .ZN(n9162) );
  AND2_X1 U5876 ( .A1(n5907), .A2(n5886), .ZN(n9138) );
  NAND2_X1 U5877 ( .A1(n5290), .A2(n7141), .ZN(n7218) );
  AND2_X1 U5878 ( .A1(n7214), .A2(n7143), .ZN(n5290) );
  AOI21_X1 U5879 ( .B1(n9075), .B2(n9076), .A(n5076), .ZN(n9150) );
  INV_X1 U5880 ( .A(n9123), .ZN(n9168) );
  INV_X1 U5881 ( .A(n9153), .ZN(n9166) );
  OAI21_X1 U5882 ( .B1(n5118), .B2(n4917), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5140) );
  INV_X1 U5883 ( .A(n5067), .ZN(n4917) );
  OAI21_X1 U5884 ( .B1(n8295), .B2(n8294), .A(n8293), .ZN(n8296) );
  AND2_X1 U5885 ( .A1(n4659), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5886 ( .A1(n5081), .A2(n5083), .ZN(n5157) );
  NOR2_X1 U5887 ( .A1(n10053), .A2(n4628), .ZN(n10066) );
  NOR2_X1 U5888 ( .A1(n6553), .A2(n6519), .ZN(n4628) );
  INV_X1 U5889 ( .A(n4612), .ZN(n6680) );
  OAI21_X1 U5890 ( .B1(n6614), .B2(n4615), .A(n4613), .ZN(n10103) );
  NAND2_X1 U5891 ( .A1(n6613), .A2(n4616), .ZN(n10105) );
  AND2_X1 U5892 ( .A1(n6526), .A2(n6525), .ZN(n6650) );
  AND2_X1 U5893 ( .A1(n6773), .A2(n6772), .ZN(n6777) );
  INV_X1 U5894 ( .A(n4621), .ZN(n10117) );
  INV_X1 U5895 ( .A(n4619), .ZN(n10115) );
  INV_X1 U5896 ( .A(n4626), .ZN(n10181) );
  INV_X1 U5897 ( .A(n4624), .ZN(n10179) );
  AOI21_X1 U5898 ( .B1(n8160), .B2(n8163), .A(n8162), .ZN(n9438) );
  AOI21_X1 U5899 ( .B1(n8451), .B2(n8163), .A(n7976), .ZN(n9443) );
  NAND2_X1 U5900 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  OR2_X1 U5901 ( .A1(n9454), .A2(n10004), .ZN(n4852) );
  AND2_X1 U5902 ( .A1(n4854), .A2(n4853), .ZN(n9453) );
  AOI22_X1 U5903 ( .A1(n9275), .A2(n9988), .B1(n9990), .B2(n9246), .ZN(n4853)
         );
  NAND2_X1 U5904 ( .A1(n9247), .A2(n9985), .ZN(n4854) );
  AND2_X1 U5905 ( .A1(n5842), .A2(n5841), .ZN(n9253) );
  NAND2_X1 U5906 ( .A1(n9281), .A2(n4912), .ZN(n9263) );
  NAND2_X1 U5907 ( .A1(n4824), .A2(n4828), .ZN(n9289) );
  NAND2_X1 U5908 ( .A1(n9321), .A2(n4830), .ZN(n4824) );
  NAND2_X1 U5909 ( .A1(n5729), .A2(n5728), .ZN(n9485) );
  NAND2_X1 U5910 ( .A1(n4834), .A2(n8125), .ZN(n9380) );
  NAND2_X1 U5911 ( .A1(n9995), .A2(n8009), .ZN(n9417) );
  INV_X1 U5912 ( .A(n10221), .ZN(n9993) );
  NAND2_X1 U5913 ( .A1(n5574), .A2(n5573), .ZN(n10009) );
  NAND2_X1 U5914 ( .A1(n4876), .A2(n7878), .ZN(n7879) );
  NAND2_X1 U5915 ( .A1(n5548), .A2(n5547), .ZN(n9169) );
  NAND2_X1 U5916 ( .A1(n5519), .A2(n5518), .ZN(n7941) );
  NAND2_X1 U5917 ( .A1(n4866), .A2(n7721), .ZN(n7844) );
  NAND2_X1 U5918 ( .A1(n10207), .A2(n7352), .ZN(n9432) );
  NAND2_X1 U5919 ( .A1(n7552), .A2(n7412), .ZN(n7527) );
  NAND2_X1 U5920 ( .A1(n5395), .A2(n5394), .ZN(n10262) );
  NAND2_X1 U5921 ( .A1(n4848), .A2(n8319), .ZN(n7423) );
  INV_X1 U5922 ( .A(n9432), .ZN(n10213) );
  NAND2_X1 U5923 ( .A1(n7450), .A2(n7449), .ZN(n7448) );
  NAND2_X1 U5924 ( .A1(n6994), .A2(n6993), .ZN(n7450) );
  AND2_X1 U5925 ( .A1(n10207), .A2(n7045), .ZN(n10212) );
  OR2_X1 U5926 ( .A1(n6853), .A2(n6832), .ZN(n10279) );
  INV_X2 U5927 ( .A(n10271), .ZN(n10273) );
  INV_X1 U5928 ( .A(n10230), .ZN(n10231) );
  AND2_X1 U5929 ( .A1(n6514), .A2(n5880), .ZN(n10234) );
  NAND2_X1 U5930 ( .A1(n5152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5150) );
  OAI21_X1 U5931 ( .B1(n5149), .B2(n5390), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5151) );
  XNOR2_X1 U5932 ( .A(n6249), .B(n6248), .ZN(n7954) );
  XNOR2_X1 U5933 ( .A(n5113), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7944) );
  INV_X1 U5934 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U5935 ( .A1(n5117), .A2(n5116), .ZN(n7927) );
  INV_X1 U5936 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7826) );
  XNOR2_X1 U5937 ( .A(n5119), .B(n5111), .ZN(n7828) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U5939 ( .A1(n4965), .A2(n5743), .ZN(n5763) );
  INV_X1 U5940 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8363) );
  OR2_X1 U5941 ( .A1(n5098), .A2(n5097), .ZN(n5099) );
  OAI21_X1 U5942 ( .B1(n5096), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5098) );
  INV_X1 U5943 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7572) );
  INV_X1 U5944 ( .A(n6844), .ZN(n8343) );
  INV_X1 U5945 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7362) );
  INV_X1 U5946 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9637) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6720) );
  INV_X1 U5948 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6624) );
  INV_X1 U5949 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9748) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6583) );
  NOR2_X1 U5951 ( .A1(n9970), .A2(n10408), .ZN(n10399) );
  AOI21_X1 U5952 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10397), .ZN(n10396) );
  NOR2_X1 U5953 ( .A1(n10396), .A2(n10395), .ZN(n10394) );
  AOI21_X1 U5954 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10394), .ZN(n10393) );
  OAI21_X1 U5955 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10391), .ZN(n10389) );
  NAND2_X1 U5956 ( .A1(n4634), .A2(n6513), .ZN(P2_U3244) );
  OAI21_X1 U5957 ( .B1(n4576), .B2(n4635), .A(n6510), .ZN(n4634) );
  NAND2_X1 U5958 ( .A1(n4557), .A2(n4554), .ZN(P2_U3264) );
  AOI21_X1 U5959 ( .B1(n8679), .B2(n4919), .A(n4555), .ZN(n4554) );
  NAND2_X1 U5960 ( .A1(n8680), .A2(n4460), .ZN(n4557) );
  NAND2_X1 U5961 ( .A1(n4556), .A2(n8681), .ZN(n4555) );
  NAND2_X1 U5962 ( .A1(n4792), .A2(n4790), .ZN(P2_U3549) );
  OR2_X1 U5963 ( .A1(n10370), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5964 ( .A1(n8991), .A2(n10370), .ZN(n4792) );
  INV_X1 U5965 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5966 ( .A1(n6546), .A2(P1_U3084), .ZN(P1_U4006) );
  OAI21_X1 U5967 ( .B1(n9453), .B2(n10216), .A(n4849), .ZN(P1_U3263) );
  AOI21_X1 U5968 ( .B1(n9450), .B2(n9428), .A(n4850), .ZN(n4849) );
  NAND2_X1 U5969 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  INV_X1 U5970 ( .A(n9248), .ZN(n4851) );
  NOR2_X1 U5971 ( .A1(n7413), .A2(n4902), .ZN(n4467) );
  AND2_X1 U5972 ( .A1(n4981), .A2(n4455), .ZN(n4468) );
  INV_X1 U5973 ( .A(n8352), .ZN(n5858) );
  AND2_X1 U5974 ( .A1(n8845), .A2(n4502), .ZN(n4469) );
  NAND2_X1 U5975 ( .A1(n8869), .A2(n8870), .ZN(n8843) );
  NAND2_X1 U5976 ( .A1(n4600), .A2(n8758), .ZN(n8759) );
  INV_X1 U5977 ( .A(n6815), .ZN(n6741) );
  NAND2_X1 U5978 ( .A1(n7762), .A2(n7761), .ZN(n4470) );
  AND2_X1 U5979 ( .A1(n5350), .A2(n4716), .ZN(n4471) );
  INV_X1 U5980 ( .A(n5895), .ZN(n5184) );
  INV_X1 U5981 ( .A(n8082), .ZN(n4843) );
  OR2_X1 U5982 ( .A1(n8136), .A2(n8158), .ZN(n4472) );
  INV_X1 U5983 ( .A(n8146), .ZN(n4826) );
  OR2_X1 U5984 ( .A1(n8567), .A2(n10323), .ZN(n4473) );
  AND2_X1 U5985 ( .A1(n6930), .A2(n6928), .ZN(n4474) );
  OR2_X1 U5986 ( .A1(n4894), .A2(n8728), .ZN(n4475) );
  NOR2_X1 U5987 ( .A1(n8741), .A2(n5021), .ZN(n5019) );
  AND2_X1 U5988 ( .A1(n6555), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5989 ( .A1(n5053), .A2(n5051), .ZN(n9083) );
  AND2_X1 U5990 ( .A1(n6373), .A2(n6098), .ZN(n7785) );
  INV_X1 U5991 ( .A(n7785), .ZN(n4642) );
  NOR2_X1 U5992 ( .A1(n10262), .A2(n9181), .ZN(n4477) );
  AND2_X1 U5993 ( .A1(n9127), .A2(n9125), .ZN(n4478) );
  OR2_X1 U5994 ( .A1(n8977), .A2(n8557), .ZN(n4479) );
  OR2_X1 U5995 ( .A1(n8921), .A2(n8750), .ZN(n8714) );
  INV_X1 U5996 ( .A(n6454), .ZN(n4856) );
  AND2_X1 U5997 ( .A1(n4735), .A2(n4504), .ZN(n4480) );
  AND2_X1 U5998 ( .A1(n4759), .A2(n4758), .ZN(n4481) );
  AND2_X1 U5999 ( .A1(n7251), .A2(n7246), .ZN(n4482) );
  AND2_X1 U6000 ( .A1(n5933), .A2(n4560), .ZN(n4483) );
  XNOR2_X1 U6001 ( .A(n6310), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6464) );
  AND2_X1 U6002 ( .A1(n4961), .A2(n5781), .ZN(n4484) );
  NOR2_X1 U6003 ( .A1(n10100), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U6004 ( .A1(n6237), .A2(n6236), .ZN(n8909) );
  INV_X1 U6005 ( .A(n8909), .ZN(n4742) );
  OR2_X1 U6006 ( .A1(n7885), .A2(n7888), .ZN(n7886) );
  NAND2_X1 U6007 ( .A1(n5024), .A2(n4469), .ZN(n8841) );
  AND2_X1 U6008 ( .A1(n10241), .A2(n10247), .ZN(n4486) );
  AND2_X1 U6009 ( .A1(n4749), .A2(n4748), .ZN(n4487) );
  AND2_X1 U6010 ( .A1(n4723), .A2(n4546), .ZN(n4488) );
  INV_X1 U6011 ( .A(n7456), .ZN(n4805) );
  OR2_X1 U6012 ( .A1(n5566), .A2(n4786), .ZN(n4489) );
  OR2_X1 U6013 ( .A1(n7868), .A2(n7880), .ZN(n4490) );
  INV_X1 U6014 ( .A(n5850), .ZN(n5298) );
  NOR2_X1 U6015 ( .A1(n7051), .A2(n5161), .ZN(n5203) );
  INV_X1 U6016 ( .A(n6419), .ZN(n4878) );
  INV_X1 U6017 ( .A(n6837), .ZN(n6838) );
  INV_X1 U6018 ( .A(n7860), .ZN(n4596) );
  AND2_X1 U6019 ( .A1(n6377), .A2(n6378), .ZN(n7858) );
  NOR2_X1 U6020 ( .A1(n9363), .A2(n9348), .ZN(n4491) );
  AND3_X1 U6021 ( .A1(n5993), .A2(n5992), .A3(n5991), .ZN(n4492) );
  AOI21_X1 U6022 ( .B1(n8374), .B2(n8878), .A(n8373), .ZN(n8902) );
  INV_X1 U6023 ( .A(n8902), .ZN(n4609) );
  NAND4_X1 U6024 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n9188)
         );
  NAND2_X1 U6025 ( .A1(n4863), .A2(n8024), .ZN(n9317) );
  NAND3_X1 U6026 ( .A1(n5955), .A2(n5954), .A3(n5953), .ZN(n6756) );
  AOI21_X1 U6027 ( .B1(n8768), .B2(n7992), .A(n5075), .ZN(n4600) );
  INV_X1 U6028 ( .A(n7652), .ZN(n4706) );
  OR3_X1 U6029 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U6030 ( .A1(n5216), .A2(n6556), .ZN(n5219) );
  INV_X1 U6031 ( .A(n5219), .ZN(n4839) );
  AND2_X1 U6032 ( .A1(n9480), .A2(n9305), .ZN(n4494) );
  OR3_X1 U6033 ( .A1(n6388), .A2(n6387), .A3(n6386), .ZN(n4495) );
  MUX2_X1 U6034 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6551), .S(n5216), .Z(n10211)
         );
  AND2_X1 U6035 ( .A1(n8234), .A2(n8315), .ZN(n4496) );
  AND2_X1 U6036 ( .A1(n5454), .A2(n5453), .ZN(n4497) );
  NAND2_X1 U6037 ( .A1(n5705), .A2(n5704), .ZN(n9489) );
  OR2_X1 U6038 ( .A1(n6382), .A2(n7860), .ZN(n4498) );
  INV_X1 U6039 ( .A(n6338), .ZN(n4682) );
  NAND2_X1 U6040 ( .A1(n4636), .A2(n6025), .ZN(n7479) );
  AND2_X1 U6041 ( .A1(n5110), .A2(n4737), .ZN(n4499) );
  OR2_X1 U6042 ( .A1(n6491), .A2(n6490), .ZN(n4500) );
  AND2_X1 U6043 ( .A1(n8900), .A2(n8444), .ZN(n6455) );
  NOR2_X1 U6044 ( .A1(n8277), .A2(n8139), .ZN(n4501) );
  NAND2_X1 U6045 ( .A1(n8964), .A2(n8556), .ZN(n4502) );
  AND2_X1 U6046 ( .A1(n6476), .A2(n7503), .ZN(n4503) );
  NAND3_X1 U6047 ( .A1(n5943), .A2(n5942), .A3(n5941), .ZN(n6317) );
  OR2_X1 U6048 ( .A1(n8414), .A2(n5085), .ZN(n8500) );
  INV_X1 U6049 ( .A(n8288), .ZN(n4664) );
  AND2_X1 U6050 ( .A1(n5077), .A2(n5622), .ZN(n4504) );
  AND2_X1 U6051 ( .A1(n4711), .A2(n5412), .ZN(n4505) );
  NOR2_X1 U6052 ( .A1(n6418), .A2(n6405), .ZN(n8777) );
  INV_X1 U6053 ( .A(n4828), .ZN(n4827) );
  AOI21_X1 U6054 ( .B1(n4830), .B2(n9318), .A(n4829), .ZN(n4828) );
  INV_X1 U6055 ( .A(n6297), .ZN(n8691) );
  NAND2_X1 U6056 ( .A1(n6280), .A2(n6279), .ZN(n6297) );
  INV_X1 U6057 ( .A(n5075), .ZN(n4603) );
  AND2_X1 U6058 ( .A1(n5025), .A2(n5921), .ZN(n5935) );
  INV_X1 U6059 ( .A(n8728), .ZN(n4899) );
  NAND2_X1 U6060 ( .A1(n8714), .A2(n6434), .ZN(n8728) );
  NOR2_X1 U6061 ( .A1(n8791), .A2(n8811), .ZN(n4506) );
  INV_X1 U6062 ( .A(n7991), .ZN(n5005) );
  AND2_X1 U6063 ( .A1(n8791), .A2(n8811), .ZN(n4507) );
  AND2_X1 U6064 ( .A1(n6458), .A2(n6449), .ZN(n4508) );
  NOR2_X1 U6065 ( .A1(n8961), .A2(n8874), .ZN(n4509) );
  INV_X1 U6066 ( .A(n4831), .ZN(n4830) );
  OAI21_X1 U6067 ( .B1(n9318), .B2(n8178), .A(n4832), .ZN(n4831) );
  AND2_X1 U6068 ( .A1(n9887), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4510) );
  INV_X1 U6069 ( .A(n5021), .ZN(n5020) );
  NOR2_X1 U6070 ( .A1(n8764), .A2(n8749), .ZN(n5021) );
  AND2_X1 U6071 ( .A1(n5644), .A2(SI_18_), .ZN(n4511) );
  INV_X1 U6072 ( .A(n4941), .ZN(n4940) );
  NAND2_X1 U6073 ( .A1(n4942), .A2(n8391), .ZN(n4941) );
  OR2_X1 U6074 ( .A1(n8944), .A2(n8821), .ZN(n6180) );
  AND2_X1 U6075 ( .A1(n5457), .A2(SI_11_), .ZN(n4512) );
  INV_X1 U6076 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U6077 ( .A1(n6451), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6078 ( .A1(n5012), .A2(n7811), .ZN(n4513) );
  OAI21_X1 U6079 ( .B1(n4689), .B2(n4692), .A(n4508), .ZN(n4687) );
  INV_X1 U6080 ( .A(n5057), .ZN(n5056) );
  OR2_X1 U6081 ( .A1(n5509), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U6082 ( .A1(n4892), .A2(n4894), .ZN(n4514) );
  OR2_X1 U6083 ( .A1(n6454), .A2(n6297), .ZN(n4515) );
  INV_X1 U6084 ( .A(n8273), .ZN(n4671) );
  NAND2_X1 U6085 ( .A1(n5599), .A2(n5598), .ZN(n9510) );
  NOR2_X1 U6086 ( .A1(n7485), .A2(n7484), .ZN(n4516) );
  AND2_X1 U6087 ( .A1(n4897), .A2(n4895), .ZN(n4517) );
  AND2_X1 U6088 ( .A1(n8159), .A2(n8034), .ZN(n4518) );
  AND2_X1 U6089 ( .A1(n7880), .A2(n7878), .ZN(n4519) );
  INV_X1 U6090 ( .A(n4907), .ZN(n4906) );
  NOR2_X1 U6091 ( .A1(n8211), .A2(n4908), .ZN(n4907) );
  AND2_X1 U6092 ( .A1(n4783), .A2(n5589), .ZN(n4520) );
  AND2_X1 U6093 ( .A1(n4688), .A2(n4695), .ZN(n4521) );
  NAND2_X1 U6094 ( .A1(n5068), .A2(n5108), .ZN(n5118) );
  INV_X1 U6095 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5139) );
  OR2_X1 U6096 ( .A1(n4714), .A2(n4471), .ZN(n4522) );
  INV_X1 U6097 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4737) );
  OR2_X1 U6098 ( .A1(n5036), .A2(n5742), .ZN(n4523) );
  INV_X1 U6099 ( .A(n5381), .ZN(n4781) );
  AND2_X1 U6100 ( .A1(n8086), .A2(n8083), .ZN(n8193) );
  INV_X1 U6101 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5093) );
  AND2_X1 U6102 ( .A1(n5027), .A2(n5026), .ZN(n4524) );
  INV_X1 U6103 ( .A(n5215), .ZN(n5848) );
  INV_X1 U6104 ( .A(n5183), .ZN(n5846) );
  AND2_X1 U6105 ( .A1(n5156), .A2(n9887), .ZN(n5183) );
  AND2_X1 U6106 ( .A1(n4657), .A2(n5156), .ZN(n5708) );
  NOR2_X1 U6107 ( .A1(n8808), .A2(n4888), .ZN(n4887) );
  INV_X1 U6108 ( .A(n7995), .ZN(n4632) );
  XNOR2_X1 U6109 ( .A(n8930), .B(n8749), .ZN(n8758) );
  INV_X1 U6110 ( .A(n8758), .ZN(n5018) );
  AND2_X1 U6111 ( .A1(n9375), .A2(n4808), .ZN(n4525) );
  OAI211_X1 U6112 ( .C1(n6902), .C2(n7077), .A(n5989), .B(n5988), .ZN(n7468)
         );
  INV_X1 U6113 ( .A(n8808), .ZN(n5002) );
  XNOR2_X1 U6114 ( .A(n5170), .B(n5171), .ZN(n6553) );
  AND2_X1 U6115 ( .A1(n5361), .A2(n5328), .ZN(n6617) );
  OAI21_X1 U6116 ( .B1(n8528), .B2(n4941), .A(n4937), .ZN(n8512) );
  NAND2_X1 U6117 ( .A1(n4643), .A2(n6088), .ZN(n7786) );
  AND2_X1 U6118 ( .A1(n9125), .A2(n5034), .ZN(n4526) );
  NAND2_X1 U6119 ( .A1(n4724), .A2(n4727), .ZN(n9092) );
  NAND2_X1 U6120 ( .A1(n4640), .A2(n4638), .ZN(n7816) );
  AND3_X2 U6121 ( .A1(n4581), .A2(n4580), .A3(n4579), .ZN(n5921) );
  NAND2_X1 U6122 ( .A1(n5053), .A2(n5564), .ZN(n9082) );
  OAI21_X1 U6123 ( .B1(n7849), .B2(n6384), .A(n6383), .ZN(n8869) );
  AND2_X1 U6124 ( .A1(n7907), .A2(n9177), .ZN(n4527) );
  NAND2_X1 U6125 ( .A1(n7981), .A2(n7980), .ZN(n9444) );
  INV_X1 U6126 ( .A(n9444), .ZN(n4796) );
  NAND2_X1 U6127 ( .A1(n5091), .A2(n5090), .ZN(n5513) );
  NAND2_X1 U6128 ( .A1(n5813), .A2(n5812), .ZN(n9460) );
  INV_X1 U6129 ( .A(n9101), .ZN(n5048) );
  NAND2_X1 U6130 ( .A1(n6211), .A2(n6210), .ZN(n8924) );
  NAND2_X1 U6131 ( .A1(n5766), .A2(n5765), .ZN(n9471) );
  NAND2_X1 U6132 ( .A1(n7979), .A2(n7978), .ZN(n9451) );
  NAND2_X1 U6133 ( .A1(n6150), .A2(n6149), .ZN(n8954) );
  NAND2_X1 U6134 ( .A1(n5627), .A2(n5626), .ZN(n9503) );
  NAND2_X1 U6135 ( .A1(n6126), .A2(n6125), .ZN(n8964) );
  NAND2_X1 U6136 ( .A1(n5497), .A2(n5496), .ZN(n7907) );
  NAND2_X1 U6137 ( .A1(n8787), .A2(n4751), .ZN(n4752) );
  NAND2_X1 U6138 ( .A1(n8888), .A2(n4746), .ZN(n4747) );
  INV_X1 U6139 ( .A(n6200), .ZN(n8775) );
  NAND2_X1 U6140 ( .A1(n6189), .A2(n6188), .ZN(n6200) );
  AND2_X1 U6141 ( .A1(n9510), .A2(n9989), .ZN(n4528) );
  AND2_X1 U6142 ( .A1(n5015), .A2(n5013), .ZN(n4529) );
  NAND2_X1 U6143 ( .A1(n7651), .A2(n7650), .ZN(n7783) );
  INV_X1 U6144 ( .A(n7783), .ZN(n5016) );
  NOR2_X1 U6145 ( .A1(n7900), .A2(n7899), .ZN(n4530) );
  AND2_X1 U6146 ( .A1(n4943), .A2(n4940), .ZN(n4531) );
  INV_X1 U6147 ( .A(n5376), .ZN(n4716) );
  OR2_X1 U6148 ( .A1(n4485), .A2(n4615), .ZN(n4532) );
  INV_X1 U6149 ( .A(n5742), .ZN(n5034) );
  NAND2_X1 U6150 ( .A1(n5921), .A2(n4955), .ZN(n4533) );
  AND2_X1 U6151 ( .A1(n5783), .A2(SI_24_), .ZN(n4534) );
  INV_X1 U6152 ( .A(n7276), .ZN(n6947) );
  AND3_X1 U6153 ( .A1(n5965), .A2(n5964), .A3(n5079), .ZN(n7276) );
  INV_X1 U6154 ( .A(n5076), .ZN(n5050) );
  NAND2_X1 U6155 ( .A1(n6253), .A2(n6252), .ZN(n8904) );
  NAND2_X1 U6156 ( .A1(n5721), .A2(n5702), .ZN(n4535) );
  AND2_X1 U6157 ( .A1(n4797), .A2(n4796), .ZN(n4536) );
  NAND2_X1 U6158 ( .A1(n8833), .A2(n8851), .ZN(n4537) );
  AND2_X1 U6159 ( .A1(n5024), .A2(n4502), .ZN(n4538) );
  AND2_X1 U6160 ( .A1(n4889), .A2(n4887), .ZN(n4539) );
  XNOR2_X1 U6161 ( .A(n6493), .B(n6492), .ZN(n6463) );
  INV_X1 U6162 ( .A(n6463), .ZN(n4920) );
  NAND2_X1 U6163 ( .A1(n5650), .A2(n5649), .ZN(n9498) );
  INV_X1 U6164 ( .A(n9498), .ZN(n4815) );
  AND2_X1 U6165 ( .A1(n4800), .A2(n7536), .ZN(n4540) );
  AND2_X1 U6166 ( .A1(n7339), .A2(n4761), .ZN(n4541) );
  NAND2_X1 U6167 ( .A1(n5858), .A2(n9342), .ZN(n8170) );
  INV_X1 U6168 ( .A(n8314), .ZN(n4844) );
  INV_X1 U6169 ( .A(n8319), .ZN(n4847) );
  AND2_X1 U6170 ( .A1(n6702), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U6171 ( .A1(n7683), .A2(n5413), .ZN(n7670) );
  NAND2_X1 U6172 ( .A1(n4835), .A2(n8315), .ZN(n7194) );
  NAND2_X1 U6173 ( .A1(n4901), .A2(n4900), .ZN(n7598) );
  NAND2_X1 U6174 ( .A1(n6219), .A2(n6218), .ZN(n8921) );
  INV_X1 U6175 ( .A(n8921), .ZN(n4748) );
  NAND2_X1 U6176 ( .A1(n5377), .A2(n7586), .ZN(n7682) );
  OAI21_X1 U6177 ( .B1(n7670), .B2(n4721), .A(n4719), .ZN(n7885) );
  AOI21_X1 U6178 ( .B1(n7365), .B2(n6472), .A(n6000), .ZN(n7127) );
  NAND2_X1 U6179 ( .A1(n4713), .A2(n5376), .ZN(n7585) );
  OR2_X1 U6180 ( .A1(n7553), .A2(n8193), .ZN(n7552) );
  NAND2_X1 U6181 ( .A1(n7128), .A2(n6343), .ZN(n7328) );
  NAND2_X1 U6182 ( .A1(n5109), .A2(n5108), .ZN(n5878) );
  INV_X1 U6183 ( .A(n5013), .ZN(n5012) );
  NOR2_X1 U6184 ( .A1(n7785), .A2(n5014), .ZN(n5013) );
  OR2_X1 U6185 ( .A1(n6501), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4543) );
  AND2_X1 U6186 ( .A1(n7186), .A2(n7185), .ZN(n4544) );
  AND2_X1 U6187 ( .A1(n4848), .A2(n4846), .ZN(n4545) );
  NAND2_X1 U6188 ( .A1(n5437), .A2(n5436), .ZN(n4546) );
  OAI21_X1 U6189 ( .B1(n6320), .B2(n6467), .A(n6324), .ZN(n6752) );
  AND2_X1 U6190 ( .A1(n5086), .A2(n6265), .ZN(n4547) );
  INV_X1 U6191 ( .A(n6786), .ZN(n7023) );
  NOR2_X1 U6192 ( .A1(n6463), .A2(n4919), .ZN(n4548) );
  AND2_X1 U6193 ( .A1(n5062), .A2(n5061), .ZN(n4549) );
  INV_X1 U6194 ( .A(n7442), .ZN(n4756) );
  INV_X1 U6195 ( .A(n7734), .ZN(n4758) );
  NAND2_X1 U6196 ( .A1(n5466), .A2(n5465), .ZN(n7894) );
  INV_X1 U6197 ( .A(n7894), .ZN(n4803) );
  INV_X1 U6198 ( .A(n6953), .ZN(n10323) );
  AND2_X1 U6199 ( .A1(n7015), .A2(n6956), .ZN(n4550) );
  INV_X1 U6200 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6309) );
  INV_X1 U6201 ( .A(n9342), .ZN(n10200) );
  XNOR2_X1 U6202 ( .A(n5155), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5156) );
  AND2_X1 U6203 ( .A1(n6462), .A2(n6461), .ZN(n4984) );
  MUX2_X1 U6204 ( .A(n6354), .B(n6353), .S(n6461), .Z(n6357) );
  NAND2_X1 U6205 ( .A1(n5302), .A2(n5301), .ZN(n4551) );
  NAND2_X1 U6206 ( .A1(n8518), .A2(n8411), .ZN(n8414) );
  NAND2_X1 U6207 ( .A1(n7404), .A2(n7403), .ZN(n7615) );
  NAND2_X1 U6208 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  XNOR2_X1 U6209 ( .A(n4552), .B(n6166), .ZN(n8678) );
  NOR2_X2 U6210 ( .A1(n4558), .A2(n5919), .ZN(n5920) );
  NAND4_X1 U6211 ( .A1(n5915), .A2(n5916), .A3(n5917), .A4(n6291), .ZN(n4558)
         );
  OAI22_X1 U6212 ( .A1(n4461), .A2(n6557), .B1(n6902), .B2(n9917), .ZN(n4605)
         );
  NAND2_X1 U6213 ( .A1(n8540), .A2(n8428), .ZN(n8457) );
  OAI22_X2 U6214 ( .A1(n8058), .A2(n8059), .B1(n6945), .B2(n4918), .ZN(n6974)
         );
  OAI21_X2 U6215 ( .B1(n7062), .B2(n7061), .A(n7060), .ZN(n7242) );
  NAND2_X1 U6216 ( .A1(n5935), .A2(n5933), .ZN(n5923) );
  NAND2_X1 U6217 ( .A1(n5935), .A2(n4483), .ZN(n4562) );
  INV_X1 U6218 ( .A(n7368), .ZN(n8566) );
  AND2_X1 U6219 ( .A1(n4581), .A2(n4585), .ZN(n4855) );
  NAND2_X1 U6220 ( .A1(n7651), .A2(n4591), .ZN(n4592) );
  OAI21_X1 U6221 ( .B1(n5009), .B2(n4592), .A(n7985), .ZN(n4595) );
  OR2_X2 U6222 ( .A1(n4605), .A2(n4604), .ZN(n6815) );
  MUX2_X1 U6223 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6519), .S(n6553), .Z(n10054)
         );
  AND2_X2 U6224 ( .A1(n4630), .A2(n4629), .ZN(n8701) );
  OR2_X2 U6225 ( .A1(n8713), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U6226 ( .A1(n7507), .A2(n4637), .ZN(n4640) );
  NAND2_X1 U6227 ( .A1(n6298), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U6228 ( .A1(n7330), .A2(n6345), .ZN(n7476) );
  NAND3_X1 U6229 ( .A1(n7128), .A2(n6343), .A3(n6035), .ZN(n7330) );
  NAND2_X1 U6230 ( .A1(n7127), .A2(n7129), .ZN(n7128) );
  OAI211_X1 U6231 ( .C1(n6874), .C2(n4654), .A(n6876), .B(n4650), .ZN(n6877)
         );
  NAND2_X1 U6232 ( .A1(n4653), .A2(n6875), .ZN(n4650) );
  INV_X1 U6233 ( .A(n8182), .ZN(n6874) );
  INV_X1 U6234 ( .A(n5156), .ZN(n4658) );
  NAND3_X1 U6235 ( .A1(n5167), .A2(n5166), .A3(n4655), .ZN(n6837) );
  NAND3_X1 U6236 ( .A1(n4658), .A2(P1_REG1_REG_1__SCAN_IN), .A3(n4657), .ZN(
        n4659) );
  AND2_X2 U6237 ( .A1(n4658), .A2(n9887), .ZN(n8046) );
  NAND2_X1 U6238 ( .A1(n4835), .A2(n4496), .ZN(n4662) );
  NAND2_X1 U6239 ( .A1(n8156), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U6240 ( .A1(n8157), .A2(n9244), .ZN(n4668) );
  NAND2_X1 U6241 ( .A1(n6441), .A2(n4521), .ZN(n4685) );
  NAND2_X1 U6242 ( .A1(n4685), .A2(n4686), .ZN(n6459) );
  INV_X1 U6243 ( .A(n4699), .ZN(n6336) );
  AND2_X1 U6244 ( .A1(n6474), .A2(n6340), .ZN(n4697) );
  NAND2_X1 U6245 ( .A1(n4699), .A2(n6461), .ZN(n4698) );
  NAND2_X1 U6246 ( .A1(n4701), .A2(n6432), .ZN(n4700) );
  NAND2_X1 U6247 ( .A1(n4473), .A2(n6474), .ZN(n4701) );
  INV_X1 U6248 ( .A(n4708), .ZN(n5143) );
  NAND2_X1 U6249 ( .A1(n5096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6250 ( .A1(n7315), .A2(n4522), .ZN(n4712) );
  NAND2_X1 U6251 ( .A1(n7670), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U6252 ( .A1(n4718), .A2(n4717), .ZN(n5055) );
  NAND2_X1 U6253 ( .A1(n9158), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U6254 ( .A1(n9111), .A2(n4732), .ZN(n4731) );
  INV_X1 U6255 ( .A(n9068), .ZN(n4734) );
  NAND2_X1 U6256 ( .A1(n9111), .A2(n5699), .ZN(n9067) );
  NAND3_X1 U6257 ( .A1(n5089), .A2(n5247), .A3(n4736), .ZN(n5464) );
  INV_X1 U6258 ( .A(n5464), .ZN(n5091) );
  INV_X1 U6259 ( .A(n5921), .ZN(n6121) );
  NOR2_X1 U6260 ( .A1(n6501), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U6261 ( .A1(n5921), .A2(n5920), .ZN(n6501) );
  NOR2_X1 U6262 ( .A1(n8719), .A2(n8909), .ZN(n8697) );
  INV_X1 U6263 ( .A(n4747), .ZN(n8853) );
  INV_X1 U6264 ( .A(n4752), .ZN(n8761) );
  NAND2_X1 U6265 ( .A1(n4970), .A2(n4766), .ZN(n4764) );
  OR2_X1 U6266 ( .A1(n4970), .A2(n5641), .ZN(n4774) );
  NAND2_X1 U6267 ( .A1(n4775), .A2(n5378), .ZN(n4777) );
  NAND2_X1 U6268 ( .A1(n5378), .A2(n5381), .ZN(n4778) );
  OAI21_X1 U6269 ( .B1(n5378), .B2(n5379), .A(n5381), .ZN(n5414) );
  NAND3_X1 U6270 ( .A1(n4777), .A2(n4975), .A3(n4776), .ZN(n5486) );
  NAND2_X1 U6271 ( .A1(n5512), .A2(n4784), .ZN(n4782) );
  NAND2_X1 U6272 ( .A1(n4782), .A2(n4520), .ZN(n5592) );
  NAND2_X1 U6273 ( .A1(n5512), .A2(n5511), .ZN(n5541) );
  INV_X1 U6274 ( .A(n10235), .ZN(n8308) );
  XNOR2_X2 U6275 ( .A(n9188), .B(n10235), .ZN(n8184) );
  AND2_X2 U6276 ( .A1(n4795), .A2(n4840), .ZN(n10235) );
  AND2_X1 U6277 ( .A1(n4837), .A2(n4836), .ZN(n4795) );
  AND2_X1 U6278 ( .A1(n9283), .A2(n4799), .ZN(n9250) );
  NAND3_X1 U6279 ( .A1(n4805), .A2(n10197), .A3(n10241), .ZN(n7189) );
  NAND2_X1 U6280 ( .A1(n5151), .A2(n5150), .ZN(n5153) );
  NAND2_X1 U6281 ( .A1(n6460), .A2(n6432), .ZN(n4982) );
  NAND2_X1 U6282 ( .A1(n4983), .A2(n4982), .ZN(n4981) );
  NOR2_X2 U6283 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6291) );
  AOI21_X1 U6284 ( .B1(n6459), .B2(n6461), .A(n4984), .ZN(n4983) );
  NAND2_X1 U6285 ( .A1(n7601), .A2(n8194), .ZN(n4816) );
  NAND2_X1 U6286 ( .A1(n7528), .A2(n8089), .ZN(n4817) );
  OAI21_X1 U6287 ( .B1(n9321), .B2(n4823), .A(n4819), .ZN(n4818) );
  INV_X1 U6288 ( .A(n4818), .ZN(n9256) );
  NAND2_X1 U6289 ( .A1(n4834), .A2(n4833), .ZN(n9361) );
  OAI21_X1 U6290 ( .B1(n7414), .B2(n4845), .A(n4842), .ZN(n7555) );
  OAI21_X2 U6291 ( .B1(n9984), .B2(n8040), .A(n8257), .ZN(n9419) );
  NAND2_X2 U6292 ( .A1(n4490), .A2(n8254), .ZN(n9984) );
  INV_X2 U6293 ( .A(n5118), .ZN(n5112) );
  NAND2_X1 U6294 ( .A1(n5112), .A2(n5066), .ZN(n5135) );
  NAND2_X1 U6295 ( .A1(n4855), .A2(n5987), .ZN(n4992) );
  INV_X1 U6296 ( .A(n6456), .ZN(n4857) );
  NAND2_X1 U6297 ( .A1(n4863), .A2(n4861), .ZN(n8026) );
  NAND2_X2 U6298 ( .A1(n4868), .A2(n4867), .ZN(n8305) );
  NAND2_X1 U6299 ( .A1(n9997), .A2(n4873), .ZN(n4872) );
  NAND2_X1 U6300 ( .A1(n4876), .A2(n4519), .ZN(n10022) );
  NAND2_X1 U6301 ( .A1(n8818), .A2(n6400), .ZN(n4886) );
  NAND2_X1 U6302 ( .A1(n7553), .A2(n4467), .ZN(n4901) );
  INV_X1 U6303 ( .A(n9298), .ZN(n4911) );
  NAND2_X1 U6304 ( .A1(n9298), .A2(n4907), .ZN(n4903) );
  NOR2_X1 U6305 ( .A1(n9298), .A2(n8027), .ZN(n9280) );
  NAND3_X1 U6306 ( .A1(n4920), .A2(n7666), .A3(n4919), .ZN(n4922) );
  INV_X1 U6307 ( .A(n4455), .ZN(n6314) );
  OAI21_X2 U6308 ( .B1(n7622), .B2(n4927), .A(n4923), .ZN(n4929) );
  INV_X1 U6309 ( .A(n4924), .ZN(n4923) );
  OR2_X1 U6310 ( .A1(n7758), .A2(n4928), .ZN(n4927) );
  INV_X1 U6311 ( .A(n4929), .ZN(n7763) );
  INV_X1 U6312 ( .A(n7017), .ZN(n4934) );
  INV_X1 U6313 ( .A(n7018), .ZN(n4935) );
  NAND2_X1 U6314 ( .A1(n7247), .A2(n4482), .ZN(n7398) );
  NAND2_X1 U6315 ( .A1(n7398), .A2(n7397), .ZN(n7404) );
  OAI21_X2 U6316 ( .B1(n7916), .B2(n4948), .A(n4945), .ZN(n8385) );
  NAND3_X1 U6317 ( .A1(n4953), .A2(n4952), .A3(n8541), .ZN(n8540) );
  INV_X1 U6318 ( .A(n8422), .ZN(n4953) );
  AND2_X1 U6319 ( .A1(n5921), .A2(n4957), .ZN(n6294) );
  NAND2_X1 U6320 ( .A1(n5745), .A2(n4484), .ZN(n4960) );
  OR2_X1 U6321 ( .A1(n5745), .A2(n5744), .ZN(n4965) );
  NAND2_X1 U6322 ( .A1(n5592), .A2(n5591), .ZN(n5621) );
  NAND2_X1 U6323 ( .A1(n5416), .A2(n5415), .ZN(n5438) );
  NAND2_X1 U6324 ( .A1(n4986), .A2(n4547), .ZN(n6278) );
  NAND3_X1 U6325 ( .A1(n4990), .A2(n4989), .A3(n5129), .ZN(n5168) );
  NAND2_X1 U6326 ( .A1(n4992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U6327 ( .A1(n4995), .A2(n4996), .ZN(n8768) );
  NAND2_X1 U6328 ( .A1(n8759), .A2(n5020), .ZN(n8740) );
  NAND2_X1 U6329 ( .A1(n8866), .A2(n4469), .ZN(n5023) );
  INV_X1 U6330 ( .A(n5024), .ZN(n8867) );
  AND2_X1 U6331 ( .A1(n5920), .A2(n4524), .ZN(n5025) );
  OAI21_X1 U6332 ( .B1(n5049), .B2(n5037), .A(n5041), .ZN(n5853) );
  OAI21_X1 U6333 ( .B1(n5049), .B2(n5038), .A(n5040), .ZN(n9075) );
  INV_X1 U6334 ( .A(n5049), .ZN(n5047) );
  NAND2_X1 U6335 ( .A1(n5055), .A2(n5054), .ZN(n7935) );
  NAND2_X1 U6336 ( .A1(n6712), .A2(n6818), .ZN(n5059) );
  NAND2_X1 U6337 ( .A1(n6713), .A2(n6818), .ZN(n5060) );
  NAND3_X1 U6338 ( .A1(n6819), .A2(n5060), .A3(n5059), .ZN(n6821) );
  NAND2_X1 U6339 ( .A1(n8071), .A2(n8070), .ZN(n8069) );
  XNOR2_X1 U6340 ( .A(n8045), .B(n8034), .ZN(n8054) );
  NAND2_X1 U6341 ( .A1(n7438), .A2(n7437), .ZN(n7436) );
  NAND2_X1 U6342 ( .A1(n6324), .A2(n6322), .ZN(n6467) );
  NAND2_X1 U6343 ( .A1(n6285), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U6344 ( .A1(n4464), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5942) );
  OR2_X1 U6345 ( .A1(n4465), .A2(n5951), .ZN(n5954) );
  NAND2_X1 U6346 ( .A1(n5923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  OAI21_X2 U6347 ( .B1(n7723), .B2(n7722), .A(n8100), .ZN(n7724) );
  NAND4_X2 U6348 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n6786)
         );
  NAND2_X1 U6349 ( .A1(n6285), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5932) );
  INV_X1 U6350 ( .A(n5708), .ZN(n5734) );
  INV_X1 U6351 ( .A(n5927), .ZN(n5926) );
  INV_X1 U6352 ( .A(n8046), .ZN(n5821) );
  OAI22_X2 U6353 ( .A1(n8495), .A2(n8494), .B1(n8387), .B2(n8386), .ZN(n8528)
         );
  NAND2_X2 U6354 ( .A1(n6893), .A2(n10306), .ZN(n8568) );
  OR4_X1 U6355 ( .A1(n10293), .A2(n6507), .A3(n6798), .A4(n8850), .ZN(n5069)
         );
  NAND2_X2 U6356 ( .A1(n7263), .A2(n8882), .ZN(n8896) );
  AND2_X1 U6357 ( .A1(n6123), .A2(n6122), .ZN(n5070) );
  AND2_X1 U6358 ( .A1(n5511), .A2(n5491), .ZN(n5071) );
  INV_X1 U6359 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6018) );
  OR2_X1 U6360 ( .A1(n5968), .A2(n7289), .ZN(n5072) );
  AND2_X1 U6361 ( .A1(n9059), .A2(n9058), .ZN(n5073) );
  AND2_X1 U6362 ( .A1(n8775), .A2(n8477), .ZN(n5075) );
  AND2_X1 U6363 ( .A1(n5804), .A2(n5803), .ZN(n5076) );
  AND2_X1 U6364 ( .A1(n5595), .A2(n5094), .ZN(n5077) );
  OR2_X1 U6365 ( .A1(n6902), .A2(n7096), .ZN(n5079) );
  INV_X1 U6366 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6066) );
  AND2_X1 U6367 ( .A1(n5439), .A2(n5420), .ZN(n5080) );
  AND2_X1 U6368 ( .A1(n5415), .A2(n5385), .ZN(n5082) );
  AND2_X1 U6369 ( .A1(n5183), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5083) );
  AOI21_X1 U6370 ( .B1(n8744), .B2(n5952), .A(n6217), .ZN(n8486) );
  INV_X1 U6371 ( .A(n6369), .ZN(n6087) );
  NOR2_X1 U6372 ( .A1(n6368), .A2(n7654), .ZN(n5084) );
  XOR2_X1 U6373 ( .A(n8930), .B(n8436), .Z(n5085) );
  NAND2_X1 U6374 ( .A1(n10221), .A2(n7418), .ZN(n10207) );
  INV_X2 U6375 ( .A(n10207), .ZN(n10216) );
  OR2_X1 U6376 ( .A1(n6276), .A2(SI_29_), .ZN(n5086) );
  INV_X1 U6377 ( .A(n8214), .ZN(n8034) );
  NAND2_X1 U6378 ( .A1(n8069), .A2(n5165), .ZN(n6670) );
  INV_X1 U6379 ( .A(n5203), .ZN(n5850) );
  INV_X1 U6380 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6381 ( .A1(n8504), .A2(n8417), .ZN(n8415) );
  NAND2_X1 U6382 ( .A1(n7555), .A2(n8193), .ZN(n7528) );
  NAND2_X1 U6383 ( .A1(n8418), .A2(n8503), .ZN(n8419) );
  INV_X1 U6384 ( .A(n6192), .ZN(n6190) );
  AND2_X1 U6385 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n6004) );
  NOR2_X1 U6386 ( .A1(n8845), .A2(n6390), .ZN(n6148) );
  INV_X1 U6387 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6155) );
  INV_X1 U6388 ( .A(n7685), .ZN(n5412) );
  INV_X1 U6389 ( .A(n5674), .ZN(n5672) );
  AND2_X1 U6390 ( .A1(n9471), .A2(n9290), .ZN(n8027) );
  INV_X1 U6391 ( .A(SI_22_), .ZN(n9816) );
  INV_X1 U6392 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5622) );
  INV_X1 U6393 ( .A(SI_15_), .ZN(n5542) );
  NAND2_X1 U6394 ( .A1(n8436), .A2(n7443), .ZN(n6794) );
  AOI21_X1 U6395 ( .B1(n8423), .B2(n8484), .A(n8483), .ZN(n8422) );
  OR2_X1 U6396 ( .A1(n6203), .A2(n8462), .ZN(n6212) );
  NAND2_X1 U6397 ( .A1(n6128), .A2(n6127), .ZN(n6141) );
  INV_X1 U6398 ( .A(n8486), .ZN(n7993) );
  OR2_X1 U6399 ( .A1(n6104), .A2(n6103), .ZN(n6130) );
  NAND2_X1 U6400 ( .A1(n5946), .A2(n10307), .ZN(n6468) );
  NOR2_X1 U6401 ( .A1(n8002), .A2(n8365), .ZN(n8001) );
  AND2_X1 U6402 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5467) );
  INV_X1 U6403 ( .A(n5686), .ZN(n5687) );
  OR2_X1 U6404 ( .A1(n5768), .A2(n5767), .ZN(n5791) );
  NAND2_X1 U6405 ( .A1(n5672), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5706) );
  INV_X1 U6406 ( .A(n5859), .ZN(n8304) );
  INV_X1 U6407 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6408 ( .A1(n5255), .A2(n9798), .ZN(n5199) );
  INV_X1 U6409 ( .A(n8552), .ZN(n8443) );
  OR2_X1 U6410 ( .A1(n6212), .A2(n9629), .ZN(n6228) );
  NAND2_X1 U6411 ( .A1(n6140), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6164) );
  OR2_X1 U6412 ( .A1(n8546), .A2(n8850), .ZN(n8531) );
  OR2_X1 U6413 ( .A1(n6254), .A2(n8441), .ZN(n6269) );
  INV_X1 U6414 ( .A(n8507), .ZN(n8744) );
  INV_X1 U6415 ( .A(n6784), .ZN(n6895) );
  AND2_X1 U6416 ( .A1(n8944), .A2(n8794), .ZN(n7991) );
  INV_X1 U6417 ( .A(n8555), .ZN(n8851) );
  OR2_X1 U6418 ( .A1(n7734), .A2(n7658), .ZN(n6478) );
  NAND2_X1 U6419 ( .A1(n6805), .A2(n6807), .ZN(n8882) );
  INV_X1 U6420 ( .A(n8560), .ZN(n7658) );
  INV_X1 U6421 ( .A(n8878), .ZN(n8847) );
  INV_X1 U6422 ( .A(n6472), .ZN(n7366) );
  OR2_X1 U6423 ( .A1(n6807), .A2(n7259), .ZN(n7034) );
  OR2_X1 U6424 ( .A1(n6048), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6060) );
  INV_X1 U6425 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  OR2_X1 U6426 ( .A1(n5652), .A2(n5651), .ZN(n5674) );
  OR2_X1 U6427 ( .A1(n5602), .A2(n5601), .ZN(n5629) );
  AND2_X1 U6428 ( .A1(n10263), .A2(n8177), .ZN(n5899) );
  NAND2_X1 U6429 ( .A1(n5815), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5890) );
  OR2_X1 U6430 ( .A1(n5706), .A2(n9069), .ZN(n5732) );
  OR2_X1 U6431 ( .A1(n8177), .A2(n6515), .ZN(n6516) );
  OR2_X1 U6432 ( .A1(n7044), .A2(n8343), .ZN(n10196) );
  AND2_X1 U6433 ( .A1(n8109), .A2(n8247), .ZN(n8199) );
  INV_X1 U6434 ( .A(n9182), .ZN(n7530) );
  NAND2_X1 U6435 ( .A1(n7960), .A2(n6871), .ZN(n6872) );
  INV_X1 U6436 ( .A(n10263), .ZN(n9511) );
  INV_X1 U6437 ( .A(n8203), .ZN(n7880) );
  OR2_X1 U6438 ( .A1(n8177), .A2(n6842), .ZN(n9425) );
  NOR2_X1 U6439 ( .A1(n7927), .A2(n7828), .ZN(n5120) );
  AND2_X1 U6440 ( .A1(n5591), .A2(n5571), .ZN(n5589) );
  OAI21_X1 U6441 ( .B1(n5255), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5199), .ZN(
        n5222) );
  INV_X1 U6442 ( .A(n8522), .ZN(n8548) );
  AND2_X1 U6443 ( .A1(n10348), .A2(n6784), .ZN(n6785) );
  AND2_X1 U6444 ( .A1(n6269), .A2(n6255), .ZN(n8440) );
  INV_X1 U6445 ( .A(n6812), .ZN(n6893) );
  INV_X1 U6446 ( .A(n10285), .ZN(n10281) );
  INV_X1 U6447 ( .A(n10282), .ZN(n9924) );
  AND2_X1 U6448 ( .A1(n6919), .A2(n6918), .ZN(n10282) );
  NAND2_X1 U6449 ( .A1(n6452), .A2(n6449), .ZN(n8369) );
  INV_X1 U6450 ( .A(n8850), .ZN(n8871) );
  OR2_X1 U6451 ( .A1(n4548), .A2(n6754), .ZN(n8878) );
  NOR2_X1 U6452 ( .A1(n7032), .A2(n7034), .ZN(n6740) );
  OR2_X1 U6453 ( .A1(n6751), .A2(n6314), .ZN(n10335) );
  AND2_X1 U6454 ( .A1(n8881), .A2(n10335), .ZN(n8981) );
  INV_X1 U6455 ( .A(n8981), .ZN(n10354) );
  AND2_X1 U6456 ( .A1(n7033), .A2(n7032), .ZN(n7260) );
  AND2_X1 U6457 ( .A1(n6024), .A2(n6048), .ZN(n8587) );
  INV_X1 U6458 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5986) );
  OAI21_X1 U6459 ( .B1(n9253), .B2(n9123), .A(n5911), .ZN(n5912) );
  AND2_X1 U6460 ( .A1(n5899), .A2(n5884), .ZN(n9115) );
  OR2_X1 U6461 ( .A1(n5890), .A2(n5889), .ZN(n8037) );
  NAND2_X1 U6462 ( .A1(n6516), .A2(n6546), .ZN(n6644) );
  INV_X1 U6463 ( .A(n10178), .ZN(n10106) );
  INV_X1 U6464 ( .A(n10190), .ZN(n10172) );
  INV_X1 U6465 ( .A(n10074), .ZN(n10184) );
  INV_X1 U6466 ( .A(n10196), .ZN(n7352) );
  AND2_X1 U6467 ( .A1(n8126), .A2(n8125), .ZN(n9394) );
  AND2_X1 U6468 ( .A1(n10207), .A2(n7354), .ZN(n7968) );
  OR2_X1 U6469 ( .A1(n8170), .A2(n6844), .ZN(n9937) );
  OR2_X1 U6470 ( .A1(n7044), .A2(n7043), .ZN(n10263) );
  AND2_X1 U6471 ( .A1(n7561), .A2(n9937), .ZN(n10016) );
  INV_X1 U6472 ( .A(n10016), .ZN(n10252) );
  OR2_X1 U6473 ( .A1(n6852), .A2(n9881), .ZN(n7040) );
  AND2_X1 U6474 ( .A1(n7744), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U6475 ( .A(n5459), .B(n5455), .ZN(n6595) );
  AND2_X1 U6476 ( .A1(n6556), .A2(P1_U3084), .ZN(n7950) );
  OAI21_X1 U6477 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10376), .ZN(n10405) );
  INV_X1 U6478 ( .A(n9913), .ZN(n10287) );
  INV_X1 U6479 ( .A(n4453), .ZN(n8551) );
  NAND2_X1 U6480 ( .A1(n6919), .A2(n6509), .ZN(n10283) );
  INV_X1 U6481 ( .A(n8891), .ZN(n8695) );
  INV_X1 U6482 ( .A(n10370), .ZN(n10368) );
  INV_X1 U6483 ( .A(n10358), .ZN(n10356) );
  NOR2_X1 U6484 ( .A1(n10293), .A2(n10292), .ZN(n10299) );
  INV_X1 U6485 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10304) );
  INV_X1 U6486 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7956) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7669) );
  INV_X1 U6488 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6622) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9741) );
  INV_X1 U6490 ( .A(n7430), .ZN(n7518) );
  AND2_X1 U6491 ( .A1(n5906), .A2(n6674), .ZN(n9153) );
  AND2_X1 U6492 ( .A1(n5883), .A2(n10221), .ZN(n9123) );
  INV_X1 U6493 ( .A(n9115), .ZN(n9172) );
  NAND2_X1 U6494 ( .A1(n5825), .A2(n5824), .ZN(n9291) );
  NAND2_X1 U6495 ( .A1(n9225), .A2(n6842), .ZN(n10178) );
  OR2_X1 U6496 ( .A1(n6644), .A2(n6544), .ZN(n10190) );
  INV_X1 U6497 ( .A(n10101), .ZN(n10193) );
  AND2_X1 U6498 ( .A1(n9992), .A2(n9991), .ZN(n10011) );
  NAND2_X1 U6499 ( .A1(n10207), .A2(n10195), .ZN(n10004) );
  OR2_X1 U6500 ( .A1(n6853), .A2(n7040), .ZN(n10271) );
  AND2_X1 U6501 ( .A1(n10234), .A2(n10222), .ZN(n10230) );
  AOI21_X1 U6502 ( .B1(n5877), .B2(n5864), .A(n5863), .ZN(n9881) );
  INV_X1 U6503 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9658) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9753) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U6506 ( .A1(n10399), .A2(n10398), .ZN(n10397) );
  OAI21_X1 U6507 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10388), .ZN(n10386) );
  INV_X1 U6508 ( .A(n8568), .ZN(P2_U3966) );
  AND2_X2 U6509 ( .A1(n5088), .A2(n5087), .ZN(n5247) );
  NAND2_X1 U6510 ( .A1(n5145), .A2(n5095), .ZN(n5096) );
  NAND2_X1 U6511 ( .A1(n5143), .A2(n5099), .ZN(n5859) );
  XNOR2_X1 U6512 ( .A(n5100), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U6513 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5104) );
  NOR2_X1 U6514 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5103) );
  NOR2_X1 U6515 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5102) );
  NOR2_X1 U6516 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5101) );
  NAND4_X1 U6517 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n5107)
         );
  NAND4_X1 U6518 ( .A1(n5093), .A2(n5622), .A3(n5595), .A4(n5105), .ZN(n5106)
         );
  NAND2_X1 U6519 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6520 ( .A1(n5116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5113) );
  INV_X1 U6521 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6522 ( .A1(n5115), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6523 ( .A1(n5118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5119) );
  INV_X1 U6524 ( .A(n6514), .ZN(n5161) );
  NAND2_X1 U6525 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  NAND2_X1 U6526 ( .A1(n5124), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5125) );
  INV_X1 U6527 ( .A(SI_0_), .ZN(n5127) );
  INV_X1 U6528 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5126) );
  OAI21_X1 U6529 ( .B1(n6555), .B2(n5127), .A(n5126), .ZN(n5130) );
  AND2_X1 U6530 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5129) );
  AND2_X1 U6531 ( .A1(n5130), .A2(n5168), .ZN(n6551) );
  NAND2_X1 U6532 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U6533 ( .A1(n5135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5136) );
  INV_X1 U6534 ( .A(n5149), .ZN(n5137) );
  NAND2_X2 U6535 ( .A1(n5138), .A2(n5137), .ZN(n5886) );
  INV_X1 U6536 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U6537 ( .A1(n6514), .A2(n10058), .ZN(n5141) );
  AOI21_X1 U6538 ( .B1(n5203), .B2(n10211), .A(n5141), .ZN(n5142) );
  INV_X1 U6539 ( .A(n5142), .ZN(n5160) );
  NAND2_X1 U6540 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6541 ( .A1(n5858), .A2(n7043), .ZN(n5148) );
  NAND2_X1 U6542 ( .A1(n5148), .A2(n5215), .ZN(n5175) );
  NAND2_X1 U6543 ( .A1(n8046), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6544 ( .A1(n5184), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5158) );
  NAND3_X1 U6545 ( .A1(n5159), .A2(n5158), .A3(n5157), .ZN(n6606) );
  NAND2_X1 U6546 ( .A1(n6606), .A2(n5203), .ZN(n5163) );
  AOI22_X1 U6547 ( .A1(n5814), .A2(n10211), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5161), .ZN(n5162) );
  NAND2_X1 U6548 ( .A1(n5163), .A2(n5162), .ZN(n8070) );
  INV_X1 U6549 ( .A(n8070), .ZN(n5164) );
  NAND2_X1 U6550 ( .A1(n5164), .A2(n5374), .ZN(n5165) );
  NAND2_X1 U6551 ( .A1(n5708), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6552 ( .A1(n5183), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5166) );
  INV_X1 U6553 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U6554 ( .A1(n6837), .A2(n5203), .ZN(n5173) );
  CLKBUF_X3 U6555 ( .A(n5255), .Z(n6556) );
  NAND3_X1 U6556 ( .A1(n5128), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5169) );
  NAND2_X1 U6557 ( .A1(n5169), .A2(n5168), .ZN(n5196) );
  XNOR2_X1 U6558 ( .A(n5196), .B(n9660), .ZN(n5195) );
  MUX2_X1 U6559 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5255), .Z(n5194) );
  XNOR2_X1 U6560 ( .A(n5195), .B(n5194), .ZN(n6558) );
  INV_X1 U6561 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6562 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5170) );
  INV_X1 U6563 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U6564 ( .A1(n5814), .A2(n8305), .ZN(n5172) );
  NAND2_X1 U6565 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  XNOR2_X1 U6566 ( .A(n5174), .B(n5828), .ZN(n5179) );
  NAND2_X1 U6567 ( .A1(n6670), .A2(n5179), .ZN(n5178) );
  NAND2_X1 U6568 ( .A1(n5298), .A2(n8305), .ZN(n5176) );
  NAND2_X1 U6569 ( .A1(n5177), .A2(n5176), .ZN(n6671) );
  NAND2_X1 U6570 ( .A1(n5178), .A2(n6671), .ZN(n5182) );
  INV_X1 U6571 ( .A(n6670), .ZN(n5180) );
  INV_X1 U6572 ( .A(n5179), .ZN(n6672) );
  NAND2_X1 U6573 ( .A1(n5180), .A2(n6672), .ZN(n5181) );
  NAND2_X1 U6574 ( .A1(n5182), .A2(n5181), .ZN(n6712) );
  NAND2_X1 U6575 ( .A1(n5708), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6576 ( .A1(n5183), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6577 ( .A1(n8046), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6578 ( .A1(n5184), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6579 ( .A1(n9188), .A2(n5203), .ZN(n5201) );
  NOR2_X1 U6580 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5191) );
  INV_X1 U6581 ( .A(n5191), .ZN(n5189) );
  NAND2_X1 U6582 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5189), .ZN(n5190) );
  INV_X1 U6583 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5192) );
  MUX2_X1 U6584 ( .A(n5190), .B(P1_IR_REG_31__SCAN_IN), .S(n5192), .Z(n5193)
         );
  NAND2_X1 U6585 ( .A1(n5192), .A2(n5191), .ZN(n5217) );
  AND2_X1 U6586 ( .A1(n5193), .A2(n5217), .ZN(n6531) );
  INV_X1 U6587 ( .A(n6531), .ZN(n10073) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U6589 ( .A1(n5195), .A2(n5194), .ZN(n5198) );
  NAND2_X1 U6590 ( .A1(n5196), .A2(SI_1_), .ZN(n5197) );
  NAND2_X1 U6591 ( .A1(n5198), .A2(n5197), .ZN(n5221) );
  INV_X1 U6592 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6560) );
  XNOR2_X1 U6593 ( .A(n5222), .B(SI_2_), .ZN(n5220) );
  XNOR2_X1 U6594 ( .A(n5221), .B(n5220), .ZN(n6559) );
  NAND2_X1 U6595 ( .A1(n5814), .A2(n8308), .ZN(n5200) );
  NAND2_X1 U6596 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  XNOR2_X1 U6597 ( .A(n5202), .B(n5828), .ZN(n5205) );
  NAND2_X1 U6598 ( .A1(n5203), .A2(n8308), .ZN(n5204) );
  AND2_X1 U6599 ( .A1(n5078), .A2(n5204), .ZN(n5206) );
  NAND2_X1 U6600 ( .A1(n5205), .A2(n5206), .ZN(n6818) );
  INV_X1 U6601 ( .A(n5205), .ZN(n5208) );
  INV_X1 U6602 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6603 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NAND2_X1 U6604 ( .A1(n6818), .A2(n5209), .ZN(n6713) );
  INV_X2 U6605 ( .A(n5734), .ZN(n5631) );
  INV_X1 U6606 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6607 ( .A1(n5631), .A2(n5210), .ZN(n5214) );
  NAND2_X1 U6608 ( .A1(n8046), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5212) );
  INV_X2 U6609 ( .A(n5895), .ZN(n6601) );
  NAND2_X1 U6610 ( .A1(n6601), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6611 ( .A1(n9187), .A2(n5298), .ZN(n5229) );
  NAND2_X1 U6612 ( .A1(n5217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6613 ( .A(n5218), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9895) );
  INV_X1 U6614 ( .A(n9895), .ZN(n6563) );
  NAND2_X1 U6615 ( .A1(n5221), .A2(n5220), .ZN(n5225) );
  INV_X1 U6616 ( .A(n5222), .ZN(n5223) );
  NAND2_X1 U6617 ( .A1(n5223), .A2(SI_2_), .ZN(n5224) );
  NAND2_X1 U6618 ( .A1(n5225), .A2(n5224), .ZN(n5250) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6568) );
  INV_X1 U6620 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U6621 ( .A(n6568), .B(n6564), .S(n5255), .Z(n5251) );
  XNOR2_X1 U6622 ( .A(n5251), .B(SI_3_), .ZN(n5249) );
  XNOR2_X1 U6623 ( .A(n5250), .B(n5249), .ZN(n6567) );
  OR2_X1 U6624 ( .A1(n5219), .A2(n6567), .ZN(n5227) );
  OR2_X1 U6625 ( .A1(n8161), .A2(n6564), .ZN(n5226) );
  OAI211_X1 U6626 ( .C1(n6640), .C2(n6563), .A(n5227), .B(n5226), .ZN(n6886)
         );
  NAND2_X1 U6627 ( .A1(n5814), .A2(n6886), .ZN(n5228) );
  NAND2_X1 U6628 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  INV_X2 U6629 ( .A(n5374), .ZN(n5828) );
  XNOR2_X1 U6630 ( .A(n5230), .B(n5828), .ZN(n5233) );
  NAND2_X1 U6631 ( .A1(n9187), .A2(n9049), .ZN(n5232) );
  NAND2_X1 U6632 ( .A1(n5298), .A2(n6886), .ZN(n5231) );
  AND2_X1 U6633 ( .A1(n5232), .A2(n5231), .ZN(n5234) );
  NAND2_X1 U6634 ( .A1(n5233), .A2(n5234), .ZN(n5238) );
  INV_X1 U6635 ( .A(n5233), .ZN(n5236) );
  INV_X1 U6636 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6637 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  AND2_X1 U6638 ( .A1(n5238), .A2(n5237), .ZN(n6819) );
  NAND2_X1 U6639 ( .A1(n6821), .A2(n5238), .ZN(n6861) );
  NAND2_X1 U6640 ( .A1(n5183), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6641 ( .A1(n6601), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5242) );
  INV_X1 U6642 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5239) );
  XNOR2_X1 U6643 ( .A(n5239), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7459) );
  NAND2_X1 U6644 ( .A1(n5892), .A2(n7459), .ZN(n5241) );
  NAND2_X1 U6645 ( .A1(n8046), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5240) );
  NAND4_X1 U6646 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n9186)
         );
  NAND2_X1 U6647 ( .A1(n9186), .A2(n5298), .ZN(n5259) );
  NOR2_X1 U6648 ( .A1(n5247), .A2(n5390), .ZN(n5244) );
  MUX2_X1 U6649 ( .A(n5390), .B(n5244), .S(P1_IR_REG_4__SCAN_IN), .Z(n5245) );
  INV_X1 U6650 ( .A(n5245), .ZN(n5248) );
  INV_X1 U6651 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6652 ( .A1(n5247), .A2(n5246), .ZN(n5299) );
  NAND2_X1 U6653 ( .A1(n5248), .A2(n5299), .ZN(n10086) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6561) );
  OR2_X1 U6655 ( .A1(n8161), .A2(n6561), .ZN(n5257) );
  NAND2_X1 U6656 ( .A1(n5250), .A2(n5249), .ZN(n5254) );
  INV_X1 U6657 ( .A(n5251), .ZN(n5252) );
  NAND2_X1 U6658 ( .A1(n5252), .A2(SI_3_), .ZN(n5253) );
  MUX2_X1 U6659 ( .A(n9741), .B(n6561), .S(n5255), .Z(n5277) );
  XNOR2_X1 U6660 ( .A(n5277), .B(SI_4_), .ZN(n5275) );
  XNOR2_X1 U6661 ( .A(n5276), .B(n5275), .ZN(n6562) );
  OR2_X1 U6662 ( .A1(n5219), .A2(n6562), .ZN(n5256) );
  OAI211_X1 U6663 ( .C1(n6640), .C2(n10086), .A(n5257), .B(n5256), .ZN(n7460)
         );
  NAND2_X1 U6664 ( .A1(n5814), .A2(n7460), .ZN(n5258) );
  NAND2_X1 U6665 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  XNOR2_X1 U6666 ( .A(n5260), .B(n5828), .ZN(n5265) );
  NAND2_X1 U6667 ( .A1(n9186), .A2(n9049), .ZN(n5262) );
  NAND2_X1 U6668 ( .A1(n5203), .A2(n7460), .ZN(n5261) );
  NAND2_X1 U6669 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  XNOR2_X1 U6670 ( .A(n5265), .B(n5263), .ZN(n6862) );
  NAND2_X1 U6671 ( .A1(n6861), .A2(n6862), .ZN(n6860) );
  INV_X1 U6672 ( .A(n5263), .ZN(n5264) );
  NAND2_X1 U6673 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6674 ( .A1(n6860), .A2(n5266), .ZN(n5289) );
  NAND2_X1 U6675 ( .A1(n6600), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6676 ( .A1(n6601), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5272) );
  NAND3_X1 U6677 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5292) );
  INV_X1 U6678 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6679 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5267) );
  NAND2_X1 U6680 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  AND2_X1 U6681 ( .A1(n5292), .A2(n5269), .ZN(n7140) );
  NAND2_X1 U6682 ( .A1(n5631), .A2(n7140), .ZN(n5271) );
  NAND2_X1 U6683 ( .A1(n8046), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5270) );
  NAND4_X1 U6684 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n9185)
         );
  NAND2_X1 U6685 ( .A1(n9185), .A2(n5298), .ZN(n5284) );
  NAND2_X1 U6686 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5274) );
  XNOR2_X1 U6687 ( .A(n5274), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6688) );
  INV_X1 U6688 ( .A(n6688), .ZN(n6565) );
  NAND2_X1 U6689 ( .A1(n5276), .A2(n5275), .ZN(n5280) );
  INV_X1 U6690 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6691 ( .A1(n5278), .A2(SI_4_), .ZN(n5279) );
  NAND2_X1 U6692 ( .A1(n5280), .A2(n5279), .ZN(n5302) );
  INV_X1 U6693 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6570) );
  INV_X1 U6694 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6566) );
  XNOR2_X1 U6695 ( .A(n5302), .B(n5301), .ZN(n6569) );
  OR2_X1 U6696 ( .A1(n5219), .A2(n6569), .ZN(n5282) );
  OR2_X1 U6697 ( .A1(n8161), .A2(n6566), .ZN(n5281) );
  OAI211_X1 U6698 ( .C1(n6640), .C2(n6565), .A(n5282), .B(n5281), .ZN(n7184)
         );
  NAND2_X1 U6699 ( .A1(n5814), .A2(n7184), .ZN(n5283) );
  NAND2_X1 U6700 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  XNOR2_X1 U6701 ( .A(n5285), .B(n5828), .ZN(n5288) );
  NAND2_X1 U6702 ( .A1(n9185), .A2(n9049), .ZN(n5287) );
  NAND2_X1 U6703 ( .A1(n9045), .A2(n7184), .ZN(n5286) );
  AND2_X1 U6704 ( .A1(n5287), .A2(n5286), .ZN(n7143) );
  OR2_X1 U6705 ( .A1(n5289), .A2(n5288), .ZN(n7141) );
  NAND2_X1 U6706 ( .A1(n7218), .A2(n7214), .ZN(n5317) );
  NAND2_X1 U6707 ( .A1(n6600), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6708 ( .A1(n8046), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5296) );
  INV_X1 U6709 ( .A(n5292), .ZN(n5291) );
  NAND2_X1 U6710 ( .A1(n5291), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5333) );
  INV_X1 U6711 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U6712 ( .A1(n5292), .A2(n6628), .ZN(n5293) );
  AND2_X1 U6713 ( .A1(n5333), .A2(n5293), .ZN(n7187) );
  NAND2_X1 U6714 ( .A1(n5631), .A2(n7187), .ZN(n5295) );
  NAND2_X1 U6715 ( .A1(n6601), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5294) );
  NAND4_X1 U6716 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n9184)
         );
  NAND2_X1 U6717 ( .A1(n9184), .A2(n5298), .ZN(n5308) );
  NOR2_X1 U6718 ( .A1(n5299), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5325) );
  OR2_X1 U6719 ( .A1(n5325), .A2(n5390), .ZN(n5300) );
  XNOR2_X1 U6720 ( .A(n5300), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6636) );
  AOI22_X1 U6721 ( .A1(n4841), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4458), .B2(
        n6636), .ZN(n5306) );
  NAND2_X1 U6722 ( .A1(n5303), .A2(SI_5_), .ZN(n5304) );
  MUX2_X1 U6723 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6556), .Z(n5321) );
  XNOR2_X1 U6724 ( .A(n5321), .B(SI_6_), .ZN(n5318) );
  XNOR2_X1 U6725 ( .A(n5320), .B(n5318), .ZN(n6571) );
  NAND2_X1 U6726 ( .A1(n6571), .A2(n4839), .ZN(n5305) );
  NAND2_X1 U6727 ( .A1(n5306), .A2(n5305), .ZN(n7225) );
  NAND2_X1 U6728 ( .A1(n7225), .A2(n5814), .ZN(n5307) );
  NAND2_X1 U6729 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  XNOR2_X1 U6730 ( .A(n5309), .B(n5828), .ZN(n5312) );
  NAND2_X1 U6731 ( .A1(n9184), .A2(n9049), .ZN(n5311) );
  NAND2_X1 U6732 ( .A1(n9045), .A2(n7225), .ZN(n5310) );
  AND2_X1 U6733 ( .A1(n5311), .A2(n5310), .ZN(n5313) );
  NAND2_X1 U6734 ( .A1(n5312), .A2(n5313), .ZN(n7311) );
  INV_X1 U6735 ( .A(n5312), .ZN(n5315) );
  INV_X1 U6736 ( .A(n5313), .ZN(n5314) );
  NAND2_X1 U6737 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  AND2_X1 U6738 ( .A1(n7311), .A2(n5316), .ZN(n7215) );
  NAND2_X1 U6739 ( .A1(n5317), .A2(n7215), .ZN(n7217) );
  NAND2_X1 U6740 ( .A1(n7217), .A2(n7311), .ZN(n5349) );
  INV_X1 U6741 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6742 ( .A1(n5320), .A2(n5319), .ZN(n5323) );
  NAND2_X1 U6743 ( .A1(n5321), .A2(SI_6_), .ZN(n5322) );
  NAND2_X1 U6744 ( .A1(n5323), .A2(n5322), .ZN(n5353) );
  MUX2_X1 U6745 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6556), .Z(n5354) );
  XNOR2_X1 U6746 ( .A(n5354), .B(SI_7_), .ZN(n5351) );
  XNOR2_X1 U6747 ( .A(n5353), .B(n5351), .ZN(n6575) );
  NAND2_X1 U6748 ( .A1(n6575), .A2(n8163), .ZN(n5330) );
  NAND2_X1 U6749 ( .A1(n5325), .A2(n5324), .ZN(n5386) );
  NAND2_X1 U6750 ( .A1(n5386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6751 ( .A1(n5327), .A2(n5326), .ZN(n5361) );
  OR2_X1 U6752 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  AOI22_X1 U6753 ( .A1(n4841), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4458), .B2(
        n6617), .ZN(n5329) );
  NAND2_X1 U6754 ( .A1(n5330), .A2(n5329), .ZN(n7430) );
  NAND2_X1 U6755 ( .A1(n7430), .A2(n5814), .ZN(n5340) );
  NAND2_X1 U6756 ( .A1(n5183), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6757 ( .A1(n8046), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5337) );
  INV_X1 U6758 ( .A(n5333), .ZN(n5331) );
  NAND2_X1 U6759 ( .A1(n5331), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5366) );
  INV_X1 U6760 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6761 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  AND2_X1 U6762 ( .A1(n5366), .A2(n5334), .ZN(n7429) );
  NAND2_X1 U6763 ( .A1(n5892), .A2(n7429), .ZN(n5336) );
  NAND2_X1 U6764 ( .A1(n6601), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5335) );
  NAND4_X1 U6765 ( .A1(n5338), .A2(n5337), .A3(n5336), .A4(n5335), .ZN(n9183)
         );
  NAND2_X1 U6766 ( .A1(n9183), .A2(n9045), .ZN(n5339) );
  NAND2_X1 U6767 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  XNOR2_X1 U6768 ( .A(n5341), .B(n5828), .ZN(n5344) );
  NAND2_X1 U6769 ( .A1(n7430), .A2(n9045), .ZN(n5343) );
  NAND2_X1 U6770 ( .A1(n9183), .A2(n9049), .ZN(n5342) );
  AND2_X1 U6771 ( .A1(n5343), .A2(n5342), .ZN(n5345) );
  NAND2_X1 U6772 ( .A1(n5344), .A2(n5345), .ZN(n5350) );
  INV_X1 U6773 ( .A(n5344), .ZN(n5347) );
  INV_X1 U6774 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6775 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  AND2_X1 U6776 ( .A1(n5350), .A2(n5348), .ZN(n7312) );
  INV_X1 U6777 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6778 ( .A1(n5353), .A2(n5352), .ZN(n5356) );
  NAND2_X1 U6779 ( .A1(n5354), .A2(SI_7_), .ZN(n5355) );
  MUX2_X1 U6780 ( .A(n6580), .B(n6583), .S(n6556), .Z(n5358) );
  INV_X1 U6781 ( .A(SI_8_), .ZN(n5357) );
  NAND2_X1 U6782 ( .A1(n5358), .A2(n5357), .ZN(n5381) );
  INV_X1 U6783 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6784 ( .A1(n5359), .A2(SI_8_), .ZN(n5360) );
  NAND2_X1 U6785 ( .A1(n5381), .A2(n5360), .ZN(n5379) );
  NAND2_X1 U6786 ( .A1(n6579), .A2(n8163), .ZN(n5364) );
  NAND2_X1 U6787 ( .A1(n5361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6788 ( .A(n5362), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U6789 ( .A1(n4841), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4458), .B2(
        n10100), .ZN(n5363) );
  NAND2_X1 U6790 ( .A1(n5364), .A2(n5363), .ZN(n7594) );
  NAND2_X1 U6791 ( .A1(n6600), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6792 ( .A1(n8046), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5370) );
  INV_X1 U6793 ( .A(n5366), .ZN(n5365) );
  NAND2_X1 U6794 ( .A1(n5365), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5397) );
  INV_X1 U6795 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U6796 ( .A1(n5366), .A2(n7589), .ZN(n5367) );
  AND2_X1 U6797 ( .A1(n5397), .A2(n5367), .ZN(n7562) );
  NAND2_X1 U6798 ( .A1(n5892), .A2(n7562), .ZN(n5369) );
  NAND2_X1 U6799 ( .A1(n6601), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5368) );
  NAND4_X1 U6800 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n9182)
         );
  AOI22_X1 U6801 ( .A1(n7594), .A2(n9045), .B1(n9049), .B2(n9182), .ZN(n5376)
         );
  NAND2_X1 U6802 ( .A1(n7594), .A2(n5814), .ZN(n5373) );
  NAND2_X1 U6803 ( .A1(n9182), .A2(n9045), .ZN(n5372) );
  NAND2_X1 U6804 ( .A1(n5373), .A2(n5372), .ZN(n5375) );
  XNOR2_X1 U6805 ( .A(n5375), .B(n5374), .ZN(n7588) );
  INV_X1 U6806 ( .A(n5379), .ZN(n5380) );
  MUX2_X1 U6807 ( .A(n6589), .B(n9748), .S(n6556), .Z(n5383) );
  INV_X1 U6808 ( .A(SI_9_), .ZN(n5382) );
  NAND2_X1 U6809 ( .A1(n5383), .A2(n5382), .ZN(n5415) );
  INV_X1 U6810 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6811 ( .A1(n5384), .A2(SI_9_), .ZN(n5385) );
  XNOR2_X1 U6812 ( .A(n5414), .B(n5082), .ZN(n6588) );
  NAND2_X1 U6813 ( .A1(n6588), .A2(n8163), .ZN(n5395) );
  INV_X1 U6814 ( .A(n5386), .ZN(n5388) );
  NOR2_X1 U6815 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5387) );
  AOI21_X1 U6816 ( .B1(n5388), .B2(n5387), .A(n5390), .ZN(n5389) );
  MUX2_X1 U6817 ( .A(n5390), .B(n5389), .S(P1_IR_REG_9__SCAN_IN), .Z(n5393) );
  INV_X1 U6818 ( .A(n5391), .ZN(n5392) );
  AOI22_X1 U6819 ( .A1(n4841), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4458), .B2(
        n6654), .ZN(n5394) );
  NAND2_X1 U6820 ( .A1(n10262), .A2(n5814), .ZN(n5404) );
  NAND2_X1 U6821 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  AND2_X1 U6822 ( .A1(n5424), .A2(n5398), .ZN(n7534) );
  NAND2_X1 U6823 ( .A1(n5631), .A2(n7534), .ZN(n5402) );
  NAND2_X1 U6824 ( .A1(n6600), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6825 ( .A1(n8046), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6826 ( .A1(n6601), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6827 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n9181)
         );
  NAND2_X1 U6828 ( .A1(n9181), .A2(n9045), .ZN(n5403) );
  NAND2_X1 U6829 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  XNOR2_X1 U6830 ( .A(n5405), .B(n5828), .ZN(n5407) );
  AND2_X1 U6831 ( .A1(n9049), .A2(n9181), .ZN(n5406) );
  AOI21_X1 U6832 ( .B1(n10262), .B2(n9045), .A(n5406), .ZN(n5408) );
  NAND2_X1 U6833 ( .A1(n5407), .A2(n5408), .ZN(n5413) );
  INV_X1 U6834 ( .A(n5407), .ZN(n5410) );
  INV_X1 U6835 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U6836 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  NAND2_X1 U6837 ( .A1(n5413), .A2(n5411), .ZN(n7685) );
  MUX2_X1 U6838 ( .A(n9602), .B(n6598), .S(n6556), .Z(n5418) );
  NAND2_X1 U6839 ( .A1(n5418), .A2(n5417), .ZN(n5439) );
  INV_X1 U6840 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6841 ( .A1(n5419), .A2(SI_10_), .ZN(n5420) );
  XNOR2_X1 U6842 ( .A(n5438), .B(n5080), .ZN(n6597) );
  NAND2_X1 U6843 ( .A1(n6597), .A2(n8163), .ZN(n5423) );
  NAND2_X1 U6844 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  XNOR2_X1 U6845 ( .A(n5421), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6702) );
  AOI22_X1 U6846 ( .A1(n4841), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4458), .B2(
        n6702), .ZN(n5422) );
  NAND2_X1 U6847 ( .A1(n5423), .A2(n5422), .ZN(n7679) );
  NAND2_X1 U6848 ( .A1(n7679), .A2(n5814), .ZN(n5431) );
  NAND2_X1 U6849 ( .A1(n6601), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6850 ( .A1(n6600), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6851 ( .A1(n5424), .A2(n6663), .ZN(n5425) );
  AND2_X1 U6852 ( .A1(n5471), .A2(n5425), .ZN(n7673) );
  NAND2_X1 U6853 ( .A1(n5631), .A2(n7673), .ZN(n5427) );
  NAND2_X1 U6854 ( .A1(n8046), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5426) );
  NAND4_X1 U6855 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9180)
         );
  NAND2_X1 U6856 ( .A1(n9180), .A2(n9045), .ZN(n5430) );
  NAND2_X1 U6857 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  XNOR2_X1 U6858 ( .A(n5432), .B(n5828), .ZN(n5437) );
  INV_X1 U6859 ( .A(n5437), .ZN(n5435) );
  AND2_X1 U6860 ( .A1(n9049), .A2(n9180), .ZN(n5433) );
  AOI21_X1 U6861 ( .B1(n7679), .B2(n9045), .A(n5433), .ZN(n5436) );
  INV_X1 U6862 ( .A(n5436), .ZN(n5434) );
  NAND2_X1 U6863 ( .A1(n5435), .A2(n5434), .ZN(n7671) );
  MUX2_X1 U6864 ( .A(n6609), .B(n5440), .S(n6556), .Z(n5456) );
  XNOR2_X1 U6865 ( .A(n5456), .B(SI_11_), .ZN(n5455) );
  NAND2_X1 U6866 ( .A1(n6595), .A2(n8163), .ZN(n5443) );
  OR2_X1 U6867 ( .A1(n5109), .A2(n5390), .ZN(n5441) );
  XNOR2_X1 U6868 ( .A(n5441), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U6869 ( .A1(n4841), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4458), .B2(
        n6765), .ZN(n5442) );
  NAND2_X1 U6870 ( .A1(n7710), .A2(n5814), .ZN(n5449) );
  NAND2_X1 U6871 ( .A1(n6601), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6872 ( .A1(n6600), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6873 ( .A(n5471), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U6874 ( .A1(n5631), .A2(n7778), .ZN(n5445) );
  NAND2_X1 U6875 ( .A1(n8046), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5444) );
  NAND4_X1 U6876 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n9179)
         );
  NAND2_X1 U6877 ( .A1(n9179), .A2(n9045), .ZN(n5448) );
  NAND2_X1 U6878 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XNOR2_X1 U6879 ( .A(n5450), .B(n5374), .ZN(n5454) );
  AND2_X1 U6880 ( .A1(n9049), .A2(n9179), .ZN(n5451) );
  AOI21_X1 U6881 ( .B1(n7710), .B2(n9045), .A(n5451), .ZN(n5452) );
  XNOR2_X1 U6882 ( .A(n5454), .B(n5452), .ZN(n7773) );
  INV_X1 U6883 ( .A(n5452), .ZN(n5453) );
  INV_X1 U6884 ( .A(n5455), .ZN(n5458) );
  INV_X1 U6885 ( .A(n5456), .ZN(n5457) );
  MUX2_X1 U6886 ( .A(n6622), .B(n6624), .S(n6556), .Z(n5461) );
  NAND2_X1 U6887 ( .A1(n5461), .A2(n5460), .ZN(n5484) );
  INV_X1 U6888 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U6889 ( .A1(n5462), .A2(SI_12_), .ZN(n5463) );
  NAND2_X1 U6890 ( .A1(n5484), .A2(n5463), .ZN(n5485) );
  XNOR2_X1 U6891 ( .A(n5486), .B(n5485), .ZN(n6621) );
  NAND2_X1 U6892 ( .A1(n6621), .A2(n8163), .ZN(n5466) );
  NAND2_X1 U6893 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5493) );
  XNOR2_X1 U6894 ( .A(n5493), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U6895 ( .A1(n4841), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4458), .B2(
        n6774), .ZN(n5465) );
  NAND2_X1 U6896 ( .A1(n7894), .A2(n5814), .ZN(n5478) );
  NAND2_X1 U6897 ( .A1(n6600), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6898 ( .A1(n6601), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5475) );
  INV_X1 U6899 ( .A(n5471), .ZN(n5468) );
  NAND2_X1 U6900 ( .A1(n5468), .A2(n5467), .ZN(n5499) );
  INV_X1 U6901 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5470) );
  INV_X1 U6902 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5469) );
  OAI21_X1 U6903 ( .B1(n5471), .B2(n5470), .A(n5469), .ZN(n5472) );
  AND2_X1 U6904 ( .A1(n5499), .A2(n5472), .ZN(n7893) );
  NAND2_X1 U6905 ( .A1(n5631), .A2(n7893), .ZN(n5474) );
  NAND2_X1 U6906 ( .A1(n8046), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5473) );
  NAND4_X1 U6907 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n9178)
         );
  NAND2_X1 U6908 ( .A1(n9178), .A2(n9045), .ZN(n5477) );
  NAND2_X1 U6909 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  XNOR2_X1 U6910 ( .A(n5479), .B(n5828), .ZN(n5482) );
  AND2_X1 U6911 ( .A1(n9049), .A2(n9178), .ZN(n5480) );
  AOI21_X1 U6912 ( .B1(n7894), .B2(n9045), .A(n5480), .ZN(n5481) );
  XNOR2_X1 U6913 ( .A(n5482), .B(n5481), .ZN(n7888) );
  NAND2_X1 U6914 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  OAI21_X1 U6915 ( .B1(n5486), .B2(n5485), .A(n5484), .ZN(n5510) );
  MUX2_X1 U6916 ( .A(n6718), .B(n5487), .S(n6556), .Z(n5489) );
  NAND2_X1 U6917 ( .A1(n5489), .A2(n5488), .ZN(n5511) );
  INV_X1 U6918 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U6919 ( .A1(n5490), .A2(SI_13_), .ZN(n5491) );
  XNOR2_X1 U6920 ( .A(n5510), .B(n5071), .ZN(n6709) );
  NAND2_X1 U6921 ( .A1(n6709), .A2(n8163), .ZN(n5497) );
  INV_X1 U6922 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6923 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  NAND2_X1 U6924 ( .A1(n5494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U6925 ( .A(n5495), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U6926 ( .A1(n4841), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4458), .B2(
        n10120), .ZN(n5496) );
  NAND2_X1 U6927 ( .A1(n7907), .A2(n5814), .ZN(n5506) );
  NAND2_X1 U6928 ( .A1(n6600), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U6929 ( .A1(n6601), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5503) );
  INV_X1 U6930 ( .A(n5499), .ZN(n5498) );
  NAND2_X1 U6931 ( .A1(n5498), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5521) );
  INV_X1 U6932 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U6933 ( .A1(n5499), .A2(n9728), .ZN(n5500) );
  AND2_X1 U6934 ( .A1(n5521), .A2(n5500), .ZN(n7902) );
  NAND2_X1 U6935 ( .A1(n5892), .A2(n7902), .ZN(n5502) );
  NAND2_X1 U6936 ( .A1(n8046), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5501) );
  NAND4_X1 U6937 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n9177)
         );
  NAND2_X1 U6938 ( .A1(n9177), .A2(n9045), .ZN(n5505) );
  NAND2_X1 U6939 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  XNOR2_X1 U6940 ( .A(n5507), .B(n5828), .ZN(n7900) );
  AND2_X1 U6941 ( .A1(n9049), .A2(n9177), .ZN(n5508) );
  AOI21_X1 U6942 ( .B1(n7907), .B2(n9045), .A(n5508), .ZN(n7899) );
  AND2_X1 U6943 ( .A1(n7900), .A2(n7899), .ZN(n5509) );
  NAND2_X1 U6944 ( .A1(n5510), .A2(n5071), .ZN(n5512) );
  MUX2_X1 U6945 ( .A(n6722), .B(n6720), .S(n6556), .Z(n5537) );
  XNOR2_X1 U6946 ( .A(n5537), .B(SI_14_), .ZN(n5536) );
  XNOR2_X1 U6947 ( .A(n5541), .B(n5536), .ZN(n6719) );
  NAND2_X1 U6948 ( .A1(n6719), .A2(n8163), .ZN(n5519) );
  NAND2_X1 U6949 ( .A1(n5513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5515) );
  MUX2_X1 U6950 ( .A(n5515), .B(P1_IR_REG_31__SCAN_IN), .S(n5514), .Z(n5517)
         );
  NAND2_X1 U6951 ( .A1(n5517), .A2(n5516), .ZN(n9210) );
  INV_X1 U6952 ( .A(n9210), .ZN(n10132) );
  AOI22_X1 U6953 ( .A1(n4841), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4458), .B2(
        n10132), .ZN(n5518) );
  NAND2_X1 U6954 ( .A1(n7941), .A2(n5814), .ZN(n5528) );
  NAND2_X1 U6955 ( .A1(n6601), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6956 ( .A1(n6600), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6957 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  AND2_X1 U6958 ( .A1(n5551), .A2(n5522), .ZN(n7936) );
  NAND2_X1 U6959 ( .A1(n5631), .A2(n7936), .ZN(n5524) );
  NAND2_X1 U6960 ( .A1(n8046), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5523) );
  NAND4_X1 U6961 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n9176)
         );
  NAND2_X1 U6962 ( .A1(n9176), .A2(n9045), .ZN(n5527) );
  NAND2_X1 U6963 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U6964 ( .A(n5529), .B(n5828), .ZN(n7933) );
  AND2_X1 U6965 ( .A1(n9049), .A2(n9176), .ZN(n5530) );
  AOI21_X1 U6966 ( .B1(n7941), .B2(n9045), .A(n5530), .ZN(n5532) );
  NAND2_X1 U6967 ( .A1(n7933), .A2(n5532), .ZN(n5531) );
  NAND2_X1 U6968 ( .A1(n7935), .A2(n5531), .ZN(n5535) );
  INV_X1 U6969 ( .A(n7933), .ZN(n5533) );
  INV_X1 U6970 ( .A(n5532), .ZN(n7932) );
  NAND2_X1 U6971 ( .A1(n5533), .A2(n7932), .ZN(n5534) );
  NAND2_X1 U6972 ( .A1(n5535), .A2(n5534), .ZN(n9158) );
  INV_X1 U6973 ( .A(n5536), .ZN(n5540) );
  INV_X1 U6974 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U6975 ( .A1(n5538), .A2(SI_14_), .ZN(n5539) );
  MUX2_X1 U6976 ( .A(n6925), .B(n9637), .S(n6556), .Z(n5543) );
  NAND2_X1 U6977 ( .A1(n5543), .A2(n5542), .ZN(n5565) );
  INV_X1 U6978 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U6979 ( .A1(n5544), .A2(SI_15_), .ZN(n5545) );
  NAND2_X1 U6980 ( .A1(n5565), .A2(n5545), .ZN(n5566) );
  XNOR2_X1 U6981 ( .A(n5567), .B(n5566), .ZN(n6924) );
  NAND2_X1 U6982 ( .A1(n6924), .A2(n8163), .ZN(n5548) );
  NAND2_X1 U6983 ( .A1(n5516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5546) );
  XNOR2_X1 U6984 ( .A(n5546), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U6985 ( .A1(n4841), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4458), .B2(
        n10146), .ZN(n5547) );
  NAND2_X1 U6986 ( .A1(n9169), .A2(n5814), .ZN(n5558) );
  NAND2_X1 U6987 ( .A1(n6601), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6988 ( .A1(n6600), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5555) );
  INV_X1 U6989 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6990 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  AND2_X1 U6991 ( .A1(n5602), .A2(n5552), .ZN(n9167) );
  NAND2_X1 U6992 ( .A1(n5892), .A2(n9167), .ZN(n5554) );
  NAND2_X1 U6993 ( .A1(n8046), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5553) );
  NAND4_X1 U6994 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n9987)
         );
  NAND2_X1 U6995 ( .A1(n9987), .A2(n9045), .ZN(n5557) );
  NAND2_X1 U6996 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  XNOR2_X1 U6997 ( .A(n5559), .B(n5828), .ZN(n9160) );
  AND2_X1 U6998 ( .A1(n9049), .A2(n9987), .ZN(n5560) );
  AOI21_X1 U6999 ( .B1(n9169), .B2(n9045), .A(n5560), .ZN(n5562) );
  NAND2_X1 U7000 ( .A1(n9160), .A2(n5562), .ZN(n5561) );
  INV_X1 U7001 ( .A(n9160), .ZN(n5563) );
  INV_X1 U7002 ( .A(n5562), .ZN(n9159) );
  NAND2_X1 U7003 ( .A1(n5563), .A2(n9159), .ZN(n5564) );
  MUX2_X1 U7004 ( .A(n9781), .B(n9753), .S(n6556), .Z(n5569) );
  NAND2_X1 U7005 ( .A1(n5569), .A2(n5568), .ZN(n5591) );
  INV_X1 U7006 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7007 ( .A1(n5570), .A2(SI_16_), .ZN(n5571) );
  XNOR2_X1 U7008 ( .A(n5590), .B(n5589), .ZN(n6940) );
  NAND2_X1 U7009 ( .A1(n6940), .A2(n8163), .ZN(n5574) );
  NAND2_X1 U7010 ( .A1(n5572), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5596) );
  XNOR2_X1 U7011 ( .A(n5596), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U7012 ( .A1(n4841), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4458), .B2(
        n10157), .ZN(n5573) );
  NAND2_X1 U7013 ( .A1(n10009), .A2(n5814), .ZN(n5580) );
  NAND2_X1 U7014 ( .A1(n6600), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7015 ( .A1(n6601), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5577) );
  XNOR2_X1 U7016 ( .A(n5602), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U7017 ( .A1(n5892), .A2(n9994), .ZN(n5576) );
  NAND2_X1 U7018 ( .A1(n8046), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5575) );
  NAND4_X1 U7019 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n9175)
         );
  NAND2_X1 U7020 ( .A1(n9175), .A2(n9045), .ZN(n5579) );
  NAND2_X1 U7021 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  XNOR2_X1 U7022 ( .A(n5581), .B(n5828), .ZN(n5583) );
  AND2_X1 U7023 ( .A1(n9049), .A2(n9175), .ZN(n5582) );
  AOI21_X1 U7024 ( .B1(n10009), .B2(n9045), .A(n5582), .ZN(n5584) );
  NAND2_X1 U7025 ( .A1(n5583), .A2(n5584), .ZN(n5588) );
  INV_X1 U7026 ( .A(n5583), .ZN(n5586) );
  INV_X1 U7027 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7028 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7029 ( .A1(n5588), .A2(n5587), .ZN(n9085) );
  MUX2_X1 U7030 ( .A(n5594), .B(n5593), .S(n6556), .Z(n5617) );
  XNOR2_X1 U7031 ( .A(n5617), .B(SI_17_), .ZN(n5616) );
  XNOR2_X1 U7032 ( .A(n5621), .B(n5616), .ZN(n6988) );
  NAND2_X1 U7033 ( .A1(n6988), .A2(n8163), .ZN(n5599) );
  NAND2_X1 U7034 ( .A1(n5596), .A2(n5595), .ZN(n5597) );
  NAND2_X1 U7035 ( .A1(n5597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5623) );
  XNOR2_X1 U7036 ( .A(n5623), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U7037 ( .A1(n4841), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4458), .B2(
        n10170), .ZN(n5598) );
  NAND2_X1 U7038 ( .A1(n9510), .A2(n5814), .ZN(n5609) );
  NAND2_X1 U7039 ( .A1(n6601), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7040 ( .A1(n6600), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5606) );
  INV_X1 U7041 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9086) );
  INV_X1 U7042 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U7043 ( .B1(n5602), .B2(n9086), .A(n5600), .ZN(n5603) );
  NAND2_X1 U7044 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5601) );
  AND2_X1 U7045 ( .A1(n5603), .A2(n5629), .ZN(n9429) );
  NAND2_X1 U7046 ( .A1(n5631), .A2(n9429), .ZN(n5605) );
  NAND2_X1 U7047 ( .A1(n8046), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5604) );
  NAND4_X1 U7048 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n9989)
         );
  NAND2_X1 U7049 ( .A1(n9989), .A2(n9045), .ZN(n5608) );
  NAND2_X1 U7050 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  XNOR2_X1 U7051 ( .A(n5610), .B(n5374), .ZN(n5612) );
  AND2_X1 U7052 ( .A1(n9049), .A2(n9989), .ZN(n5611) );
  AOI21_X1 U7053 ( .B1(n9510), .B2(n9045), .A(n5611), .ZN(n5613) );
  XNOR2_X1 U7054 ( .A(n5612), .B(n5613), .ZN(n9094) );
  INV_X1 U7055 ( .A(n5612), .ZN(n5614) );
  NAND2_X1 U7056 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U7057 ( .A1(n9092), .A2(n5615), .ZN(n5685) );
  INV_X1 U7058 ( .A(n5616), .ZN(n5620) );
  INV_X1 U7059 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7060 ( .A1(n5618), .A2(SI_17_), .ZN(n5619) );
  MUX2_X1 U7061 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6556), .Z(n5644) );
  XNOR2_X1 U7062 ( .A(n5644), .B(SI_18_), .ZN(n5641) );
  XNOR2_X1 U7063 ( .A(n5643), .B(n5641), .ZN(n7308) );
  NAND2_X1 U7064 ( .A1(n7308), .A2(n8163), .ZN(n5627) );
  NAND2_X1 U7065 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  NAND2_X1 U7066 ( .A1(n5624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  XNOR2_X1 U7067 ( .A(n5625), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U7068 ( .A1(n4841), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10185), 
        .B2(n4458), .ZN(n5626) );
  NAND2_X1 U7069 ( .A1(n9503), .A2(n5814), .ZN(n5637) );
  NAND2_X1 U7070 ( .A1(n6601), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7071 ( .A1(n6600), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5634) );
  INV_X1 U7072 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U7073 ( .A1(n5629), .A2(n9824), .ZN(n5630) );
  AND2_X1 U7074 ( .A1(n5652), .A2(n5630), .ZN(n9405) );
  NAND2_X1 U7075 ( .A1(n5631), .A2(n9405), .ZN(n5633) );
  NAND2_X1 U7076 ( .A1(n8046), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5632) );
  NAND4_X1 U7077 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n9395)
         );
  NAND2_X1 U7078 ( .A1(n9395), .A2(n9045), .ZN(n5636) );
  NAND2_X1 U7079 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  XNOR2_X1 U7080 ( .A(n5638), .B(n5828), .ZN(n5686) );
  NAND2_X1 U7081 ( .A1(n5685), .A2(n5686), .ZN(n9134) );
  NAND2_X1 U7082 ( .A1(n9503), .A2(n9045), .ZN(n5640) );
  NAND2_X1 U7083 ( .A1(n9395), .A2(n9049), .ZN(n5639) );
  NAND2_X1 U7084 ( .A1(n5640), .A2(n5639), .ZN(n9137) );
  NAND2_X1 U7085 ( .A1(n9134), .A2(n9137), .ZN(n9034) );
  INV_X1 U7086 ( .A(n5641), .ZN(n5642) );
  MUX2_X1 U7087 ( .A(n8361), .B(n7362), .S(n6556), .Z(n5646) );
  NAND2_X1 U7088 ( .A1(n5646), .A2(n5645), .ZN(n5663) );
  INV_X1 U7089 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7090 ( .A1(n5647), .A2(SI_19_), .ZN(n5648) );
  NAND2_X1 U7091 ( .A1(n5663), .A2(n5648), .ZN(n5664) );
  XNOR2_X1 U7092 ( .A(n5665), .B(n5664), .ZN(n7361) );
  NAND2_X1 U7093 ( .A1(n7361), .A2(n8163), .ZN(n5650) );
  AOI22_X1 U7094 ( .A1(n4841), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9342), .B2(
        n4458), .ZN(n5649) );
  NAND2_X1 U7095 ( .A1(n9498), .A2(n5814), .ZN(n5659) );
  NAND2_X1 U7096 ( .A1(n6601), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5657) );
  INV_X1 U7097 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7098 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  AND2_X1 U7099 ( .A1(n5674), .A2(n5653), .ZN(n9391) );
  NAND2_X1 U7100 ( .A1(n9391), .A2(n5892), .ZN(n5656) );
  NAND2_X1 U7101 ( .A1(n6600), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7102 ( .A1(n8046), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5654) );
  NAND4_X1 U7103 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n9412)
         );
  NAND2_X1 U7104 ( .A1(n9412), .A2(n9045), .ZN(n5658) );
  NAND2_X1 U7105 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  XNOR2_X1 U7106 ( .A(n5660), .B(n5374), .ZN(n5693) );
  NAND2_X1 U7107 ( .A1(n9498), .A2(n9045), .ZN(n5662) );
  NAND2_X1 U7108 ( .A1(n9412), .A2(n9049), .ZN(n5661) );
  NAND2_X1 U7109 ( .A1(n5662), .A2(n5661), .ZN(n5694) );
  AND2_X1 U7110 ( .A1(n5693), .A2(n5694), .ZN(n9036) );
  MUX2_X1 U7111 ( .A(n7669), .B(n7572), .S(n6556), .Z(n5667) );
  INV_X1 U7112 ( .A(SI_20_), .ZN(n5666) );
  NAND2_X1 U7113 ( .A1(n5667), .A2(n5666), .ZN(n5702) );
  INV_X1 U7114 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U7115 ( .A1(n5668), .A2(SI_20_), .ZN(n5669) );
  XNOR2_X1 U7116 ( .A(n5701), .B(n5700), .ZN(n7571) );
  NAND2_X1 U7117 ( .A1(n7571), .A2(n8163), .ZN(n5671) );
  OR2_X1 U7118 ( .A1(n8161), .A2(n7572), .ZN(n5670) );
  NAND2_X1 U7119 ( .A1(n9493), .A2(n5814), .ZN(n5682) );
  INV_X1 U7120 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5680) );
  INV_X1 U7121 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7122 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U7123 ( .A1(n5706), .A2(n5675), .ZN(n9117) );
  OR2_X1 U7124 ( .A1(n9117), .A2(n5734), .ZN(n5679) );
  NAND2_X1 U7125 ( .A1(n6600), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7126 ( .A1(n8046), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5676) );
  AND2_X1 U7127 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  OAI211_X1 U7128 ( .C1(n5895), .C2(n5680), .A(n5679), .B(n5678), .ZN(n9396)
         );
  NAND2_X1 U7129 ( .A1(n9396), .A2(n9045), .ZN(n5681) );
  NAND2_X1 U7130 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  XNOR2_X1 U7131 ( .A(n5683), .B(n5374), .ZN(n5690) );
  AND2_X1 U7132 ( .A1(n9396), .A2(n9049), .ZN(n5684) );
  AOI21_X1 U7133 ( .B1(n9493), .B2(n9045), .A(n5684), .ZN(n5691) );
  XNOR2_X1 U7134 ( .A(n5690), .B(n5691), .ZN(n9114) );
  INV_X1 U7135 ( .A(n9114), .ZN(n5697) );
  NOR2_X1 U7136 ( .A1(n9036), .A2(n5697), .ZN(n5689) );
  INV_X1 U7137 ( .A(n5685), .ZN(n5688) );
  NAND2_X1 U7138 ( .A1(n5688), .A2(n5687), .ZN(n9135) );
  NAND3_X1 U7139 ( .A1(n9034), .A2(n5689), .A3(n9135), .ZN(n9111) );
  INV_X1 U7140 ( .A(n5690), .ZN(n5692) );
  NAND2_X1 U7141 ( .A1(n5692), .A2(n5691), .ZN(n5698) );
  INV_X1 U7142 ( .A(n5693), .ZN(n5696) );
  INV_X1 U7143 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7144 ( .A1(n5696), .A2(n5695), .ZN(n9108) );
  OR2_X1 U7145 ( .A1(n5697), .A2(n9108), .ZN(n9110) );
  AND2_X1 U7146 ( .A1(n5698), .A2(n9110), .ZN(n5699) );
  MUX2_X1 U7147 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6556), .Z(n5722) );
  XNOR2_X1 U7148 ( .A(n5722), .B(n5703), .ZN(n5721) );
  XNOR2_X1 U7149 ( .A(n5720), .B(n5721), .ZN(n7665) );
  NAND2_X1 U7150 ( .A1(n7665), .A2(n8163), .ZN(n5705) );
  INV_X1 U7151 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8383) );
  OR2_X1 U7152 ( .A1(n8161), .A2(n8383), .ZN(n5704) );
  NAND2_X1 U7153 ( .A1(n9489), .A2(n5814), .ZN(n5712) );
  INV_X1 U7154 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U7155 ( .A1(n5706), .A2(n9069), .ZN(n5707) );
  NAND2_X1 U7156 ( .A1(n5732), .A2(n5707), .ZN(n9356) );
  AOI22_X1 U7157 ( .A1(n6600), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n6601), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7158 ( .A1(n8046), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U7159 ( .C1(n9356), .C2(n5734), .A(n5710), .B(n5709), .ZN(n9381)
         );
  NAND2_X1 U7160 ( .A1(n9381), .A2(n9045), .ZN(n5711) );
  NAND2_X1 U7161 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  XNOR2_X1 U7162 ( .A(n5713), .B(n5374), .ZN(n5715) );
  AND2_X1 U7163 ( .A1(n9381), .A2(n9049), .ZN(n5714) );
  AOI21_X1 U7164 ( .B1(n9489), .B2(n9045), .A(n5714), .ZN(n5716) );
  XNOR2_X1 U7165 ( .A(n5715), .B(n5716), .ZN(n9068) );
  INV_X1 U7166 ( .A(n5715), .ZN(n5717) );
  NAND2_X1 U7167 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U7168 ( .A1(n5722), .A2(SI_21_), .ZN(n5723) );
  NAND2_X1 U7169 ( .A1(n5724), .A2(n5723), .ZN(n5745) );
  MUX2_X1 U7170 ( .A(n8068), .B(n8363), .S(n6556), .Z(n5725) );
  NAND2_X1 U7171 ( .A1(n5725), .A2(n9816), .ZN(n5743) );
  INV_X1 U7172 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U7173 ( .A1(n5726), .A2(SI_22_), .ZN(n5727) );
  NAND2_X1 U7174 ( .A1(n5743), .A2(n5727), .ZN(n5744) );
  XNOR2_X1 U7175 ( .A(n5745), .B(n5744), .ZN(n8067) );
  NAND2_X1 U7176 ( .A1(n8067), .A2(n8163), .ZN(n5729) );
  OR2_X1 U7177 ( .A1(n8161), .A2(n8363), .ZN(n5728) );
  INV_X1 U7178 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7179 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  NAND2_X1 U7180 ( .A1(n5752), .A2(n5733), .ZN(n9341) );
  OR2_X1 U7181 ( .A1(n9341), .A2(n5734), .ZN(n5739) );
  INV_X1 U7182 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U7183 ( .A1(n5184), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7184 ( .A1(n6600), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5735) );
  OAI211_X1 U7185 ( .C1(n9800), .C2(n5821), .A(n5736), .B(n5735), .ZN(n5737)
         );
  INV_X1 U7186 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7187 ( .A1(n5739), .A2(n5738), .ZN(n9365) );
  AND2_X1 U7188 ( .A1(n9365), .A2(n9049), .ZN(n5740) );
  AOI21_X1 U7189 ( .B1(n9485), .B2(n9045), .A(n5740), .ZN(n5742) );
  AOI22_X1 U7190 ( .A1(n9485), .A2(n5814), .B1(n9045), .B2(n9365), .ZN(n5741)
         );
  XOR2_X1 U7191 ( .A(n5374), .B(n5741), .Z(n9125) );
  MUX2_X1 U7192 ( .A(n7751), .B(n7746), .S(n6556), .Z(n5747) );
  INV_X1 U7193 ( .A(SI_23_), .ZN(n5746) );
  NAND2_X1 U7194 ( .A1(n5747), .A2(n5746), .ZN(n5764) );
  INV_X1 U7195 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7196 ( .A1(n5748), .A2(SI_23_), .ZN(n5749) );
  XNOR2_X1 U7197 ( .A(n5763), .B(n5762), .ZN(n7748) );
  NAND2_X1 U7198 ( .A1(n7748), .A2(n8163), .ZN(n5751) );
  OR2_X1 U7199 ( .A1(n8161), .A2(n7746), .ZN(n5750) );
  INV_X1 U7200 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U7201 ( .A1(n5752), .A2(n9028), .ZN(n5753) );
  NAND2_X1 U7202 ( .A1(n5768), .A2(n5753), .ZN(n9326) );
  OR2_X1 U7203 ( .A1(n9326), .A2(n5734), .ZN(n5759) );
  INV_X1 U7204 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7205 ( .A1(n6600), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7206 ( .A1(n5184), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U7207 ( .C1(n5756), .C2(n5821), .A(n5755), .B(n5754), .ZN(n5757)
         );
  INV_X1 U7208 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7209 ( .A1(n5759), .A2(n5758), .ZN(n9305) );
  AOI22_X1 U7210 ( .A1(n9480), .A2(n5814), .B1(n9045), .B2(n9305), .ZN(n5760)
         );
  XOR2_X1 U7211 ( .A(n5374), .B(n5760), .Z(n5761) );
  NOR2_X1 U7212 ( .A1(n9124), .A2(n5761), .ZN(n9023) );
  AOI22_X1 U7213 ( .A1(n9480), .A2(n9045), .B1(n9049), .B2(n9305), .ZN(n9026)
         );
  NAND2_X1 U7214 ( .A1(n9124), .A2(n5761), .ZN(n9024) );
  MUX2_X1 U7215 ( .A(n7824), .B(n7826), .S(n6556), .Z(n5782) );
  XNOR2_X1 U7216 ( .A(n5782), .B(SI_24_), .ZN(n5781) );
  NAND2_X1 U7217 ( .A1(n7823), .A2(n8163), .ZN(n5766) );
  OR2_X1 U7218 ( .A1(n8161), .A2(n7826), .ZN(n5765) );
  INV_X1 U7219 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7220 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  AND2_X1 U7221 ( .A1(n5791), .A2(n5769), .ZN(n9311) );
  NAND2_X1 U7222 ( .A1(n9311), .A2(n5892), .ZN(n5775) );
  INV_X1 U7223 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7224 ( .A1(n5184), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7225 ( .A1(n6600), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5770) );
  OAI211_X1 U7226 ( .C1(n5772), .C2(n5821), .A(n5771), .B(n5770), .ZN(n5773)
         );
  INV_X1 U7227 ( .A(n5773), .ZN(n5774) );
  NAND2_X1 U7228 ( .A1(n5775), .A2(n5774), .ZN(n9290) );
  AOI22_X1 U7229 ( .A1(n9471), .A2(n5814), .B1(n9045), .B2(n9290), .ZN(n5776)
         );
  XNOR2_X1 U7230 ( .A(n5776), .B(n5374), .ZN(n5778) );
  AOI22_X1 U7231 ( .A1(n9471), .A2(n9045), .B1(n9049), .B2(n9290), .ZN(n5777)
         );
  XNOR2_X1 U7232 ( .A(n5778), .B(n5777), .ZN(n9101) );
  INV_X1 U7233 ( .A(n5777), .ZN(n5780) );
  INV_X1 U7234 ( .A(n5778), .ZN(n5779) );
  INV_X1 U7235 ( .A(n5782), .ZN(n5783) );
  MUX2_X1 U7236 ( .A(n7931), .B(n7928), .S(n6556), .Z(n5784) );
  INV_X1 U7237 ( .A(SI_25_), .ZN(n9662) );
  NAND2_X1 U7238 ( .A1(n5784), .A2(n9662), .ZN(n5805) );
  INV_X1 U7239 ( .A(n5784), .ZN(n5785) );
  NAND2_X1 U7240 ( .A1(n5785), .A2(SI_25_), .ZN(n5786) );
  NAND2_X1 U7241 ( .A1(n5805), .A2(n5786), .ZN(n5806) );
  XNOR2_X1 U7242 ( .A(n5807), .B(n5806), .ZN(n7926) );
  NAND2_X1 U7243 ( .A1(n7926), .A2(n8163), .ZN(n5788) );
  OR2_X1 U7244 ( .A1(n8161), .A2(n7928), .ZN(n5787) );
  NAND2_X1 U7245 ( .A1(n9465), .A2(n5814), .ZN(n5800) );
  INV_X1 U7246 ( .A(n5791), .ZN(n5789) );
  NAND2_X1 U7247 ( .A1(n5789), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5817) );
  INV_X1 U7248 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7249 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U7250 ( .A1(n5817), .A2(n5792), .ZN(n9284) );
  INV_X1 U7251 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7252 ( .A1(n5184), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7253 ( .A1(n6600), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5793) );
  OAI211_X1 U7254 ( .C1(n5795), .C2(n5821), .A(n5794), .B(n5793), .ZN(n5796)
         );
  INV_X1 U7255 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U7256 ( .A1(n9306), .A2(n9045), .ZN(n5799) );
  NAND2_X1 U7257 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  XNOR2_X1 U7258 ( .A(n5801), .B(n5374), .ZN(n5802) );
  AOI22_X1 U7259 ( .A1(n9465), .A2(n9045), .B1(n9049), .B2(n9306), .ZN(n5803)
         );
  XNOR2_X1 U7260 ( .A(n5802), .B(n5803), .ZN(n9076) );
  INV_X1 U7261 ( .A(n5802), .ZN(n5804) );
  INV_X1 U7262 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7947) );
  MUX2_X1 U7263 ( .A(n7947), .B(n9658), .S(n6556), .Z(n5809) );
  INV_X1 U7264 ( .A(SI_26_), .ZN(n5808) );
  NAND2_X1 U7265 ( .A1(n5809), .A2(n5808), .ZN(n5835) );
  INV_X1 U7266 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U7267 ( .A1(n5810), .A2(SI_26_), .ZN(n5811) );
  XNOR2_X1 U7268 ( .A(n5834), .B(n5833), .ZN(n7945) );
  NAND2_X1 U7269 ( .A1(n7945), .A2(n8163), .ZN(n5813) );
  OR2_X1 U7270 ( .A1(n8161), .A2(n9658), .ZN(n5812) );
  NAND2_X1 U7271 ( .A1(n9460), .A2(n5814), .ZN(n5827) );
  INV_X1 U7272 ( .A(n5817), .ZN(n5815) );
  INV_X1 U7273 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7274 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U7275 ( .A1(n5890), .A2(n5818), .ZN(n9267) );
  OR2_X1 U7276 ( .A1(n9267), .A2(n5734), .ZN(n5825) );
  INV_X1 U7277 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7278 ( .A1(n6600), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7279 ( .A1(n6601), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5819) );
  OAI211_X1 U7280 ( .C1(n5822), .C2(n5821), .A(n5820), .B(n5819), .ZN(n5823)
         );
  INV_X1 U7281 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7282 ( .A1(n9291), .A2(n9045), .ZN(n5826) );
  NAND2_X1 U7283 ( .A1(n5827), .A2(n5826), .ZN(n5829) );
  XNOR2_X1 U7284 ( .A(n5829), .B(n5828), .ZN(n5832) );
  AND2_X1 U7285 ( .A1(n9291), .A2(n9049), .ZN(n5830) );
  AOI21_X1 U7286 ( .B1(n9460), .B2(n9045), .A(n5830), .ZN(n5831) );
  NOR2_X1 U7287 ( .A1(n5832), .A2(n5831), .ZN(n9148) );
  NAND2_X1 U7288 ( .A1(n5832), .A2(n5831), .ZN(n9146) );
  NAND2_X1 U7289 ( .A1(n5834), .A2(n5833), .ZN(n5836) );
  INV_X1 U7290 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7953) );
  MUX2_X1 U7291 ( .A(n7956), .B(n7953), .S(n6556), .Z(n5838) );
  INV_X1 U7292 ( .A(SI_27_), .ZN(n5837) );
  NAND2_X1 U7293 ( .A1(n5838), .A2(n5837), .ZN(n6250) );
  INV_X1 U7294 ( .A(n5838), .ZN(n5839) );
  NAND2_X1 U7295 ( .A1(n5839), .A2(SI_27_), .ZN(n5840) );
  NAND2_X1 U7296 ( .A1(n7954), .A2(n8163), .ZN(n5842) );
  OR2_X1 U7297 ( .A1(n8161), .A2(n7953), .ZN(n5841) );
  XNOR2_X1 U7298 ( .A(n5890), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9251) );
  INV_X1 U7299 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7300 ( .A1(n8046), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7301 ( .A1(n6601), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5843) );
  OAI211_X1 U7302 ( .C1(n5846), .C2(n5845), .A(n5844), .B(n5843), .ZN(n5847)
         );
  AOI21_X1 U7303 ( .B1(n9251), .B2(n5892), .A(n5847), .ZN(n9151) );
  OAI22_X1 U7304 ( .A1(n9253), .A2(n5848), .B1(n9151), .B2(n5850), .ZN(n5849)
         );
  XNOR2_X1 U7305 ( .A(n5849), .B(n5374), .ZN(n5852) );
  OAI22_X1 U7306 ( .A1(n9253), .A2(n5850), .B1(n9151), .B2(n5175), .ZN(n5851)
         );
  NOR2_X1 U7307 ( .A1(n5852), .A2(n5851), .ZN(n9061) );
  AOI21_X1 U7308 ( .B1(n5852), .B2(n5851), .A(n9061), .ZN(n5854) );
  NAND2_X1 U7309 ( .A1(n5853), .A2(n5854), .ZN(n9060) );
  INV_X1 U7310 ( .A(n5853), .ZN(n5856) );
  INV_X1 U7311 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U7312 ( .A1(n5856), .A2(n5855), .ZN(n5857) );
  NAND2_X1 U7313 ( .A1(n9060), .A2(n5857), .ZN(n5881) );
  NAND2_X1 U7314 ( .A1(n5858), .A2(n5859), .ZN(n7044) );
  NAND2_X1 U7315 ( .A1(n7927), .A2(P1_B_REG_SCAN_IN), .ZN(n5860) );
  MUX2_X1 U7316 ( .A(P1_B_REG_SCAN_IN), .B(n5860), .S(n7828), .Z(n5861) );
  NAND2_X1 U7317 ( .A1(n5861), .A2(n7944), .ZN(n10222) );
  INV_X1 U7318 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5864) );
  INV_X1 U7319 ( .A(n7828), .ZN(n5862) );
  NOR2_X1 U7320 ( .A1(n7944), .A2(n5862), .ZN(n5863) );
  INV_X1 U7321 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10233) );
  INV_X1 U7322 ( .A(n7927), .ZN(n5865) );
  NOR2_X1 U7323 ( .A1(n7944), .A2(n5865), .ZN(n5866) );
  AOI21_X1 U7324 ( .B1(n5877), .B2(n10233), .A(n5866), .ZN(n7039) );
  NOR4_X1 U7325 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5875) );
  NOR4_X1 U7326 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5874) );
  INV_X1 U7327 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10228) );
  INV_X1 U7328 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10225) );
  INV_X1 U7329 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10229) );
  INV_X1 U7330 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U7331 ( .A1(n10228), .A2(n10225), .A3(n10229), .A4(n10224), .ZN(
        n5872) );
  NOR4_X1 U7332 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5870) );
  NOR4_X1 U7333 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5869) );
  NOR4_X1 U7334 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n5868) );
  NOR4_X1 U7335 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5867) );
  NAND4_X1 U7336 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n5871)
         );
  NOR4_X1 U7337 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5872), .A4(n5871), .ZN(n5873) );
  NAND3_X1 U7338 ( .A1(n5875), .A2(n5874), .A3(n5873), .ZN(n5876) );
  NAND2_X1 U7339 ( .A1(n5877), .A2(n5876), .ZN(n6851) );
  AND3_X1 U7340 ( .A1(n9881), .A2(n7039), .A3(n6851), .ZN(n6676) );
  NAND2_X1 U7341 ( .A1(n5878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7342 ( .A1(n5881), .A2(n9115), .ZN(n5914) );
  NAND2_X1 U7343 ( .A1(n7352), .A2(n5884), .ZN(n5883) );
  NAND2_X1 U7344 ( .A1(n5859), .A2(n10234), .ZN(n5882) );
  OR2_X1 U7345 ( .A1(n7051), .A2(n6833), .ZN(n8350) );
  INV_X1 U7346 ( .A(n5884), .ZN(n5885) );
  NOR2_X1 U7347 ( .A1(n8350), .A2(n5885), .ZN(n5907) );
  INV_X1 U7348 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5888) );
  INV_X1 U7349 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5887) );
  OAI21_X1 U7350 ( .B1(n5890), .B2(n5888), .A(n5887), .ZN(n5891) );
  NAND2_X1 U7351 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5889) );
  NAND2_X1 U7352 ( .A1(n9239), .A2(n5892), .ZN(n5898) );
  INV_X1 U7353 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U7354 ( .A1(n6600), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7355 ( .A1(n8046), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5893) );
  OAI211_X1 U7356 ( .C1(n9793), .C2(n5895), .A(n5894), .B(n5893), .ZN(n5896)
         );
  INV_X1 U7357 ( .A(n5896), .ZN(n5897) );
  INV_X1 U7358 ( .A(n5899), .ZN(n5901) );
  AND3_X1 U7359 ( .A1(n7042), .A2(n6514), .A3(n7744), .ZN(n5900) );
  OAI21_X1 U7360 ( .B1(n5901), .B2(n6676), .A(n5900), .ZN(n5902) );
  NAND2_X1 U7361 ( .A1(n5902), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7362 ( .A1(n8350), .A2(n10196), .ZN(n5905) );
  INV_X1 U7363 ( .A(n6676), .ZN(n5903) );
  AND2_X1 U7364 ( .A1(n5903), .A2(n10234), .ZN(n5904) );
  NAND2_X1 U7365 ( .A1(n5905), .A2(n5904), .ZN(n6674) );
  INV_X1 U7366 ( .A(n9251), .ZN(n5909) );
  AOI22_X1 U7367 ( .A1(n9291), .A2(n9162), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n5908) );
  OAI21_X1 U7368 ( .B1(n9153), .B2(n5909), .A(n5908), .ZN(n5910) );
  AOI21_X1 U7369 ( .B1(n9138), .B2(n9257), .A(n5910), .ZN(n5911) );
  INV_X1 U7370 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7371 ( .A1(n5914), .A2(n5913), .ZN(P1_U3212) );
  NOR2_X1 U7372 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5917) );
  NOR2_X1 U7373 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5916) );
  NOR2_X1 U7374 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5915) );
  NOR2_X1 U7375 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5918) );
  NAND2_X1 U7376 ( .A1(n6123), .A2(n5918), .ZN(n5919) );
  INV_X1 U7377 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6898) );
  NAND2_X2 U7378 ( .A1(n5926), .A2(n5925), .ZN(n5968) );
  INV_X1 U7379 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9912) );
  OR2_X1 U7380 ( .A1(n4463), .A2(n9912), .ZN(n5930) );
  NAND2_X1 U7381 ( .A1(n4464), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5929) );
  XNOR2_X2 U7382 ( .A(n5934), .B(n5933), .ZN(n6508) );
  NAND2_X1 U7383 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5936) );
  MUX2_X1 U7384 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5936), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5938) );
  INV_X1 U7385 ( .A(n5956), .ZN(n5937) );
  NAND2_X1 U7386 ( .A1(n5938), .A2(n5937), .ZN(n9917) );
  INV_X1 U7387 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7388 ( .A1(n7023), .A2(n6815), .ZN(n6470) );
  INV_X1 U7389 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7289) );
  INV_X1 U7390 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5939) );
  INV_X1 U7391 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10359) );
  INV_X1 U7392 ( .A(n6317), .ZN(n5946) );
  INV_X1 U7393 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U7394 ( .A1(n6555), .A2(SI_0_), .ZN(n5945) );
  INV_X1 U7395 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5944) );
  XNOR2_X1 U7396 ( .A(n5945), .B(n5944), .ZN(n9021) );
  MUX2_X1 U7397 ( .A(n10290), .B(n9021), .S(n6902), .Z(n7443) );
  INV_X1 U7398 ( .A(n7443), .ZN(n10307) );
  NAND2_X1 U7399 ( .A1(n6470), .A2(n6468), .ZN(n5947) );
  NAND2_X1 U7400 ( .A1(n6786), .A2(n6741), .ZN(n6469) );
  NAND2_X1 U7401 ( .A1(n5947), .A2(n6469), .ZN(n6320) );
  INV_X1 U7402 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9734) );
  AND2_X1 U7403 ( .A1(n5950), .A2(n5949), .ZN(n5955) );
  INV_X1 U7404 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5951) );
  INV_X2 U7405 ( .A(n5968), .ZN(n5952) );
  OR2_X1 U7406 ( .A1(n5956), .A2(n6156), .ZN(n5958) );
  INV_X1 U7407 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5957) );
  XNOR2_X1 U7408 ( .A(n5958), .B(n5957), .ZN(n6912) );
  NAND2_X1 U7409 ( .A1(n6756), .A2(n4457), .ZN(n6322) );
  OR2_X1 U7410 ( .A1(n4465), .A2(n9010), .ZN(n5961) );
  OR2_X1 U7411 ( .A1(n5968), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5960) );
  INV_X1 U7412 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6897) );
  OR2_X1 U7413 ( .A1(n5969), .A2(n6897), .ZN(n5959) );
  INV_X1 U7414 ( .A(n6946), .ZN(n6927) );
  OR2_X1 U7415 ( .A1(n5976), .A2(n6568), .ZN(n5965) );
  OR2_X1 U7416 ( .A1(n5975), .A2(n6567), .ZN(n5964) );
  NAND2_X1 U7417 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4493), .ZN(n5963) );
  XNOR2_X1 U7418 ( .A(n5963), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6913) );
  INV_X1 U7419 ( .A(n6913), .ZN(n7096) );
  NAND2_X1 U7420 ( .A1(n6927), .A2(n6947), .ZN(n6330) );
  NAND2_X1 U7421 ( .A1(n6752), .A2(n6753), .ZN(n5966) );
  NAND2_X1 U7422 ( .A1(n5966), .A2(n6330), .ZN(n7387) );
  INV_X1 U7423 ( .A(n7387), .ZN(n5979) );
  NAND2_X1 U7424 ( .A1(n5928), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5973) );
  INV_X1 U7425 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5967) );
  OR2_X1 U7426 ( .A1(n6258), .A2(n5967), .ZN(n5972) );
  NAND2_X1 U7427 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5982) );
  OAI21_X1 U7428 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n5982), .ZN(n7379) );
  OR2_X1 U7429 ( .A1(n5968), .A2(n7379), .ZN(n5971) );
  INV_X1 U7430 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6900) );
  OR2_X1 U7431 ( .A1(n6287), .A2(n6900), .ZN(n5970) );
  OR2_X1 U7432 ( .A1(n5987), .A2(n6156), .ZN(n5974) );
  XNOR2_X1 U7433 ( .A(n5974), .B(n5986), .ZN(n6916) );
  OR2_X1 U7434 ( .A1(n5975), .A2(n6562), .ZN(n5978) );
  OR2_X1 U7435 ( .A1(n5976), .A2(n9741), .ZN(n5977) );
  OAI211_X1 U7436 ( .C1(n6902), .C2(n6916), .A(n5978), .B(n5977), .ZN(n6953)
         );
  NAND2_X1 U7437 ( .A1(n5979), .A2(n4473), .ZN(n6933) );
  NAND2_X1 U7438 ( .A1(n5928), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5985) );
  INV_X1 U7439 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6901) );
  OR2_X1 U7440 ( .A1(n6287), .A2(n6901), .ZN(n5984) );
  INV_X1 U7441 ( .A(n5982), .ZN(n5980) );
  NAND2_X1 U7442 ( .A1(n5980), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6003) );
  INV_X1 U7443 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7444 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  NAND2_X1 U7445 ( .A1(n6003), .A2(n5983), .ZN(n7011) );
  INV_X1 U7446 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U7447 ( .A1(n5987), .A2(n5986), .ZN(n6020) );
  NAND2_X1 U7448 ( .A1(n6020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7449 ( .A(n5996), .B(n6018), .ZN(n7077) );
  OR2_X1 U7450 ( .A1(n6569), .A2(n5975), .ZN(n5989) );
  OR2_X1 U7451 ( .A1(n5976), .A2(n6570), .ZN(n5988) );
  INV_X1 U7452 ( .A(n7468), .ZN(n7122) );
  NAND2_X1 U7453 ( .A1(n8567), .A2(n10323), .ZN(n6934) );
  NAND2_X1 U7454 ( .A1(n6933), .A2(n6336), .ZN(n5990) );
  NAND2_X1 U7455 ( .A1(n5990), .A2(n6474), .ZN(n7365) );
  NAND2_X1 U7456 ( .A1(n5928), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5993) );
  INV_X1 U7457 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U7458 ( .A(n6003), .B(n6002), .ZN(n7373) );
  OR2_X1 U7459 ( .A1(n5968), .A2(n7373), .ZN(n5992) );
  INV_X1 U7460 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7078) );
  OR2_X1 U7461 ( .A1(n6287), .A2(n7078), .ZN(n5991) );
  INV_X1 U7462 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7463 ( .A1(n6258), .A2(n5994), .ZN(n5995) );
  INV_X2 U7464 ( .A(n5975), .ZN(n6171) );
  NAND2_X1 U7465 ( .A1(n6571), .A2(n6171), .ZN(n5999) );
  NAND2_X1 U7466 ( .A1(n5996), .A2(n6018), .ZN(n5997) );
  NAND2_X1 U7467 ( .A1(n5997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U7468 ( .A(n6011), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7108) );
  AOI22_X1 U7469 ( .A1(n6159), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6584), .B2(
        n7108), .ZN(n5998) );
  NAND2_X1 U7470 ( .A1(n5999), .A2(n5998), .ZN(n7132) );
  NAND2_X1 U7471 ( .A1(n10329), .A2(n8565), .ZN(n6338) );
  INV_X1 U7472 ( .A(n6340), .ZN(n6000) );
  NAND2_X1 U7473 ( .A1(n5928), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6010) );
  INV_X1 U7474 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7107) );
  OR2_X1 U7475 ( .A1(n6287), .A2(n7107), .ZN(n6009) );
  INV_X1 U7476 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U7477 ( .B1(n6003), .B2(n6002), .A(n6001), .ZN(n6006) );
  INV_X1 U7478 ( .A(n6003), .ZN(n6005) );
  NAND2_X1 U7479 ( .A1(n6005), .A2(n6004), .ZN(n6029) );
  NAND2_X1 U7480 ( .A1(n6006), .A2(n6029), .ZN(n7543) );
  OR2_X1 U7481 ( .A1(n5968), .A2(n7543), .ZN(n6008) );
  INV_X1 U7482 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7544) );
  OR2_X1 U7483 ( .A1(n6258), .A2(n7544), .ZN(n6007) );
  NAND4_X1 U7484 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n8564)
         );
  INV_X1 U7485 ( .A(n8564), .ZN(n7369) );
  NAND2_X1 U7486 ( .A1(n6575), .A2(n6171), .ZN(n6015) );
  INV_X1 U7487 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7488 ( .A1(n6011), .A2(n6017), .ZN(n6012) );
  NAND2_X1 U7489 ( .A1(n6012), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U7490 ( .A(n6013), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U7491 ( .A1(n6159), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6584), .B2(
        n7234), .ZN(n6014) );
  NAND2_X1 U7492 ( .A1(n6015), .A2(n6014), .ZN(n7323) );
  OR2_X1 U7493 ( .A1(n7369), .A2(n7323), .ZN(n6343) );
  NAND2_X1 U7494 ( .A1(n7323), .A2(n7369), .ZN(n6358) );
  INV_X1 U7495 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6016) );
  NAND3_X1 U7496 ( .A1(n6018), .A2(n6017), .A3(n6016), .ZN(n6019) );
  NOR2_X1 U7497 ( .A1(n6020), .A2(n6019), .ZN(n6023) );
  OR2_X1 U7498 ( .A1(n6023), .A2(n6156), .ZN(n6021) );
  MUX2_X1 U7499 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6021), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6024) );
  INV_X1 U7500 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7501 ( .A1(n6023), .A2(n6022), .ZN(n6048) );
  AOI22_X1 U7502 ( .A1(n6159), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6584), .B2(
        n8587), .ZN(n6025) );
  NAND2_X1 U7503 ( .A1(n6285), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6034) );
  INV_X1 U7504 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7113) );
  OR2_X1 U7505 ( .A1(n6287), .A2(n7113), .ZN(n6033) );
  INV_X1 U7506 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7507 ( .A1(n4465), .A2(n6027), .ZN(n6032) );
  INV_X1 U7508 ( .A(n6029), .ZN(n6028) );
  NAND2_X1 U7509 ( .A1(n6028), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6041) );
  INV_X1 U7510 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U7511 ( .A1(n6029), .A2(n8588), .ZN(n6030) );
  NAND2_X1 U7512 ( .A1(n6041), .A2(n6030), .ZN(n7337) );
  OR2_X1 U7513 ( .A1(n5968), .A2(n7337), .ZN(n6031) );
  NAND4_X1 U7514 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n8563)
         );
  INV_X1 U7515 ( .A(n8563), .ZN(n7478) );
  OR2_X1 U7516 ( .A1(n7479), .A2(n7478), .ZN(n6348) );
  NAND2_X1 U7517 ( .A1(n7479), .A2(n7478), .ZN(n6345) );
  NAND2_X1 U7518 ( .A1(n6348), .A2(n6345), .ZN(n7483) );
  INV_X1 U7519 ( .A(n7483), .ZN(n6035) );
  NAND2_X1 U7520 ( .A1(n6588), .A2(n6171), .ZN(n6038) );
  NAND2_X1 U7521 ( .A1(n6048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7522 ( .A(n6036), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8602) );
  AOI22_X1 U7523 ( .A1(n6159), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6584), .B2(
        n8602), .ZN(n6037) );
  NAND2_X1 U7524 ( .A1(n6285), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6046) );
  INV_X1 U7525 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6039) );
  OR2_X1 U7526 ( .A1(n4465), .A2(n6039), .ZN(n6045) );
  INV_X1 U7527 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7106) );
  OR2_X1 U7528 ( .A1(n6287), .A2(n7106), .ZN(n6044) );
  NAND2_X1 U7529 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7530 ( .A1(n6053), .A2(n6042), .ZN(n7495) );
  OR2_X1 U7531 ( .A1(n5968), .A2(n7495), .ZN(n6043) );
  NAND4_X1 U7532 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n8562)
         );
  INV_X1 U7533 ( .A(n8562), .ZN(n7347) );
  OR2_X1 U7534 ( .A1(n7630), .A2(n7347), .ZN(n6347) );
  NAND2_X1 U7535 ( .A1(n7630), .A2(n7347), .ZN(n6355) );
  NAND2_X1 U7536 ( .A1(n7476), .A2(n7490), .ZN(n6047) );
  NAND2_X1 U7537 ( .A1(n6597), .A2(n6171), .ZN(n6051) );
  NAND2_X1 U7538 ( .A1(n6060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6049) );
  XNOR2_X1 U7539 ( .A(n6049), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7151) );
  AOI22_X1 U7540 ( .A1(n6159), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6584), .B2(
        n7151), .ZN(n6050) );
  NAND2_X1 U7541 ( .A1(n5928), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6058) );
  INV_X1 U7542 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7511) );
  OR2_X1 U7543 ( .A1(n6258), .A2(n7511), .ZN(n6057) );
  INV_X1 U7544 ( .A(n6053), .ZN(n6052) );
  NAND2_X1 U7545 ( .A1(n6052), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6067) );
  INV_X1 U7546 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U7547 ( .A1(n6053), .A2(n7346), .ZN(n6054) );
  NAND2_X1 U7548 ( .A1(n6067), .A2(n6054), .ZN(n7510) );
  OR2_X1 U7549 ( .A1(n5968), .A2(n7510), .ZN(n6056) );
  INV_X1 U7550 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7115) );
  OR2_X1 U7551 ( .A1(n6287), .A2(n7115), .ZN(n6055) );
  NAND4_X1 U7552 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n8561)
         );
  INV_X1 U7553 ( .A(n8561), .ZN(n7477) );
  OR2_X1 U7554 ( .A1(n7647), .A2(n7477), .ZN(n7694) );
  NAND2_X1 U7555 ( .A1(n7647), .A2(n7477), .ZN(n6362) );
  NAND2_X1 U7556 ( .A1(n7694), .A2(n6362), .ZN(n6476) );
  INV_X1 U7557 ( .A(n6476), .ZN(n6059) );
  NAND2_X1 U7558 ( .A1(n4454), .A2(n6059), .ZN(n7507) );
  NAND2_X1 U7559 ( .A1(n6595), .A2(n6171), .ZN(n6065) );
  OAI21_X1 U7560 ( .B1(n6060), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6062) );
  INV_X1 U7561 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7562 ( .A(n6062), .B(n6061), .ZN(n7174) );
  INV_X1 U7563 ( .A(n7174), .ZN(n6063) );
  AOI22_X1 U7564 ( .A1(n6159), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6584), .B2(
        n6063), .ZN(n6064) );
  NAND2_X1 U7565 ( .A1(n5928), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6072) );
  INV_X1 U7566 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7173) );
  OR2_X1 U7567 ( .A1(n6258), .A2(n7173), .ZN(n6071) );
  NAND2_X1 U7568 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  NAND2_X1 U7569 ( .A1(n6079), .A2(n6068), .ZN(n7735) );
  OR2_X1 U7570 ( .A1(n4463), .A2(n7735), .ZN(n6070) );
  INV_X1 U7571 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7157) );
  OR2_X1 U7572 ( .A1(n6287), .A2(n7157), .ZN(n6069) );
  NAND4_X1 U7573 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n8560)
         );
  AND2_X1 U7574 ( .A1(n7694), .A2(n6478), .ZN(n7653) );
  NAND2_X1 U7575 ( .A1(n6621), .A2(n6171), .ZN(n6075) );
  XNOR2_X1 U7576 ( .A(n6073), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7206) );
  AOI22_X1 U7577 ( .A1(n6159), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6584), .B2(
        n7206), .ZN(n6074) );
  NAND2_X1 U7578 ( .A1(n6075), .A2(n6074), .ZN(n7781) );
  NAND2_X1 U7579 ( .A1(n5928), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6085) );
  INV_X1 U7580 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7581 ( .A1(n6287), .A2(n6076), .ZN(n6084) );
  INV_X1 U7582 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7583 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7584 ( .A1(n6092), .A2(n6080), .ZN(n7624) );
  OR2_X1 U7585 ( .A1(n5968), .A2(n7624), .ZN(n6083) );
  INV_X1 U7586 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6081) );
  OR2_X1 U7587 ( .A1(n6258), .A2(n6081), .ZN(n6082) );
  NAND4_X1 U7588 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n8559)
         );
  INV_X1 U7589 ( .A(n8559), .ZN(n7640) );
  NOR2_X1 U7590 ( .A1(n7781), .A2(n7640), .ZN(n6368) );
  INV_X1 U7591 ( .A(n6368), .ZN(n6367) );
  AND2_X1 U7592 ( .A1(n7653), .A2(n6367), .ZN(n6086) );
  NAND2_X1 U7593 ( .A1(n7781), .A2(n7640), .ZN(n6369) );
  NAND2_X1 U7594 ( .A1(n7734), .A2(n7658), .ZN(n7654) );
  NOR2_X1 U7595 ( .A1(n6087), .A2(n5084), .ZN(n6088) );
  NAND2_X1 U7596 ( .A1(n6709), .A2(n6171), .ZN(n6090) );
  NAND2_X1 U7597 ( .A1(n6121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7598 ( .A(n6099), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7295) );
  AOI22_X1 U7599 ( .A1(n6159), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6584), .B2(
        n7295), .ZN(n6089) );
  NAND2_X1 U7600 ( .A1(n5928), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6097) );
  INV_X1 U7601 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7795) );
  OR2_X1 U7602 ( .A1(n6258), .A2(n7795), .ZN(n6096) );
  NAND2_X1 U7603 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  NAND2_X1 U7604 ( .A1(n6104), .A2(n6093), .ZN(n7794) );
  OR2_X1 U7605 ( .A1(n4463), .A2(n7794), .ZN(n6095) );
  INV_X1 U7606 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9616) );
  OR2_X1 U7607 ( .A1(n6287), .A2(n9616), .ZN(n6094) );
  NAND4_X1 U7608 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n8558)
         );
  OR2_X1 U7609 ( .A1(n8984), .A2(n7767), .ZN(n6373) );
  NAND2_X1 U7610 ( .A1(n8984), .A2(n7767), .ZN(n6098) );
  INV_X1 U7611 ( .A(n6098), .ZN(n6375) );
  NAND2_X1 U7612 ( .A1(n6719), .A2(n6171), .ZN(n6102) );
  NAND2_X1 U7613 ( .A1(n6099), .A2(n6122), .ZN(n6100) );
  NAND2_X1 U7614 ( .A1(n6100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6112) );
  XNOR2_X1 U7615 ( .A(n6112), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7574) );
  AOI22_X1 U7616 ( .A1(n6159), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6584), .B2(
        n7574), .ZN(n6101) );
  NAND2_X1 U7617 ( .A1(n5928), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6110) );
  INV_X1 U7618 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9680) );
  OR2_X1 U7619 ( .A1(n6287), .A2(n9680), .ZN(n6109) );
  NAND2_X1 U7620 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  NAND2_X1 U7621 ( .A1(n6130), .A2(n6105), .ZN(n7766) );
  OR2_X1 U7622 ( .A1(n5968), .A2(n7766), .ZN(n6108) );
  INV_X1 U7623 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7624 ( .A1(n6258), .A2(n6106), .ZN(n6107) );
  NAND4_X1 U7625 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n8557)
         );
  INV_X1 U7626 ( .A(n8557), .ZN(n7805) );
  NAND2_X1 U7627 ( .A1(n8977), .A2(n7805), .ZN(n6378) );
  NAND2_X1 U7628 ( .A1(n6924), .A2(n6171), .ZN(n6116) );
  INV_X1 U7629 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7630 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  NAND2_X1 U7631 ( .A1(n6113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7632 ( .A(n6114), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8611) );
  AOI22_X1 U7633 ( .A1(n6159), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6584), .B2(
        n8611), .ZN(n6115) );
  NAND2_X1 U7634 ( .A1(n5928), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6120) );
  INV_X1 U7635 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9651) );
  OR2_X1 U7636 ( .A1(n6287), .A2(n9651), .ZN(n6119) );
  INV_X1 U7637 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7804) );
  XNOR2_X1 U7638 ( .A(n6130), .B(n7804), .ZN(n7854) );
  OR2_X1 U7639 ( .A1(n4463), .A2(n7854), .ZN(n6118) );
  INV_X1 U7640 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7855) );
  OR2_X1 U7641 ( .A1(n6258), .A2(n7855), .ZN(n6117) );
  NAND4_X1 U7642 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n8872)
         );
  INV_X1 U7643 ( .A(n8872), .ZN(n7921) );
  NOR2_X1 U7644 ( .A1(n8972), .A2(n7921), .ZN(n6384) );
  NAND2_X1 U7645 ( .A1(n8972), .A2(n7921), .ZN(n6383) );
  NAND2_X1 U7646 ( .A1(n6940), .A2(n6171), .ZN(n6126) );
  NAND2_X1 U7647 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7648 ( .A(n6124), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8631) );
  AOI22_X1 U7649 ( .A1(n6159), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6584), .B2(
        n8631), .ZN(n6125) );
  NAND2_X1 U7650 ( .A1(n5928), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6135) );
  INV_X1 U7651 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8884) );
  OR2_X1 U7652 ( .A1(n6258), .A2(n8884), .ZN(n6134) );
  AND2_X1 U7653 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6127) );
  INV_X1 U7654 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7655 ( .B1(n6130), .B2(n7804), .A(n6129), .ZN(n6131) );
  NAND2_X1 U7656 ( .A1(n6141), .A2(n6131), .ZN(n8883) );
  OR2_X1 U7657 ( .A1(n5968), .A2(n8883), .ZN(n6133) );
  INV_X1 U7658 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9810) );
  OR2_X1 U7659 ( .A1(n6287), .A2(n9810), .ZN(n6132) );
  NAND4_X1 U7660 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n8556)
         );
  INV_X1 U7661 ( .A(n8556), .ZN(n8849) );
  OR2_X1 U7662 ( .A1(n8964), .A2(n8849), .ZN(n6389) );
  NAND2_X1 U7663 ( .A1(n8964), .A2(n8849), .ZN(n8844) );
  NAND2_X1 U7664 ( .A1(n6988), .A2(n6171), .ZN(n6139) );
  NAND2_X1 U7665 ( .A1(n4533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7666 ( .A(n6137), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8659) );
  AOI22_X1 U7667 ( .A1(n6159), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6584), .B2(
        n8659), .ZN(n6138) );
  NAND2_X1 U7668 ( .A1(n5928), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6146) );
  INV_X1 U7669 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8630) );
  OR2_X1 U7670 ( .A1(n6287), .A2(n8630), .ZN(n6145) );
  INV_X1 U7671 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U7672 ( .A1(n6141), .A2(n8629), .ZN(n6142) );
  NAND2_X1 U7673 ( .A1(n6164), .A2(n6142), .ZN(n8855) );
  OR2_X1 U7674 ( .A1(n4463), .A2(n8855), .ZN(n6144) );
  INV_X1 U7675 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8642) );
  OR2_X1 U7676 ( .A1(n6258), .A2(n8642), .ZN(n6143) );
  NAND4_X1 U7677 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n8874)
         );
  INV_X1 U7678 ( .A(n8874), .ZN(n8532) );
  NAND2_X1 U7679 ( .A1(n8961), .A2(n8532), .ZN(n6394) );
  NAND2_X1 U7680 ( .A1(n6393), .A2(n6394), .ZN(n8845) );
  INV_X1 U7681 ( .A(n8844), .ZN(n6390) );
  INV_X1 U7682 ( .A(n6393), .ZN(n6147) );
  NAND2_X1 U7683 ( .A1(n7308), .A2(n6171), .ZN(n6150) );
  XNOR2_X1 U7684 ( .A(n6158), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8671) );
  AOI22_X1 U7685 ( .A1(n6159), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6584), .B2(
        n8671), .ZN(n6149) );
  XNOR2_X1 U7686 ( .A(n6164), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U7687 ( .A1(n8831), .A2(n5952), .ZN(n6154) );
  NAND2_X1 U7688 ( .A1(n4466), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7689 ( .A1(n5928), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7690 ( .A1(n6285), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6151) );
  NAND4_X1 U7691 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n8555)
         );
  AND2_X1 U7692 ( .A1(n8954), .A2(n8851), .ZN(n6399) );
  OR2_X1 U7693 ( .A1(n8954), .A2(n8851), .ZN(n6466) );
  NAND2_X1 U7694 ( .A1(n7361), .A2(n6171), .ZN(n6161) );
  AOI22_X1 U7695 ( .A1(n6159), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4460), .B2(
        n6584), .ZN(n6160) );
  INV_X1 U7696 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8529) );
  INV_X1 U7697 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U7698 ( .B1(n6164), .B2(n8529), .A(n6162), .ZN(n6165) );
  NAND2_X1 U7699 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6163) );
  NAND2_X1 U7700 ( .A1(n6165), .A2(n6175), .ZN(n8823) );
  INV_X1 U7701 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9828) );
  OR2_X1 U7702 ( .A1(n4465), .A2(n9828), .ZN(n6168) );
  INV_X1 U7703 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7704 ( .A1(n6258), .A2(n6166), .ZN(n6167) );
  AND2_X1 U7705 ( .A1(n6168), .A2(n6167), .ZN(n6170) );
  NAND2_X1 U7706 ( .A1(n4466), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6169) );
  OAI211_X1 U7707 ( .C1(n8823), .C2(n4463), .A(n6170), .B(n6169), .ZN(n8836)
         );
  INV_X1 U7708 ( .A(n8836), .ZN(n8810) );
  OR2_X1 U7709 ( .A1(n8951), .A2(n8810), .ZN(n6411) );
  NAND2_X1 U7710 ( .A1(n8951), .A2(n8810), .ZN(n6400) );
  NAND2_X1 U7711 ( .A1(n6411), .A2(n6400), .ZN(n8818) );
  NAND2_X1 U7712 ( .A1(n7571), .A2(n6171), .ZN(n6173) );
  OR2_X1 U7713 ( .A1(n5976), .A2(n7669), .ZN(n6172) );
  INV_X1 U7714 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6179) );
  INV_X1 U7715 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U7716 ( .A1(n6175), .A2(n9626), .ZN(n6176) );
  NAND2_X1 U7717 ( .A1(n6183), .A2(n6176), .ZN(n8804) );
  OR2_X1 U7718 ( .A1(n8804), .A2(n5968), .ZN(n6178) );
  AOI22_X1 U7719 ( .A1(n4466), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5928), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7720 ( .C1(n6258), .C2(n6179), .A(n6178), .B(n6177), .ZN(n8794)
         );
  INV_X1 U7721 ( .A(n8794), .ZN(n8821) );
  NAND2_X1 U7722 ( .A1(n8944), .A2(n8821), .ZN(n6416) );
  NAND2_X1 U7723 ( .A1(n6180), .A2(n6416), .ZN(n8808) );
  INV_X1 U7724 ( .A(n6180), .ZN(n6401) );
  NAND2_X1 U7725 ( .A1(n7665), .A2(n6171), .ZN(n6182) );
  INV_X1 U7726 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7667) );
  OR2_X1 U7727 ( .A1(n5976), .A2(n7667), .ZN(n6181) );
  INV_X1 U7728 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U7729 ( .A1(n6183), .A2(n8476), .ZN(n6184) );
  NAND2_X1 U7730 ( .A1(n6192), .A2(n6184), .ZN(n8788) );
  AOI22_X1 U7731 ( .A1(n4466), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5928), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6187) );
  INV_X1 U7732 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6185) );
  OR2_X1 U7733 ( .A1(n6258), .A2(n6185), .ZN(n6186) );
  OAI211_X1 U7734 ( .C1(n8788), .C2(n4463), .A(n6187), .B(n6186), .ZN(n8779)
         );
  XNOR2_X1 U7735 ( .A(n8939), .B(n8779), .ZN(n8792) );
  INV_X1 U7736 ( .A(n8939), .ZN(n8791) );
  NOR2_X1 U7737 ( .A1(n8791), .A2(n8779), .ZN(n6419) );
  NAND2_X1 U7738 ( .A1(n8067), .A2(n6171), .ZN(n6189) );
  OR2_X1 U7739 ( .A1(n5976), .A2(n8068), .ZN(n6188) );
  INV_X1 U7740 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7741 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  NAND2_X1 U7742 ( .A1(n6203), .A2(n6193), .ZN(n8772) );
  OR2_X1 U7743 ( .A1(n8772), .A2(n5968), .ZN(n6199) );
  INV_X1 U7744 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7745 ( .A1(n4466), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7746 ( .A1(n5928), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7747 ( .C1(n6196), .C2(n6258), .A(n6195), .B(n6194), .ZN(n6197)
         );
  INV_X1 U7748 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7749 ( .A1(n6199), .A2(n6198), .ZN(n8795) );
  INV_X1 U7750 ( .A(n8795), .ZN(n8477) );
  NOR2_X1 U7751 ( .A1(n6200), .A2(n8477), .ZN(n6405) );
  NAND2_X1 U7752 ( .A1(n8778), .A2(n8777), .ZN(n8776) );
  INV_X1 U7753 ( .A(n6405), .ZN(n6421) );
  NAND2_X1 U7754 ( .A1(n8776), .A2(n6421), .ZN(n8756) );
  NAND2_X1 U7755 ( .A1(n7748), .A2(n6171), .ZN(n6202) );
  OR2_X1 U7756 ( .A1(n5976), .A2(n7751), .ZN(n6201) );
  INV_X1 U7757 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U7758 ( .A1(n6203), .A2(n8462), .ZN(n6204) );
  AND2_X1 U7759 ( .A1(n6212), .A2(n6204), .ZN(n8762) );
  NAND2_X1 U7760 ( .A1(n8762), .A2(n5952), .ZN(n6209) );
  INV_X1 U7761 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U7762 ( .A1(n6285), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7763 ( .A1(n4466), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7764 ( .C1(n4465), .C2(n9743), .A(n6206), .B(n6205), .ZN(n6207)
         );
  INV_X1 U7765 ( .A(n6207), .ZN(n6208) );
  NAND2_X1 U7766 ( .A1(n6209), .A2(n6208), .ZN(n8780) );
  NAND2_X1 U7767 ( .A1(n8930), .A2(n8749), .ZN(n6424) );
  OR2_X1 U7768 ( .A1(n5976), .A2(n7824), .ZN(n6210) );
  INV_X1 U7769 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U7770 ( .A1(n6212), .A2(n9629), .ZN(n6213) );
  NAND2_X1 U7771 ( .A1(n6228), .A2(n6213), .ZN(n8507) );
  INV_X1 U7772 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7773 ( .A1(n5928), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7774 ( .A1(n4466), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6214) );
  OAI211_X1 U7775 ( .C1(n6258), .C2(n6216), .A(n6215), .B(n6214), .ZN(n6217)
         );
  OR2_X1 U7776 ( .A1(n8924), .A2(n8486), .ZN(n6426) );
  NAND2_X1 U7777 ( .A1(n8924), .A2(n8486), .ZN(n6430) );
  NAND2_X1 U7778 ( .A1(n6426), .A2(n6430), .ZN(n8747) );
  INV_X1 U7779 ( .A(n6426), .ZN(n6409) );
  NAND2_X1 U7780 ( .A1(n7926), .A2(n6171), .ZN(n6219) );
  OR2_X1 U7781 ( .A1(n5976), .A2(n7931), .ZN(n6218) );
  XNOR2_X1 U7782 ( .A(n6228), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8734) );
  INV_X1 U7783 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7784 ( .A1(n4466), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7785 ( .A1(n5928), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6220) );
  OAI211_X1 U7786 ( .C1(n6222), .C2(n6258), .A(n6221), .B(n6220), .ZN(n6223)
         );
  AOI21_X1 U7787 ( .B1(n8734), .B2(n5952), .A(n6223), .ZN(n8750) );
  NAND2_X1 U7788 ( .A1(n8921), .A2(n8750), .ZN(n6434) );
  NAND2_X1 U7789 ( .A1(n7945), .A2(n6171), .ZN(n6225) );
  OR2_X1 U7790 ( .A1(n5976), .A2(n7947), .ZN(n6224) );
  INV_X1 U7791 ( .A(n6228), .ZN(n6227) );
  AND2_X1 U7792 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n6226) );
  NAND2_X1 U7793 ( .A1(n6227), .A2(n6226), .ZN(n6239) );
  INV_X1 U7794 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8489) );
  INV_X1 U7795 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8545) );
  OAI21_X1 U7796 ( .B1(n6228), .B2(n8489), .A(n8545), .ZN(n6229) );
  AND2_X1 U7797 ( .A1(n6239), .A2(n6229), .ZN(n8722) );
  NAND2_X1 U7798 ( .A1(n8722), .A2(n5952), .ZN(n6235) );
  INV_X1 U7799 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7800 ( .A1(n4466), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7801 ( .A1(n5928), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6230) );
  OAI211_X1 U7802 ( .C1(n6232), .C2(n6258), .A(n6231), .B(n6230), .ZN(n6233)
         );
  INV_X1 U7803 ( .A(n6233), .ZN(n6234) );
  NAND2_X1 U7804 ( .A1(n6235), .A2(n6234), .ZN(n8553) );
  NAND2_X1 U7805 ( .A1(n8725), .A2(n8553), .ZN(n6437) );
  INV_X1 U7806 ( .A(n8553), .ZN(n8704) );
  NAND2_X1 U7807 ( .A1(n8916), .A2(n8704), .ZN(n6438) );
  NAND2_X1 U7808 ( .A1(n6437), .A2(n6438), .ZN(n7995) );
  INV_X1 U7809 ( .A(n6438), .ZN(n8703) );
  NAND2_X1 U7810 ( .A1(n7954), .A2(n6171), .ZN(n6237) );
  OR2_X1 U7811 ( .A1(n5976), .A2(n7956), .ZN(n6236) );
  INV_X1 U7812 ( .A(n6239), .ZN(n6238) );
  NAND2_X1 U7813 ( .A1(n6238), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6254) );
  INV_X1 U7814 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U7815 ( .A1(n6239), .A2(n9811), .ZN(n6240) );
  NAND2_X1 U7816 ( .A1(n6254), .A2(n6240), .ZN(n8698) );
  INV_X1 U7817 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7818 ( .A1(n4466), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7819 ( .A1(n5928), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6241) );
  OAI211_X1 U7820 ( .C1(n6243), .C2(n6258), .A(n6242), .B(n6241), .ZN(n6244)
         );
  INV_X1 U7821 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7822 ( .A1(n6246), .A2(n6245), .ZN(n8552) );
  NAND2_X1 U7823 ( .A1(n8909), .A2(n8443), .ZN(n6442) );
  INV_X1 U7824 ( .A(n6247), .ZN(n6444) );
  NOR2_X1 U7825 ( .A1(n8701), .A2(n6444), .ZN(n8002) );
  NAND2_X1 U7826 ( .A1(n6249), .A2(n6248), .ZN(n6251) );
  NAND2_X1 U7827 ( .A1(n6251), .A2(n6250), .ZN(n6263) );
  MUX2_X1 U7828 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6555), .Z(n6264) );
  XNOR2_X1 U7829 ( .A(n6264), .B(n9735), .ZN(n6262) );
  NAND2_X1 U7830 ( .A1(n8449), .A2(n6171), .ZN(n6253) );
  INV_X1 U7831 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8450) );
  OR2_X1 U7832 ( .A1(n5976), .A2(n8450), .ZN(n6252) );
  INV_X1 U7833 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U7834 ( .A1(n6254), .A2(n8441), .ZN(n6255) );
  INV_X1 U7835 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7836 ( .A1(n4466), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7837 ( .A1(n5928), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6256) );
  OAI211_X1 U7838 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n6256), .ZN(n6260)
         );
  AOI21_X1 U7839 ( .B1(n8440), .B2(n5952), .A(n6260), .ZN(n8705) );
  NAND2_X1 U7840 ( .A1(n8904), .A2(n8705), .ZN(n6446) );
  INV_X1 U7841 ( .A(n6261), .ZN(n6447) );
  NOR2_X1 U7842 ( .A1(n8001), .A2(n6447), .ZN(n8368) );
  OR2_X1 U7843 ( .A1(n6264), .A2(SI_28_), .ZN(n6265) );
  INV_X1 U7844 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9889) );
  INV_X1 U7845 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9019) );
  MUX2_X1 U7846 ( .A(n9889), .B(n9019), .S(n6555), .Z(n6275) );
  XNOR2_X1 U7847 ( .A(n6275), .B(SI_29_), .ZN(n6266) );
  NAND2_X1 U7848 ( .A1(n9017), .A2(n6171), .ZN(n6268) );
  OR2_X1 U7849 ( .A1(n5976), .A2(n9019), .ZN(n6267) );
  INV_X1 U7850 ( .A(n6269), .ZN(n8376) );
  INV_X1 U7851 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7852 ( .A1(n4466), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7853 ( .A1(n6285), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U7854 ( .C1(n4465), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6273)
         );
  AOI21_X1 U7855 ( .B1(n8376), .B2(n5952), .A(n6273), .ZN(n8444) );
  AOI21_X1 U7856 ( .B1(n8368), .B2(n6452), .A(n6455), .ZN(n6298) );
  INV_X1 U7857 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U7858 ( .A1(n6276), .A2(SI_29_), .ZN(n6277) );
  NAND2_X1 U7859 ( .A1(n6278), .A2(n6277), .ZN(n6302) );
  MUX2_X1 U7860 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6555), .Z(n6301) );
  NAND2_X1 U7861 ( .A1(n8451), .A2(n6171), .ZN(n6280) );
  INV_X1 U7862 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9639) );
  OR2_X1 U7863 ( .A1(n5976), .A2(n9639), .ZN(n6279) );
  NAND2_X1 U7864 ( .A1(n5928), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7865 ( .A1(n6285), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6283) );
  INV_X1 U7866 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6281) );
  OR2_X1 U7867 ( .A1(n6287), .A2(n6281), .ZN(n6282) );
  AND3_X1 U7868 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(n8372) );
  OR2_X1 U7869 ( .A1(n6297), .A2(n8372), .ZN(n6456) );
  NAND2_X1 U7870 ( .A1(n6285), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7871 ( .A1(n5928), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6289) );
  INV_X1 U7872 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6286) );
  OR2_X1 U7873 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  AND3_X1 U7874 ( .A1(n6290), .A2(n6289), .A3(n6288), .ZN(n8685) );
  INV_X1 U7875 ( .A(n6291), .ZN(n6292) );
  NOR2_X1 U7876 ( .A1(n6292), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7877 ( .A1(n8685), .A2(n6747), .ZN(n6299) );
  NAND2_X1 U7878 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  MUX2_X1 U7879 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6555), .Z(n6304) );
  XNOR2_X1 U7880 ( .A(n6304), .B(SI_31_), .ZN(n6305) );
  NAND2_X1 U7881 ( .A1(n8160), .A2(n6171), .ZN(n6307) );
  INV_X1 U7882 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9013) );
  OR2_X1 U7883 ( .A1(n4462), .A2(n9013), .ZN(n6306) );
  NAND2_X1 U7884 ( .A1(n6307), .A2(n6306), .ZN(n8683) );
  NAND2_X1 U7885 ( .A1(n6297), .A2(n8372), .ZN(n6458) );
  NAND2_X1 U7886 ( .A1(n6315), .A2(n6458), .ZN(n6454) );
  NAND2_X1 U7887 ( .A1(n8683), .A2(n8685), .ZN(n6457) );
  XNOR2_X1 U7888 ( .A(n6308), .B(n4919), .ZN(n6491) );
  NAND2_X1 U7889 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  AND2_X1 U7890 ( .A1(n6314), .A2(n6747), .ZN(n6754) );
  NOR2_X1 U7891 ( .A1(n7025), .A2(n6754), .ZN(n6490) );
  INV_X1 U7892 ( .A(n6315), .ZN(n6462) );
  NOR2_X1 U7893 ( .A1(n4919), .A2(n7666), .ZN(n6316) );
  NAND2_X1 U7894 ( .A1(n6316), .A2(n6463), .ZN(n6461) );
  INV_X1 U7895 ( .A(n6461), .ZN(n6432) );
  NOR2_X1 U7896 ( .A1(n8795), .A2(n6461), .ZN(n6410) );
  NAND2_X1 U7897 ( .A1(n8569), .A2(n7443), .ZN(n7024) );
  NAND2_X1 U7898 ( .A1(n7024), .A2(n6469), .ZN(n6318) );
  NAND3_X1 U7899 ( .A1(n6324), .A2(n6470), .A3(n6318), .ZN(n6319) );
  NAND2_X1 U7900 ( .A1(n6319), .A2(n6322), .ZN(n6327) );
  NAND3_X1 U7901 ( .A1(n7024), .A2(n6469), .A3(n6747), .ZN(n6321) );
  NAND2_X1 U7902 ( .A1(n6320), .A2(n6321), .ZN(n6323) );
  NAND2_X1 U7903 ( .A1(n6323), .A2(n6322), .ZN(n6325) );
  NAND2_X1 U7904 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  MUX2_X1 U7905 ( .A(n6327), .B(n6326), .S(n6461), .Z(n6329) );
  INV_X1 U7906 ( .A(n6337), .ZN(n6328) );
  NAND3_X1 U7907 ( .A1(n6329), .A2(n6753), .A3(n6328), .ZN(n6334) );
  AND2_X1 U7908 ( .A1(n4473), .A2(n6330), .ZN(n6331) );
  NAND2_X1 U7909 ( .A1(n6332), .A2(n6461), .ZN(n6333) );
  AOI22_X1 U7910 ( .A1(n6337), .A2(n6473), .B1(n6336), .B2(n6335), .ZN(n6339)
         );
  OAI21_X1 U7911 ( .B1(n6339), .B2(n4682), .A(n6432), .ZN(n6342) );
  OAI21_X1 U7912 ( .B1(n6461), .B2(n6340), .A(n7129), .ZN(n6341) );
  INV_X1 U7913 ( .A(n6343), .ZN(n6344) );
  INV_X1 U7914 ( .A(n6345), .ZN(n6346) );
  INV_X1 U7915 ( .A(n6347), .ZN(n6352) );
  INV_X1 U7916 ( .A(n6348), .ZN(n6349) );
  NOR2_X1 U7917 ( .A1(n6352), .A2(n6349), .ZN(n6350) );
  MUX2_X1 U7918 ( .A(n6351), .B(n6350), .S(n6461), .Z(n6356) );
  OR2_X1 U7919 ( .A1(n6476), .A2(n6352), .ZN(n6354) );
  NAND2_X1 U7920 ( .A1(n6362), .A2(n6355), .ZN(n6353) );
  AOI21_X1 U7921 ( .B1(n6356), .B2(n6355), .A(n6357), .ZN(n6366) );
  INV_X1 U7922 ( .A(n6357), .ZN(n6360) );
  NAND4_X1 U7923 ( .A1(n6360), .A2(n6035), .A3(n6359), .A4(n6358), .ZN(n6361)
         );
  NAND3_X1 U7924 ( .A1(n6361), .A2(n7694), .A3(n6478), .ZN(n6364) );
  NAND2_X1 U7925 ( .A1(n7654), .A2(n6362), .ZN(n6363) );
  NAND2_X1 U7926 ( .A1(n6367), .A2(n6369), .ZN(n7652) );
  AOI21_X1 U7927 ( .B1(n6478), .B2(n6367), .A(n6087), .ZN(n6371) );
  AOI21_X1 U7928 ( .B1(n7654), .B2(n6369), .A(n6368), .ZN(n6370) );
  MUX2_X1 U7929 ( .A(n6371), .B(n6370), .S(n6461), .Z(n6372) );
  INV_X1 U7930 ( .A(n6373), .ZN(n6374) );
  MUX2_X1 U7931 ( .A(n6375), .B(n6374), .S(n6461), .Z(n6376) );
  INV_X1 U7932 ( .A(n7858), .ZN(n7811) );
  INV_X1 U7933 ( .A(n6377), .ZN(n6380) );
  INV_X1 U7934 ( .A(n6378), .ZN(n6379) );
  MUX2_X1 U7935 ( .A(n6380), .B(n6379), .S(n6461), .Z(n6382) );
  INV_X1 U7936 ( .A(n6384), .ZN(n6381) );
  NAND2_X1 U7937 ( .A1(n6381), .A2(n6383), .ZN(n7860) );
  INV_X1 U7938 ( .A(n6383), .ZN(n6385) );
  MUX2_X1 U7939 ( .A(n6385), .B(n6384), .S(n6461), .Z(n6387) );
  INV_X1 U7940 ( .A(n8870), .ZN(n6386) );
  INV_X1 U7941 ( .A(n6389), .ZN(n6391) );
  MUX2_X1 U7942 ( .A(n6391), .B(n6390), .S(n6461), .Z(n6392) );
  NAND2_X1 U7943 ( .A1(n6466), .A2(n6393), .ZN(n6396) );
  INV_X1 U7944 ( .A(n6394), .ZN(n6395) );
  MUX2_X1 U7945 ( .A(n6396), .B(n6395), .S(n6432), .Z(n6397) );
  INV_X1 U7946 ( .A(n6466), .ZN(n6398) );
  INV_X1 U7947 ( .A(n6399), .ZN(n6465) );
  NAND2_X1 U7948 ( .A1(n6400), .A2(n6465), .ZN(n6412) );
  INV_X1 U7949 ( .A(n8779), .ZN(n8811) );
  NOR2_X1 U7950 ( .A1(n8939), .A2(n8811), .ZN(n6402) );
  NOR2_X1 U7951 ( .A1(n6402), .A2(n6401), .ZN(n6414) );
  INV_X1 U7952 ( .A(n6416), .ZN(n6404) );
  INV_X1 U7953 ( .A(n6402), .ZN(n6403) );
  OAI21_X1 U7954 ( .B1(n6419), .B2(n6404), .A(n6403), .ZN(n6406) );
  AOI211_X1 U7955 ( .C1(n6407), .C2(n6406), .A(n6405), .B(n6461), .ZN(n6408)
         );
  AOI211_X1 U7956 ( .C1(n6410), .C2(n6200), .A(n6409), .B(n6408), .ZN(n6429)
         );
  OAI21_X1 U7957 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(n6417) );
  INV_X1 U7958 ( .A(n6414), .ZN(n6415) );
  AOI21_X1 U7959 ( .B1(n6417), .B2(n6416), .A(n6415), .ZN(n6423) );
  INV_X1 U7960 ( .A(n6418), .ZN(n6420) );
  NAND3_X1 U7961 ( .A1(n6420), .A2(n6461), .A3(n4878), .ZN(n6422) );
  OAI22_X1 U7962 ( .A1(n6423), .A2(n6422), .B1(n6432), .B2(n6421), .ZN(n6425)
         );
  OAI22_X1 U7963 ( .A1(n6425), .A2(n8758), .B1(n6432), .B2(n6424), .ZN(n6428)
         );
  OAI21_X1 U7964 ( .B1(n8749), .B2(n8930), .A(n6426), .ZN(n6427) );
  AOI22_X1 U7965 ( .A1(n6429), .A2(n6428), .B1(n6432), .B2(n6427), .ZN(n6431)
         );
  NAND2_X1 U7966 ( .A1(n6437), .A2(n8714), .ZN(n6436) );
  NAND2_X1 U7967 ( .A1(n6438), .A2(n6434), .ZN(n6435) );
  MUX2_X1 U7968 ( .A(n6436), .B(n6435), .S(n6461), .Z(n6440) );
  INV_X1 U7969 ( .A(n8702), .ZN(n7996) );
  MUX2_X1 U7970 ( .A(n6438), .B(n6437), .S(n6461), .Z(n6439) );
  INV_X1 U7971 ( .A(n6442), .ZN(n6443) );
  MUX2_X1 U7972 ( .A(n6444), .B(n6443), .S(n6461), .Z(n6445) );
  NOR2_X1 U7973 ( .A1(n8365), .A2(n6445), .ZN(n6451) );
  INV_X1 U7974 ( .A(n6446), .ZN(n6448) );
  MUX2_X1 U7975 ( .A(n6448), .B(n6447), .S(n6461), .Z(n6450) );
  INV_X1 U7976 ( .A(n6455), .ZN(n6449) );
  INV_X1 U7977 ( .A(n6452), .ZN(n6453) );
  NAND2_X1 U7978 ( .A1(n6457), .A2(n6456), .ZN(n6486) );
  INV_X1 U7979 ( .A(n6804), .ZN(n10308) );
  INV_X1 U7980 ( .A(n8365), .ZN(n7997) );
  NAND2_X1 U7981 ( .A1(n6466), .A2(n6465), .ZN(n8834) );
  NAND2_X1 U7982 ( .A1(n6468), .A2(n7024), .ZN(n10309) );
  NOR4_X1 U7983 ( .A1(n7284), .A2(n10309), .A3(n7438), .A4(n4455), .ZN(n6471)
         );
  AND2_X1 U7984 ( .A1(n4473), .A2(n6934), .ZN(n7388) );
  NAND3_X1 U7985 ( .A1(n6471), .A2(n6753), .A3(n7388), .ZN(n6475) );
  NAND2_X1 U7986 ( .A1(n6474), .A2(n6473), .ZN(n6936) );
  NOR4_X1 U7987 ( .A1(n6475), .A2(n7480), .A3(n7366), .A4(n6936), .ZN(n6477)
         );
  NAND4_X1 U7988 ( .A1(n6477), .A2(n6059), .A3(n6035), .A4(n7490), .ZN(n6479)
         );
  NAND2_X1 U7989 ( .A1(n6478), .A2(n7654), .ZN(n7695) );
  NOR4_X1 U7990 ( .A1(n4642), .A2(n7652), .A3(n6479), .A4(n7695), .ZN(n6480)
         );
  NAND4_X1 U7991 ( .A1(n8870), .A2(n7858), .A3(n4596), .A4(n6480), .ZN(n6481)
         );
  NOR4_X1 U7992 ( .A1(n8818), .A2(n8834), .A3(n8845), .A4(n6481), .ZN(n6482)
         );
  NAND4_X1 U7993 ( .A1(n8777), .A2(n5002), .A3(n6482), .A4(n8792), .ZN(n6483)
         );
  NOR4_X1 U7994 ( .A1(n8728), .A2(n6483), .A3(n8747), .A4(n8758), .ZN(n6484)
         );
  NAND4_X1 U7995 ( .A1(n7997), .A2(n7996), .A3(n4632), .A4(n6484), .ZN(n6485)
         );
  NOR4_X1 U7996 ( .A1(n6454), .A2(n6486), .A3(n8369), .A4(n6485), .ZN(n6487)
         );
  XNOR2_X1 U7997 ( .A(n6487), .B(n4919), .ZN(n6488) );
  AOI22_X1 U7998 ( .A1(n6488), .A2(n7666), .B1(n4548), .B2(n4455), .ZN(n6489)
         );
  OR2_X1 U7999 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  NAND2_X1 U8000 ( .A1(n6498), .A2(n6497), .ZN(n6811) );
  NOR2_X1 U8001 ( .A1(n6811), .A2(P2_U3152), .ZN(n6510) );
  NAND2_X1 U8002 ( .A1(n6501), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6502) );
  MUX2_X1 U8003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6502), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6503) );
  NAND2_X1 U8004 ( .A1(n6503), .A2(n4543), .ZN(n7929) );
  NAND2_X1 U8005 ( .A1(n4543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6504) );
  MUX2_X1 U8006 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6504), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6506) );
  NAND2_X1 U8007 ( .A1(n6506), .A2(n6505), .ZN(n7949) );
  INV_X1 U8008 ( .A(n6510), .ZN(n7749) );
  OAI21_X1 U8009 ( .B1(n7749), .B2(n4920), .A(P2_B_REG_SCAN_IN), .ZN(n6511) );
  INV_X1 U8010 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U8011 ( .A1(n5069), .A2(n6512), .ZN(n6513) );
  INV_X1 U8012 ( .A(n7744), .ZN(n6515) );
  OR2_X1 U8013 ( .A1(n6644), .A2(n4458), .ZN(n6517) );
  NAND2_X1 U8014 ( .A1(n6517), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8015 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7686) );
  INV_X1 U8016 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9785) );
  INV_X1 U8017 ( .A(n10100), .ZN(n6581) );
  AOI22_X1 U8018 ( .A1(n10100), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9785), .B2(
        n6581), .ZN(n10104) );
  NOR2_X1 U8019 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6617), .ZN(n6518) );
  AOI21_X1 U8020 ( .B1(n6617), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6518), .ZN(
        n6615) );
  INV_X1 U8021 ( .A(n6553), .ZN(n10056) );
  NAND2_X1 U8022 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10076) );
  INV_X1 U8023 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6519) );
  INV_X1 U8024 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6520) );
  MUX2_X1 U8025 ( .A(n6520), .B(P1_REG2_REG_2__SCAN_IN), .S(n6531), .Z(n10067)
         );
  NOR2_X1 U8026 ( .A1(n10066), .A2(n10067), .ZN(n10065) );
  AOI21_X1 U8027 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6531), .A(n10065), .ZN(
        n9897) );
  NAND2_X1 U8028 ( .A1(n9895), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6521) );
  OAI21_X1 U8029 ( .B1(n9895), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6521), .ZN(
        n9898) );
  NOR2_X1 U8030 ( .A1(n9897), .A2(n9898), .ZN(n9896) );
  XNOR2_X1 U8031 ( .A(n10086), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10087) );
  INV_X1 U8032 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6522) );
  AND2_X1 U8033 ( .A1(n10086), .A2(n6522), .ZN(n6523) );
  AOI21_X1 U8034 ( .B1(n10088), .B2(n10087), .A(n6523), .ZN(n6681) );
  INV_X1 U8035 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10209) );
  MUX2_X1 U8036 ( .A(n10209), .B(P1_REG2_REG_5__SCAN_IN), .S(n6688), .Z(n6682)
         );
  NAND2_X1 U8037 ( .A1(n6636), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6524) );
  OAI21_X1 U8038 ( .B1(n6636), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6524), .ZN(
        n6632) );
  INV_X1 U8039 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7535) );
  XNOR2_X1 U8040 ( .A(n6654), .B(n7535), .ZN(n6525) );
  OR2_X1 U8041 ( .A1(n8349), .A2(P1_U3084), .ZN(n7951) );
  NOR2_X1 U8042 ( .A1(n6644), .A2(n7951), .ZN(n9225) );
  OAI21_X1 U8043 ( .B1(n6526), .B2(n6525), .A(n10106), .ZN(n6527) );
  NOR2_X1 U8044 ( .A1(n6527), .A2(n6650), .ZN(n6550) );
  NAND2_X1 U8045 ( .A1(n10100), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6540) );
  INV_X1 U8046 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8047 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6528), .S(n10100), .Z(n10109) );
  NOR2_X1 U8048 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6617), .ZN(n6539) );
  NOR2_X1 U8049 ( .A1(n6636), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8050 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6688), .ZN(n6536) );
  INV_X1 U8051 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6529) );
  MUX2_X1 U8052 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6529), .S(n6688), .Z(n6684)
         );
  INV_X1 U8053 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6535) );
  MUX2_X1 U8054 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6535), .S(n10086), .Z(n10092) );
  NAND2_X1 U8055 ( .A1(n9895), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6534) );
  INV_X1 U8056 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8057 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6530), .S(n9895), .Z(n9901)
         );
  INV_X1 U8058 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10274) );
  MUX2_X1 U8059 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10274), .S(n6531), .Z(n10070) );
  OR2_X1 U8060 ( .A1(n6553), .A2(n6532), .ZN(n6533) );
  MUX2_X1 U8061 ( .A(n6532), .B(P1_REG1_REG_1__SCAN_IN), .S(n6553), .Z(n10060)
         );
  NAND3_X1 U8062 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n10060), .ZN(n10059) );
  NAND2_X1 U8063 ( .A1(n6533), .A2(n10059), .ZN(n10069) );
  NAND2_X1 U8064 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  OAI21_X1 U8065 ( .B1(n10073), .B2(n10274), .A(n10068), .ZN(n9902) );
  NAND2_X1 U8066 ( .A1(n9901), .A2(n9902), .ZN(n9900) );
  NAND2_X1 U8067 ( .A1(n6534), .A2(n9900), .ZN(n10093) );
  NOR2_X1 U8068 ( .A1(n10092), .A2(n10093), .ZN(n10091) );
  AOI21_X1 U8069 ( .B1(n10086), .B2(n6535), .A(n10091), .ZN(n6685) );
  NAND2_X1 U8070 ( .A1(n6684), .A2(n6685), .ZN(n6683) );
  NAND2_X1 U8071 ( .A1(n6536), .A2(n6683), .ZN(n6627) );
  INV_X1 U8072 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8073 ( .A(n6537), .B(P1_REG1_REG_6__SCAN_IN), .S(n6636), .Z(n6626)
         );
  NOR2_X1 U8074 ( .A1(n6627), .A2(n6626), .ZN(n6625) );
  NOR2_X1 U8075 ( .A1(n6538), .A2(n6625), .ZN(n6612) );
  INV_X1 U8076 ( .A(n6617), .ZN(n6577) );
  INV_X1 U8077 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7526) );
  AOI22_X1 U8078 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6577), .B1(n6617), .B2(
        n7526), .ZN(n6611) );
  NOR2_X1 U8079 ( .A1(n6612), .A2(n6611), .ZN(n6610) );
  NOR2_X1 U8080 ( .A1(n6539), .A2(n6610), .ZN(n10110) );
  NAND2_X1 U8081 ( .A1(n10109), .A2(n10110), .ZN(n10108) );
  NAND2_X1 U8082 ( .A1(n6540), .A2(n10108), .ZN(n6543) );
  INV_X1 U8083 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6541) );
  MUX2_X1 U8084 ( .A(n6541), .B(P1_REG1_REG_9__SCAN_IN), .S(n6654), .Z(n6542)
         );
  NOR2_X1 U8085 ( .A1(n6543), .A2(n6542), .ZN(n6655) );
  AOI21_X1 U8086 ( .B1(n6543), .B2(n6542), .A(n6655), .ZN(n6545) );
  NOR2_X1 U8087 ( .A1(n5886), .A2(P1_U3084), .ZN(n9891) );
  NAND2_X1 U8088 ( .A1(n9891), .A2(n8349), .ZN(n6544) );
  NOR2_X1 U8089 ( .A1(n6545), .A2(n10190), .ZN(n6549) );
  INV_X1 U8090 ( .A(n6546), .ZN(n6547) );
  NOR2_X1 U8091 ( .A1(P1_U3083), .A2(n6547), .ZN(n10101) );
  INV_X1 U8092 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10410) );
  INV_X1 U8093 ( .A(n6654), .ZN(n6591) );
  NAND2_X1 U8094 ( .A1(n9225), .A2(n5886), .ZN(n10074) );
  OAI22_X1 U8095 ( .A1(n10193), .A2(n10410), .B1(n6591), .B2(n10074), .ZN(
        n6548) );
  OR4_X1 U8096 ( .A1(n7686), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(P1_U3250)
         );
  OR2_X1 U8097 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_U3084), .ZN(n6639) );
  OAI21_X1 U8098 ( .B1(n6551), .B2(P1_STATE_REG_SCAN_IN), .A(n6639), .ZN(n6552) );
  INV_X1 U8099 ( .A(n6552), .ZN(P1_U3353) );
  NAND2_X2 U8100 ( .A1(n6555), .A2(P1_U3084), .ZN(n9890) );
  OAI222_X1 U8101 ( .A1(n9890), .A2(n6554), .B1(n4459), .B2(n6558), .C1(
        P1_U3084), .C2(n6553), .ZN(P1_U3352) );
  OAI222_X1 U8102 ( .A1(n9890), .A2(n9798), .B1(n4459), .B2(n6559), .C1(
        P1_U3084), .C2(n10073), .ZN(P1_U3351) );
  NAND2_X2 U8103 ( .A1(n6555), .A2(P2_U3152), .ZN(n8454) );
  AND2_X1 U8104 ( .A1(n6556), .A2(P2_U3152), .ZN(n6989) );
  INV_X2 U8105 ( .A(n6989), .ZN(n9018) );
  OAI222_X1 U8106 ( .A1(P2_U3152), .A2(n9917), .B1(n8454), .B2(n6558), .C1(
        n6557), .C2(n9018), .ZN(P2_U3357) );
  OAI222_X1 U8107 ( .A1(n9018), .A2(n6560), .B1(n8454), .B2(n6559), .C1(
        P2_U3152), .C2(n6912), .ZN(P2_U3356) );
  OAI222_X1 U8108 ( .A1(n9890), .A2(n6561), .B1(n4459), .B2(n6562), .C1(
        P1_U3084), .C2(n10086), .ZN(P1_U3349) );
  OAI222_X1 U8109 ( .A1(n9018), .A2(n9741), .B1(n8454), .B2(n6562), .C1(
        P2_U3152), .C2(n6916), .ZN(P2_U3354) );
  OAI222_X1 U8110 ( .A1(n9890), .A2(n6564), .B1(n4459), .B2(n6567), .C1(
        P1_U3084), .C2(n6563), .ZN(P1_U3350) );
  OAI222_X1 U8111 ( .A1(n9890), .A2(n6566), .B1(n4459), .B2(n6569), .C1(
        P1_U3084), .C2(n6565), .ZN(P1_U3348) );
  INV_X1 U8112 ( .A(n8454), .ZN(n7747) );
  OAI222_X1 U8113 ( .A1(n9018), .A2(n6568), .B1(n8454), .B2(n6567), .C1(
        P2_U3152), .C2(n7096), .ZN(P2_U3355) );
  OAI222_X1 U8114 ( .A1(n9018), .A2(n6570), .B1(n8454), .B2(n6569), .C1(
        P2_U3152), .C2(n7077), .ZN(P2_U3353) );
  INV_X1 U8115 ( .A(n6571), .ZN(n6573) );
  INV_X1 U8116 ( .A(n9890), .ZN(n9892) );
  AOI22_X1 U8117 ( .A1(n6636), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9892), .ZN(n6572) );
  OAI21_X1 U8118 ( .B1(n6573), .B2(n4459), .A(n6572), .ZN(P1_U3347) );
  INV_X1 U8119 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6574) );
  INV_X1 U8120 ( .A(n7108), .ZN(n7083) );
  OAI222_X1 U8121 ( .A1(n9018), .A2(n6574), .B1(n8454), .B2(n6573), .C1(
        P2_U3152), .C2(n7083), .ZN(P2_U3352) );
  INV_X1 U8122 ( .A(n6575), .ZN(n6578) );
  AOI22_X1 U8123 ( .A1(n7234), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n6989), .ZN(n6576) );
  OAI21_X1 U8124 ( .B1(n6578), .B2(n8454), .A(n6576), .ZN(P2_U3351) );
  INV_X1 U8125 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9815) );
  OAI222_X1 U8126 ( .A1(n9890), .A2(n9815), .B1(n4459), .B2(n6578), .C1(
        P1_U3084), .C2(n6577), .ZN(P1_U3346) );
  INV_X1 U8127 ( .A(n6579), .ZN(n6582) );
  INV_X1 U8128 ( .A(n8587), .ZN(n7112) );
  OAI222_X1 U8129 ( .A1(n9018), .A2(n6580), .B1(n8454), .B2(n6582), .C1(
        P2_U3152), .C2(n7112), .ZN(P2_U3350) );
  OAI222_X1 U8130 ( .A1(n9890), .A2(n6583), .B1(n4459), .B2(n6582), .C1(
        P1_U3084), .C2(n6581), .ZN(P1_U3345) );
  INV_X1 U8131 ( .A(n10293), .ZN(n6805) );
  NAND2_X1 U8132 ( .A1(n6805), .A2(n6895), .ZN(n6587) );
  NAND2_X1 U8133 ( .A1(n10293), .A2(n7749), .ZN(n6585) );
  NAND2_X1 U8134 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  AND2_X1 U8135 ( .A1(n6587), .A2(n6586), .ZN(n9913) );
  NOR2_X1 U8136 ( .A1(n10287), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8137 ( .A(n6588), .ZN(n6590) );
  INV_X1 U8138 ( .A(n8602), .ZN(n7114) );
  OAI222_X1 U8139 ( .A1(n9018), .A2(n6589), .B1(n8454), .B2(n6590), .C1(n7114), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8140 ( .A1(P1_U3084), .A2(n6591), .B1(n4459), .B2(n6590), .C1(
        n9748), .C2(n9890), .ZN(P1_U3344) );
  INV_X1 U8141 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6594) );
  INV_X1 U8142 ( .A(n8685), .ZN(n6592) );
  NAND2_X1 U8143 ( .A1(n6592), .A2(P2_U3966), .ZN(n6593) );
  OAI21_X1 U8144 ( .B1(n6594), .B2(P2_U3966), .A(n6593), .ZN(P2_U3583) );
  INV_X1 U8145 ( .A(n6595), .ZN(n6608) );
  AOI22_X1 U8146 ( .A1(n6765), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9892), .ZN(n6596) );
  OAI21_X1 U8147 ( .B1(n6608), .B2(n4459), .A(n6596), .ZN(P1_U3342) );
  INV_X1 U8148 ( .A(n6597), .ZN(n6599) );
  INV_X1 U8149 ( .A(n6702), .ZN(n6695) );
  OAI222_X1 U8150 ( .A1(n9890), .A2(n6598), .B1(n4459), .B2(n6599), .C1(n6695), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8151 ( .A(n7151), .ZN(n7156) );
  OAI222_X1 U8152 ( .A1(n9018), .A2(n9602), .B1(n8454), .B2(n6599), .C1(n7156), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  CLKBUF_X2 U8153 ( .A(P1_U4006), .Z(n10079) );
  NAND2_X1 U8154 ( .A1(n8046), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U8155 ( .A1(n6600), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8156 ( .A1(n6601), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6602) );
  NAND3_X1 U8157 ( .A1(n6604), .A2(n6603), .A3(n6602), .ZN(n8173) );
  NAND2_X1 U8158 ( .A1(n8173), .A2(n10079), .ZN(n6605) );
  OAI21_X1 U8159 ( .B1(n10079), .B2(n9013), .A(n6605), .ZN(P1_U3586) );
  NAND2_X1 U8160 ( .A1(n6606), .A2(n10079), .ZN(n6607) );
  OAI21_X1 U8161 ( .B1(n10079), .B2(n5944), .A(n6607), .ZN(P1_U3555) );
  OAI222_X1 U8162 ( .A1(n9018), .A2(n6609), .B1(n8454), .B2(n6608), .C1(n7174), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  AOI21_X1 U8163 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(n6620) );
  OAI21_X1 U8164 ( .B1(n6615), .B2(n6614), .A(n6613), .ZN(n6616) );
  AOI22_X1 U8165 ( .A1(n10106), .A2(n6616), .B1(n10101), .B2(
        P1_ADDR_REG_7__SCAN_IN), .ZN(n6619) );
  AND2_X1 U8166 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7318) );
  AOI21_X1 U8167 ( .B1(n10184), .B2(n6617), .A(n7318), .ZN(n6618) );
  OAI211_X1 U8168 ( .C1(n6620), .C2(n10190), .A(n6619), .B(n6618), .ZN(
        P1_U3248) );
  INV_X1 U8169 ( .A(n6621), .ZN(n6623) );
  INV_X1 U8170 ( .A(n7206), .ZN(n7166) );
  OAI222_X1 U8171 ( .A1(n9018), .A2(n6622), .B1(n8454), .B2(n6623), .C1(
        P2_U3152), .C2(n7166), .ZN(P2_U3346) );
  INV_X1 U8172 ( .A(n6774), .ZN(n9203) );
  OAI222_X1 U8173 ( .A1(n9890), .A2(n6624), .B1(n4459), .B2(n6623), .C1(
        P1_U3084), .C2(n9203), .ZN(P1_U3341) );
  INV_X1 U8174 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6638) );
  AOI21_X1 U8175 ( .B1(n6627), .B2(n6626), .A(n6625), .ZN(n6630) );
  NOR2_X1 U8176 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6628), .ZN(n7220) );
  INV_X1 U8177 ( .A(n7220), .ZN(n6629) );
  OAI21_X1 U8178 ( .B1(n10190), .B2(n6630), .A(n6629), .ZN(n6635) );
  AOI211_X1 U8179 ( .C1(n6633), .C2(n6632), .A(n6631), .B(n10178), .ZN(n6634)
         );
  AOI211_X1 U8180 ( .C1(n10184), .C2(n6636), .A(n6635), .B(n6634), .ZN(n6637)
         );
  OAI21_X1 U8181 ( .B1(n10193), .B2(n6638), .A(n6637), .ZN(P1_U3247) );
  INV_X1 U8182 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6648) );
  INV_X1 U8183 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10057) );
  AOI21_X1 U8184 ( .B1(n8349), .B2(n10057), .A(n6639), .ZN(n6642) );
  OAI21_X1 U8185 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n8349), .A(n6842), .ZN(
        n6641) );
  OAI21_X1 U8186 ( .B1(P1_U3084), .B2(n10058), .A(n6641), .ZN(n10078) );
  OAI211_X1 U8187 ( .C1(n6642), .C2(n6641), .A(n10078), .B(n6640), .ZN(n6643)
         );
  NOR2_X1 U8188 ( .A1(n6644), .A2(n6643), .ZN(n6645) );
  AOI21_X1 U8189 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6645), .ZN(
        n6647) );
  NAND3_X1 U8190 ( .A1(n10172), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10057), .ZN(
        n6646) );
  OAI211_X1 U8191 ( .C1(n10193), .C2(n6648), .A(n6647), .B(n6646), .ZN(
        P1_U3241) );
  INV_X1 U8192 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6669) );
  INV_X1 U8193 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9791) );
  NOR2_X1 U8194 ( .A1(n6702), .A2(n9791), .ZN(n6649) );
  AOI21_X1 U8195 ( .B1(n9791), .B2(n6702), .A(n6649), .ZN(n6652) );
  AOI211_X1 U8196 ( .C1(n6652), .C2(n6651), .A(n10178), .B(n6701), .ZN(n6653)
         );
  INV_X1 U8197 ( .A(n6653), .ZN(n6668) );
  OR2_X1 U8198 ( .A1(n6654), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6657) );
  INV_X1 U8199 ( .A(n6655), .ZN(n6656) );
  AND2_X1 U8200 ( .A1(n6657), .A2(n6656), .ZN(n6662) );
  INV_X1 U8201 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6658) );
  OR2_X1 U8202 ( .A1(n6702), .A2(n6658), .ZN(n6660) );
  NAND2_X1 U8203 ( .A1(n6702), .A2(n6658), .ZN(n6659) );
  AND2_X1 U8204 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  NOR2_X1 U8205 ( .A1(n6662), .A2(n6661), .ZN(n6694) );
  AOI21_X1 U8206 ( .B1(n6662), .B2(n6661), .A(n6694), .ZN(n6665) );
  NOR2_X1 U8207 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6663), .ZN(n7674) );
  INV_X1 U8208 ( .A(n7674), .ZN(n6664) );
  OAI21_X1 U8209 ( .B1(n10190), .B2(n6665), .A(n6664), .ZN(n6666) );
  AOI21_X1 U8210 ( .B1(n10184), .B2(n6702), .A(n6666), .ZN(n6667) );
  OAI211_X1 U8211 ( .C1(n10193), .C2(n6669), .A(n6668), .B(n6667), .ZN(
        P1_U3251) );
  XNOR2_X1 U8212 ( .A(n6670), .B(n6671), .ZN(n6673) );
  XNOR2_X1 U8213 ( .A(n6673), .B(n6672), .ZN(n6679) );
  AOI22_X1 U8214 ( .A1(n9162), .A2(n6606), .B1(n9138), .B2(n9188), .ZN(n6678)
         );
  NAND2_X1 U8215 ( .A1(n7042), .A2(n10234), .ZN(n6830) );
  INV_X1 U8216 ( .A(n6830), .ZN(n6675) );
  OAI211_X1 U8217 ( .C1(n9511), .C2(n6676), .A(n6675), .B(n6674), .ZN(n8074)
         );
  AOI22_X1 U8218 ( .A1(n9168), .A2(n8305), .B1(n8074), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6677) );
  OAI211_X1 U8219 ( .C1(n6679), .C2(n9172), .A(n6678), .B(n6677), .ZN(P1_U3220) );
  AOI21_X1 U8220 ( .B1(n6682), .B2(n6681), .A(n6680), .ZN(n6691) );
  AND2_X1 U8221 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7147) );
  OAI211_X1 U8222 ( .C1(n6685), .C2(n6684), .A(n10172), .B(n6683), .ZN(n6686)
         );
  INV_X1 U8223 ( .A(n6686), .ZN(n6687) );
  AOI211_X1 U8224 ( .C1(n10184), .C2(n6688), .A(n7147), .B(n6687), .ZN(n6690)
         );
  NAND2_X1 U8225 ( .A1(n10101), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6689) );
  OAI211_X1 U8226 ( .C1(n6691), .C2(n10178), .A(n6690), .B(n6689), .ZN(
        P1_U3246) );
  NAND2_X1 U8227 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8568), .ZN(n6692) );
  OAI21_X1 U8228 ( .B1(n8372), .B2(n8568), .A(n6692), .ZN(P2_U3582) );
  INV_X1 U8229 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6708) );
  AND2_X1 U8230 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7774) );
  INV_X1 U8231 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U8232 ( .A1(n6765), .A2(n10042), .ZN(n6693) );
  AOI21_X1 U8233 ( .B1(n6765), .B2(n10042), .A(n6693), .ZN(n6697) );
  AOI21_X1 U8234 ( .B1(n6695), .B2(n6658), .A(n6694), .ZN(n6696) );
  NOR2_X1 U8235 ( .A1(n6697), .A2(n6696), .ZN(n6766) );
  AOI21_X1 U8236 ( .B1(n6697), .B2(n6696), .A(n6766), .ZN(n6698) );
  NOR2_X1 U8237 ( .A1(n10190), .A2(n6698), .ZN(n6699) );
  AOI211_X1 U8238 ( .C1(n10184), .C2(n6765), .A(n7774), .B(n6699), .ZN(n6707)
         );
  OR2_X1 U8239 ( .A1(n6765), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U8240 ( .A1(n6765), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6700) );
  AND2_X1 U8241 ( .A1(n6772), .A2(n6700), .ZN(n6704) );
  OAI21_X1 U8242 ( .B1(n6704), .B2(n6703), .A(n6773), .ZN(n6705) );
  NAND2_X1 U8243 ( .A1(n10106), .A2(n6705), .ZN(n6706) );
  OAI211_X1 U8244 ( .C1(n6708), .C2(n10193), .A(n6707), .B(n6706), .ZN(
        P1_U3252) );
  INV_X1 U8245 ( .A(n6709), .ZN(n6717) );
  AOI22_X1 U8246 ( .A1(n10120), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9892), .ZN(n6710) );
  OAI21_X1 U8247 ( .B1(n6717), .B2(n4459), .A(n6710), .ZN(P1_U3340) );
  NAND2_X1 U8248 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8568), .ZN(n6711) );
  OAI21_X1 U8249 ( .B1(n8444), .B2(n8568), .A(n6711), .ZN(P2_U3581) );
  AOI21_X1 U8250 ( .B1(n6713), .B2(n6712), .A(n4549), .ZN(n6716) );
  AOI22_X1 U8251 ( .A1(n9162), .A2(n6837), .B1(n9138), .B2(n9187), .ZN(n6715)
         );
  AOI22_X1 U8252 ( .A1(n9168), .A2(n8308), .B1(n8074), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6714) );
  OAI211_X1 U8253 ( .C1(n6716), .C2(n9172), .A(n6715), .B(n6714), .ZN(P1_U3235) );
  INV_X1 U8254 ( .A(n7295), .ZN(n7300) );
  OAI222_X1 U8255 ( .A1(n9018), .A2(n6718), .B1(n8454), .B2(n6717), .C1(n7300), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8256 ( .A(n6719), .ZN(n6721) );
  OAI222_X1 U8257 ( .A1(n9890), .A2(n6720), .B1(n4459), .B2(n6721), .C1(n9210), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8258 ( .A(n7574), .ZN(n7577) );
  OAI222_X1 U8259 ( .A1(n9018), .A2(n6722), .B1(n8454), .B2(n6721), .C1(n7577), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NOR4_X1 U8260 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6726) );
  NOR4_X1 U8261 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6725) );
  NOR4_X1 U8262 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6724) );
  NOR4_X1 U8263 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6723) );
  NAND4_X1 U8264 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6735)
         );
  NOR2_X1 U8265 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .ZN(
        n6730) );
  NOR4_X1 U8266 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6729) );
  NOR4_X1 U8267 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6728) );
  NOR4_X1 U8268 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6727) );
  NAND4_X1 U8269 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6734)
         );
  INV_X1 U8270 ( .A(n7949), .ZN(n6733) );
  XNOR2_X1 U8271 ( .A(n7825), .B(P2_B_REG_SCAN_IN), .ZN(n6731) );
  NAND2_X1 U8272 ( .A1(n7929), .A2(n6731), .ZN(n6732) );
  OAI21_X1 U8273 ( .B1(n6735), .B2(n6734), .A(n10292), .ZN(n6783) );
  NAND2_X1 U8274 ( .A1(n6798), .A2(n6895), .ZN(n6810) );
  INV_X1 U8275 ( .A(n6810), .ZN(n6736) );
  NOR2_X1 U8276 ( .A1(n10293), .A2(n6736), .ZN(n6737) );
  AND2_X1 U8277 ( .A1(n7825), .A2(n7949), .ZN(n10301) );
  INV_X1 U8278 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10300) );
  AND2_X1 U8279 ( .A1(n10292), .A2(n10300), .ZN(n6738) );
  NAND2_X1 U8280 ( .A1(n10292), .A2(n10304), .ZN(n6739) );
  NAND2_X1 U8281 ( .A1(n7949), .A2(n7929), .ZN(n10302) );
  NAND2_X1 U8282 ( .A1(n6739), .A2(n10302), .ZN(n6781) );
  NAND2_X1 U8283 ( .A1(n6317), .A2(n10307), .ZN(n7437) );
  NAND2_X1 U8284 ( .A1(n7023), .A2(n6741), .ZN(n6742) );
  NAND2_X1 U8285 ( .A1(n7436), .A2(n6742), .ZN(n7285) );
  NAND2_X1 U8286 ( .A1(n6743), .A2(n4457), .ZN(n6744) );
  INV_X1 U8287 ( .A(n6753), .ZN(n6745) );
  OAI21_X1 U8288 ( .B1(n6746), .B2(n6745), .A(n6929), .ZN(n7273) );
  INV_X1 U8289 ( .A(n7273), .ZN(n6763) );
  AND2_X1 U8290 ( .A1(n6784), .A2(n4919), .ZN(n6750) );
  NAND2_X1 U8291 ( .A1(n7270), .A2(n6463), .ZN(n6749) );
  NAND2_X1 U8292 ( .A1(n6750), .A2(n6749), .ZN(n8881) );
  NAND2_X1 U8293 ( .A1(n4460), .A2(n6463), .ZN(n6751) );
  XNOR2_X1 U8294 ( .A(n6753), .B(n6752), .ZN(n6755) );
  NAND2_X1 U8295 ( .A1(n6755), .A2(n8878), .ZN(n6759) );
  INV_X1 U8296 ( .A(n6509), .ZN(n6757) );
  AOI22_X1 U8297 ( .A1(n8871), .A2(n6756), .B1(n8567), .B2(n8873), .ZN(n6758)
         );
  NAND2_X1 U8298 ( .A1(n6759), .A2(n6758), .ZN(n7264) );
  INV_X1 U8299 ( .A(n7264), .ZN(n6762) );
  NAND2_X1 U8300 ( .A1(n6741), .A2(n7443), .ZN(n7442) );
  AND2_X1 U8301 ( .A1(n7280), .A2(n6947), .ZN(n6760) );
  NOR2_X1 U8302 ( .A1(n7381), .A2(n6760), .ZN(n7269) );
  AOI22_X1 U8303 ( .A1(n7269), .A2(n8985), .B1(n9980), .B2(n6947), .ZN(n6761)
         );
  OAI211_X1 U8304 ( .C1(n6763), .C2(n8981), .A(n6762), .B(n6761), .ZN(n9011)
         );
  NAND2_X1 U8305 ( .A1(n9011), .A2(n10370), .ZN(n6764) );
  OAI21_X1 U8306 ( .B1(n10370), .B2(n6897), .A(n6764), .ZN(P2_U3523) );
  INV_X1 U8307 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6780) );
  INV_X1 U8308 ( .A(n6765), .ZN(n6767) );
  AOI21_X1 U8309 ( .B1(n10042), .B2(n6767), .A(n6766), .ZN(n6769) );
  INV_X1 U8310 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9202) );
  AOI22_X1 U8311 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9203), .B1(n6774), .B2(
        n9202), .ZN(n6768) );
  NOR2_X1 U8312 ( .A1(n6769), .A2(n6768), .ZN(n9201) );
  AOI21_X1 U8313 ( .B1(n6769), .B2(n6768), .A(n9201), .ZN(n6770) );
  NAND2_X1 U8314 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7889) );
  OAI21_X1 U8315 ( .B1(n10190), .B2(n6770), .A(n7889), .ZN(n6771) );
  AOI21_X1 U8316 ( .B1(n10184), .B2(n6774), .A(n6771), .ZN(n6779) );
  OR2_X1 U8317 ( .A1(n6774), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8318 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6774), .ZN(n9189) );
  AND2_X1 U8319 ( .A1(n6775), .A2(n9189), .ZN(n6776) );
  NAND2_X1 U8320 ( .A1(n6777), .A2(n6776), .ZN(n9190) );
  OAI211_X1 U8321 ( .C1(n6777), .C2(n6776), .A(n10106), .B(n9190), .ZN(n6778)
         );
  OAI211_X1 U8322 ( .C1(n10193), .C2(n6780), .A(n6779), .B(n6778), .ZN(
        P1_U3253) );
  NOR2_X1 U8323 ( .A1(n7032), .A2(n6781), .ZN(n6782) );
  NAND2_X1 U8324 ( .A1(n6783), .A2(n6782), .ZN(n6809) );
  XNOR2_X1 U8325 ( .A(n6815), .B(n6793), .ZN(n6789) );
  INV_X1 U8326 ( .A(n6789), .ZN(n6787) );
  NAND2_X1 U8327 ( .A1(n6786), .A2(n6944), .ZN(n6788) );
  NAND2_X1 U8328 ( .A1(n6787), .A2(n6788), .ZN(n6942) );
  INV_X1 U8329 ( .A(n6788), .ZN(n6790) );
  NAND2_X1 U8330 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  NAND2_X1 U8331 ( .A1(n6317), .A2(n6944), .ZN(n6792) );
  NAND2_X1 U8332 ( .A1(n6792), .A2(n10307), .ZN(n6795) );
  NAND2_X1 U8333 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  NAND2_X1 U8334 ( .A1(n6797), .A2(n6796), .ZN(n6943) );
  OAI21_X1 U8335 ( .B1(n6797), .B2(n6796), .A(n6943), .ZN(n6802) );
  INV_X1 U8336 ( .A(n6798), .ZN(n6799) );
  NAND2_X1 U8337 ( .A1(n6803), .A2(n6799), .ZN(n8546) );
  INV_X1 U8338 ( .A(n8546), .ZN(n7010) );
  NAND2_X1 U8339 ( .A1(n8569), .A2(n8871), .ZN(n6801) );
  NAND2_X1 U8340 ( .A1(n6756), .A2(n8873), .ZN(n6800) );
  NAND2_X1 U8341 ( .A1(n6801), .A2(n6800), .ZN(n7439) );
  AOI22_X1 U8342 ( .A1(n8539), .A2(n6802), .B1(n7010), .B2(n7439), .ZN(n6817)
         );
  INV_X1 U8343 ( .A(n6803), .ZN(n6806) );
  OR2_X1 U8344 ( .A1(n4455), .A2(n6804), .ZN(n7261) );
  INV_X1 U8345 ( .A(n6807), .ZN(n6808) );
  NAND2_X1 U8346 ( .A1(n6809), .A2(n6808), .ZN(n6814) );
  AND3_X1 U8347 ( .A1(n6812), .A2(n6811), .A3(n6810), .ZN(n6813) );
  NAND2_X1 U8348 ( .A1(n6814), .A2(n6813), .ZN(n6967) );
  OR2_X1 U8349 ( .A1(n6967), .A2(P2_U3152), .ZN(n8062) );
  AOI22_X1 U8350 ( .A1(n4453), .A2(n6815), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8062), .ZN(n6816) );
  NAND2_X1 U8351 ( .A1(n6817), .A2(n6816), .ZN(P2_U3224) );
  INV_X1 U8352 ( .A(n6818), .ZN(n6820) );
  NOR3_X1 U8353 ( .A1(n4549), .A2(n6820), .A3(n6819), .ZN(n6823) );
  INV_X1 U8354 ( .A(n6821), .ZN(n6822) );
  OAI21_X1 U8355 ( .B1(n6823), .B2(n6822), .A(n9115), .ZN(n6827) );
  NAND2_X1 U8356 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9905) );
  INV_X1 U8357 ( .A(n9905), .ZN(n6825) );
  INV_X1 U8358 ( .A(n9186), .ZN(n7145) );
  INV_X1 U8359 ( .A(n6886), .ZN(n7047) );
  OAI22_X1 U8360 ( .A1(n9164), .A2(n7145), .B1(n7047), .B2(n9123), .ZN(n6824)
         );
  AOI211_X1 U8361 ( .C1(n9162), .C2(n9188), .A(n6825), .B(n6824), .ZN(n6826)
         );
  OAI211_X1 U8362 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9153), .A(n6827), .B(
        n6826), .ZN(P1_U3216) );
  NAND2_X1 U8363 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8568), .ZN(n6828) );
  OAI21_X1 U8364 ( .B1(n8705), .B2(n8568), .A(n6828), .ZN(P2_U3580) );
  INV_X1 U8365 ( .A(n7039), .ZN(n6829) );
  OAI21_X1 U8366 ( .B1(n9937), .B2(n8304), .A(n6829), .ZN(n6831) );
  NAND2_X1 U8367 ( .A1(n9881), .A2(n6851), .ZN(n6832) );
  INV_X1 U8368 ( .A(n7051), .ZN(n6834) );
  OR2_X1 U8369 ( .A1(n6834), .A2(n6833), .ZN(n6836) );
  NAND3_X1 U8370 ( .A1(n5858), .A2(n8304), .A3(n7043), .ZN(n6835) );
  AND2_X1 U8371 ( .A1(n6836), .A2(n6835), .ZN(n7561) );
  NAND2_X1 U8372 ( .A1(n6606), .A2(n10211), .ZN(n6839) );
  NAND2_X1 U8373 ( .A1(n6839), .A2(n8182), .ZN(n6870) );
  OAI21_X1 U8374 ( .B1(n8182), .B2(n6839), .A(n6870), .ZN(n7353) );
  INV_X1 U8375 ( .A(n7353), .ZN(n6846) );
  OR2_X1 U8376 ( .A1(n5858), .A2(n10200), .ZN(n6841) );
  OR2_X1 U8377 ( .A1(n5859), .A2(n8343), .ZN(n6840) );
  INV_X1 U8378 ( .A(n10211), .ZN(n8072) );
  XNOR2_X1 U8379 ( .A(n6874), .B(n6873), .ZN(n6843) );
  AOI222_X1 U8380 ( .A1(n9985), .A2(n6843), .B1(n9188), .B2(n9990), .C1(n6606), 
        .C2(n9988), .ZN(n7357) );
  AOI211_X1 U8381 ( .C1(n10211), .C2(n8305), .A(n10265), .B(n7965), .ZN(n7358)
         );
  AOI21_X1 U8382 ( .B1(n9511), .B2(n8305), .A(n7358), .ZN(n6845) );
  OAI211_X1 U8383 ( .C1(n10016), .C2(n6846), .A(n7357), .B(n6845), .ZN(n6857)
         );
  NAND2_X1 U8384 ( .A1(n6857), .A2(n4456), .ZN(n6847) );
  OAI21_X1 U8385 ( .B1(n4456), .B2(n6532), .A(n6847), .ZN(P1_U3524) );
  AND2_X1 U8386 ( .A1(n6606), .A2(n8072), .ZN(n8302) );
  OR2_X1 U8387 ( .A1(n8302), .A2(n6873), .ZN(n8183) );
  AND2_X1 U8388 ( .A1(n8350), .A2(n7044), .ZN(n6849) );
  AND2_X1 U8389 ( .A1(n9990), .A2(n6837), .ZN(n6848) );
  AOI21_X1 U8390 ( .B1(n8183), .B2(n6849), .A(n6848), .ZN(n10217) );
  OAI21_X1 U8391 ( .B1(n8072), .B2(n7044), .A(n10217), .ZN(n6854) );
  NAND2_X1 U8392 ( .A1(n6854), .A2(n4456), .ZN(n6850) );
  OAI21_X1 U8393 ( .B1(n4456), .B2(n10057), .A(n6850), .ZN(P1_U3523) );
  INV_X1 U8394 ( .A(n6851), .ZN(n6852) );
  INV_X1 U8395 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8396 ( .A1(n6854), .A2(n10273), .ZN(n6855) );
  OAI21_X1 U8397 ( .B1(n10273), .B2(n6856), .A(n6855), .ZN(P1_U3454) );
  INV_X1 U8398 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8399 ( .A1(n6857), .A2(n10273), .ZN(n6858) );
  OAI21_X1 U8400 ( .B1(n10273), .B2(n6859), .A(n6858), .ZN(P1_U3457) );
  INV_X1 U8401 ( .A(n7459), .ZN(n6867) );
  OAI21_X1 U8402 ( .B1(n6862), .B2(n6861), .A(n6860), .ZN(n6863) );
  NAND2_X1 U8403 ( .A1(n6863), .A2(n9115), .ZN(n6866) );
  AND2_X1 U8404 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10096) );
  INV_X1 U8405 ( .A(n9185), .ZN(n7451) );
  INV_X1 U8406 ( .A(n7460), .ZN(n10241) );
  OAI22_X1 U8407 ( .A1(n9164), .A2(n7451), .B1(n10241), .B2(n9123), .ZN(n6864)
         );
  AOI211_X1 U8408 ( .C1(n9162), .C2(n9187), .A(n10096), .B(n6864), .ZN(n6865)
         );
  OAI211_X1 U8409 ( .C1(n9153), .C2(n6867), .A(n6866), .B(n6865), .ZN(P1_U3228) );
  INV_X1 U8410 ( .A(n8305), .ZN(n6868) );
  NAND2_X1 U8411 ( .A1(n6838), .A2(n6868), .ZN(n6869) );
  NAND2_X1 U8412 ( .A1(n6870), .A2(n6869), .ZN(n7958) );
  NAND2_X1 U8413 ( .A1(n7958), .A2(n8184), .ZN(n7960) );
  INV_X1 U8414 ( .A(n9188), .ZN(n8309) );
  NAND2_X1 U8415 ( .A1(n8309), .A2(n10235), .ZN(n6871) );
  INV_X1 U8416 ( .A(n9187), .ZN(n7452) );
  NAND2_X1 U8417 ( .A1(n7452), .A2(n6886), .ZN(n8312) );
  NAND2_X1 U8418 ( .A1(n9187), .A2(n7047), .ZN(n8181) );
  NAND2_X1 U8419 ( .A1(n8312), .A2(n8181), .ZN(n6879) );
  OAI21_X1 U8420 ( .B1(n6872), .B2(n6879), .A(n6994), .ZN(n7052) );
  INV_X1 U8421 ( .A(n7052), .ZN(n6888) );
  INV_X1 U8422 ( .A(n7561), .ZN(n7961) );
  OAI22_X1 U8423 ( .A1(n8309), .A2(n9423), .B1(n7145), .B2(n9425), .ZN(n6884)
         );
  NAND2_X1 U8424 ( .A1(n6838), .A2(n8305), .ZN(n6875) );
  INV_X1 U8425 ( .A(n8184), .ZN(n6876) );
  NAND2_X1 U8426 ( .A1(n8309), .A2(n8308), .ZN(n8306) );
  NAND2_X1 U8427 ( .A1(n6877), .A2(n8306), .ZN(n6881) );
  INV_X1 U8428 ( .A(n6881), .ZN(n6878) );
  NAND2_X1 U8429 ( .A1(n6878), .A2(n6879), .ZN(n6882) );
  INV_X1 U8430 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U8431 ( .A1(n6881), .A2(n6880), .ZN(n6998) );
  AOI21_X1 U8432 ( .B1(n6882), .B2(n6998), .A(n9421), .ZN(n6883) );
  AOI211_X1 U8433 ( .C1(n7961), .C2(n7052), .A(n6884), .B(n6883), .ZN(n7055)
         );
  INV_X1 U8434 ( .A(n7967), .ZN(n6885) );
  NAND2_X1 U8435 ( .A1(n7967), .A2(n7047), .ZN(n7456) );
  AOI21_X1 U8436 ( .B1(n6886), .B2(n6885), .A(n4805), .ZN(n7050) );
  AOI22_X1 U8437 ( .A1(n7050), .A2(n9999), .B1(n9511), .B2(n6886), .ZN(n6887)
         );
  OAI211_X1 U8438 ( .C1(n6888), .C2(n9937), .A(n7055), .B(n6887), .ZN(n6890)
         );
  NAND2_X1 U8439 ( .A1(n6890), .A2(n4456), .ZN(n6889) );
  OAI21_X1 U8440 ( .B1(n4456), .B2(n6530), .A(n6889), .ZN(P1_U3526) );
  INV_X1 U8441 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8442 ( .A1(n6890), .A2(n10273), .ZN(n6891) );
  OAI21_X1 U8443 ( .B1(n10273), .B2(n6892), .A(n6891), .ZN(P1_U3463) );
  NAND2_X1 U8444 ( .A1(n6893), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6894) );
  OAI211_X1 U8445 ( .C1(n10293), .C2(n6895), .A(n7749), .B(n6894), .ZN(n6904)
         );
  NAND2_X1 U8446 ( .A1(n6904), .A2(n6902), .ZN(n6896) );
  NAND2_X1 U8447 ( .A1(n6896), .A2(n8568), .ZN(n6919) );
  AND2_X1 U8448 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8449 ( .A1(n6913), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6899) );
  MUX2_X1 U8450 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6897), .S(n6913), .Z(n7092)
         );
  INV_X1 U8451 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10362) );
  MUX2_X1 U8452 ( .A(n10362), .B(P2_REG1_REG_2__SCAN_IN), .S(n6912), .Z(n9932)
         );
  MUX2_X1 U8453 ( .A(n6898), .B(P2_REG1_REG_1__SCAN_IN), .S(n9917), .Z(n9920)
         );
  NAND3_X1 U8454 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9920), .ZN(n9919) );
  OAI21_X1 U8455 ( .B1(n9917), .B2(n6898), .A(n9919), .ZN(n9933) );
  NAND2_X1 U8456 ( .A1(n9932), .A2(n9933), .ZN(n9931) );
  OAI21_X1 U8457 ( .B1(n6912), .B2(n10362), .A(n9931), .ZN(n7093) );
  NAND2_X1 U8458 ( .A1(n7092), .A2(n7093), .ZN(n7091) );
  NAND2_X1 U8459 ( .A1(n6899), .A2(n7091), .ZN(n8578) );
  MUX2_X1 U8460 ( .A(n6900), .B(P2_REG1_REG_4__SCAN_IN), .S(n6916), .Z(n8577)
         );
  NAND2_X1 U8461 ( .A1(n8578), .A2(n8577), .ZN(n8576) );
  OAI21_X1 U8462 ( .B1(n6900), .B2(n6916), .A(n8576), .ZN(n6906) );
  MUX2_X1 U8463 ( .A(n6901), .B(P2_REG1_REG_5__SCAN_IN), .S(n7077), .Z(n6905)
         );
  AND2_X1 U8464 ( .A1(n6902), .A2(n6507), .ZN(n6903) );
  NAND2_X1 U8465 ( .A1(n6904), .A2(n6903), .ZN(n10285) );
  NAND2_X1 U8466 ( .A1(n6905), .A2(n6906), .ZN(n7076) );
  OAI211_X1 U8467 ( .C1(n6906), .C2(n6905), .A(n10281), .B(n7076), .ZN(n6907)
         );
  INV_X1 U8468 ( .A(n6907), .ZN(n6908) );
  AOI211_X1 U8469 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10287), .A(n6909), .B(
        n6908), .ZN(n6923) );
  MUX2_X1 U8470 ( .A(n7067), .B(P2_REG2_REG_5__SCAN_IN), .S(n7077), .Z(n6921)
         );
  XNOR2_X1 U8471 ( .A(n6916), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U8472 ( .A1(n6913), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6915) );
  INV_X1 U8473 ( .A(n6912), .ZN(n9929) );
  INV_X1 U8474 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6910) );
  MUX2_X1 U8475 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6910), .S(n9917), .Z(n9909)
         );
  NOR2_X1 U8476 ( .A1(n9917), .A2(n6910), .ZN(n6911) );
  NOR2_X1 U8477 ( .A1(n9907), .A2(n6911), .ZN(n9927) );
  XNOR2_X1 U8478 ( .A(n6912), .B(n9734), .ZN(n9926) );
  NOR2_X1 U8479 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  AOI21_X1 U8480 ( .B1(n9929), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9925), .ZN(
        n7088) );
  OAI21_X1 U8481 ( .B1(n6913), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6915), .ZN(
        n7087) );
  INV_X1 U8482 ( .A(n7086), .ZN(n6914) );
  NAND2_X1 U8483 ( .A1(n6915), .A2(n6914), .ZN(n8572) );
  NAND2_X1 U8484 ( .A1(n8573), .A2(n8572), .ZN(n8571) );
  INV_X1 U8485 ( .A(n6916), .ZN(n8570) );
  NAND2_X1 U8486 ( .A1(n8570), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8487 ( .A1(n8571), .A2(n6917), .ZN(n6920) );
  NOR2_X1 U8488 ( .A1(n6509), .A2(n6507), .ZN(n6918) );
  NAND2_X1 U8489 ( .A1(n6920), .A2(n6921), .ZN(n7069) );
  OAI211_X1 U8490 ( .C1(n6921), .C2(n6920), .A(n10282), .B(n7069), .ZN(n6922)
         );
  OAI211_X1 U8491 ( .C1(n10283), .C2(n7077), .A(n6923), .B(n6922), .ZN(
        P2_U3250) );
  INV_X1 U8492 ( .A(n6924), .ZN(n6926) );
  INV_X1 U8493 ( .A(n8611), .ZN(n8617) );
  OAI222_X1 U8494 ( .A1(n9018), .A2(n6925), .B1(n8454), .B2(n6926), .C1(
        P2_U3152), .C2(n8617), .ZN(P2_U3343) );
  INV_X1 U8495 ( .A(n10146), .ZN(n9212) );
  OAI222_X1 U8496 ( .A1(n9890), .A2(n9637), .B1(n4459), .B2(n6926), .C1(
        P1_U3084), .C2(n9212), .ZN(P1_U3338) );
  NAND2_X1 U8497 ( .A1(n6927), .A2(n7276), .ZN(n6928) );
  INV_X1 U8498 ( .A(n7388), .ZN(n7385) );
  INV_X1 U8499 ( .A(n8567), .ZN(n6975) );
  NAND2_X1 U8500 ( .A1(n6975), .A2(n10323), .ZN(n6930) );
  OAI21_X1 U8501 ( .B1(n6931), .B2(n6936), .A(n7124), .ZN(n7474) );
  INV_X1 U8502 ( .A(n7380), .ZN(n6932) );
  OAI211_X1 U8503 ( .C1(n6932), .C2(n7122), .A(n8985), .B(n7370), .ZN(n7470)
         );
  OAI21_X1 U8504 ( .B1(n7122), .B2(n10348), .A(n7470), .ZN(n6938) );
  NAND2_X1 U8505 ( .A1(n6933), .A2(n6934), .ZN(n6935) );
  XOR2_X1 U8506 ( .A(n6936), .B(n6935), .Z(n6937) );
  AOI22_X1 U8507 ( .A1(n8871), .A2(n8567), .B1(n8565), .B2(n8873), .ZN(n7008)
         );
  OAI21_X1 U8508 ( .B1(n6937), .B2(n8847), .A(n7008), .ZN(n7466) );
  AOI211_X1 U8509 ( .C1(n10354), .C2(n7474), .A(n6938), .B(n7466), .ZN(n7036)
         );
  NAND2_X1 U8510 ( .A1(n10368), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6939) );
  OAI21_X1 U8511 ( .B1(n7036), .B2(n10368), .A(n6939), .ZN(P2_U3525) );
  INV_X1 U8512 ( .A(n6940), .ZN(n6941) );
  INV_X1 U8513 ( .A(n10157), .ZN(n9214) );
  OAI222_X1 U8514 ( .A1(n9890), .A2(n9753), .B1(n4459), .B2(n6941), .C1(n9214), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8515 ( .A(n8631), .ZN(n8624) );
  OAI222_X1 U8516 ( .A1(n9018), .A2(n9781), .B1(n8454), .B2(n6941), .C1(n8624), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  NAND2_X1 U8517 ( .A1(n6943), .A2(n6942), .ZN(n8058) );
  NAND2_X1 U8518 ( .A1(n6756), .A2(n6944), .ZN(n6945) );
  NAND2_X1 U8519 ( .A1(n6946), .A2(n8430), .ZN(n6948) );
  XNOR2_X1 U8520 ( .A(n6947), .B(n8436), .ZN(n6949) );
  XNOR2_X1 U8521 ( .A(n6948), .B(n6949), .ZN(n6973) );
  NAND2_X1 U8522 ( .A1(n6974), .A2(n6973), .ZN(n6952) );
  INV_X1 U8523 ( .A(n6948), .ZN(n6950) );
  NAND2_X1 U8524 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  NAND2_X1 U8525 ( .A1(n6952), .A2(n6951), .ZN(n7018) );
  NAND2_X1 U8526 ( .A1(n8567), .A2(n8430), .ZN(n6955) );
  XNOR2_X1 U8527 ( .A(n8429), .B(n6953), .ZN(n6954) );
  NAND2_X1 U8528 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  OAI21_X1 U8529 ( .B1(n6955), .B2(n6954), .A(n6956), .ZN(n7017) );
  XNOR2_X1 U8530 ( .A(n7468), .B(n8436), .ZN(n6957) );
  INV_X4 U8531 ( .A(n7025), .ZN(n8430) );
  NAND2_X1 U8532 ( .A1(n8566), .A2(n8430), .ZN(n6958) );
  XNOR2_X1 U8533 ( .A(n6957), .B(n6958), .ZN(n7007) );
  INV_X1 U8534 ( .A(n6957), .ZN(n6959) );
  NOR2_X1 U8535 ( .A1(n6959), .A2(n6958), .ZN(n6960) );
  XNOR2_X1 U8536 ( .A(n7132), .B(n8429), .ZN(n6961) );
  NAND2_X1 U8537 ( .A1(n8565), .A2(n8430), .ZN(n6962) );
  NAND2_X1 U8538 ( .A1(n6961), .A2(n6962), .ZN(n6966) );
  INV_X1 U8539 ( .A(n6961), .ZN(n6964) );
  INV_X1 U8540 ( .A(n6962), .ZN(n6963) );
  NAND2_X1 U8541 ( .A1(n6964), .A2(n6963), .ZN(n6965) );
  AND2_X1 U8542 ( .A1(n6966), .A2(n6965), .ZN(n6982) );
  NAND2_X1 U8543 ( .A1(n6980), .A2(n6966), .ZN(n7062) );
  XNOR2_X1 U8544 ( .A(n7323), .B(n8429), .ZN(n7056) );
  NAND2_X1 U8545 ( .A1(n8564), .A2(n8430), .ZN(n7057) );
  XNOR2_X1 U8546 ( .A(n7056), .B(n7057), .ZN(n7061) );
  XNOR2_X1 U8547 ( .A(n7062), .B(n7061), .ZN(n6972) );
  INV_X1 U8548 ( .A(n8531), .ZN(n8061) );
  AND2_X1 U8549 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7235) );
  INV_X1 U8550 ( .A(n7235), .ZN(n6968) );
  OAI21_X1 U8551 ( .B1(n8522), .B2(n7543), .A(n6968), .ZN(n6970) );
  INV_X1 U8552 ( .A(n7323), .ZN(n7545) );
  OAI22_X1 U8553 ( .A1(n8551), .A2(n7545), .B1(n8530), .B2(n7478), .ZN(n6969)
         );
  AOI211_X1 U8554 ( .C1(n8061), .C2(n8565), .A(n6970), .B(n6969), .ZN(n6971)
         );
  OAI21_X1 U8555 ( .B1(n6972), .B2(n8537), .A(n6971), .ZN(P2_U3215) );
  XNOR2_X1 U8556 ( .A(n6974), .B(n6973), .ZN(n6979) );
  MUX2_X1 U8557 ( .A(n8548), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n6977) );
  OAI22_X1 U8558 ( .A1(n8551), .A2(n7276), .B1(n8530), .B2(n6975), .ZN(n6976)
         );
  AOI211_X1 U8559 ( .C1(n8061), .C2(n6756), .A(n6977), .B(n6976), .ZN(n6978)
         );
  OAI21_X1 U8560 ( .B1(n8537), .B2(n6979), .A(n6978), .ZN(P2_U3220) );
  OAI21_X1 U8561 ( .B1(n6982), .B2(n6981), .A(n6980), .ZN(n6986) );
  OAI22_X1 U8562 ( .A1(n8551), .A2(n10329), .B1(n8530), .B2(n7369), .ZN(n6985)
         );
  NAND2_X1 U8563 ( .A1(n8061), .A2(n8566), .ZN(n6983) );
  NAND2_X1 U8564 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7074) );
  OAI211_X1 U8565 ( .C1(n8522), .C2(n7373), .A(n6983), .B(n7074), .ZN(n6984)
         );
  AOI211_X1 U8566 ( .C1(n6986), .C2(n8539), .A(n6985), .B(n6984), .ZN(n6987)
         );
  INV_X1 U8567 ( .A(n6987), .ZN(P2_U3241) );
  INV_X1 U8568 ( .A(n6988), .ZN(n6992) );
  AOI22_X1 U8569 ( .A1(n8659), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6989), .ZN(n6990) );
  OAI21_X1 U8570 ( .B1(n6992), .B2(n8454), .A(n6990), .ZN(P2_U3341) );
  AOI22_X1 U8571 ( .A1(n10170), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9892), .ZN(n6991) );
  OAI21_X1 U8572 ( .B1(n6992), .B2(n4459), .A(n6991), .ZN(P1_U3336) );
  NAND2_X1 U8573 ( .A1(n7452), .A2(n7047), .ZN(n6993) );
  NAND2_X1 U8574 ( .A1(n7145), .A2(n7460), .ZN(n8315) );
  NAND2_X1 U8575 ( .A1(n9186), .A2(n10241), .ZN(n8231) );
  NAND2_X1 U8576 ( .A1(n8315), .A2(n8231), .ZN(n7449) );
  NAND2_X1 U8577 ( .A1(n7145), .A2(n10241), .ZN(n6995) );
  NAND2_X1 U8578 ( .A1(n7451), .A2(n7184), .ZN(n8234) );
  INV_X1 U8579 ( .A(n7184), .ZN(n10197) );
  NAND2_X1 U8580 ( .A1(n9185), .A2(n10197), .ZN(n8232) );
  INV_X1 U8581 ( .A(n8186), .ZN(n6996) );
  OAI21_X1 U8582 ( .B1(n6997), .B2(n6996), .A(n7186), .ZN(n10204) );
  INV_X1 U8583 ( .A(n7449), .ZN(n6999) );
  XNOR2_X1 U8584 ( .A(n7194), .B(n8186), .ZN(n7000) );
  AOI222_X1 U8585 ( .A1(n9985), .A2(n7000), .B1(n9184), .B2(n9990), .C1(n9186), 
        .C2(n9988), .ZN(n10203) );
  AOI21_X1 U8586 ( .B1(n7458), .B2(n7184), .A(n10265), .ZN(n7001) );
  AND2_X1 U8587 ( .A1(n7189), .A2(n7001), .ZN(n10201) );
  AOI21_X1 U8588 ( .B1(n9511), .B2(n7184), .A(n10201), .ZN(n7002) );
  OAI211_X1 U8589 ( .C1(n10016), .C2(n10204), .A(n10203), .B(n7002), .ZN(n7004) );
  NAND2_X1 U8590 ( .A1(n7004), .A2(n4456), .ZN(n7003) );
  OAI21_X1 U8591 ( .B1(n4456), .B2(n6529), .A(n7003), .ZN(P1_U3528) );
  INV_X1 U8592 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U8593 ( .A1(n7004), .A2(n10273), .ZN(n7005) );
  OAI21_X1 U8594 ( .B1(n10273), .B2(n7006), .A(n7005), .ZN(P1_U3469) );
  XNOR2_X1 U8595 ( .A(n4550), .B(n7007), .ZN(n7014) );
  INV_X1 U8596 ( .A(n7008), .ZN(n7009) );
  AOI22_X1 U8597 ( .A1(n7010), .A2(n7009), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7013) );
  INV_X1 U8598 ( .A(n7011), .ZN(n7467) );
  AOI22_X1 U8599 ( .A1(n4453), .A2(n7468), .B1(n8548), .B2(n7467), .ZN(n7012)
         );
  OAI211_X1 U8600 ( .C1(n7014), .C2(n8537), .A(n7013), .B(n7012), .ZN(P2_U3229) );
  INV_X1 U8601 ( .A(n7015), .ZN(n7016) );
  AOI21_X1 U8602 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7022) );
  NAND2_X1 U8603 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8574) );
  OAI21_X1 U8604 ( .B1(n8522), .B2(n7379), .A(n8574), .ZN(n7020) );
  OAI22_X1 U8605 ( .A1(n8551), .A2(n10323), .B1(n8530), .B2(n7368), .ZN(n7019)
         );
  AOI211_X1 U8606 ( .C1(n8061), .C2(n6946), .A(n7020), .B(n7019), .ZN(n7021)
         );
  OAI21_X1 U8607 ( .B1(n7022), .B2(n8537), .A(n7021), .ZN(P2_U3232) );
  INV_X1 U8608 ( .A(n8062), .ZN(n7031) );
  INV_X1 U8609 ( .A(n8530), .ZN(n8060) );
  AOI22_X1 U8610 ( .A1(n8060), .A2(n6786), .B1(n10307), .B2(n4453), .ZN(n7030)
         );
  INV_X1 U8611 ( .A(n6468), .ZN(n7028) );
  INV_X1 U8612 ( .A(n7024), .ZN(n7026) );
  MUX2_X1 U8613 ( .A(n7026), .B(n10307), .S(n7025), .Z(n7027) );
  OAI21_X1 U8614 ( .B1(n7028), .B2(n7027), .A(n8539), .ZN(n7029) );
  OAI211_X1 U8615 ( .C1(n7031), .C2(n7289), .A(n7030), .B(n7029), .ZN(P2_U3234) );
  INV_X1 U8616 ( .A(n7034), .ZN(n7035) );
  INV_X1 U8617 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7038) );
  OR2_X1 U8618 ( .A1(n7036), .A2(n10356), .ZN(n7037) );
  OAI21_X1 U8619 ( .B1(n10358), .B2(n7038), .A(n7037), .ZN(P2_U3466) );
  NAND2_X1 U8620 ( .A1(n7039), .A2(n10234), .ZN(n10232) );
  NOR2_X1 U8621 ( .A1(n7040), .A2(n10232), .ZN(n7041) );
  NAND2_X1 U8622 ( .A1(n7042), .A2(n7041), .ZN(n7418) );
  INV_X1 U8623 ( .A(n7043), .ZN(n8346) );
  NOR2_X1 U8624 ( .A1(n7044), .A2(n8346), .ZN(n7045) );
  INV_X1 U8625 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7046) );
  OAI22_X1 U8626 ( .A1(n10207), .A2(n7046), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10221), .ZN(n7049) );
  NOR2_X1 U8627 ( .A1(n9432), .A2(n7047), .ZN(n7048) );
  AOI211_X1 U8628 ( .C1(n7050), .C2(n10212), .A(n7049), .B(n7048), .ZN(n7054)
         );
  NOR2_X1 U8629 ( .A1(n7051), .A2(n10200), .ZN(n7354) );
  NAND2_X1 U8630 ( .A1(n7052), .A2(n7968), .ZN(n7053) );
  OAI211_X1 U8631 ( .C1(n7055), .C2(n10216), .A(n7054), .B(n7053), .ZN(
        P1_U3288) );
  INV_X1 U8632 ( .A(n7056), .ZN(n7059) );
  INV_X1 U8633 ( .A(n7057), .ZN(n7058) );
  NAND2_X1 U8634 ( .A1(n7059), .A2(n7058), .ZN(n7060) );
  XNOR2_X1 U8635 ( .A(n7479), .B(n8436), .ZN(n7245) );
  NAND2_X1 U8636 ( .A1(n8563), .A2(n8430), .ZN(n7243) );
  XNOR2_X1 U8637 ( .A(n7245), .B(n7243), .ZN(n7241) );
  XNOR2_X1 U8638 ( .A(n7242), .B(n7241), .ZN(n7066) );
  OAI22_X1 U8639 ( .A1(n8522), .A2(n7337), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8588), .ZN(n7064) );
  OAI22_X1 U8640 ( .A1(n7369), .A2(n8531), .B1(n8530), .B2(n7347), .ZN(n7063)
         );
  AOI211_X1 U8641 ( .C1(n7479), .C2(n4453), .A(n7064), .B(n7063), .ZN(n7065)
         );
  OAI21_X1 U8642 ( .B1(n7066), .B2(n8537), .A(n7065), .ZN(P2_U3223) );
  OR2_X1 U8643 ( .A1(n7077), .A2(n7067), .ZN(n7068) );
  AND2_X1 U8644 ( .A1(n7069), .A2(n7068), .ZN(n7073) );
  OR2_X1 U8645 ( .A1(n7108), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U8646 ( .A1(n7108), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7070) );
  NAND2_X1 U8647 ( .A1(n7071), .A2(n7070), .ZN(n7072) );
  AOI211_X1 U8648 ( .C1(n7073), .C2(n7072), .A(n7099), .B(n9924), .ZN(n7085)
         );
  INV_X1 U8649 ( .A(n7074), .ZN(n7075) );
  AOI21_X1 U8650 ( .B1(n10287), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7075), .ZN(
        n7082) );
  OAI21_X1 U8651 ( .B1(n7077), .B2(n6901), .A(n7076), .ZN(n7080) );
  MUX2_X1 U8652 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7078), .S(n7108), .Z(n7079)
         );
  NAND2_X1 U8653 ( .A1(n7079), .A2(n7080), .ZN(n7109) );
  OAI211_X1 U8654 ( .C1(n7080), .C2(n7079), .A(n10281), .B(n7109), .ZN(n7081)
         );
  OAI211_X1 U8655 ( .C1(n10283), .C2(n7083), .A(n7082), .B(n7081), .ZN(n7084)
         );
  OR2_X1 U8656 ( .A1(n7085), .A2(n7084), .ZN(P2_U3251) );
  AOI211_X1 U8657 ( .C1(n7088), .C2(n7087), .A(n7086), .B(n9924), .ZN(n7098)
         );
  INV_X1 U8658 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7089) );
  NOR2_X1 U8659 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7089), .ZN(n7090) );
  AOI21_X1 U8660 ( .B1(n10287), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7090), .ZN(
        n7095) );
  OAI211_X1 U8661 ( .C1(n7093), .C2(n7092), .A(n10281), .B(n7091), .ZN(n7094)
         );
  OAI211_X1 U8662 ( .C1(n10283), .C2(n7096), .A(n7095), .B(n7094), .ZN(n7097)
         );
  OR2_X1 U8663 ( .A1(n7098), .A2(n7097), .ZN(P2_U3248) );
  AOI21_X1 U8664 ( .B1(n7108), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7099), .ZN(
        n7230) );
  NAND2_X1 U8665 ( .A1(n7234), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7100) );
  OAI21_X1 U8666 ( .B1(n7234), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7100), .ZN(
        n7229) );
  NOR2_X1 U8667 ( .A1(n7230), .A2(n7229), .ZN(n7228) );
  AOI21_X1 U8668 ( .B1(n7234), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7228), .ZN(
        n8585) );
  XNOR2_X1 U8669 ( .A(n8587), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n8584) );
  AOI21_X1 U8670 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n8587), .A(n8583), .ZN(
        n8598) );
  NAND2_X1 U8671 ( .A1(n8602), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7101) );
  OAI21_X1 U8672 ( .B1(n8602), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7101), .ZN(
        n8597) );
  AOI21_X1 U8673 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8602), .A(n8596), .ZN(
        n7104) );
  NAND2_X1 U8674 ( .A1(n7151), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7102) );
  OAI21_X1 U8675 ( .B1(n7151), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7102), .ZN(
        n7103) );
  AOI211_X1 U8676 ( .C1(n7104), .C2(n7103), .A(n7150), .B(n9924), .ZN(n7121)
         );
  NOR2_X1 U8677 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7346), .ZN(n7105) );
  AOI21_X1 U8678 ( .B1(n10287), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7105), .ZN(
        n7119) );
  MUX2_X1 U8679 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7106), .S(n8602), .Z(n8604)
         );
  NAND2_X1 U8680 ( .A1(n7234), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7111) );
  MUX2_X1 U8681 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7107), .S(n7234), .Z(n7232)
         );
  NAND2_X1 U8682 ( .A1(n7108), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U8683 ( .A1(n7110), .A2(n7109), .ZN(n7233) );
  NAND2_X1 U8684 ( .A1(n7232), .A2(n7233), .ZN(n7231) );
  NAND2_X1 U8685 ( .A1(n7111), .A2(n7231), .ZN(n8592) );
  MUX2_X1 U8686 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7113), .S(n8587), .Z(n8591)
         );
  NAND2_X1 U8687 ( .A1(n8592), .A2(n8591), .ZN(n8590) );
  OAI21_X1 U8688 ( .B1(n7113), .B2(n7112), .A(n8590), .ZN(n8605) );
  NAND2_X1 U8689 ( .A1(n8604), .A2(n8605), .ZN(n8603) );
  OAI21_X1 U8690 ( .B1(n7114), .B2(n7106), .A(n8603), .ZN(n7117) );
  MUX2_X1 U8691 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7115), .S(n7151), .Z(n7116)
         );
  NAND2_X1 U8692 ( .A1(n7116), .A2(n7117), .ZN(n7155) );
  OAI211_X1 U8693 ( .C1(n7117), .C2(n7116), .A(n10281), .B(n7155), .ZN(n7118)
         );
  OAI211_X1 U8694 ( .C1(n10283), .C2(n7156), .A(n7119), .B(n7118), .ZN(n7120)
         );
  OR2_X1 U8695 ( .A1(n7121), .A2(n7120), .ZN(P2_U3255) );
  INV_X1 U8696 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8697 ( .A1(n7368), .A2(n7122), .ZN(n7123) );
  NAND2_X1 U8698 ( .A1(n7124), .A2(n7123), .ZN(n7364) );
  NAND2_X1 U8699 ( .A1(n7364), .A2(n7366), .ZN(n7363) );
  NAND2_X1 U8700 ( .A1(n7125), .A2(n10329), .ZN(n7126) );
  NAND2_X1 U8701 ( .A1(n7363), .A2(n7126), .ZN(n7487) );
  NAND2_X1 U8702 ( .A1(n7487), .A2(n7480), .ZN(n7324) );
  OAI21_X1 U8703 ( .B1(n7487), .B2(n7480), .A(n7324), .ZN(n7542) );
  INV_X1 U8704 ( .A(n7542), .ZN(n7135) );
  OAI211_X1 U8705 ( .C1(n7127), .C2(n7129), .A(n7128), .B(n8878), .ZN(n7131)
         );
  AOI22_X1 U8706 ( .A1(n8871), .A2(n8565), .B1(n8563), .B2(n8873), .ZN(n7130)
         );
  AND2_X1 U8707 ( .A1(n7131), .A2(n7130), .ZN(n7551) );
  NOR2_X1 U8708 ( .A1(n7370), .A2(n7132), .ZN(n7133) );
  INV_X1 U8709 ( .A(n7133), .ZN(n7371) );
  AOI21_X1 U8710 ( .B1(n7323), .B2(n7371), .A(n7339), .ZN(n7548) );
  AOI22_X1 U8711 ( .A1(n7548), .A2(n8985), .B1(n9980), .B2(n7323), .ZN(n7134)
         );
  OAI211_X1 U8712 ( .C1(n7135), .C2(n8981), .A(n7551), .B(n7134), .ZN(n7138)
         );
  NAND2_X1 U8713 ( .A1(n7138), .A2(n10358), .ZN(n7136) );
  OAI21_X1 U8714 ( .B1(n10358), .B2(n7137), .A(n7136), .ZN(P2_U3472) );
  NAND2_X1 U8715 ( .A1(n7138), .A2(n10370), .ZN(n7139) );
  OAI21_X1 U8716 ( .B1(n10370), .B2(n7107), .A(n7139), .ZN(P2_U3527) );
  INV_X1 U8717 ( .A(n7140), .ZN(n10198) );
  AND2_X1 U8718 ( .A1(n7141), .A2(n7214), .ZN(n7142) );
  OAI21_X1 U8719 ( .B1(n7143), .B2(n7142), .A(n7218), .ZN(n7144) );
  NAND2_X1 U8720 ( .A1(n7144), .A2(n9115), .ZN(n7149) );
  INV_X1 U8721 ( .A(n9162), .ZN(n9141) );
  OAI22_X1 U8722 ( .A1(n9141), .A2(n7145), .B1(n10197), .B2(n9123), .ZN(n7146)
         );
  AOI211_X1 U8723 ( .C1(n9138), .C2(n9184), .A(n7147), .B(n7146), .ZN(n7148)
         );
  OAI211_X1 U8724 ( .C1(n9153), .C2(n10198), .A(n7149), .B(n7148), .ZN(
        P1_U3225) );
  MUX2_X1 U8725 ( .A(n7173), .B(P2_REG2_REG_11__SCAN_IN), .S(n7174), .Z(n7153)
         );
  NAND2_X1 U8726 ( .A1(n7152), .A2(n7153), .ZN(n7175) );
  OAI21_X1 U8727 ( .B1(n7153), .B2(n7152), .A(n7175), .ZN(n7163) );
  NOR2_X1 U8728 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6066), .ZN(n7154) );
  AOI21_X1 U8729 ( .B1(n10287), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7154), .ZN(
        n7161) );
  OAI21_X1 U8730 ( .B1(n7156), .B2(n7115), .A(n7155), .ZN(n7159) );
  MUX2_X1 U8731 ( .A(n7157), .B(P2_REG1_REG_11__SCAN_IN), .S(n7174), .Z(n7158)
         );
  NAND2_X1 U8732 ( .A1(n7158), .A2(n7159), .ZN(n7165) );
  OAI211_X1 U8733 ( .C1(n7159), .C2(n7158), .A(n10281), .B(n7165), .ZN(n7160)
         );
  OAI211_X1 U8734 ( .C1(n10283), .C2(n7174), .A(n7161), .B(n7160), .ZN(n7162)
         );
  AOI21_X1 U8735 ( .B1(n10282), .B2(n7163), .A(n7162), .ZN(n7164) );
  INV_X1 U8736 ( .A(n7164), .ZN(P2_U3256) );
  OAI21_X1 U8737 ( .B1(n7157), .B2(n7174), .A(n7165), .ZN(n7204) );
  AOI22_X1 U8738 ( .A1(n7206), .A2(n6076), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7166), .ZN(n7203) );
  NOR2_X1 U8739 ( .A1(n7204), .A2(n7203), .ZN(n7202) );
  NOR2_X1 U8740 ( .A1(n7206), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7167) );
  NOR2_X1 U8741 ( .A1(n7202), .A2(n7167), .ZN(n7169) );
  XNOR2_X1 U8742 ( .A(n7295), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n7168) );
  NOR2_X1 U8743 ( .A1(n7169), .A2(n7168), .ZN(n7299) );
  AOI21_X1 U8744 ( .B1(n7169), .B2(n7168), .A(n7299), .ZN(n7183) );
  OR2_X1 U8745 ( .A1(n7295), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8746 ( .A1(n7295), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7170) );
  AND2_X1 U8747 ( .A1(n7171), .A2(n7170), .ZN(n7178) );
  NAND2_X1 U8748 ( .A1(n7206), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7172) );
  OAI21_X1 U8749 ( .B1(n7206), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7172), .ZN(
        n7208) );
  NAND2_X1 U8750 ( .A1(n7174), .A2(n7173), .ZN(n7176) );
  NAND2_X1 U8751 ( .A1(n7176), .A2(n7175), .ZN(n7209) );
  AOI21_X1 U8752 ( .B1(n7206), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7207), .ZN(
        n7177) );
  NAND2_X1 U8753 ( .A1(n7178), .A2(n7177), .ZN(n7294) );
  OAI21_X1 U8754 ( .B1(n7178), .B2(n7177), .A(n7294), .ZN(n7181) );
  AND2_X1 U8755 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7642) );
  AOI21_X1 U8756 ( .B1(n10287), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7642), .ZN(
        n7179) );
  OAI21_X1 U8757 ( .B1(n10283), .B2(n7300), .A(n7179), .ZN(n7180) );
  AOI21_X1 U8758 ( .B1(n10282), .B2(n7181), .A(n7180), .ZN(n7182) );
  OAI21_X1 U8759 ( .B1(n7183), .B2(n10285), .A(n7182), .ZN(P2_U3258) );
  NAND2_X1 U8760 ( .A1(n9185), .A2(n7184), .ZN(n7185) );
  INV_X1 U8761 ( .A(n9184), .ZN(n7425) );
  NAND2_X1 U8762 ( .A1(n7425), .A2(n7225), .ZN(n8314) );
  INV_X1 U8763 ( .A(n7225), .ZN(n10247) );
  NAND2_X1 U8764 ( .A1(n9184), .A2(n10247), .ZN(n8319) );
  INV_X1 U8765 ( .A(n8187), .ZN(n7195) );
  OAI21_X1 U8766 ( .B1(n4544), .B2(n7195), .A(n7410), .ZN(n10251) );
  INV_X1 U8767 ( .A(n10251), .ZN(n7201) );
  AND2_X1 U8768 ( .A1(n8350), .A2(n5374), .ZN(n10195) );
  INV_X1 U8769 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7188) );
  INV_X1 U8770 ( .A(n7187), .ZN(n7223) );
  OAI22_X1 U8771 ( .A1(n10207), .A2(n7188), .B1(n7223), .B2(n10221), .ZN(n7193) );
  INV_X1 U8772 ( .A(n7189), .ZN(n7191) );
  INV_X1 U8773 ( .A(n7428), .ZN(n7190) );
  OAI21_X1 U8774 ( .B1(n10247), .B2(n7191), .A(n7190), .ZN(n10248) );
  INV_X1 U8775 ( .A(n10212), .ZN(n7973) );
  NOR2_X1 U8776 ( .A1(n10248), .A2(n7973), .ZN(n7192) );
  AOI211_X1 U8777 ( .C1(n10213), .C2(n7225), .A(n7193), .B(n7192), .ZN(n7200)
         );
  INV_X1 U8778 ( .A(n8234), .ZN(n8317) );
  XNOR2_X1 U8779 ( .A(n7414), .B(n7195), .ZN(n7196) );
  NAND2_X1 U8780 ( .A1(n7196), .A2(n9985), .ZN(n7198) );
  AOI22_X1 U8781 ( .A1(n9988), .A2(n9185), .B1(n9990), .B2(n9183), .ZN(n7197)
         );
  NAND2_X1 U8782 ( .A1(n7198), .A2(n7197), .ZN(n10249) );
  NAND2_X1 U8783 ( .A1(n10249), .A2(n10207), .ZN(n7199) );
  OAI211_X1 U8784 ( .C1(n7201), .C2(n10004), .A(n7200), .B(n7199), .ZN(
        P1_U3285) );
  AOI21_X1 U8785 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7213) );
  INV_X1 U8786 ( .A(n10283), .ZN(n9930) );
  INV_X1 U8787 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U8788 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7625) );
  OAI21_X1 U8789 ( .B1(n9913), .B2(n9787), .A(n7625), .ZN(n7205) );
  AOI21_X1 U8790 ( .B1(n9930), .B2(n7206), .A(n7205), .ZN(n7212) );
  AOI21_X1 U8791 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n7210) );
  NAND2_X1 U8792 ( .A1(n10282), .A2(n7210), .ZN(n7211) );
  OAI211_X1 U8793 ( .C1(n7213), .C2(n10285), .A(n7212), .B(n7211), .ZN(
        P2_U3257) );
  INV_X1 U8794 ( .A(n7214), .ZN(n7216) );
  NOR2_X1 U8795 ( .A1(n7216), .A2(n7215), .ZN(n7219) );
  INV_X1 U8796 ( .A(n7217), .ZN(n7314) );
  AOI21_X1 U8797 ( .B1(n7219), .B2(n7218), .A(n7314), .ZN(n7227) );
  AOI21_X1 U8798 ( .B1(n9138), .B2(n9183), .A(n7220), .ZN(n7222) );
  NAND2_X1 U8799 ( .A1(n9162), .A2(n9185), .ZN(n7221) );
  OAI211_X1 U8800 ( .C1(n9153), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7224)
         );
  AOI21_X1 U8801 ( .B1(n7225), .B2(n9168), .A(n7224), .ZN(n7226) );
  OAI21_X1 U8802 ( .B1(n7227), .B2(n9172), .A(n7226), .ZN(P1_U3237) );
  AOI211_X1 U8803 ( .C1(n7230), .C2(n7229), .A(n7228), .B(n9924), .ZN(n7240)
         );
  OAI21_X1 U8804 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7238) );
  NAND2_X1 U8805 ( .A1(n9930), .A2(n7234), .ZN(n7237) );
  AOI21_X1 U8806 ( .B1(n10287), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7235), .ZN(
        n7236) );
  OAI211_X1 U8807 ( .C1(n10285), .C2(n7238), .A(n7237), .B(n7236), .ZN(n7239)
         );
  OR2_X1 U8808 ( .A1(n7240), .A2(n7239), .ZN(P2_U3252) );
  NAND2_X1 U8809 ( .A1(n7242), .A2(n7241), .ZN(n7247) );
  INV_X1 U8810 ( .A(n7243), .ZN(n7244) );
  NAND2_X1 U8811 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  XNOR2_X1 U8812 ( .A(n7630), .B(n8429), .ZN(n7248) );
  NAND2_X1 U8813 ( .A1(n8562), .A2(n8430), .ZN(n7249) );
  NAND2_X1 U8814 ( .A1(n7248), .A2(n7249), .ZN(n7395) );
  NAND2_X1 U8815 ( .A1(n7395), .A2(n7250), .ZN(n7253) );
  INV_X1 U8816 ( .A(n7253), .ZN(n7251) );
  INV_X1 U8817 ( .A(n7398), .ZN(n7252) );
  AOI21_X1 U8818 ( .B1(n7254), .B2(n7253), .A(n7252), .ZN(n7258) );
  NAND2_X1 U8819 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8600) );
  OAI21_X1 U8820 ( .B1(n8522), .B2(n7495), .A(n8600), .ZN(n7256) );
  OAI22_X1 U8821 ( .A1(n7478), .A2(n8531), .B1(n8530), .B2(n7477), .ZN(n7255)
         );
  AOI211_X1 U8822 ( .C1(n7630), .C2(n4453), .A(n7256), .B(n7255), .ZN(n7257)
         );
  OAI21_X1 U8823 ( .B1(n7258), .B2(n8537), .A(n7257), .ZN(P2_U3233) );
  INV_X1 U8824 ( .A(n7261), .ZN(n7262) );
  NAND2_X2 U8825 ( .A1(n8896), .A2(n7262), .ZN(n8861) );
  NOR2_X2 U8826 ( .A1(n7263), .A2(n8430), .ZN(n8891) );
  NOR2_X1 U8827 ( .A1(n8882), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7268) );
  INV_X1 U8828 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U8829 ( .A1(n8896), .A2(n7264), .ZN(n7265) );
  OAI21_X1 U8830 ( .B1(n8896), .B2(n7266), .A(n7265), .ZN(n7267) );
  AOI211_X1 U8831 ( .C1(n8891), .C2(n7269), .A(n7268), .B(n7267), .ZN(n7275)
         );
  NOR2_X1 U8832 ( .A1(n7270), .A2(n4919), .ZN(n7271) );
  NAND2_X1 U8833 ( .A1(n8896), .A2(n7271), .ZN(n8894) );
  INV_X1 U8834 ( .A(n8881), .ZN(n7790) );
  NAND2_X1 U8835 ( .A1(n8896), .A2(n7790), .ZN(n7272) );
  NAND2_X1 U8836 ( .A1(n8760), .A2(n7273), .ZN(n7274) );
  OAI211_X1 U8837 ( .C1(n7276), .C2(n8861), .A(n7275), .B(n7274), .ZN(P2_U3293) );
  XNOR2_X1 U8838 ( .A(n6320), .B(n7284), .ZN(n7277) );
  NAND2_X1 U8839 ( .A1(n7277), .A2(n8878), .ZN(n7279) );
  AOI22_X1 U8840 ( .A1(n8871), .A2(n6786), .B1(n6946), .B2(n8873), .ZN(n7278)
         );
  NAND2_X1 U8841 ( .A1(n7279), .A2(n7278), .ZN(n10320) );
  INV_X1 U8842 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9779) );
  OAI22_X1 U8843 ( .A1(n8882), .A2(n9779), .B1(n9734), .B2(n8896), .ZN(n7282)
         );
  OAI21_X1 U8844 ( .B1(n4756), .B2(n4457), .A(n7280), .ZN(n10319) );
  NOR2_X1 U8845 ( .A1(n8695), .A2(n10319), .ZN(n7281) );
  AOI211_X1 U8846 ( .C1(n8896), .C2(n10320), .A(n7282), .B(n7281), .ZN(n7287)
         );
  OAI21_X1 U8847 ( .B1(n7285), .B2(n7284), .A(n7283), .ZN(n10322) );
  NAND2_X1 U8848 ( .A1(n8760), .A2(n10322), .ZN(n7286) );
  OAI211_X1 U8849 ( .C1(n4457), .C2(n8861), .A(n7287), .B(n7286), .ZN(P2_U3294) );
  INV_X1 U8850 ( .A(n10309), .ZN(n7293) );
  INV_X2 U8851 ( .A(n8896), .ZN(n8858) );
  AND2_X1 U8852 ( .A1(n6786), .A2(n8873), .ZN(n7288) );
  AOI21_X1 U8853 ( .B1(n10309), .B2(n8878), .A(n7288), .ZN(n10311) );
  OAI22_X1 U8854 ( .A1(n8858), .A2(n10311), .B1(n7289), .B2(n8882), .ZN(n7291)
         );
  AOI21_X1 U8855 ( .B1(n8695), .B2(n8861), .A(n7443), .ZN(n7290) );
  AOI211_X1 U8856 ( .C1(n8858), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7291), .B(
        n7290), .ZN(n7292) );
  OAI21_X1 U8857 ( .B1(n7293), .B2(n8865), .A(n7292), .ZN(P2_U3296) );
  AOI22_X1 U8858 ( .A1(n7574), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6106), .B2(
        n7577), .ZN(n7297) );
  OAI21_X1 U8859 ( .B1(n7295), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7294), .ZN(
        n7296) );
  OAI21_X1 U8860 ( .B1(n7297), .B2(n7296), .A(n7573), .ZN(n7306) );
  AND2_X1 U8861 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7769) );
  AOI21_X1 U8862 ( .B1(n10287), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7769), .ZN(
        n7298) );
  OAI21_X1 U8863 ( .B1(n10283), .B2(n7577), .A(n7298), .ZN(n7305) );
  AOI21_X1 U8864 ( .B1(n7300), .B2(n9616), .A(n7299), .ZN(n7302) );
  AOI22_X1 U8865 ( .A1(n7574), .A2(n9680), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7577), .ZN(n7301) );
  NOR2_X1 U8866 ( .A1(n7302), .A2(n7301), .ZN(n7576) );
  AOI21_X1 U8867 ( .B1(n7302), .B2(n7301), .A(n7576), .ZN(n7303) );
  NOR2_X1 U8868 ( .A1(n7303), .A2(n10285), .ZN(n7304) );
  AOI211_X1 U8869 ( .C1(n7306), .C2(n10282), .A(n7305), .B(n7304), .ZN(n7307)
         );
  INV_X1 U8870 ( .A(n7307), .ZN(P2_U3259) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9813) );
  INV_X1 U8872 ( .A(n7308), .ZN(n7309) );
  INV_X1 U8873 ( .A(n8671), .ZN(n8667) );
  OAI222_X1 U8874 ( .A1(n9018), .A2(n9813), .B1(n8454), .B2(n7309), .C1(
        P2_U3152), .C2(n8667), .ZN(P2_U3340) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7310) );
  INV_X1 U8876 ( .A(n10185), .ZN(n9217) );
  OAI222_X1 U8877 ( .A1(n9890), .A2(n7310), .B1(n4459), .B2(n7309), .C1(
        P1_U3084), .C2(n9217), .ZN(P1_U3335) );
  INV_X1 U8878 ( .A(n7311), .ZN(n7313) );
  NOR3_X1 U8879 ( .A1(n7314), .A2(n7313), .A3(n7312), .ZN(n7317) );
  INV_X1 U8880 ( .A(n7315), .ZN(n7316) );
  OAI21_X1 U8881 ( .B1(n7317), .B2(n7316), .A(n9115), .ZN(n7322) );
  AOI21_X1 U8882 ( .B1(n9162), .B2(n9184), .A(n7318), .ZN(n7319) );
  OAI21_X1 U8883 ( .B1(n9164), .B2(n7530), .A(n7319), .ZN(n7320) );
  AOI21_X1 U8884 ( .B1(n7429), .B2(n9166), .A(n7320), .ZN(n7321) );
  OAI211_X1 U8885 ( .C1(n7518), .C2(n9123), .A(n7322), .B(n7321), .ZN(P1_U3211) );
  OR2_X1 U8886 ( .A1(n7323), .A2(n8564), .ZN(n7482) );
  NAND2_X1 U8887 ( .A1(n7324), .A2(n7482), .ZN(n7325) );
  OR2_X1 U8888 ( .A1(n7325), .A2(n6035), .ZN(n7327) );
  NAND2_X1 U8889 ( .A1(n7325), .A2(n6035), .ZN(n7326) );
  NAND2_X1 U8890 ( .A1(n7327), .A2(n7326), .ZN(n10336) );
  OR2_X1 U8891 ( .A1(n10336), .A2(n8881), .ZN(n7336) );
  NAND2_X1 U8892 ( .A1(n7328), .A2(n7483), .ZN(n7329) );
  NAND2_X1 U8893 ( .A1(n7330), .A2(n7329), .ZN(n7334) );
  NAND2_X1 U8894 ( .A1(n8564), .A2(n8871), .ZN(n7332) );
  NAND2_X1 U8895 ( .A1(n8562), .A2(n8873), .ZN(n7331) );
  NAND2_X1 U8896 ( .A1(n7332), .A2(n7331), .ZN(n7333) );
  AOI21_X1 U8897 ( .B1(n7334), .B2(n8878), .A(n7333), .ZN(n7335) );
  NAND2_X1 U8898 ( .A1(n7336), .A2(n7335), .ZN(n10341) );
  NAND2_X1 U8899 ( .A1(n10341), .A2(n8896), .ZN(n7344) );
  INV_X1 U8900 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7338) );
  OAI22_X1 U8901 ( .A1(n8896), .A2(n7338), .B1(n7337), .B2(n8882), .ZN(n7342)
         );
  INV_X1 U8902 ( .A(n7479), .ZN(n10337) );
  OR2_X1 U8903 ( .A1(n7339), .A2(n10337), .ZN(n7340) );
  NAND2_X1 U8904 ( .A1(n7494), .A2(n7340), .ZN(n10338) );
  NOR2_X1 U8905 ( .A1(n8695), .A2(n10338), .ZN(n7341) );
  AOI211_X1 U8906 ( .C1(n8886), .C2(n7479), .A(n7342), .B(n7341), .ZN(n7343)
         );
  OAI211_X1 U8907 ( .C1(n10336), .C2(n8894), .A(n7344), .B(n7343), .ZN(
        P2_U3288) );
  NAND2_X1 U8908 ( .A1(n7398), .A2(n7395), .ZN(n7345) );
  XNOR2_X1 U8909 ( .A(n7647), .B(n8429), .ZN(n7399) );
  NAND2_X1 U8910 ( .A1(n8561), .A2(n8430), .ZN(n7400) );
  XNOR2_X1 U8911 ( .A(n7399), .B(n7400), .ZN(n7394) );
  XNOR2_X1 U8912 ( .A(n7345), .B(n7394), .ZN(n7351) );
  OAI22_X1 U8913 ( .A1(n8522), .A2(n7510), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7346), .ZN(n7349) );
  OAI22_X1 U8914 ( .A1(n7347), .A2(n8531), .B1(n8530), .B2(n7658), .ZN(n7348)
         );
  AOI211_X1 U8915 ( .C1(n7647), .C2(n4453), .A(n7349), .B(n7348), .ZN(n7350)
         );
  OAI21_X1 U8916 ( .B1(n7351), .B2(n8537), .A(n7350), .ZN(P2_U3219) );
  AOI22_X1 U8917 ( .A1(n9993), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7352), .B2(
        n8305), .ZN(n7356) );
  OAI21_X1 U8918 ( .B1(n7354), .B2(n7961), .A(n7353), .ZN(n7355) );
  AND3_X1 U8919 ( .A1(n7357), .A2(n7356), .A3(n7355), .ZN(n7360) );
  NOR2_X1 U8920 ( .A1(n10216), .A2(n9342), .ZN(n9428) );
  AOI22_X1 U8921 ( .A1(n9428), .A2(n7358), .B1(n10216), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7359) );
  OAI21_X1 U8922 ( .B1(n7360), .B2(n10216), .A(n7359), .ZN(P1_U3290) );
  INV_X1 U8923 ( .A(n7361), .ZN(n8360) );
  OAI222_X1 U8924 ( .A1(n9890), .A2(n7362), .B1(n4459), .B2(n8360), .C1(
        P1_U3084), .C2(n10200), .ZN(P1_U3334) );
  OAI21_X1 U8925 ( .B1(n7364), .B2(n7366), .A(n7363), .ZN(n10333) );
  INV_X1 U8926 ( .A(n10333), .ZN(n7378) );
  XNOR2_X1 U8927 ( .A(n7365), .B(n7366), .ZN(n7367) );
  OAI222_X1 U8928 ( .A1(n8852), .A2(n7369), .B1(n8850), .B2(n7368), .C1(n7367), 
        .C2(n8847), .ZN(n10331) );
  INV_X1 U8929 ( .A(n7370), .ZN(n7372) );
  OAI21_X1 U8930 ( .B1(n10329), .B2(n7372), .A(n7371), .ZN(n10330) );
  OAI22_X1 U8931 ( .A1(n8695), .A2(n10330), .B1(n7373), .B2(n8882), .ZN(n7374)
         );
  AOI21_X1 U8932 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n8858), .A(n7374), .ZN(
        n7375) );
  OAI21_X1 U8933 ( .B1(n10329), .B2(n8861), .A(n7375), .ZN(n7376) );
  AOI21_X1 U8934 ( .B1(n8896), .B2(n10331), .A(n7376), .ZN(n7377) );
  OAI21_X1 U8935 ( .B1(n8865), .B2(n7378), .A(n7377), .ZN(P2_U3290) );
  NOR2_X1 U8936 ( .A1(n8882), .A2(n7379), .ZN(n7383) );
  OAI21_X1 U8937 ( .B1(n7381), .B2(n10323), .A(n7380), .ZN(n10324) );
  NOR2_X1 U8938 ( .A1(n8695), .A2(n10324), .ZN(n7382) );
  AOI211_X1 U8939 ( .C1(n8858), .C2(P2_REG2_REG_4__SCAN_IN), .A(n7383), .B(
        n7382), .ZN(n7393) );
  OAI21_X1 U8940 ( .B1(n7386), .B2(n7385), .A(n7384), .ZN(n10327) );
  XNOR2_X1 U8941 ( .A(n7388), .B(n7387), .ZN(n7389) );
  NAND2_X1 U8942 ( .A1(n7389), .A2(n8878), .ZN(n7391) );
  AOI22_X1 U8943 ( .A1(n8871), .A2(n6946), .B1(n8566), .B2(n8873), .ZN(n7390)
         );
  NAND2_X1 U8944 ( .A1(n7391), .A2(n7390), .ZN(n10325) );
  AOI22_X1 U8945 ( .A1(n8760), .A2(n10327), .B1(n8896), .B2(n10325), .ZN(n7392) );
  OAI211_X1 U8946 ( .C1(n10323), .C2(n8861), .A(n7393), .B(n7392), .ZN(
        P2_U3292) );
  INV_X1 U8947 ( .A(n7394), .ZN(n7396) );
  AND2_X1 U8948 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  INV_X1 U8949 ( .A(n7399), .ZN(n7402) );
  INV_X1 U8950 ( .A(n7400), .ZN(n7401) );
  NAND2_X1 U8951 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  XNOR2_X1 U8952 ( .A(n7734), .B(n8436), .ZN(n7612) );
  NAND2_X1 U8953 ( .A1(n8560), .A2(n8430), .ZN(n7610) );
  XNOR2_X1 U8954 ( .A(n7612), .B(n7610), .ZN(n7614) );
  XNOR2_X1 U8955 ( .A(n7615), .B(n7614), .ZN(n7408) );
  OAI22_X1 U8956 ( .A1(n8522), .A2(n7735), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6066), .ZN(n7406) );
  OAI22_X1 U8957 ( .A1(n7477), .A2(n8531), .B1(n8530), .B2(n7640), .ZN(n7405)
         );
  AOI211_X1 U8958 ( .C1(n7734), .C2(n4453), .A(n7406), .B(n7405), .ZN(n7407)
         );
  OAI21_X1 U8959 ( .B1(n7408), .B2(n8537), .A(n7407), .ZN(P2_U3238) );
  NAND2_X1 U8960 ( .A1(n7425), .A2(n10247), .ZN(n7409) );
  NAND2_X1 U8961 ( .A1(n7518), .A2(n9183), .ZN(n8081) );
  INV_X1 U8962 ( .A(n9183), .ZN(n7557) );
  NAND2_X1 U8963 ( .A1(n7557), .A2(n7430), .ZN(n8082) );
  NAND2_X1 U8964 ( .A1(n8081), .A2(n8082), .ZN(n8189) );
  NAND2_X1 U8965 ( .A1(n7427), .A2(n8189), .ZN(n7426) );
  NAND2_X1 U8966 ( .A1(n7518), .A2(n7557), .ZN(n7411) );
  NAND2_X1 U8967 ( .A1(n7426), .A2(n7411), .ZN(n7553) );
  OR2_X1 U8968 ( .A1(n7594), .A2(n7530), .ZN(n8086) );
  NAND2_X1 U8969 ( .A1(n7594), .A2(n7530), .ZN(n8083) );
  NAND2_X1 U8970 ( .A1(n7594), .A2(n9182), .ZN(n7412) );
  AND2_X1 U8971 ( .A1(n10262), .A2(n9181), .ZN(n7413) );
  OR2_X1 U8972 ( .A1(n7679), .A2(n7776), .ZN(n8241) );
  NAND2_X1 U8973 ( .A1(n7679), .A2(n7776), .ZN(n8223) );
  NAND2_X1 U8974 ( .A1(n8241), .A2(n8223), .ZN(n7597) );
  XNOR2_X1 U8975 ( .A(n7598), .B(n7597), .ZN(n9941) );
  INV_X1 U8976 ( .A(n9181), .ZN(n7556) );
  NAND2_X1 U8977 ( .A1(n10262), .A2(n7556), .ZN(n8222) );
  AND2_X1 U8978 ( .A1(n8222), .A2(n8083), .ZN(n8089) );
  OR2_X1 U8979 ( .A1(n10262), .A2(n7556), .ZN(n8091) );
  INV_X1 U8980 ( .A(n7597), .ZN(n8194) );
  XNOR2_X1 U8981 ( .A(n7601), .B(n8194), .ZN(n7416) );
  AOI22_X1 U8982 ( .A1(n9988), .A2(n9181), .B1(n9990), .B2(n9179), .ZN(n7415)
         );
  OAI21_X1 U8983 ( .B1(n7416), .B2(n9421), .A(n7415), .ZN(n7417) );
  AOI21_X1 U8984 ( .B1(n9941), .B2(n7961), .A(n7417), .ZN(n9943) );
  INV_X1 U8985 ( .A(n7679), .ZN(n9939) );
  OAI211_X1 U8986 ( .C1(n7536), .C2(n9939), .A(n9999), .B(n7603), .ZN(n9938)
         );
  OR2_X1 U8987 ( .A1(n7418), .A2(n9342), .ZN(n10003) );
  AOI22_X1 U8988 ( .A1(n10216), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7673), .B2(
        n9993), .ZN(n7420) );
  NAND2_X1 U8989 ( .A1(n7679), .A2(n10213), .ZN(n7419) );
  OAI211_X1 U8990 ( .C1(n9938), .C2(n10003), .A(n7420), .B(n7419), .ZN(n7421)
         );
  AOI21_X1 U8991 ( .B1(n9941), .B2(n7968), .A(n7421), .ZN(n7422) );
  OAI21_X1 U8992 ( .B1(n9943), .B2(n10216), .A(n7422), .ZN(P1_U3281) );
  AOI21_X1 U8993 ( .B1(n8189), .B2(n7423), .A(n4545), .ZN(n7424) );
  OAI222_X1 U8994 ( .A1(n9425), .A2(n7530), .B1(n9423), .B2(n7425), .C1(n9421), 
        .C2(n7424), .ZN(n7519) );
  INV_X1 U8995 ( .A(n7519), .ZN(n7435) );
  OAI21_X1 U8996 ( .B1(n7427), .B2(n8189), .A(n7426), .ZN(n7521) );
  INV_X1 U8997 ( .A(n10004), .ZN(n7881) );
  OAI211_X1 U8998 ( .C1(n7428), .C2(n7518), .A(n7563), .B(n9999), .ZN(n7517)
         );
  AOI22_X1 U8999 ( .A1(n10216), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7429), .B2(
        n9993), .ZN(n7432) );
  NAND2_X1 U9000 ( .A1(n10213), .A2(n7430), .ZN(n7431) );
  OAI211_X1 U9001 ( .C1(n7517), .C2(n10003), .A(n7432), .B(n7431), .ZN(n7433)
         );
  AOI21_X1 U9002 ( .B1(n7521), .B2(n7881), .A(n7433), .ZN(n7434) );
  OAI21_X1 U9003 ( .B1(n7435), .B2(n10216), .A(n7434), .ZN(P1_U3284) );
  OAI21_X1 U9004 ( .B1(n7438), .B2(n7437), .A(n7436), .ZN(n10317) );
  XNOR2_X1 U9005 ( .A(n6468), .B(n7438), .ZN(n7440) );
  AOI21_X1 U9006 ( .B1(n7440), .B2(n8878), .A(n7439), .ZN(n10314) );
  OAI21_X1 U9007 ( .B1(n9912), .B2(n8882), .A(n10314), .ZN(n7441) );
  MUX2_X1 U9008 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7441), .S(n8896), .Z(n7445)
         );
  OAI21_X1 U9009 ( .B1(n6741), .B2(n7443), .A(n7442), .ZN(n10313) );
  OAI22_X1 U9010 ( .A1(n8695), .A2(n10313), .B1(n6741), .B2(n8861), .ZN(n7444)
         );
  AOI211_X1 U9011 ( .C1(n8760), .C2(n10317), .A(n7445), .B(n7444), .ZN(n7446)
         );
  INV_X1 U9012 ( .A(n7446), .ZN(P2_U3295) );
  XNOR2_X1 U9013 ( .A(n7447), .B(n7449), .ZN(n7455) );
  OAI21_X1 U9014 ( .B1(n7450), .B2(n7449), .A(n7448), .ZN(n10245) );
  OAI22_X1 U9015 ( .A1(n7452), .A2(n9423), .B1(n7451), .B2(n9425), .ZN(n7453)
         );
  AOI21_X1 U9016 ( .B1(n10245), .B2(n7961), .A(n7453), .ZN(n7454) );
  OAI21_X1 U9017 ( .B1(n9421), .B2(n7455), .A(n7454), .ZN(n10243) );
  INV_X1 U9018 ( .A(n10243), .ZN(n7465) );
  NAND2_X1 U9019 ( .A1(n7456), .A2(n7460), .ZN(n7457) );
  NAND2_X1 U9020 ( .A1(n7458), .A2(n7457), .ZN(n10242) );
  AOI22_X1 U9021 ( .A1(n10216), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7459), .B2(
        n9993), .ZN(n7462) );
  NAND2_X1 U9022 ( .A1(n10213), .A2(n7460), .ZN(n7461) );
  OAI211_X1 U9023 ( .C1(n7973), .C2(n10242), .A(n7462), .B(n7461), .ZN(n7463)
         );
  AOI21_X1 U9024 ( .B1(n10245), .B2(n7968), .A(n7463), .ZN(n7464) );
  OAI21_X1 U9025 ( .B1(n7465), .B2(n10216), .A(n7464), .ZN(P1_U3287) );
  MUX2_X1 U9026 ( .A(n7466), .B(P2_REG2_REG_5__SCAN_IN), .S(n8858), .Z(n7473)
         );
  NOR2_X1 U9027 ( .A1(n8858), .A2(n4460), .ZN(n8854) );
  INV_X1 U9028 ( .A(n8854), .ZN(n7471) );
  INV_X1 U9029 ( .A(n8882), .ZN(n8856) );
  AOI22_X1 U9030 ( .A1(n8886), .A2(n7468), .B1(n8856), .B2(n7467), .ZN(n7469)
         );
  OAI21_X1 U9031 ( .B1(n7471), .B2(n7470), .A(n7469), .ZN(n7472) );
  AOI211_X1 U9032 ( .C1(n8760), .C2(n7474), .A(n7473), .B(n7472), .ZN(n7475)
         );
  INV_X1 U9033 ( .A(n7475), .ZN(P2_U3291) );
  XNOR2_X1 U9034 ( .A(n7476), .B(n7490), .ZN(n7493) );
  OAI22_X1 U9035 ( .A1(n7478), .A2(n8850), .B1(n7477), .B2(n8852), .ZN(n7492)
         );
  NAND2_X1 U9036 ( .A1(n7479), .A2(n8563), .ZN(n7481) );
  AND2_X1 U9037 ( .A1(n7480), .A2(n7481), .ZN(n7486) );
  INV_X1 U9038 ( .A(n7481), .ZN(n7485) );
  AND2_X1 U9039 ( .A1(n7483), .A2(n7482), .ZN(n7484) );
  AOI21_X1 U9040 ( .B1(n7487), .B2(n7486), .A(n4516), .ZN(n7489) );
  INV_X1 U9041 ( .A(n7504), .ZN(n7488) );
  AOI21_X1 U9042 ( .B1(n7490), .B2(n7489), .A(n7488), .ZN(n7634) );
  NOR2_X1 U9043 ( .A1(n7634), .A2(n8881), .ZN(n7491) );
  AOI211_X1 U9044 ( .C1(n7493), .C2(n8878), .A(n7492), .B(n7491), .ZN(n7633)
         );
  AOI21_X1 U9045 ( .B1(n7630), .B2(n7494), .A(n4541), .ZN(n7631) );
  INV_X1 U9046 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7496) );
  OAI22_X1 U9047 ( .A1(n8896), .A2(n7496), .B1(n7495), .B2(n8882), .ZN(n7499)
         );
  INV_X1 U9048 ( .A(n7630), .ZN(n7497) );
  NOR2_X1 U9049 ( .A1(n8861), .A2(n7497), .ZN(n7498) );
  AOI211_X1 U9050 ( .C1(n7631), .C2(n8891), .A(n7499), .B(n7498), .ZN(n7502)
         );
  INV_X1 U9051 ( .A(n7634), .ZN(n7500) );
  INV_X1 U9052 ( .A(n8894), .ZN(n7798) );
  NAND2_X1 U9053 ( .A1(n7500), .A2(n7798), .ZN(n7501) );
  OAI211_X1 U9054 ( .C1(n7633), .C2(n8858), .A(n7502), .B(n7501), .ZN(P2_U3287) );
  OR2_X1 U9055 ( .A1(n7630), .A2(n8562), .ZN(n7503) );
  INV_X1 U9056 ( .A(n7649), .ZN(n7505) );
  AOI21_X1 U9057 ( .B1(n6059), .B2(n7506), .A(n7505), .ZN(n10346) );
  INV_X1 U9058 ( .A(n10346), .ZN(n7516) );
  OAI211_X1 U9059 ( .C1(n4454), .C2(n6059), .A(n8878), .B(n7507), .ZN(n7509)
         );
  AOI22_X1 U9060 ( .A1(n8871), .A2(n8562), .B1(n8560), .B2(n8873), .ZN(n7508)
         );
  NAND2_X1 U9061 ( .A1(n7509), .A2(n7508), .ZN(n10345) );
  INV_X1 U9062 ( .A(n7647), .ZN(n10342) );
  OAI21_X1 U9063 ( .B1(n4541), .B2(n10342), .A(n7699), .ZN(n10343) );
  OAI22_X1 U9064 ( .A1(n8896), .A2(n7511), .B1(n7510), .B2(n8882), .ZN(n7512)
         );
  AOI21_X1 U9065 ( .B1(n8886), .B2(n7647), .A(n7512), .ZN(n7513) );
  OAI21_X1 U9066 ( .B1(n10343), .B2(n8695), .A(n7513), .ZN(n7514) );
  AOI21_X1 U9067 ( .B1(n10345), .B2(n8896), .A(n7514), .ZN(n7515) );
  OAI21_X1 U9068 ( .B1(n7516), .B2(n8865), .A(n7515), .ZN(P2_U3286) );
  INV_X1 U9069 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9070 ( .B1(n7518), .B2(n10263), .A(n7517), .ZN(n7520) );
  AOI211_X1 U9071 ( .C1(n10252), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7524)
         );
  OR2_X1 U9072 ( .A1(n7524), .A2(n10271), .ZN(n7522) );
  OAI21_X1 U9073 ( .B1(n10273), .B2(n7523), .A(n7522), .ZN(P1_U3475) );
  OR2_X1 U9074 ( .A1(n7524), .A2(n10279), .ZN(n7525) );
  OAI21_X1 U9075 ( .B1(n4456), .B2(n7526), .A(n7525), .ZN(P1_U3530) );
  XNOR2_X1 U9076 ( .A(n10262), .B(n9181), .ZN(n8191) );
  XOR2_X1 U9077 ( .A(n8191), .B(n7527), .Z(n10261) );
  INV_X1 U9078 ( .A(n7968), .ZN(n7570) );
  NAND2_X1 U9079 ( .A1(n7528), .A2(n8083), .ZN(n7529) );
  XNOR2_X1 U9080 ( .A(n7529), .B(n8191), .ZN(n7532) );
  OAI22_X1 U9081 ( .A1(n7530), .A2(n9423), .B1(n7776), .B2(n9425), .ZN(n7531)
         );
  AOI21_X1 U9082 ( .B1(n7532), .B2(n9985), .A(n7531), .ZN(n7533) );
  OAI21_X1 U9083 ( .B1(n10261), .B2(n7561), .A(n7533), .ZN(n10267) );
  NAND2_X1 U9084 ( .A1(n10267), .A2(n10207), .ZN(n7541) );
  INV_X1 U9085 ( .A(n7534), .ZN(n7689) );
  OAI22_X1 U9086 ( .A1(n10207), .A2(n7535), .B1(n7689), .B2(n10221), .ZN(n7539) );
  AND2_X1 U9087 ( .A1(n7564), .A2(n10262), .ZN(n7537) );
  OR2_X1 U9088 ( .A1(n7537), .A2(n7536), .ZN(n10266) );
  NOR2_X1 U9089 ( .A1(n10266), .A2(n7973), .ZN(n7538) );
  AOI211_X1 U9090 ( .C1(n10213), .C2(n10262), .A(n7539), .B(n7538), .ZN(n7540)
         );
  OAI211_X1 U9091 ( .C1(n10261), .C2(n7570), .A(n7541), .B(n7540), .ZN(
        P1_U3282) );
  NAND2_X1 U9092 ( .A1(n7542), .A2(n8760), .ZN(n7550) );
  OAI22_X1 U9093 ( .A1(n8896), .A2(n7544), .B1(n7543), .B2(n8882), .ZN(n7547)
         );
  NOR2_X1 U9094 ( .A1(n8861), .A2(n7545), .ZN(n7546) );
  AOI211_X1 U9095 ( .C1(n7548), .C2(n8891), .A(n7547), .B(n7546), .ZN(n7549)
         );
  OAI211_X1 U9096 ( .C1(n8858), .C2(n7551), .A(n7550), .B(n7549), .ZN(P2_U3289) );
  NAND2_X1 U9097 ( .A1(n7553), .A2(n8193), .ZN(n7554) );
  NAND2_X1 U9098 ( .A1(n7552), .A2(n7554), .ZN(n10254) );
  OAI21_X1 U9099 ( .B1(n8193), .B2(n7555), .A(n7528), .ZN(n7559) );
  OAI22_X1 U9100 ( .A1(n7557), .A2(n9423), .B1(n7556), .B2(n9425), .ZN(n7558)
         );
  AOI21_X1 U9101 ( .B1(n7559), .B2(n9985), .A(n7558), .ZN(n7560) );
  OAI21_X1 U9102 ( .B1(n10254), .B2(n7561), .A(n7560), .ZN(n10257) );
  NAND2_X1 U9103 ( .A1(n10257), .A2(n10207), .ZN(n7569) );
  INV_X1 U9104 ( .A(n7562), .ZN(n7592) );
  OAI22_X1 U9105 ( .A1(n10207), .A2(n9785), .B1(n7592), .B2(n10221), .ZN(n7567) );
  INV_X1 U9106 ( .A(n7563), .ZN(n7565) );
  INV_X1 U9107 ( .A(n7594), .ZN(n10256) );
  OAI211_X1 U9108 ( .C1(n7565), .C2(n10256), .A(n9999), .B(n7564), .ZN(n10255)
         );
  INV_X1 U9109 ( .A(n9428), .ZN(n7874) );
  NOR2_X1 U9110 ( .A1(n10255), .A2(n7874), .ZN(n7566) );
  AOI211_X1 U9111 ( .C1(n10213), .C2(n7594), .A(n7567), .B(n7566), .ZN(n7568)
         );
  OAI211_X1 U9112 ( .C1(n10254), .C2(n7570), .A(n7569), .B(n7568), .ZN(
        P1_U3283) );
  INV_X1 U9113 ( .A(n7571), .ZN(n7668) );
  OAI222_X1 U9114 ( .A1(n9890), .A2(n7572), .B1(n4459), .B2(n7668), .C1(n8343), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  XNOR2_X1 U9115 ( .A(n8616), .B(n8611), .ZN(n7575) );
  NAND2_X1 U9116 ( .A1(n7575), .A2(n7855), .ZN(n8618) );
  OAI21_X1 U9117 ( .B1(n7575), .B2(n7855), .A(n8618), .ZN(n7583) );
  AOI21_X1 U9118 ( .B1(n7577), .B2(n9680), .A(n7576), .ZN(n8610) );
  XNOR2_X1 U9119 ( .A(n8610), .B(n8617), .ZN(n7578) );
  NAND2_X1 U9120 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7578), .ZN(n8612) );
  OAI211_X1 U9121 ( .C1(n7578), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10281), .B(
        n8612), .ZN(n7581) );
  AND2_X1 U9122 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7579) );
  AOI21_X1 U9123 ( .B1(n10287), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7579), .ZN(
        n7580) );
  OAI211_X1 U9124 ( .C1(n10283), .C2(n8617), .A(n7581), .B(n7580), .ZN(n7582)
         );
  AOI21_X1 U9125 ( .B1(n10282), .B2(n7583), .A(n7582), .ZN(n7584) );
  INV_X1 U9126 ( .A(n7584), .ZN(P2_U3260) );
  NAND2_X1 U9127 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  XOR2_X1 U9128 ( .A(n7588), .B(n7587), .Z(n7596) );
  NOR2_X1 U9129 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7589), .ZN(n10102) );
  AOI21_X1 U9130 ( .B1(n9162), .B2(n9183), .A(n10102), .ZN(n7591) );
  NAND2_X1 U9131 ( .A1(n9138), .A2(n9181), .ZN(n7590) );
  OAI211_X1 U9132 ( .C1(n9153), .C2(n7592), .A(n7591), .B(n7590), .ZN(n7593)
         );
  AOI21_X1 U9133 ( .B1(n7594), .B2(n9168), .A(n7593), .ZN(n7595) );
  OAI21_X1 U9134 ( .B1(n7596), .B2(n9172), .A(n7595), .ZN(P1_U3219) );
  NAND2_X1 U9135 ( .A1(n7598), .A2(n7597), .ZN(n7600) );
  OR2_X1 U9136 ( .A1(n7679), .A2(n9180), .ZN(n7599) );
  XNOR2_X1 U9137 ( .A(n7710), .B(n9179), .ZN(n8197) );
  XOR2_X1 U9138 ( .A(n7707), .B(n8197), .Z(n10041) );
  INV_X1 U9139 ( .A(n10041), .ZN(n7609) );
  INV_X1 U9140 ( .A(n9178), .ZN(n7708) );
  XNOR2_X1 U9141 ( .A(n7709), .B(n8197), .ZN(n7602) );
  OAI222_X1 U9142 ( .A1(n9425), .A2(n7708), .B1(n9423), .B2(n7776), .C1(n7602), 
        .C2(n9421), .ZN(n10039) );
  INV_X1 U9143 ( .A(n7603), .ZN(n7604) );
  INV_X1 U9144 ( .A(n7710), .ZN(n10037) );
  OAI21_X1 U9145 ( .B1(n7604), .B2(n10037), .A(n7714), .ZN(n10038) );
  AOI22_X1 U9146 ( .A1(n10216), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7778), .B2(
        n9993), .ZN(n7606) );
  NAND2_X1 U9147 ( .A1(n7710), .A2(n10213), .ZN(n7605) );
  OAI211_X1 U9148 ( .C1(n10038), .C2(n7973), .A(n7606), .B(n7605), .ZN(n7607)
         );
  AOI21_X1 U9149 ( .B1(n10039), .B2(n10207), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9150 ( .B1(n7609), .B2(n10004), .A(n7608), .ZN(P1_U3280) );
  INV_X1 U9151 ( .A(n7781), .ZN(n10349) );
  INV_X1 U9152 ( .A(n7610), .ZN(n7611) );
  AND2_X1 U9153 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  AOI21_X2 U9154 ( .B1(n7615), .B2(n7614), .A(n7613), .ZN(n7622) );
  XNOR2_X1 U9155 ( .A(n7781), .B(n8429), .ZN(n7616) );
  NAND2_X1 U9156 ( .A1(n8559), .A2(n8430), .ZN(n7617) );
  NAND2_X1 U9157 ( .A1(n7616), .A2(n7617), .ZN(n7638) );
  INV_X1 U9158 ( .A(n7616), .ZN(n7619) );
  INV_X1 U9159 ( .A(n7617), .ZN(n7618) );
  NAND2_X1 U9160 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  AND2_X1 U9161 ( .A1(n7638), .A2(n7620), .ZN(n7621) );
  OAI21_X1 U9162 ( .B1(n7622), .B2(n7621), .A(n7639), .ZN(n7623) );
  NAND2_X1 U9163 ( .A1(n7623), .A2(n8539), .ZN(n7629) );
  INV_X1 U9164 ( .A(n7624), .ZN(n7659) );
  INV_X1 U9165 ( .A(n7625), .ZN(n7627) );
  OAI22_X1 U9166 ( .A1(n7658), .A2(n8531), .B1(n8530), .B2(n7767), .ZN(n7626)
         );
  AOI211_X1 U9167 ( .C1(n7659), .C2(n8548), .A(n7627), .B(n7626), .ZN(n7628)
         );
  OAI211_X1 U9168 ( .C1(n10349), .C2(n8551), .A(n7629), .B(n7628), .ZN(
        P2_U3226) );
  AOI22_X1 U9169 ( .A1(n7631), .A2(n8985), .B1(n9980), .B2(n7630), .ZN(n7632)
         );
  OAI211_X1 U9170 ( .C1(n7634), .C2(n10335), .A(n7633), .B(n7632), .ZN(n7636)
         );
  NAND2_X1 U9171 ( .A1(n7636), .A2(n10358), .ZN(n7635) );
  OAI21_X1 U9172 ( .B1(n10358), .B2(n6039), .A(n7635), .ZN(P2_U3478) );
  NAND2_X1 U9173 ( .A1(n7636), .A2(n10370), .ZN(n7637) );
  OAI21_X1 U9174 ( .B1(n10370), .B2(n7106), .A(n7637), .ZN(P2_U3529) );
  XNOR2_X1 U9175 ( .A(n8984), .B(n8429), .ZN(n7759) );
  NAND2_X1 U9176 ( .A1(n8558), .A2(n8430), .ZN(n7760) );
  XNOR2_X1 U9177 ( .A(n7759), .B(n7760), .ZN(n7758) );
  XNOR2_X1 U9178 ( .A(n7757), .B(n7758), .ZN(n7646) );
  INV_X1 U9179 ( .A(n7794), .ZN(n7643) );
  OAI22_X1 U9180 ( .A1(n7640), .A2(n8531), .B1(n8530), .B2(n7805), .ZN(n7641)
         );
  AOI211_X1 U9181 ( .C1(n8548), .C2(n7643), .A(n7642), .B(n7641), .ZN(n7645)
         );
  NAND2_X1 U9182 ( .A1(n8984), .A2(n4453), .ZN(n7644) );
  OAI211_X1 U9183 ( .C1(n7646), .C2(n8537), .A(n7645), .B(n7644), .ZN(P2_U3236) );
  NAND2_X1 U9184 ( .A1(n7647), .A2(n8561), .ZN(n7648) );
  NAND2_X1 U9185 ( .A1(n7693), .A2(n7695), .ZN(n7651) );
  NAND2_X1 U9186 ( .A1(n7734), .A2(n8560), .ZN(n7650) );
  XNOR2_X1 U9187 ( .A(n7783), .B(n4706), .ZN(n10355) );
  INV_X1 U9188 ( .A(n10355), .ZN(n7664) );
  NAND2_X1 U9189 ( .A1(n7507), .A2(n7653), .ZN(n7655) );
  AND2_X1 U9190 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  XNOR2_X1 U9191 ( .A(n7656), .B(n4706), .ZN(n7657) );
  OAI222_X1 U9192 ( .A1(n8852), .A2(n7767), .B1(n8850), .B2(n7658), .C1(n8847), 
        .C2(n7657), .ZN(n10352) );
  NAND2_X1 U9193 ( .A1(n7698), .A2(n10349), .ZN(n7792) );
  OAI21_X1 U9194 ( .B1(n7698), .B2(n10349), .A(n7792), .ZN(n10351) );
  AOI22_X1 U9195 ( .A1(n8858), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7659), .B2(
        n8856), .ZN(n7661) );
  NAND2_X1 U9196 ( .A1(n8886), .A2(n7781), .ZN(n7660) );
  OAI211_X1 U9197 ( .C1(n10351), .C2(n8695), .A(n7661), .B(n7660), .ZN(n7662)
         );
  AOI21_X1 U9198 ( .B1(n10352), .B2(n8896), .A(n7662), .ZN(n7663) );
  OAI21_X1 U9199 ( .B1(n8865), .B2(n7664), .A(n7663), .ZN(P2_U3284) );
  INV_X1 U9200 ( .A(n7665), .ZN(n8382) );
  OAI222_X1 U9201 ( .A1(n9018), .A2(n7667), .B1(P2_U3152), .B2(n7666), .C1(
        n8454), .C2(n8382), .ZN(P2_U3337) );
  OAI222_X1 U9202 ( .A1(n9018), .A2(n7669), .B1(P2_U3152), .B2(n4455), .C1(
        n8454), .C2(n7668), .ZN(P2_U3338) );
  NAND2_X1 U9203 ( .A1(n4546), .A2(n7671), .ZN(n7672) );
  XNOR2_X1 U9204 ( .A(n7670), .B(n7672), .ZN(n7681) );
  INV_X1 U9205 ( .A(n7673), .ZN(n7677) );
  AOI21_X1 U9206 ( .B1(n9138), .B2(n9179), .A(n7674), .ZN(n7676) );
  NAND2_X1 U9207 ( .A1(n9162), .A2(n9181), .ZN(n7675) );
  OAI211_X1 U9208 ( .C1(n9153), .C2(n7677), .A(n7676), .B(n7675), .ZN(n7678)
         );
  AOI21_X1 U9209 ( .B1(n7679), .B2(n9168), .A(n7678), .ZN(n7680) );
  OAI21_X1 U9210 ( .B1(n7681), .B2(n9172), .A(n7680), .ZN(P1_U3215) );
  INV_X1 U9211 ( .A(n7683), .ZN(n7684) );
  AOI21_X1 U9212 ( .B1(n7685), .B2(n7682), .A(n7684), .ZN(n7692) );
  AOI21_X1 U9213 ( .B1(n9162), .B2(n9182), .A(n7686), .ZN(n7688) );
  NAND2_X1 U9214 ( .A1(n9138), .A2(n9180), .ZN(n7687) );
  OAI211_X1 U9215 ( .C1(n9153), .C2(n7689), .A(n7688), .B(n7687), .ZN(n7690)
         );
  AOI21_X1 U9216 ( .B1(n10262), .B2(n9168), .A(n7690), .ZN(n7691) );
  OAI21_X1 U9217 ( .B1(n7692), .B2(n9172), .A(n7691), .ZN(P1_U3229) );
  INV_X1 U9218 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U9219 ( .A(n7693), .B(n7695), .ZN(n7743) );
  NAND2_X1 U9220 ( .A1(n7507), .A2(n7694), .ZN(n7696) );
  XNOR2_X1 U9221 ( .A(n7696), .B(n7695), .ZN(n7697) );
  AOI222_X1 U9222 ( .A1(n8878), .A2(n7697), .B1(n8559), .B2(n8873), .C1(n8561), 
        .C2(n8871), .ZN(n7738) );
  AOI21_X1 U9223 ( .B1(n7734), .B2(n7699), .A(n7698), .ZN(n7741) );
  AOI22_X1 U9224 ( .A1(n7741), .A2(n8985), .B1(n9980), .B2(n7734), .ZN(n7700)
         );
  OAI211_X1 U9225 ( .C1(n8981), .C2(n7743), .A(n7738), .B(n7700), .ZN(n7703)
         );
  NAND2_X1 U9226 ( .A1(n7703), .A2(n10358), .ZN(n7701) );
  OAI21_X1 U9227 ( .B1(n10358), .B2(n7702), .A(n7701), .ZN(P2_U3484) );
  NAND2_X1 U9228 ( .A1(n7703), .A2(n10370), .ZN(n7704) );
  OAI21_X1 U9229 ( .B1(n10370), .B2(n7157), .A(n7704), .ZN(P2_U3531) );
  NOR2_X1 U9230 ( .A1(n7710), .A2(n9179), .ZN(n7706) );
  NAND2_X1 U9231 ( .A1(n7710), .A2(n9179), .ZN(n7705) );
  OAI21_X1 U9232 ( .B1(n7707), .B2(n7706), .A(n7705), .ZN(n7720) );
  OR2_X1 U9233 ( .A1(n7894), .A2(n7708), .ZN(n8099) );
  NAND2_X1 U9234 ( .A1(n7894), .A2(n7708), .ZN(n8100) );
  NAND2_X1 U9235 ( .A1(n8099), .A2(n8100), .ZN(n8196) );
  XNOR2_X1 U9236 ( .A(n7720), .B(n8196), .ZN(n7832) );
  INV_X1 U9237 ( .A(n9177), .ZN(n7891) );
  INV_X1 U9238 ( .A(n9179), .ZN(n7713) );
  NAND2_X1 U9239 ( .A1(n7710), .A2(n7713), .ZN(n8096) );
  NAND2_X1 U9240 ( .A1(n7709), .A2(n8096), .ZN(n7711) );
  OR2_X1 U9241 ( .A1(n7710), .A2(n7713), .ZN(n8098) );
  NAND2_X1 U9242 ( .A1(n7711), .A2(n8098), .ZN(n7723) );
  XOR2_X1 U9243 ( .A(n7723), .B(n8196), .Z(n7712) );
  OAI222_X1 U9244 ( .A1(n9425), .A2(n7891), .B1(n9423), .B2(n7713), .C1(n9421), 
        .C2(n7712), .ZN(n7829) );
  AOI211_X1 U9245 ( .C1(n7894), .C2(n7714), .A(n10265), .B(n4540), .ZN(n7830)
         );
  INV_X1 U9246 ( .A(n10003), .ZN(n7715) );
  NAND2_X1 U9247 ( .A1(n7830), .A2(n7715), .ZN(n7717) );
  AOI22_X1 U9248 ( .A1(n10216), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7893), .B2(
        n9993), .ZN(n7716) );
  OAI211_X1 U9249 ( .C1(n4803), .C2(n9432), .A(n7717), .B(n7716), .ZN(n7718)
         );
  AOI21_X1 U9250 ( .B1(n7829), .B2(n10207), .A(n7718), .ZN(n7719) );
  OAI21_X1 U9251 ( .B1(n10004), .B2(n7832), .A(n7719), .ZN(P1_U3279) );
  NAND2_X1 U9252 ( .A1(n7894), .A2(n9178), .ZN(n7721) );
  OR2_X1 U9253 ( .A1(n7907), .A2(n7891), .ZN(n8109) );
  NAND2_X1 U9254 ( .A1(n7907), .A2(n7891), .ZN(n8247) );
  XNOR2_X1 U9255 ( .A(n7844), .B(n8199), .ZN(n10034) );
  INV_X1 U9256 ( .A(n8099), .ZN(n7722) );
  NAND2_X1 U9257 ( .A1(n7724), .A2(n8199), .ZN(n7866) );
  OAI21_X1 U9258 ( .B1(n8199), .B2(n7724), .A(n7866), .ZN(n7725) );
  NAND2_X1 U9259 ( .A1(n7725), .A2(n9985), .ZN(n7727) );
  AOI22_X1 U9260 ( .A1(n9988), .A2(n9178), .B1(n9990), .B2(n9176), .ZN(n7726)
         );
  NAND2_X1 U9261 ( .A1(n7727), .A2(n7726), .ZN(n7728) );
  AOI21_X1 U9262 ( .B1(n10034), .B2(n7961), .A(n7728), .ZN(n10036) );
  INV_X1 U9263 ( .A(n7907), .ZN(n10031) );
  NOR2_X1 U9264 ( .A1(n4540), .A2(n10031), .ZN(n7729) );
  OR2_X1 U9265 ( .A1(n7841), .A2(n7729), .ZN(n10032) );
  AOI22_X1 U9266 ( .A1(n10216), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7902), .B2(
        n9993), .ZN(n7731) );
  NAND2_X1 U9267 ( .A1(n7907), .A2(n10213), .ZN(n7730) );
  OAI211_X1 U9268 ( .C1(n10032), .C2(n7973), .A(n7731), .B(n7730), .ZN(n7732)
         );
  AOI21_X1 U9269 ( .B1(n10034), .B2(n7968), .A(n7732), .ZN(n7733) );
  OAI21_X1 U9270 ( .B1(n10036), .B2(n10216), .A(n7733), .ZN(P1_U3278) );
  INV_X1 U9271 ( .A(n7735), .ZN(n7736) );
  AOI22_X1 U9272 ( .A1(n8858), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7736), .B2(
        n8856), .ZN(n7737) );
  OAI21_X1 U9273 ( .B1(n4758), .B2(n8861), .A(n7737), .ZN(n7740) );
  NOR2_X1 U9274 ( .A1(n7738), .A2(n8858), .ZN(n7739) );
  AOI211_X1 U9275 ( .C1(n7741), .C2(n8891), .A(n7740), .B(n7739), .ZN(n7742)
         );
  OAI21_X1 U9276 ( .B1(n8865), .B2(n7743), .A(n7742), .ZN(P2_U3285) );
  NAND2_X1 U9277 ( .A1(n7748), .A2(n7950), .ZN(n7745) );
  OR2_X1 U9278 ( .A1(n7744), .A2(P1_U3084), .ZN(n8351) );
  OAI211_X1 U9279 ( .C1(n7746), .C2(n9890), .A(n7745), .B(n8351), .ZN(P1_U3330) );
  NAND2_X1 U9280 ( .A1(n7748), .A2(n7747), .ZN(n7750) );
  OAI211_X1 U9281 ( .C1(n7751), .C2(n9018), .A(n7750), .B(n7749), .ZN(P2_U3335) );
  INV_X1 U9282 ( .A(n8977), .ZN(n7815) );
  XNOR2_X1 U9283 ( .A(n8977), .B(n8429), .ZN(n7752) );
  NAND2_X1 U9284 ( .A1(n8557), .A2(n8430), .ZN(n7753) );
  NAND2_X1 U9285 ( .A1(n7752), .A2(n7753), .ZN(n7801) );
  INV_X1 U9286 ( .A(n7752), .ZN(n7755) );
  INV_X1 U9287 ( .A(n7753), .ZN(n7754) );
  NAND2_X1 U9288 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  AND2_X1 U9289 ( .A1(n7801), .A2(n7756), .ZN(n7764) );
  INV_X1 U9290 ( .A(n7759), .ZN(n7762) );
  INV_X1 U9291 ( .A(n7760), .ZN(n7761) );
  OAI21_X1 U9292 ( .B1(n7764), .B2(n7763), .A(n7802), .ZN(n7765) );
  NAND2_X1 U9293 ( .A1(n7765), .A2(n8539), .ZN(n7771) );
  INV_X1 U9294 ( .A(n7766), .ZN(n7813) );
  OAI22_X1 U9295 ( .A1(n7921), .A2(n8530), .B1(n8531), .B2(n7767), .ZN(n7768)
         );
  AOI211_X1 U9296 ( .C1(n8548), .C2(n7813), .A(n7769), .B(n7768), .ZN(n7770)
         );
  OAI211_X1 U9297 ( .C1(n7815), .C2(n8551), .A(n7771), .B(n7770), .ZN(P2_U3217) );
  OAI211_X1 U9298 ( .C1(n4488), .C2(n7773), .A(n7772), .B(n9115), .ZN(n7780)
         );
  AOI21_X1 U9299 ( .B1(n9138), .B2(n9178), .A(n7774), .ZN(n7775) );
  OAI21_X1 U9300 ( .B1(n9141), .B2(n7776), .A(n7775), .ZN(n7777) );
  AOI21_X1 U9301 ( .B1(n7778), .B2(n9166), .A(n7777), .ZN(n7779) );
  OAI211_X1 U9302 ( .C1(n10037), .C2(n9123), .A(n7780), .B(n7779), .ZN(
        P1_U3234) );
  OR2_X1 U9303 ( .A1(n7781), .A2(n8559), .ZN(n7782) );
  AOI21_X1 U9304 ( .B1(n7785), .B2(n7784), .A(n4529), .ZN(n8983) );
  XNOR2_X1 U9305 ( .A(n7786), .B(n4642), .ZN(n7788) );
  AOI22_X1 U9306 ( .A1(n8871), .A2(n8559), .B1(n8557), .B2(n8873), .ZN(n7787)
         );
  OAI21_X1 U9307 ( .B1(n7788), .B2(n8847), .A(n7787), .ZN(n7789) );
  AOI21_X1 U9308 ( .B1(n8983), .B2(n7790), .A(n7789), .ZN(n8988) );
  INV_X1 U9309 ( .A(n7812), .ZN(n7791) );
  AOI21_X1 U9310 ( .B1(n8984), .B2(n7792), .A(n7791), .ZN(n8986) );
  INV_X1 U9311 ( .A(n8984), .ZN(n7793) );
  NOR2_X1 U9312 ( .A1(n7793), .A2(n8861), .ZN(n7797) );
  OAI22_X1 U9313 ( .A1(n8896), .A2(n7795), .B1(n7794), .B2(n8882), .ZN(n7796)
         );
  AOI211_X1 U9314 ( .C1(n8986), .C2(n8891), .A(n7797), .B(n7796), .ZN(n7800)
         );
  NAND2_X1 U9315 ( .A1(n8983), .A2(n7798), .ZN(n7799) );
  OAI211_X1 U9316 ( .C1(n8988), .C2(n8858), .A(n7800), .B(n7799), .ZN(P2_U3283) );
  AND2_X1 U9317 ( .A1(n8872), .A2(n8430), .ZN(n7915) );
  XNOR2_X1 U9318 ( .A(n8972), .B(n8429), .ZN(n7917) );
  XOR2_X1 U9319 ( .A(n7915), .B(n7917), .Z(n7803) );
  XNOR2_X1 U9320 ( .A(n7916), .B(n7803), .ZN(n7809) );
  OAI22_X1 U9321 ( .A1(n8522), .A2(n7854), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7804), .ZN(n7807) );
  OAI22_X1 U9322 ( .A1(n7805), .A2(n8531), .B1(n8530), .B2(n8849), .ZN(n7806)
         );
  AOI211_X1 U9323 ( .C1(n8972), .C2(n4453), .A(n7807), .B(n7806), .ZN(n7808)
         );
  OAI21_X1 U9324 ( .B1(n7809), .B2(n8537), .A(n7808), .ZN(P2_U3243) );
  NAND2_X1 U9325 ( .A1(n8984), .A2(n8558), .ZN(n7810) );
  XNOR2_X1 U9326 ( .A(n7859), .B(n7811), .ZN(n8982) );
  AOI21_X1 U9327 ( .B1(n8977), .B2(n7812), .A(n7851), .ZN(n8978) );
  AOI22_X1 U9328 ( .A1(n8858), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7813), .B2(
        n8856), .ZN(n7814) );
  OAI21_X1 U9329 ( .B1(n7815), .B2(n8861), .A(n7814), .ZN(n7821) );
  OAI211_X1 U9330 ( .C1(n7817), .C2(n7858), .A(n7816), .B(n8878), .ZN(n7819)
         );
  AOI22_X1 U9331 ( .A1(n8873), .A2(n8872), .B1(n8558), .B2(n8871), .ZN(n7818)
         );
  AND2_X1 U9332 ( .A1(n7819), .A2(n7818), .ZN(n8980) );
  NOR2_X1 U9333 ( .A1(n8980), .A2(n8858), .ZN(n7820) );
  AOI211_X1 U9334 ( .C1(n8978), .C2(n8891), .A(n7821), .B(n7820), .ZN(n7822)
         );
  OAI21_X1 U9335 ( .B1(n8865), .B2(n8982), .A(n7822), .ZN(P2_U3282) );
  INV_X1 U9336 ( .A(n7823), .ZN(n7827) );
  OAI222_X1 U9337 ( .A1(P2_U3152), .A2(n7825), .B1(n8454), .B2(n7827), .C1(
        n7824), .C2(n9018), .ZN(P2_U3334) );
  OAI222_X1 U9338 ( .A1(P1_U3084), .A2(n7828), .B1(n4459), .B2(n7827), .C1(
        n7826), .C2(n9890), .ZN(P1_U3329) );
  AOI211_X1 U9339 ( .C1(n9511), .C2(n7894), .A(n7830), .B(n7829), .ZN(n7831)
         );
  OAI21_X1 U9340 ( .B1(n10016), .B2(n7832), .A(n7831), .ZN(n7834) );
  NAND2_X1 U9341 ( .A1(n7834), .A2(n4456), .ZN(n7833) );
  OAI21_X1 U9342 ( .B1(n4456), .B2(n9202), .A(n7833), .ZN(P1_U3535) );
  INV_X1 U9343 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U9344 ( .A1(n7834), .A2(n10273), .ZN(n7835) );
  OAI21_X1 U9345 ( .B1(n10273), .B2(n7836), .A(n7835), .ZN(P1_U3490) );
  INV_X1 U9346 ( .A(n9176), .ZN(n7905) );
  NAND2_X1 U9347 ( .A1(n7941), .A2(n7905), .ZN(n8252) );
  NAND2_X1 U9348 ( .A1(n8250), .A2(n8252), .ZN(n8201) );
  NAND2_X1 U9349 ( .A1(n7866), .A2(n8247), .ZN(n7837) );
  XOR2_X1 U9350 ( .A(n8201), .B(n7837), .Z(n7838) );
  AOI222_X1 U9351 ( .A1(n9985), .A2(n7838), .B1(n9987), .B2(n9990), .C1(n9177), 
        .C2(n9988), .ZN(n10026) );
  INV_X1 U9352 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7840) );
  INV_X1 U9353 ( .A(n7936), .ZN(n7839) );
  OAI22_X1 U9354 ( .A1(n10207), .A2(n7840), .B1(n7839), .B2(n10221), .ZN(n7843) );
  INV_X1 U9355 ( .A(n7941), .ZN(n10027) );
  NAND2_X1 U9356 ( .A1(n7841), .A2(n10027), .ZN(n7872) );
  OAI211_X1 U9357 ( .C1(n7841), .C2(n10027), .A(n9999), .B(n7872), .ZN(n10025)
         );
  NOR2_X1 U9358 ( .A1(n10025), .A2(n10003), .ZN(n7842) );
  AOI211_X1 U9359 ( .C1(n10213), .C2(n7941), .A(n7843), .B(n7842), .ZN(n7848)
         );
  OR2_X1 U9360 ( .A1(n7907), .A2(n9177), .ZN(n7845) );
  XNOR2_X1 U9361 ( .A(n7877), .B(n8201), .ZN(n10029) );
  NAND2_X1 U9362 ( .A1(n10029), .A2(n7881), .ZN(n7847) );
  OAI211_X1 U9363 ( .C1(n10026), .C2(n10216), .A(n7848), .B(n7847), .ZN(
        P1_U3277) );
  XNOR2_X1 U9364 ( .A(n7849), .B(n7860), .ZN(n7850) );
  AOI222_X1 U9365 ( .A1(n8878), .A2(n7850), .B1(n8556), .B2(n8873), .C1(n8557), 
        .C2(n8871), .ZN(n8975) );
  INV_X1 U9366 ( .A(n7851), .ZN(n7852) );
  INV_X1 U9367 ( .A(n8972), .ZN(n7853) );
  AOI21_X1 U9368 ( .B1(n8972), .B2(n7852), .A(n8888), .ZN(n8973) );
  NOR2_X1 U9369 ( .A1(n7853), .A2(n8861), .ZN(n7857) );
  OAI22_X1 U9370 ( .A1(n8896), .A2(n7855), .B1(n7854), .B2(n8882), .ZN(n7856)
         );
  AOI211_X1 U9371 ( .C1(n8973), .C2(n8891), .A(n7857), .B(n7856), .ZN(n7863)
         );
  OAI21_X1 U9372 ( .B1(n7861), .B2(n7860), .A(n7986), .ZN(n8971) );
  NAND2_X1 U9373 ( .A1(n8971), .A2(n8760), .ZN(n7862) );
  OAI211_X1 U9374 ( .C1(n8975), .C2(n8858), .A(n7863), .B(n7862), .ZN(P2_U3281) );
  INV_X1 U9375 ( .A(n8247), .ZN(n7864) );
  NOR2_X1 U9376 ( .A1(n8201), .A2(n7864), .ZN(n7865) );
  NAND2_X1 U9377 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U9378 ( .A1(n7867), .A2(n8250), .ZN(n7868) );
  INV_X1 U9379 ( .A(n7868), .ZN(n7869) );
  INV_X1 U9380 ( .A(n9987), .ZN(n7939) );
  OR2_X1 U9381 ( .A1(n9169), .A2(n7939), .ZN(n8256) );
  NAND2_X1 U9382 ( .A1(n9169), .A2(n7939), .ZN(n8254) );
  OAI21_X1 U9383 ( .B1(n7869), .B2(n8203), .A(n4490), .ZN(n7870) );
  AOI222_X1 U9384 ( .A1(n9985), .A2(n7870), .B1(n9175), .B2(n9990), .C1(n9176), 
        .C2(n9988), .ZN(n10019) );
  INV_X1 U9385 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10142) );
  INV_X1 U9386 ( .A(n9167), .ZN(n7871) );
  OAI22_X1 U9387 ( .A1(n10207), .A2(n10142), .B1(n7871), .B2(n10221), .ZN(
        n7876) );
  INV_X1 U9388 ( .A(n7872), .ZN(n7873) );
  INV_X1 U9389 ( .A(n9169), .ZN(n10020) );
  OAI211_X1 U9390 ( .C1(n7873), .C2(n10020), .A(n9999), .B(n9998), .ZN(n10018)
         );
  NOR2_X1 U9391 ( .A1(n10018), .A2(n7874), .ZN(n7875) );
  AOI211_X1 U9392 ( .C1(n10213), .C2(n9169), .A(n7876), .B(n7875), .ZN(n7884)
         );
  OR2_X1 U9393 ( .A1(n7941), .A2(n9176), .ZN(n7878) );
  AND2_X1 U9394 ( .A1(n7879), .A2(n8203), .ZN(n10017) );
  INV_X1 U9395 ( .A(n10017), .ZN(n7882) );
  NAND3_X1 U9396 ( .A1(n7882), .A2(n7881), .A3(n10022), .ZN(n7883) );
  OAI211_X1 U9397 ( .C1(n10019), .C2(n10216), .A(n7884), .B(n7883), .ZN(
        P1_U3276) );
  INV_X1 U9398 ( .A(n7886), .ZN(n7887) );
  AOI21_X1 U9399 ( .B1(n7888), .B2(n7885), .A(n7887), .ZN(n7897) );
  NAND2_X1 U9400 ( .A1(n9162), .A2(n9179), .ZN(n7890) );
  OAI211_X1 U9401 ( .C1(n9164), .C2(n7891), .A(n7890), .B(n7889), .ZN(n7892)
         );
  AOI21_X1 U9402 ( .B1(n7893), .B2(n9166), .A(n7892), .ZN(n7896) );
  NAND2_X1 U9403 ( .A1(n7894), .A2(n9168), .ZN(n7895) );
  OAI211_X1 U9404 ( .C1(n7897), .C2(n9172), .A(n7896), .B(n7895), .ZN(P1_U3222) );
  XNOR2_X1 U9405 ( .A(n7900), .B(n7899), .ZN(n7901) );
  XNOR2_X1 U9406 ( .A(n7898), .B(n7901), .ZN(n7909) );
  NAND2_X1 U9407 ( .A1(n9166), .A2(n7902), .ZN(n7904) );
  NOR2_X1 U9408 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9728), .ZN(n10119) );
  AOI21_X1 U9409 ( .B1(n9162), .B2(n9178), .A(n10119), .ZN(n7903) );
  OAI211_X1 U9410 ( .C1(n7905), .C2(n9164), .A(n7904), .B(n7903), .ZN(n7906)
         );
  AOI21_X1 U9411 ( .B1(n7907), .B2(n9168), .A(n7906), .ZN(n7908) );
  OAI21_X1 U9412 ( .B1(n7909), .B2(n9172), .A(n7908), .ZN(P1_U3232) );
  INV_X1 U9413 ( .A(n8964), .ZN(n8887) );
  XNOR2_X1 U9414 ( .A(n8964), .B(n8429), .ZN(n7910) );
  NAND2_X1 U9415 ( .A1(n8556), .A2(n8430), .ZN(n7911) );
  NAND2_X1 U9416 ( .A1(n7910), .A2(n7911), .ZN(n8384) );
  INV_X1 U9417 ( .A(n7910), .ZN(n7913) );
  INV_X1 U9418 ( .A(n7911), .ZN(n7912) );
  NAND2_X1 U9419 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  AND2_X1 U9420 ( .A1(n8384), .A2(n7914), .ZN(n7919) );
  OAI21_X1 U9421 ( .B1(n7919), .B2(n7918), .A(n8385), .ZN(n7920) );
  NAND2_X1 U9422 ( .A1(n7920), .A2(n8539), .ZN(n7925) );
  INV_X1 U9423 ( .A(n8883), .ZN(n7923) );
  AND2_X1 U9424 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8622) );
  OAI22_X1 U9425 ( .A1(n7921), .A2(n8531), .B1(n8530), .B2(n8532), .ZN(n7922)
         );
  AOI211_X1 U9426 ( .C1(n7923), .C2(n8548), .A(n8622), .B(n7922), .ZN(n7924)
         );
  OAI211_X1 U9427 ( .C1(n8887), .C2(n8551), .A(n7925), .B(n7924), .ZN(P2_U3228) );
  INV_X1 U9428 ( .A(n7926), .ZN(n7930) );
  OAI222_X1 U9429 ( .A1(n9890), .A2(n7928), .B1(n4459), .B2(n7930), .C1(
        P1_U3084), .C2(n7927), .ZN(P1_U3328) );
  OAI222_X1 U9430 ( .A1(n9018), .A2(n7931), .B1(n8454), .B2(n7930), .C1(
        P2_U3152), .C2(n7929), .ZN(P2_U3333) );
  XNOR2_X1 U9431 ( .A(n7933), .B(n7932), .ZN(n7934) );
  XNOR2_X1 U9432 ( .A(n7935), .B(n7934), .ZN(n7943) );
  NAND2_X1 U9433 ( .A1(n9166), .A2(n7936), .ZN(n7938) );
  AND2_X1 U9434 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10131) );
  AOI21_X1 U9435 ( .B1(n9162), .B2(n9177), .A(n10131), .ZN(n7937) );
  OAI211_X1 U9436 ( .C1(n7939), .C2(n9164), .A(n7938), .B(n7937), .ZN(n7940)
         );
  AOI21_X1 U9437 ( .B1(n7941), .B2(n9168), .A(n7940), .ZN(n7942) );
  OAI21_X1 U9438 ( .B1(n7943), .B2(n9172), .A(n7942), .ZN(P1_U3213) );
  INV_X1 U9439 ( .A(n7944), .ZN(n7946) );
  INV_X1 U9440 ( .A(n7945), .ZN(n7948) );
  OAI222_X1 U9441 ( .A1(P1_U3084), .A2(n7946), .B1(n4459), .B2(n7948), .C1(
        n9658), .C2(n9890), .ZN(P1_U3327) );
  OAI222_X1 U9442 ( .A1(P2_U3152), .A2(n7949), .B1(n8454), .B2(n7948), .C1(
        n7947), .C2(n9018), .ZN(P2_U3332) );
  NAND2_X1 U9443 ( .A1(n7954), .A2(n7950), .ZN(n7952) );
  OAI211_X1 U9444 ( .C1(n9890), .C2(n7953), .A(n7952), .B(n7951), .ZN(P1_U3326) );
  INV_X1 U9445 ( .A(n7954), .ZN(n7955) );
  OAI222_X1 U9446 ( .A1(n9018), .A2(n7956), .B1(n8454), .B2(n7955), .C1(n6507), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  XNOR2_X1 U9447 ( .A(n7957), .B(n8184), .ZN(n7964) );
  OR2_X1 U9448 ( .A1(n7958), .A2(n8184), .ZN(n7959) );
  NAND2_X1 U9449 ( .A1(n7960), .A2(n7959), .ZN(n10239) );
  NAND2_X1 U9450 ( .A1(n10239), .A2(n7961), .ZN(n7963) );
  AOI22_X1 U9451 ( .A1(n9988), .A2(n6837), .B1(n9990), .B2(n9187), .ZN(n7962)
         );
  OAI211_X1 U9452 ( .C1(n7964), .C2(n9421), .A(n7963), .B(n7962), .ZN(n10237)
         );
  MUX2_X1 U9453 ( .A(n10237), .B(P1_REG2_REG_2__SCAN_IN), .S(n10216), .Z(n7975) );
  NOR2_X1 U9454 ( .A1(n7965), .A2(n10235), .ZN(n7966) );
  OR2_X1 U9455 ( .A1(n7967), .A2(n7966), .ZN(n10236) );
  NAND2_X1 U9456 ( .A1(n10239), .A2(n7968), .ZN(n7972) );
  INV_X1 U9457 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7969) );
  OAI22_X1 U9458 ( .A1(n9432), .A2(n10235), .B1(n7969), .B2(n10221), .ZN(n7970) );
  INV_X1 U9459 ( .A(n7970), .ZN(n7971) );
  OAI211_X1 U9460 ( .C1(n7973), .C2(n10236), .A(n7972), .B(n7971), .ZN(n7974)
         );
  OR2_X1 U9461 ( .A1(n7975), .A2(n7974), .ZN(P1_U3289) );
  INV_X1 U9462 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8452) );
  NOR2_X1 U9463 ( .A1(n8161), .A2(n8452), .ZN(n7976) );
  INV_X1 U9464 ( .A(n9443), .ZN(n8078) );
  INV_X1 U9465 ( .A(n9460), .ZN(n9270) );
  INV_X1 U9466 ( .A(n9471), .ZN(n9310) );
  INV_X1 U9467 ( .A(n9510), .ZN(n9433) );
  INV_X1 U9468 ( .A(n9503), .ZN(n9407) );
  INV_X1 U9469 ( .A(n9489), .ZN(n9359) );
  NAND2_X1 U9470 ( .A1(n8449), .A2(n8163), .ZN(n7979) );
  INV_X1 U9471 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7977) );
  OR2_X1 U9472 ( .A1(n8161), .A2(n7977), .ZN(n7978) );
  INV_X1 U9473 ( .A(n9451), .ZN(n9241) );
  NAND2_X1 U9474 ( .A1(n9017), .A2(n8163), .ZN(n7981) );
  OR2_X1 U9475 ( .A1(n8161), .A2(n9889), .ZN(n7980) );
  INV_X1 U9476 ( .A(n8036), .ZN(n7982) );
  NAND2_X1 U9477 ( .A1(n8078), .A2(n7982), .ZN(n9440) );
  NAND2_X1 U9478 ( .A1(n9443), .A2(n8036), .ZN(n9439) );
  NAND3_X1 U9479 ( .A1(n9440), .A2(n10212), .A3(n9439), .ZN(n7984) );
  INV_X1 U9480 ( .A(n8349), .ZN(n10075) );
  AOI21_X1 U9481 ( .B1(n10075), .B2(P1_B_REG_SCAN_IN), .A(n9425), .ZN(n8050)
         );
  NAND2_X1 U9482 ( .A1(n8050), .A2(n8173), .ZN(n9441) );
  NOR2_X1 U9483 ( .A1(n9441), .A2(n10216), .ZN(n8357) );
  AOI21_X1 U9484 ( .B1(n10216), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8357), .ZN(
        n7983) );
  OAI211_X1 U9485 ( .C1(n9443), .C2(n9432), .A(n7984), .B(n7983), .ZN(P1_U3262) );
  INV_X1 U9486 ( .A(n8930), .ZN(n8764) );
  OR2_X1 U9487 ( .A1(n8972), .A2(n8872), .ZN(n7985) );
  NAND2_X1 U9488 ( .A1(n8954), .A2(n8555), .ZN(n7987) );
  INV_X1 U9489 ( .A(n8954), .ZN(n8833) );
  INV_X1 U9490 ( .A(n8951), .ZN(n7989) );
  INV_X1 U9491 ( .A(n8777), .ZN(n7992) );
  INV_X1 U9492 ( .A(n8747), .ZN(n8741) );
  INV_X1 U9493 ( .A(n8924), .ZN(n8746) );
  INV_X1 U9494 ( .A(n8750), .ZN(n8554) );
  AOI22_X1 U9495 ( .A1(n8712), .A2(n7995), .B1(n8725), .B2(n8704), .ZN(n8696)
         );
  OAI22_X1 U9496 ( .A1(n8696), .A2(n7996), .B1(n8909), .B2(n8552), .ZN(n8366)
         );
  XNOR2_X1 U9497 ( .A(n8366), .B(n7997), .ZN(n8908) );
  INV_X1 U9498 ( .A(n8944), .ZN(n8807) );
  NAND2_X1 U9499 ( .A1(n8822), .A2(n8807), .ZN(n8801) );
  NAND2_X1 U9500 ( .A1(n8725), .A2(n8733), .ZN(n8719) );
  INV_X1 U9501 ( .A(n8697), .ZN(n7999) );
  INV_X1 U9502 ( .A(n8904), .ZN(n8364) );
  INV_X1 U9503 ( .A(n8375), .ZN(n7998) );
  AOI21_X1 U9504 ( .B1(n8904), .B2(n7999), .A(n7998), .ZN(n8905) );
  AOI22_X1 U9505 ( .A1(n8858), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8440), .B2(
        n8856), .ZN(n8000) );
  OAI21_X1 U9506 ( .B1(n8364), .B2(n8861), .A(n8000), .ZN(n8006) );
  AOI211_X1 U9507 ( .C1(n8002), .C2(n8365), .A(n8847), .B(n8001), .ZN(n8004)
         );
  OAI22_X1 U9508 ( .A1(n8444), .A2(n8852), .B1(n8443), .B2(n8850), .ZN(n8003)
         );
  NOR2_X1 U9509 ( .A1(n8004), .A2(n8003), .ZN(n8907) );
  NOR2_X1 U9510 ( .A1(n8907), .A2(n8858), .ZN(n8005) );
  AOI211_X1 U9511 ( .C1(n8891), .C2(n8905), .A(n8006), .B(n8005), .ZN(n8007)
         );
  OAI21_X1 U9512 ( .B1(n8908), .B2(n8865), .A(n8007), .ZN(P2_U3268) );
  NAND2_X1 U9513 ( .A1(n9169), .A2(n9987), .ZN(n8008) );
  NAND2_X1 U9514 ( .A1(n10022), .A2(n8008), .ZN(n9997) );
  INV_X1 U9515 ( .A(n9175), .ZN(n9422) );
  NAND2_X1 U9516 ( .A1(n10009), .A2(n9422), .ZN(n8259) );
  NAND2_X1 U9517 ( .A1(n8257), .A2(n8259), .ZN(n9996) );
  NAND2_X1 U9518 ( .A1(n10009), .A2(n9175), .ZN(n8009) );
  OR2_X1 U9519 ( .A1(n9510), .A2(n9989), .ZN(n8010) );
  INV_X1 U9520 ( .A(n9395), .ZN(n9424) );
  OR2_X1 U9521 ( .A1(n9503), .A2(n9424), .ZN(n8122) );
  NAND2_X1 U9522 ( .A1(n9503), .A2(n9424), .ZN(n8262) );
  NAND2_X1 U9523 ( .A1(n8122), .A2(n8262), .ZN(n9410) );
  AND2_X1 U9524 ( .A1(n9493), .A2(n9396), .ZN(n8015) );
  OR2_X1 U9525 ( .A1(n9498), .A2(n9412), .ZN(n9371) );
  OR2_X1 U9526 ( .A1(n8015), .A2(n9371), .ZN(n8013) );
  AND2_X1 U9527 ( .A1(n9410), .A2(n8013), .ZN(n8011) );
  OR2_X1 U9528 ( .A1(n9493), .A2(n9396), .ZN(n8012) );
  AND2_X1 U9529 ( .A1(n8011), .A2(n8012), .ZN(n9347) );
  INV_X1 U9530 ( .A(n9381), .ZN(n9337) );
  OR2_X1 U9531 ( .A1(n9489), .A2(n9337), .ZN(n8268) );
  NAND2_X1 U9532 ( .A1(n9489), .A2(n9337), .ZN(n8133) );
  INV_X1 U9533 ( .A(n9363), .ZN(n9351) );
  AND2_X1 U9534 ( .A1(n9347), .A2(n9351), .ZN(n8021) );
  INV_X1 U9535 ( .A(n8012), .ZN(n8020) );
  INV_X1 U9536 ( .A(n8013), .ZN(n8018) );
  NAND2_X1 U9537 ( .A1(n9503), .A2(n9395), .ZN(n9386) );
  NAND2_X1 U9538 ( .A1(n9498), .A2(n9412), .ZN(n8014) );
  AND2_X1 U9539 ( .A1(n9386), .A2(n8014), .ZN(n9370) );
  INV_X1 U9540 ( .A(n8015), .ZN(n8016) );
  AND2_X1 U9541 ( .A1(n9370), .A2(n8016), .ZN(n8017) );
  OR2_X1 U9542 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  NAND2_X1 U9543 ( .A1(n9489), .A2(n9381), .ZN(n8022) );
  NAND2_X1 U9544 ( .A1(n9350), .A2(n8022), .ZN(n9333) );
  OR2_X1 U9545 ( .A1(n9485), .A2(n9365), .ZN(n8023) );
  NAND2_X1 U9546 ( .A1(n9485), .A2(n9365), .ZN(n8024) );
  OR2_X1 U9547 ( .A1(n9480), .A2(n9305), .ZN(n8025) );
  NAND2_X1 U9548 ( .A1(n8026), .A2(n8025), .ZN(n9296) );
  INV_X1 U9549 ( .A(n9290), .ZN(n9325) );
  NAND2_X1 U9550 ( .A1(n9471), .A2(n9325), .ZN(n8141) );
  NOR2_X1 U9551 ( .A1(n9296), .A2(n9302), .ZN(n9298) );
  INV_X1 U9552 ( .A(n9306), .ZN(n9104) );
  NAND2_X1 U9553 ( .A1(n9465), .A2(n9104), .ZN(n8146) );
  NAND2_X1 U9554 ( .A1(n9271), .A2(n8146), .ZN(n9288) );
  NOR2_X1 U9555 ( .A1(n9460), .A2(n9291), .ZN(n8211) );
  NAND2_X1 U9556 ( .A1(n9460), .A2(n9291), .ZN(n8209) );
  OR2_X1 U9557 ( .A1(n9253), .A2(n9275), .ZN(n8283) );
  NAND2_X1 U9558 ( .A1(n9253), .A2(n9275), .ZN(n9242) );
  OAI22_X1 U9559 ( .A1(n9249), .A2(n9255), .B1(n9455), .B2(n9275), .ZN(n9234)
         );
  INV_X1 U9560 ( .A(n9257), .ZN(n8028) );
  OR2_X1 U9561 ( .A1(n9451), .A2(n8028), .ZN(n8286) );
  NAND2_X1 U9562 ( .A1(n9451), .A2(n8028), .ZN(n8284) );
  NOR2_X1 U9563 ( .A1(n9234), .A2(n9244), .ZN(n9233) );
  AOI21_X1 U9564 ( .B1(n9257), .B2(n9451), .A(n9233), .ZN(n8035) );
  NAND2_X1 U9565 ( .A1(n8046), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U9566 ( .A1(n6600), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U9567 ( .A1(n5184), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8029) );
  AND3_X1 U9568 ( .A1(n8031), .A2(n8030), .A3(n8029), .ZN(n8032) );
  OAI21_X1 U9569 ( .B1(n8037), .B2(n5734), .A(n8032), .ZN(n9246) );
  INV_X1 U9570 ( .A(n9246), .ZN(n8033) );
  NAND2_X1 U9571 ( .A1(n9444), .A2(n8033), .ZN(n8299) );
  NAND2_X1 U9572 ( .A1(n8287), .A2(n8299), .ZN(n8214) );
  XNOR2_X1 U9573 ( .A(n8035), .B(n8034), .ZN(n9449) );
  AOI21_X1 U9574 ( .B1(n9444), .B2(n9236), .A(n8036), .ZN(n9445) );
  INV_X1 U9575 ( .A(n8037), .ZN(n8038) );
  AOI22_X1 U9576 ( .A1(n8038), .A2(n9993), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10216), .ZN(n8039) );
  OAI21_X1 U9577 ( .B1(n4796), .B2(n9432), .A(n8039), .ZN(n8056) );
  INV_X1 U9578 ( .A(n8259), .ZN(n8040) );
  INV_X1 U9579 ( .A(n9989), .ZN(n9142) );
  NAND2_X1 U9580 ( .A1(n9510), .A2(n9142), .ZN(n8260) );
  OR2_X1 U9581 ( .A1(n9510), .A2(n9142), .ZN(n9408) );
  AND2_X1 U9582 ( .A1(n8122), .A2(n9408), .ZN(n8271) );
  NAND2_X1 U9583 ( .A1(n9409), .A2(n8271), .ZN(n8041) );
  NAND2_X1 U9584 ( .A1(n8041), .A2(n8262), .ZN(n9393) );
  INV_X1 U9585 ( .A(n9412), .ZN(n9119) );
  OR2_X1 U9586 ( .A1(n9498), .A2(n9119), .ZN(n8126) );
  NAND2_X1 U9587 ( .A1(n9498), .A2(n9119), .ZN(n8125) );
  INV_X1 U9588 ( .A(n9396), .ZN(n9041) );
  AND2_X1 U9589 ( .A1(n9493), .A2(n9041), .ZN(n8179) );
  NOR2_X1 U9590 ( .A1(n9493), .A2(n9041), .ZN(n8180) );
  NOR2_X1 U9591 ( .A1(n9351), .A2(n8180), .ZN(n8042) );
  NAND2_X1 U9592 ( .A1(n9361), .A2(n8042), .ZN(n9362) );
  NAND2_X1 U9593 ( .A1(n9362), .A2(n8133), .ZN(n9335) );
  INV_X1 U9594 ( .A(n9365), .ZN(n9324) );
  NAND2_X1 U9595 ( .A1(n9335), .A2(n8274), .ZN(n9321) );
  NAND2_X1 U9596 ( .A1(n9485), .A2(n9324), .ZN(n8178) );
  INV_X1 U9597 ( .A(n9305), .ZN(n9338) );
  XNOR2_X1 U9598 ( .A(n9480), .B(n9338), .ZN(n9318) );
  NAND2_X1 U9599 ( .A1(n9480), .A2(n9338), .ZN(n9300) );
  NAND2_X1 U9600 ( .A1(n8141), .A2(n9300), .ZN(n8139) );
  INV_X1 U9601 ( .A(n9291), .ZN(n8044) );
  OR2_X1 U9602 ( .A1(n9460), .A2(n8044), .ZN(n8043) );
  AND2_X1 U9603 ( .A1(n8043), .A2(n9271), .ZN(n8329) );
  AND2_X1 U9604 ( .A1(n9460), .A2(n8044), .ZN(n8281) );
  NAND2_X1 U9605 ( .A1(n9256), .A2(n9255), .ZN(n9254) );
  NAND3_X1 U9606 ( .A1(n9254), .A2(n9244), .A3(n9242), .ZN(n9243) );
  NAND2_X1 U9607 ( .A1(n9243), .A2(n8284), .ZN(n8045) );
  NAND2_X1 U9608 ( .A1(n9257), .A2(n9988), .ZN(n8052) );
  NAND2_X1 U9609 ( .A1(n5184), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9610 ( .A1(n6600), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U9611 ( .A1(n8046), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8047) );
  NAND3_X1 U9612 ( .A1(n8049), .A2(n8048), .A3(n8047), .ZN(n9174) );
  NAND2_X1 U9613 ( .A1(n8050), .A2(n9174), .ZN(n8051) );
  NOR2_X1 U9614 ( .A1(n9447), .A2(n10216), .ZN(n8055) );
  OAI21_X1 U9615 ( .B1(n9449), .B2(n10004), .A(n8057), .ZN(P1_U3355) );
  XNOR2_X1 U9616 ( .A(n8058), .B(n8059), .ZN(n8066) );
  AOI22_X1 U9617 ( .A1(n8061), .A2(n6786), .B1(n8060), .B2(n6946), .ZN(n8065)
         );
  AOI22_X1 U9618 ( .A1(n4453), .A2(n8063), .B1(n8062), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8064) );
  OAI211_X1 U9619 ( .C1(n8066), .C2(n8537), .A(n8065), .B(n8064), .ZN(P2_U3239) );
  INV_X1 U9620 ( .A(n8067), .ZN(n8362) );
  OAI222_X1 U9621 ( .A1(n9018), .A2(n8068), .B1(n8454), .B2(n8362), .C1(n6463), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI21_X1 U9622 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n10077) );
  INV_X1 U9623 ( .A(n10077), .ZN(n8076) );
  OAI22_X1 U9624 ( .A1(n9164), .A2(n6838), .B1(n9123), .B2(n8072), .ZN(n8073)
         );
  AOI21_X1 U9625 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8074), .A(n8073), .ZN(
        n8075) );
  OAI21_X1 U9626 ( .B1(n8076), .B2(n9172), .A(n8075), .ZN(P1_U3230) );
  NAND2_X1 U9627 ( .A1(n9174), .A2(n8173), .ZN(n8077) );
  NAND2_X1 U9628 ( .A1(n8078), .A2(n8077), .ZN(n8288) );
  INV_X1 U9629 ( .A(n8170), .ZN(n8158) );
  NAND2_X1 U9630 ( .A1(n8084), .A2(n8314), .ZN(n8080) );
  INV_X1 U9631 ( .A(n8232), .ZN(n8079) );
  NAND2_X1 U9632 ( .A1(n8314), .A2(n8079), .ZN(n8229) );
  AND2_X1 U9633 ( .A1(n8229), .A2(n8081), .ZN(n8320) );
  AND2_X1 U9634 ( .A1(n8081), .A2(n8319), .ZN(n8236) );
  NAND2_X1 U9635 ( .A1(n8083), .A2(n8082), .ZN(n8224) );
  AOI21_X1 U9636 ( .B1(n8084), .B2(n8236), .A(n8224), .ZN(n8085) );
  AND2_X1 U9637 ( .A1(n8091), .A2(n8086), .ZN(n8242) );
  NAND2_X1 U9638 ( .A1(n8090), .A2(n8242), .ZN(n8087) );
  NAND3_X1 U9639 ( .A1(n8087), .A2(n8194), .A3(n8222), .ZN(n8088) );
  NAND3_X1 U9640 ( .A1(n8088), .A2(n8099), .A3(n8241), .ZN(n8095) );
  NAND2_X1 U9641 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  NAND3_X1 U9642 ( .A1(n8092), .A2(n8194), .A3(n8091), .ZN(n8093) );
  NAND2_X1 U9643 ( .A1(n8093), .A2(n8223), .ZN(n8094) );
  NAND2_X1 U9644 ( .A1(n8100), .A2(n8197), .ZN(n8107) );
  NAND2_X1 U9645 ( .A1(n8252), .A2(n8247), .ZN(n8226) );
  NAND2_X1 U9646 ( .A1(n8100), .A2(n8096), .ZN(n8246) );
  AND2_X1 U9647 ( .A1(n8246), .A2(n8099), .ZN(n8097) );
  OR2_X1 U9648 ( .A1(n8226), .A2(n8097), .ZN(n8104) );
  NAND2_X1 U9649 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  NAND2_X1 U9650 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  AND2_X1 U9651 ( .A1(n8109), .A2(n8102), .ZN(n8240) );
  NAND2_X1 U9652 ( .A1(n8250), .A2(n8240), .ZN(n8103) );
  MUX2_X1 U9653 ( .A(n8104), .B(n8103), .S(n8170), .Z(n8105) );
  INV_X1 U9654 ( .A(n8105), .ZN(n8106) );
  NAND2_X1 U9655 ( .A1(n8250), .A2(n8109), .ZN(n8110) );
  NAND2_X1 U9656 ( .A1(n8110), .A2(n8252), .ZN(n8112) );
  NAND2_X1 U9657 ( .A1(n8226), .A2(n8250), .ZN(n8111) );
  MUX2_X1 U9658 ( .A(n8112), .B(n8111), .S(n8170), .Z(n8113) );
  NAND3_X1 U9659 ( .A1(n8114), .A2(n8203), .A3(n8113), .ZN(n8116) );
  INV_X1 U9660 ( .A(n9996), .ZN(n9983) );
  MUX2_X1 U9661 ( .A(n8256), .B(n8254), .S(n8158), .Z(n8115) );
  NAND3_X1 U9662 ( .A1(n8116), .A2(n9983), .A3(n8115), .ZN(n8118) );
  MUX2_X1 U9663 ( .A(n8257), .B(n8259), .S(n8170), .Z(n8117) );
  NAND3_X1 U9664 ( .A1(n8118), .A2(n9418), .A3(n8117), .ZN(n8121) );
  AND2_X1 U9665 ( .A1(n8262), .A2(n8260), .ZN(n8119) );
  MUX2_X1 U9666 ( .A(n8271), .B(n8119), .S(n8158), .Z(n8120) );
  NAND2_X1 U9667 ( .A1(n8121), .A2(n8120), .ZN(n8128) );
  AND2_X1 U9668 ( .A1(n8126), .A2(n8122), .ZN(n8124) );
  INV_X1 U9669 ( .A(n8125), .ZN(n8221) );
  OR2_X1 U9670 ( .A1(n8179), .A2(n8221), .ZN(n8123) );
  AOI21_X1 U9671 ( .B1(n8128), .B2(n8124), .A(n8123), .ZN(n8130) );
  AND2_X1 U9672 ( .A1(n8125), .A2(n8262), .ZN(n8266) );
  INV_X1 U9673 ( .A(n8126), .ZN(n8127) );
  OR2_X1 U9674 ( .A1(n8180), .A2(n8127), .ZN(n8267) );
  AOI21_X1 U9675 ( .B1(n8128), .B2(n8266), .A(n8267), .ZN(n8129) );
  INV_X1 U9676 ( .A(n8180), .ZN(n9360) );
  NAND2_X1 U9677 ( .A1(n9360), .A2(n8268), .ZN(n8131) );
  INV_X1 U9678 ( .A(n8178), .ZN(n9319) );
  NAND2_X1 U9679 ( .A1(n8268), .A2(n8179), .ZN(n8134) );
  AND2_X1 U9680 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  AND2_X1 U9681 ( .A1(n8178), .A2(n8135), .ZN(n8273) );
  INV_X1 U9682 ( .A(n8274), .ZN(n8136) );
  OR2_X1 U9683 ( .A1(n9480), .A2(n9338), .ZN(n8137) );
  NAND2_X1 U9684 ( .A1(n8138), .A2(n8137), .ZN(n8277) );
  NAND2_X1 U9685 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  NAND2_X1 U9686 ( .A1(n8146), .A2(n8140), .ZN(n8330) );
  NAND2_X1 U9687 ( .A1(n8277), .A2(n8141), .ZN(n8142) );
  NAND2_X1 U9688 ( .A1(n9271), .A2(n8142), .ZN(n8143) );
  MUX2_X1 U9689 ( .A(n8330), .B(n8143), .S(n8170), .Z(n8144) );
  INV_X1 U9690 ( .A(n8144), .ZN(n8145) );
  MUX2_X1 U9691 ( .A(n9291), .B(n9460), .S(n8158), .Z(n8152) );
  INV_X1 U9692 ( .A(n9271), .ZN(n8147) );
  MUX2_X1 U9693 ( .A(n8147), .B(n4826), .S(n8170), .Z(n8150) );
  MUX2_X1 U9694 ( .A(n9291), .B(n9460), .S(n8170), .Z(n8148) );
  AOI21_X1 U9695 ( .B1(n8150), .B2(n8211), .A(n8148), .ZN(n8149) );
  OAI21_X1 U9696 ( .B1(n8153), .B2(n8152), .A(n8149), .ZN(n8155) );
  INV_X1 U9697 ( .A(n8150), .ZN(n8151) );
  NAND3_X1 U9698 ( .A1(n8153), .A2(n8152), .A3(n8151), .ZN(n8154) );
  NAND2_X1 U9699 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  MUX2_X1 U9700 ( .A(n9242), .B(n8283), .S(n8158), .Z(n8157) );
  MUX2_X1 U9701 ( .A(n8284), .B(n8286), .S(n8158), .Z(n8159) );
  INV_X1 U9702 ( .A(n8167), .ZN(n8164) );
  NAND2_X1 U9703 ( .A1(n9443), .A2(n9174), .ZN(n8216) );
  NOR2_X1 U9704 ( .A1(n8161), .A2(n6594), .ZN(n8162) );
  AOI21_X1 U9705 ( .B1(n8173), .B2(n8216), .A(n9438), .ZN(n8220) );
  AOI21_X1 U9706 ( .B1(n8164), .B2(n8299), .A(n8220), .ZN(n8172) );
  INV_X1 U9707 ( .A(n9438), .ZN(n8166) );
  INV_X1 U9708 ( .A(n8173), .ZN(n8165) );
  NAND2_X1 U9709 ( .A1(n8166), .A2(n8165), .ZN(n8215) );
  INV_X1 U9710 ( .A(n8287), .ZN(n8168) );
  NOR3_X1 U9711 ( .A1(n8220), .A2(n8168), .A3(n8167), .ZN(n8169) );
  INV_X1 U9712 ( .A(n8176), .ZN(n8175) );
  NAND2_X1 U9713 ( .A1(n5858), .A2(n8304), .ZN(n8174) );
  AOI21_X1 U9714 ( .B1(n8175), .B2(n8174), .A(n8339), .ZN(n8298) );
  OAI21_X1 U9715 ( .B1(n10200), .B2(n8177), .A(n8176), .ZN(n8297) );
  NOR2_X1 U9716 ( .A1(n9443), .A2(n9174), .ZN(n8337) );
  NAND2_X1 U9717 ( .A1(n8274), .A2(n8178), .ZN(n9334) );
  INV_X1 U9718 ( .A(n9373), .ZN(n9379) );
  NAND2_X1 U9719 ( .A1(n8231), .A2(n8181), .ZN(n8311) );
  NOR3_X1 U9720 ( .A1(n8183), .A2(n8182), .A3(n8311), .ZN(n8188) );
  NAND2_X1 U9721 ( .A1(n8315), .A2(n8312), .ZN(n8233) );
  NOR2_X1 U9722 ( .A1(n8233), .A2(n8184), .ZN(n8185) );
  NAND4_X1 U9723 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n8190)
         );
  NOR2_X1 U9724 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  NAND4_X1 U9725 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8195)
         );
  NOR2_X1 U9726 ( .A1(n8196), .A2(n8195), .ZN(n8198) );
  NAND3_X1 U9727 ( .A1(n8199), .A2(n8198), .A3(n8197), .ZN(n8200) );
  NOR2_X1 U9728 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  NAND4_X1 U9729 ( .A1(n9418), .A2(n9983), .A3(n8203), .A4(n8202), .ZN(n8204)
         );
  NOR2_X1 U9730 ( .A1(n9410), .A2(n8204), .ZN(n8205) );
  NAND4_X1 U9731 ( .A1(n9363), .A2(n9394), .A3(n9379), .A4(n8205), .ZN(n8206)
         );
  NOR2_X1 U9732 ( .A1(n9334), .A2(n8206), .ZN(n8207) );
  INV_X1 U9733 ( .A(n9318), .ZN(n9320) );
  NAND3_X1 U9734 ( .A1(n9302), .A2(n8207), .A3(n9320), .ZN(n8208) );
  NOR2_X1 U9735 ( .A1(n9288), .A2(n8208), .ZN(n8212) );
  INV_X1 U9736 ( .A(n8209), .ZN(n8210) );
  NAND4_X1 U9737 ( .A1(n9244), .A2(n9255), .A3(n8212), .A4(n9274), .ZN(n8213)
         );
  NOR4_X1 U9738 ( .A1(n8339), .A2(n8337), .A3(n8214), .A4(n8213), .ZN(n8219)
         );
  INV_X1 U9739 ( .A(n8215), .ZN(n8218) );
  INV_X1 U9740 ( .A(n8216), .ZN(n8217) );
  NOR2_X1 U9741 ( .A1(n8218), .A2(n8217), .ZN(n8338) );
  AOI21_X1 U9742 ( .B1(n8219), .B2(n8338), .A(n8304), .ZN(n8295) );
  INV_X1 U9743 ( .A(n8220), .ZN(n8291) );
  OR2_X1 U9744 ( .A1(n4671), .A2(n8221), .ZN(n8301) );
  NAND2_X1 U9745 ( .A1(n8223), .A2(n8222), .ZN(n8243) );
  OR3_X1 U9746 ( .A1(n8246), .A2(n8224), .A3(n8243), .ZN(n8225) );
  NOR2_X1 U9747 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  AND4_X1 U9748 ( .A1(n8260), .A2(n8227), .A3(n8259), .A4(n8254), .ZN(n8228)
         );
  NAND2_X1 U9749 ( .A1(n8262), .A2(n8228), .ZN(n8325) );
  INV_X1 U9750 ( .A(n8311), .ZN(n8230) );
  NAND3_X1 U9751 ( .A1(n6881), .A2(n8230), .A3(n8229), .ZN(n8239) );
  NAND3_X1 U9752 ( .A1(n8233), .A2(n8232), .A3(n8231), .ZN(n8235) );
  AND3_X1 U9753 ( .A1(n8235), .A2(n8314), .A3(n8234), .ZN(n8238) );
  INV_X1 U9754 ( .A(n8236), .ZN(n8237) );
  AOI21_X1 U9755 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8263) );
  INV_X1 U9756 ( .A(n8240), .ZN(n8249) );
  OAI21_X1 U9757 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8244) );
  INV_X1 U9758 ( .A(n8244), .ZN(n8245) );
  NOR2_X1 U9759 ( .A1(n8246), .A2(n8245), .ZN(n8248) );
  OAI21_X1 U9760 ( .B1(n8249), .B2(n8248), .A(n8247), .ZN(n8251) );
  NAND2_X1 U9761 ( .A1(n8251), .A2(n8250), .ZN(n8253) );
  NAND3_X1 U9762 ( .A1(n8254), .A2(n8253), .A3(n8252), .ZN(n8255) );
  NAND3_X1 U9763 ( .A1(n8257), .A2(n8256), .A3(n8255), .ZN(n8258) );
  AND3_X1 U9764 ( .A1(n8260), .A2(n8259), .A3(n8258), .ZN(n8261) );
  NAND2_X1 U9765 ( .A1(n8262), .A2(n8261), .ZN(n8323) );
  OAI21_X1 U9766 ( .B1(n8325), .B2(n8263), .A(n8323), .ZN(n8264) );
  INV_X1 U9767 ( .A(n8264), .ZN(n8265) );
  NOR2_X1 U9768 ( .A1(n8301), .A2(n8265), .ZN(n8279) );
  INV_X1 U9769 ( .A(n8266), .ZN(n8270) );
  INV_X1 U9770 ( .A(n8267), .ZN(n8269) );
  OAI211_X1 U9771 ( .C1(n8271), .C2(n8270), .A(n8269), .B(n8268), .ZN(n8272)
         );
  NAND2_X1 U9772 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  NAND2_X1 U9773 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  OR2_X1 U9774 ( .A1(n8277), .A2(n8276), .ZN(n8326) );
  INV_X1 U9775 ( .A(n8330), .ZN(n8278) );
  OAI21_X1 U9776 ( .B1(n8279), .B2(n8326), .A(n8278), .ZN(n8280) );
  AND2_X1 U9777 ( .A1(n8329), .A2(n8280), .ZN(n8285) );
  NAND2_X1 U9778 ( .A1(n9242), .A2(n8281), .ZN(n8282) );
  NAND3_X1 U9779 ( .A1(n8284), .A2(n8283), .A3(n8282), .ZN(n8300) );
  AOI21_X1 U9780 ( .B1(n8285), .B2(n9242), .A(n8300), .ZN(n8289) );
  NAND2_X1 U9781 ( .A1(n8287), .A2(n8286), .ZN(n8332) );
  OAI211_X1 U9782 ( .C1(n8289), .C2(n8332), .A(n8288), .B(n8299), .ZN(n8290)
         );
  AOI211_X1 U9783 ( .C1(n8291), .C2(n8290), .A(n5859), .B(n8339), .ZN(n8292)
         );
  AOI211_X1 U9784 ( .C1(n8298), .C2(n8297), .A(n8343), .B(n8296), .ZN(n8356)
         );
  INV_X1 U9785 ( .A(n8299), .ZN(n8336) );
  INV_X1 U9786 ( .A(n8300), .ZN(n8334) );
  INV_X1 U9787 ( .A(n8301), .ZN(n8328) );
  INV_X1 U9788 ( .A(n8302), .ZN(n8303) );
  OAI211_X1 U9789 ( .C1(n6838), .C2(n8305), .A(n8304), .B(n8303), .ZN(n8307)
         );
  NAND2_X1 U9790 ( .A1(n8307), .A2(n8306), .ZN(n8310) );
  OAI22_X1 U9791 ( .A1(n7957), .A2(n8310), .B1(n8309), .B2(n8308), .ZN(n8313)
         );
  AOI21_X1 U9792 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8318) );
  INV_X1 U9793 ( .A(n8315), .ZN(n8316) );
  NOR4_X1 U9794 ( .A1(n8318), .A2(n4844), .A3(n8317), .A4(n8316), .ZN(n8322)
         );
  INV_X1 U9795 ( .A(n8320), .ZN(n8321) );
  NOR3_X1 U9796 ( .A1(n8322), .A2(n4847), .A3(n8321), .ZN(n8324) );
  OAI21_X1 U9797 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8327) );
  AOI21_X1 U9798 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n8331) );
  OAI211_X1 U9799 ( .C1(n8331), .C2(n8330), .A(n9255), .B(n8329), .ZN(n8333)
         );
  AOI21_X1 U9800 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8335) );
  NOR3_X1 U9801 ( .A1(n8337), .A2(n8336), .A3(n8335), .ZN(n8342) );
  INV_X1 U9802 ( .A(n8338), .ZN(n8341) );
  INV_X1 U9803 ( .A(n8339), .ZN(n8340) );
  OAI21_X1 U9804 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8347) );
  NAND3_X1 U9805 ( .A1(n8347), .A2(n9342), .A3(n8343), .ZN(n8345) );
  INV_X1 U9806 ( .A(n8351), .ZN(n8344) );
  OAI211_X1 U9807 ( .C1(n8347), .C2(n8346), .A(n8345), .B(n8344), .ZN(n8355)
         );
  INV_X1 U9808 ( .A(n10234), .ZN(n8348) );
  NOR4_X1 U9809 ( .A1(n8350), .A2(n5886), .A3(n8349), .A4(n8348), .ZN(n8354)
         );
  OAI21_X1 U9810 ( .B1(n8352), .B2(n8351), .A(P1_B_REG_SCAN_IN), .ZN(n8353) );
  OAI22_X1 U9811 ( .A1(n8356), .A2(n8355), .B1(n8354), .B2(n8353), .ZN(
        P1_U3240) );
  XNOR2_X1 U9812 ( .A(n9438), .B(n9439), .ZN(n9436) );
  NAND2_X1 U9813 ( .A1(n9436), .A2(n10212), .ZN(n8359) );
  AOI21_X1 U9814 ( .B1(n10216), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8357), .ZN(
        n8358) );
  OAI211_X1 U9815 ( .C1(n9438), .C2(n9432), .A(n8359), .B(n8358), .ZN(P1_U3261) );
  OAI222_X1 U9816 ( .A1(n9018), .A2(n8361), .B1(n8454), .B2(n8360), .C1(n4919), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U9817 ( .A1(n9890), .A2(n8363), .B1(n4459), .B2(n8362), .C1(
        P1_U3084), .C2(n5858), .ZN(P1_U3331) );
  AOI22_X1 U9818 ( .A1(n8366), .A2(n8365), .B1(n8364), .B2(n8705), .ZN(n8367)
         );
  XOR2_X1 U9819 ( .A(n8369), .B(n8368), .Z(n8374) );
  INV_X1 U9820 ( .A(n6507), .ZN(n8370) );
  NAND2_X1 U9821 ( .A1(n8370), .A2(P2_B_REG_SCAN_IN), .ZN(n8371) );
  NAND2_X1 U9822 ( .A1(n8873), .A2(n8371), .ZN(n8684) );
  OAI22_X1 U9823 ( .A1(n8705), .A2(n8850), .B1(n8372), .B2(n8684), .ZN(n8373)
         );
  NAND2_X1 U9824 ( .A1(n4609), .A2(n8896), .ZN(n8381) );
  AOI21_X1 U9825 ( .B1(n8900), .B2(n8375), .A(n8690), .ZN(n8901) );
  INV_X1 U9826 ( .A(n8900), .ZN(n8378) );
  AOI22_X1 U9827 ( .A1(n8858), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8376), .B2(
        n8856), .ZN(n8377) );
  OAI21_X1 U9828 ( .B1(n8378), .B2(n8861), .A(n8377), .ZN(n8379) );
  AOI21_X1 U9829 ( .B1(n8901), .B2(n8891), .A(n8379), .ZN(n8380) );
  OAI211_X1 U9830 ( .C1(n8903), .C2(n8865), .A(n8381), .B(n8380), .ZN(P2_U3267) );
  OAI222_X1 U9831 ( .A1(n9890), .A2(n8383), .B1(n4459), .B2(n8382), .C1(n5859), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  NAND2_X1 U9832 ( .A1(n8385), .A2(n8384), .ZN(n8495) );
  XNOR2_X1 U9833 ( .A(n8961), .B(n8429), .ZN(n8387) );
  NAND2_X1 U9834 ( .A1(n8874), .A2(n8430), .ZN(n8386) );
  XNOR2_X1 U9835 ( .A(n8387), .B(n8386), .ZN(n8494) );
  XNOR2_X1 U9836 ( .A(n8954), .B(n8436), .ZN(n8390) );
  NAND2_X1 U9837 ( .A1(n8555), .A2(n8430), .ZN(n8388) );
  XNOR2_X1 U9838 ( .A(n8390), .B(n8388), .ZN(n8527) );
  INV_X1 U9839 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U9840 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  XNOR2_X1 U9841 ( .A(n8951), .B(n8429), .ZN(n8392) );
  NAND2_X1 U9842 ( .A1(n8836), .A2(n8430), .ZN(n8393) );
  NAND2_X1 U9843 ( .A1(n8392), .A2(n8393), .ZN(n8397) );
  INV_X1 U9844 ( .A(n8392), .ZN(n8395) );
  INV_X1 U9845 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U9846 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  NAND2_X1 U9847 ( .A1(n8397), .A2(n8396), .ZN(n8468) );
  XNOR2_X1 U9848 ( .A(n8944), .B(n8429), .ZN(n8398) );
  NAND2_X1 U9849 ( .A1(n8794), .A2(n8430), .ZN(n8399) );
  XNOR2_X1 U9850 ( .A(n8398), .B(n8399), .ZN(n8513) );
  INV_X1 U9851 ( .A(n8398), .ZN(n8401) );
  INV_X1 U9852 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U9853 ( .A1(n8401), .A2(n8400), .ZN(n8402) );
  OAI21_X2 U9854 ( .B1(n8512), .B2(n8513), .A(n8402), .ZN(n8475) );
  XNOR2_X1 U9855 ( .A(n8939), .B(n8436), .ZN(n8405) );
  NAND2_X1 U9856 ( .A1(n8779), .A2(n8430), .ZN(n8403) );
  XNOR2_X1 U9857 ( .A(n8405), .B(n8403), .ZN(n8474) );
  NAND2_X1 U9858 ( .A1(n8475), .A2(n8474), .ZN(n8407) );
  INV_X1 U9859 ( .A(n8403), .ZN(n8404) );
  NAND2_X1 U9860 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  XNOR2_X1 U9861 ( .A(n6200), .B(n8429), .ZN(n8409) );
  XNOR2_X1 U9862 ( .A(n8408), .B(n8409), .ZN(n8520) );
  NAND2_X1 U9863 ( .A1(n8795), .A2(n8430), .ZN(n8519) );
  NAND2_X1 U9864 ( .A1(n8520), .A2(n8519), .ZN(n8518) );
  INV_X1 U9865 ( .A(n8408), .ZN(n8410) );
  NAND2_X1 U9866 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  XOR2_X1 U9867 ( .A(n8436), .B(n8924), .Z(n8504) );
  NAND2_X1 U9868 ( .A1(n8504), .A2(n8486), .ZN(n8413) );
  NAND2_X1 U9869 ( .A1(n8780), .A2(n8430), .ZN(n8501) );
  INV_X1 U9870 ( .A(n8501), .ZN(n8412) );
  NAND2_X1 U9871 ( .A1(n8413), .A2(n8412), .ZN(n8421) );
  INV_X1 U9872 ( .A(n8500), .ZN(n8416) );
  NAND2_X1 U9873 ( .A1(n7993), .A2(n8430), .ZN(n8417) );
  NAND2_X1 U9874 ( .A1(n8416), .A2(n8415), .ZN(n8420) );
  INV_X1 U9875 ( .A(n8504), .ZN(n8418) );
  INV_X1 U9876 ( .A(n8417), .ZN(n8503) );
  OAI211_X1 U9877 ( .C1(n8502), .C2(n8421), .A(n8420), .B(n8419), .ZN(n8423)
         );
  XNOR2_X1 U9878 ( .A(n8921), .B(n8436), .ZN(n8484) );
  NOR2_X1 U9879 ( .A1(n8750), .A2(n7025), .ZN(n8483) );
  INV_X1 U9880 ( .A(n8423), .ZN(n8482) );
  INV_X1 U9881 ( .A(n8484), .ZN(n8424) );
  XNOR2_X1 U9882 ( .A(n8916), .B(n8429), .ZN(n8426) );
  NAND2_X1 U9883 ( .A1(n8553), .A2(n8430), .ZN(n8425) );
  NOR2_X1 U9884 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  AOI21_X1 U9885 ( .B1(n8426), .B2(n8425), .A(n8427), .ZN(n8541) );
  INV_X1 U9886 ( .A(n8427), .ZN(n8428) );
  XNOR2_X1 U9887 ( .A(n8909), .B(n8429), .ZN(n8432) );
  NAND2_X1 U9888 ( .A1(n8552), .A2(n8430), .ZN(n8431) );
  NOR2_X1 U9889 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  AOI21_X1 U9890 ( .B1(n8432), .B2(n8431), .A(n8433), .ZN(n8456) );
  NAND2_X1 U9891 ( .A1(n8457), .A2(n8456), .ZN(n8455) );
  INV_X1 U9892 ( .A(n8433), .ZN(n8434) );
  NAND2_X1 U9893 ( .A1(n8455), .A2(n8434), .ZN(n8439) );
  NOR2_X1 U9894 ( .A1(n8705), .A2(n7025), .ZN(n8435) );
  XOR2_X1 U9895 ( .A(n8436), .B(n8435), .Z(n8437) );
  XNOR2_X1 U9896 ( .A(n8904), .B(n8437), .ZN(n8438) );
  XNOR2_X1 U9897 ( .A(n8439), .B(n8438), .ZN(n8448) );
  INV_X1 U9898 ( .A(n8440), .ZN(n8442) );
  OAI22_X1 U9899 ( .A1(n8522), .A2(n8442), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8441), .ZN(n8446) );
  OAI22_X1 U9900 ( .A1(n8444), .A2(n8530), .B1(n8531), .B2(n8443), .ZN(n8445)
         );
  AOI211_X1 U9901 ( .C1(n8904), .C2(n4453), .A(n8446), .B(n8445), .ZN(n8447)
         );
  OAI21_X1 U9902 ( .B1(n8448), .B2(n8537), .A(n8447), .ZN(P2_U3222) );
  INV_X1 U9903 ( .A(n8449), .ZN(n9894) );
  OAI222_X1 U9904 ( .A1(n9018), .A2(n8450), .B1(P2_U3152), .B2(n6509), .C1(
        n8454), .C2(n9894), .ZN(P2_U3330) );
  INV_X1 U9905 ( .A(n8451), .ZN(n8453) );
  OAI222_X1 U9906 ( .A1(n9890), .A2(n8452), .B1(n4459), .B2(n8453), .C1(n4658), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  OAI222_X1 U9907 ( .A1(n9018), .A2(n9639), .B1(n8454), .B2(n8453), .C1(n5927), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  OAI211_X1 U9908 ( .C1(n8457), .C2(n8456), .A(n8455), .B(n8539), .ZN(n8461)
         );
  OAI22_X1 U9909 ( .A1(n8522), .A2(n8698), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9811), .ZN(n8459) );
  OAI22_X1 U9910 ( .A1(n8705), .A2(n8530), .B1(n8531), .B2(n8704), .ZN(n8458)
         );
  AOI211_X1 U9911 ( .C1(n8909), .C2(n4453), .A(n8459), .B(n8458), .ZN(n8460)
         );
  NAND2_X1 U9912 ( .A1(n8461), .A2(n8460), .ZN(P2_U3216) );
  XNOR2_X1 U9913 ( .A(n8502), .B(n8501), .ZN(n8467) );
  INV_X1 U9914 ( .A(n8762), .ZN(n8463) );
  OAI22_X1 U9915 ( .A1(n8522), .A2(n8463), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8462), .ZN(n8465) );
  OAI22_X1 U9916 ( .A1(n8486), .A2(n8530), .B1(n8531), .B2(n8477), .ZN(n8464)
         );
  AOI211_X1 U9917 ( .C1(n8930), .C2(n4453), .A(n8465), .B(n8464), .ZN(n8466)
         );
  OAI21_X1 U9918 ( .B1(n8467), .B2(n8537), .A(n8466), .ZN(P2_U3218) );
  AOI21_X1 U9919 ( .B1(n8469), .B2(n8468), .A(n4531), .ZN(n8473) );
  NAND2_X1 U9920 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8681) );
  OAI21_X1 U9921 ( .B1(n8522), .B2(n8823), .A(n8681), .ZN(n8471) );
  OAI22_X1 U9922 ( .A1(n8851), .A2(n8531), .B1(n8530), .B2(n8821), .ZN(n8470)
         );
  AOI211_X1 U9923 ( .C1(n8951), .C2(n4453), .A(n8471), .B(n8470), .ZN(n8472)
         );
  OAI21_X1 U9924 ( .B1(n8473), .B2(n8537), .A(n8472), .ZN(P2_U3221) );
  XNOR2_X1 U9925 ( .A(n8475), .B(n8474), .ZN(n8481) );
  OAI22_X1 U9926 ( .A1(n8522), .A2(n8788), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8476), .ZN(n8479) );
  OAI22_X1 U9927 ( .A1(n8821), .A2(n8531), .B1(n8530), .B2(n8477), .ZN(n8478)
         );
  AOI211_X1 U9928 ( .C1(n8939), .C2(n4453), .A(n8479), .B(n8478), .ZN(n8480)
         );
  OAI21_X1 U9929 ( .B1(n8481), .B2(n8537), .A(n8480), .ZN(P2_U3225) );
  XNOR2_X1 U9930 ( .A(n8484), .B(n8483), .ZN(n8485) );
  XNOR2_X1 U9931 ( .A(n8482), .B(n8485), .ZN(n8493) );
  NAND2_X1 U9932 ( .A1(n8553), .A2(n8873), .ZN(n8488) );
  OR2_X1 U9933 ( .A1(n8486), .A2(n8850), .ZN(n8487) );
  AND2_X1 U9934 ( .A1(n8488), .A2(n8487), .ZN(n8731) );
  OAI22_X1 U9935 ( .A1(n8731), .A2(n8546), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8489), .ZN(n8490) );
  AOI21_X1 U9936 ( .B1(n8734), .B2(n8548), .A(n8490), .ZN(n8492) );
  NAND2_X1 U9937 ( .A1(n8921), .A2(n4453), .ZN(n8491) );
  OAI211_X1 U9938 ( .C1(n8493), .C2(n8537), .A(n8492), .B(n8491), .ZN(P2_U3227) );
  XNOR2_X1 U9939 ( .A(n8495), .B(n8494), .ZN(n8499) );
  OAI22_X1 U9940 ( .A1(n8522), .A2(n8855), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8629), .ZN(n8497) );
  OAI22_X1 U9941 ( .A1(n8849), .A2(n8531), .B1(n8530), .B2(n8851), .ZN(n8496)
         );
  AOI211_X1 U9942 ( .C1(n8961), .C2(n4453), .A(n8497), .B(n8496), .ZN(n8498)
         );
  OAI21_X1 U9943 ( .B1(n8499), .B2(n8537), .A(n8498), .ZN(P2_U3230) );
  OAI21_X1 U9944 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8506) );
  XNOR2_X1 U9945 ( .A(n8504), .B(n8503), .ZN(n8505) );
  XNOR2_X1 U9946 ( .A(n8506), .B(n8505), .ZN(n8511) );
  OAI22_X1 U9947 ( .A1(n8522), .A2(n8507), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9629), .ZN(n8509) );
  OAI22_X1 U9948 ( .A1(n8749), .A2(n8531), .B1(n8530), .B2(n8750), .ZN(n8508)
         );
  AOI211_X1 U9949 ( .C1(n8924), .C2(n4453), .A(n8509), .B(n8508), .ZN(n8510)
         );
  OAI21_X1 U9950 ( .B1(n8511), .B2(n8537), .A(n8510), .ZN(P2_U3231) );
  XNOR2_X1 U9951 ( .A(n8512), .B(n8513), .ZN(n8517) );
  OAI22_X1 U9952 ( .A1(n8522), .A2(n8804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9626), .ZN(n8515) );
  OAI22_X1 U9953 ( .A1(n8810), .A2(n8531), .B1(n8530), .B2(n8811), .ZN(n8514)
         );
  AOI211_X1 U9954 ( .C1(n8944), .C2(n4453), .A(n8515), .B(n8514), .ZN(n8516)
         );
  OAI21_X1 U9955 ( .B1(n8517), .B2(n8537), .A(n8516), .ZN(P2_U3235) );
  OAI21_X1 U9956 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8521) );
  NAND2_X1 U9957 ( .A1(n8521), .A2(n8539), .ZN(n8526) );
  NOR2_X1 U9958 ( .A1(n8522), .A2(n8772), .ZN(n8524) );
  OAI22_X1 U9959 ( .A1(n8749), .A2(n8530), .B1(n8531), .B2(n8811), .ZN(n8523)
         );
  AOI211_X1 U9960 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8524), 
        .B(n8523), .ZN(n8525) );
  OAI211_X1 U9961 ( .C1(n8775), .C2(n8551), .A(n8526), .B(n8525), .ZN(P2_U3237) );
  XNOR2_X1 U9962 ( .A(n8528), .B(n8527), .ZN(n8538) );
  NOR2_X1 U9963 ( .A1(n8529), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8658) );
  OAI22_X1 U9964 ( .A1(n8532), .A2(n8531), .B1(n8530), .B2(n8810), .ZN(n8533)
         );
  AOI211_X1 U9965 ( .C1(n8548), .C2(n8831), .A(n8658), .B(n8533), .ZN(n8536)
         );
  NAND2_X1 U9966 ( .A1(n8954), .A2(n4453), .ZN(n8535) );
  OAI211_X1 U9967 ( .C1(n8538), .C2(n8537), .A(n8536), .B(n8535), .ZN(P2_U3240) );
  OAI211_X1 U9968 ( .C1(n8542), .C2(n8541), .A(n8540), .B(n8539), .ZN(n8550)
         );
  NAND2_X1 U9969 ( .A1(n8552), .A2(n8873), .ZN(n8544) );
  OR2_X1 U9970 ( .A1(n8750), .A2(n8850), .ZN(n8543) );
  AND2_X1 U9971 ( .A1(n8544), .A2(n8543), .ZN(n8717) );
  OAI22_X1 U9972 ( .A1(n8717), .A2(n8546), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8545), .ZN(n8547) );
  AOI21_X1 U9973 ( .B1(n8722), .B2(n8548), .A(n8547), .ZN(n8549) );
  OAI211_X1 U9974 ( .C1(n8725), .C2(n8551), .A(n8550), .B(n8549), .ZN(P2_U3242) );
  MUX2_X1 U9975 ( .A(n8552), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8568), .Z(
        P2_U3579) );
  MUX2_X1 U9976 ( .A(n8553), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8568), .Z(
        P2_U3578) );
  MUX2_X1 U9977 ( .A(n8554), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8568), .Z(
        P2_U3577) );
  MUX2_X1 U9978 ( .A(n7993), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8568), .Z(
        P2_U3576) );
  MUX2_X1 U9979 ( .A(n8780), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8568), .Z(
        P2_U3575) );
  MUX2_X1 U9980 ( .A(n8795), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8568), .Z(
        P2_U3574) );
  MUX2_X1 U9981 ( .A(n8779), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8568), .Z(
        P2_U3573) );
  MUX2_X1 U9982 ( .A(n8794), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8568), .Z(
        P2_U3572) );
  MUX2_X1 U9983 ( .A(n8836), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8568), .Z(
        P2_U3571) );
  MUX2_X1 U9984 ( .A(n8555), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8568), .Z(
        P2_U3570) );
  MUX2_X1 U9985 ( .A(n8874), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8568), .Z(
        P2_U3569) );
  MUX2_X1 U9986 ( .A(n8556), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8568), .Z(
        P2_U3568) );
  MUX2_X1 U9987 ( .A(n8872), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8568), .Z(
        P2_U3567) );
  MUX2_X1 U9988 ( .A(n8557), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8568), .Z(
        P2_U3566) );
  MUX2_X1 U9989 ( .A(n8558), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8568), .Z(
        P2_U3565) );
  MUX2_X1 U9990 ( .A(n8559), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8568), .Z(
        P2_U3564) );
  MUX2_X1 U9991 ( .A(n8560), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8568), .Z(
        P2_U3563) );
  MUX2_X1 U9992 ( .A(n8561), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8568), .Z(
        P2_U3562) );
  MUX2_X1 U9993 ( .A(n8562), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8568), .Z(
        P2_U3561) );
  MUX2_X1 U9994 ( .A(n8563), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8568), .Z(
        P2_U3560) );
  MUX2_X1 U9995 ( .A(n8564), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8568), .Z(
        P2_U3559) );
  MUX2_X1 U9996 ( .A(n8565), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8568), .Z(
        P2_U3558) );
  MUX2_X1 U9997 ( .A(n8566), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8568), .Z(
        P2_U3557) );
  MUX2_X1 U9998 ( .A(n8567), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8568), .Z(
        P2_U3556) );
  MUX2_X1 U9999 ( .A(n6946), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8568), .Z(
        P2_U3555) );
  MUX2_X1 U10000 ( .A(n6756), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8568), .Z(
        P2_U3554) );
  MUX2_X1 U10001 ( .A(n6786), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8568), .Z(
        P2_U3553) );
  MUX2_X1 U10002 ( .A(n8569), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8568), .Z(
        P2_U3552) );
  NAND2_X1 U10003 ( .A1(n9930), .A2(n8570), .ZN(n8582) );
  OAI211_X1 U10004 ( .C1(n8573), .C2(n8572), .A(n10282), .B(n8571), .ZN(n8581)
         );
  INV_X1 U10005 ( .A(n8574), .ZN(n8575) );
  AOI21_X1 U10006 ( .B1(n10287), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8575), .ZN(
        n8580) );
  OAI211_X1 U10007 ( .C1(n8578), .C2(n8577), .A(n10281), .B(n8576), .ZN(n8579)
         );
  NAND4_X1 U10008 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(
        P2_U3249) );
  AOI211_X1 U10009 ( .C1(n8585), .C2(n8584), .A(n8583), .B(n9924), .ZN(n8586)
         );
  AOI21_X1 U10010 ( .B1(n9930), .B2(n8587), .A(n8586), .ZN(n8595) );
  NOR2_X1 U10011 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8588), .ZN(n8589) );
  AOI21_X1 U10012 ( .B1(n10287), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8589), .ZN(
        n8594) );
  OAI211_X1 U10013 ( .C1(n8592), .C2(n8591), .A(n8590), .B(n10281), .ZN(n8593)
         );
  NAND3_X1 U10014 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(P2_U3253) );
  AOI211_X1 U10015 ( .C1(n8598), .C2(n8597), .A(n8596), .B(n9924), .ZN(n8599)
         );
  INV_X1 U10016 ( .A(n8599), .ZN(n8609) );
  INV_X1 U10017 ( .A(n8600), .ZN(n8601) );
  AOI21_X1 U10018 ( .B1(n10287), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8601), .ZN(
        n8608) );
  NAND2_X1 U10019 ( .A1(n9930), .A2(n8602), .ZN(n8607) );
  OAI211_X1 U10020 ( .C1(n8605), .C2(n8604), .A(n10281), .B(n8603), .ZN(n8606)
         );
  NAND4_X1 U10021 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(
        P2_U3254) );
  NAND2_X1 U10022 ( .A1(n8611), .A2(n8610), .ZN(n8613) );
  NAND2_X1 U10023 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  XNOR2_X1 U10024 ( .A(n8631), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8614) );
  NOR2_X1 U10025 ( .A1(n8614), .A2(n8615), .ZN(n8632) );
  AOI21_X1 U10026 ( .B1(n8615), .B2(n8614), .A(n8632), .ZN(n8628) );
  NAND2_X1 U10027 ( .A1(n8617), .A2(n8616), .ZN(n8619) );
  NAND2_X1 U10028 ( .A1(n8619), .A2(n8618), .ZN(n8621) );
  NAND2_X1 U10029 ( .A1(n8631), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8645) );
  OAI21_X1 U10030 ( .B1(n8631), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8645), .ZN(
        n8620) );
  AOI211_X1 U10031 ( .C1(n8621), .C2(n8620), .A(n8643), .B(n9924), .ZN(n8626)
         );
  AOI21_X1 U10032 ( .B1(n10287), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8622), .ZN(
        n8623) );
  OAI21_X1 U10033 ( .B1(n10283), .B2(n8624), .A(n8623), .ZN(n8625) );
  NOR2_X1 U10034 ( .A1(n8626), .A2(n8625), .ZN(n8627) );
  OAI21_X1 U10035 ( .B1(n8628), .B2(n10285), .A(n8627), .ZN(P2_U3261) );
  INV_X1 U10036 ( .A(n8659), .ZN(n8650) );
  NOR2_X1 U10037 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8629), .ZN(n8641) );
  XNOR2_X1 U10038 ( .A(n8659), .B(n8630), .ZN(n8636) );
  INV_X1 U10039 ( .A(n8636), .ZN(n8639) );
  OR2_X1 U10040 ( .A1(n8631), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8634) );
  INV_X1 U10041 ( .A(n8632), .ZN(n8633) );
  NAND2_X1 U10042 ( .A1(n8634), .A2(n8633), .ZN(n8638) );
  INV_X1 U10043 ( .A(n8638), .ZN(n8635) );
  NAND2_X1 U10044 ( .A1(n8636), .A2(n8635), .ZN(n8654) );
  INV_X1 U10045 ( .A(n8654), .ZN(n8637) );
  AOI211_X1 U10046 ( .C1(n8639), .C2(n8638), .A(n8637), .B(n10285), .ZN(n8640)
         );
  AOI211_X1 U10047 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n10287), .A(n8641), .B(
        n8640), .ZN(n8649) );
  XNOR2_X1 U10048 ( .A(n8659), .B(n8642), .ZN(n8647) );
  INV_X1 U10049 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U10050 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U10051 ( .A1(n8647), .A2(n8646), .ZN(n8661) );
  OAI211_X1 U10052 ( .C1(n8647), .C2(n8646), .A(n10282), .B(n8661), .ZN(n8648)
         );
  OAI211_X1 U10053 ( .C1(n10283), .C2(n8650), .A(n8649), .B(n8648), .ZN(
        P2_U3262) );
  OR2_X1 U10054 ( .A1(n8671), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8668) );
  NAND2_X1 U10055 ( .A1(n8671), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8651) );
  AND2_X1 U10056 ( .A1(n8668), .A2(n8651), .ZN(n8652) );
  NAND2_X1 U10057 ( .A1(n8659), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8653) );
  NAND3_X1 U10058 ( .A1(n8652), .A2(n8654), .A3(n8653), .ZN(n8669) );
  AOI21_X1 U10059 ( .B1(n8654), .B2(n8653), .A(n8652), .ZN(n8655) );
  INV_X1 U10060 ( .A(n8655), .ZN(n8656) );
  AOI21_X1 U10061 ( .B1(n8669), .B2(n8656), .A(n10285), .ZN(n8657) );
  AOI211_X1 U10062 ( .C1(n10287), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8658), .B(
        n8657), .ZN(n8666) );
  NAND2_X1 U10063 ( .A1(n8659), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10064 ( .A1(n8661), .A2(n8660), .ZN(n8672) );
  XNOR2_X1 U10065 ( .A(n8672), .B(n8667), .ZN(n8663) );
  INV_X1 U10066 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U10067 ( .A1(n8663), .A2(n8662), .ZN(n8673) );
  OAI21_X1 U10068 ( .B1(n8663), .B2(n8662), .A(n8673), .ZN(n8664) );
  NAND2_X1 U10069 ( .A1(n10282), .A2(n8664), .ZN(n8665) );
  OAI211_X1 U10070 ( .C1(n10283), .C2(n8667), .A(n8666), .B(n8665), .ZN(
        P2_U3263) );
  INV_X1 U10071 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U10072 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  XNOR2_X1 U10073 ( .A(n8670), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8676) );
  OR2_X1 U10074 ( .A1(n8672), .A2(n8671), .ZN(n8674) );
  NAND2_X1 U10075 ( .A1(n8678), .A2(n10282), .ZN(n8675) );
  OAI211_X1 U10076 ( .C1(n8676), .C2(n10285), .A(n8675), .B(n10283), .ZN(n8680) );
  INV_X1 U10077 ( .A(n8676), .ZN(n8677) );
  OAI22_X1 U10078 ( .A1(n8678), .A2(n9924), .B1(n8677), .B2(n10285), .ZN(n8679) );
  XNOR2_X1 U10079 ( .A(n8689), .B(n8683), .ZN(n8899) );
  NOR2_X1 U10080 ( .A1(n8685), .A2(n8684), .ZN(n9979) );
  INV_X1 U10081 ( .A(n9979), .ZN(n8686) );
  NOR2_X1 U10082 ( .A1(n8858), .A2(n8686), .ZN(n8693) );
  AOI21_X1 U10083 ( .B1(n8858), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8693), .ZN(
        n8688) );
  NAND2_X1 U10084 ( .A1(n8683), .A2(n8886), .ZN(n8687) );
  OAI211_X1 U10085 ( .C1(n8899), .C2(n8695), .A(n8688), .B(n8687), .ZN(
        P2_U3265) );
  OAI21_X1 U10086 ( .B1(n8691), .B2(n8690), .A(n8689), .ZN(n9977) );
  NOR2_X1 U10087 ( .A1(n8691), .A2(n8861), .ZN(n8692) );
  AOI211_X1 U10088 ( .C1(n8858), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8693), .B(
        n8692), .ZN(n8694) );
  OAI21_X1 U10089 ( .B1(n8695), .B2(n9977), .A(n8694), .ZN(P2_U3266) );
  XNOR2_X1 U10090 ( .A(n8696), .B(n8702), .ZN(n8913) );
  AOI21_X1 U10091 ( .B1(n8909), .B2(n8719), .A(n8697), .ZN(n8910) );
  INV_X1 U10092 ( .A(n8698), .ZN(n8699) );
  AOI22_X1 U10093 ( .A1(n8858), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8699), .B2(
        n8856), .ZN(n8700) );
  OAI21_X1 U10094 ( .B1(n4742), .B2(n8861), .A(n8700), .ZN(n8710) );
  NOR2_X1 U10095 ( .A1(n8701), .A2(n8847), .ZN(n8708) );
  OAI21_X1 U10096 ( .B1(n8716), .B2(n8703), .A(n8702), .ZN(n8707) );
  OAI22_X1 U10097 ( .A1(n8705), .A2(n8852), .B1(n8704), .B2(n8850), .ZN(n8706)
         );
  AOI21_X1 U10098 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8912) );
  NOR2_X1 U10099 ( .A1(n8912), .A2(n8858), .ZN(n8709) );
  AOI211_X1 U10100 ( .C1(n8891), .C2(n8910), .A(n8710), .B(n8709), .ZN(n8711)
         );
  OAI21_X1 U10101 ( .B1(n8913), .B2(n8865), .A(n8711), .ZN(P2_U3269) );
  XNOR2_X1 U10102 ( .A(n8712), .B(n4632), .ZN(n8918) );
  INV_X1 U10103 ( .A(n8713), .ZN(n8730) );
  AOI21_X1 U10104 ( .B1(n8730), .B2(n8714), .A(n4632), .ZN(n8715) );
  OAI21_X1 U10105 ( .B1(n8716), .B2(n8715), .A(n8878), .ZN(n8718) );
  NAND2_X1 U10106 ( .A1(n8718), .A2(n8717), .ZN(n8914) );
  INV_X1 U10107 ( .A(n8733), .ZN(n8721) );
  INV_X1 U10108 ( .A(n8719), .ZN(n8720) );
  AOI211_X1 U10109 ( .C1(n8916), .C2(n8721), .A(n10350), .B(n8720), .ZN(n8915)
         );
  NAND2_X1 U10110 ( .A1(n8915), .A2(n8854), .ZN(n8724) );
  AOI22_X1 U10111 ( .A1(n8858), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8722), .B2(
        n8856), .ZN(n8723) );
  OAI211_X1 U10112 ( .C1(n8725), .C2(n8861), .A(n8724), .B(n8723), .ZN(n8726)
         );
  AOI21_X1 U10113 ( .B1(n8914), .B2(n8896), .A(n8726), .ZN(n8727) );
  OAI21_X1 U10114 ( .B1(n8918), .B2(n8865), .A(n8727), .ZN(P2_U3270) );
  XNOR2_X1 U10115 ( .A(n8729), .B(n8728), .ZN(n8923) );
  OAI211_X1 U10116 ( .C1(n4899), .C2(n4514), .A(n8730), .B(n8878), .ZN(n8732)
         );
  NAND2_X1 U10117 ( .A1(n8732), .A2(n8731), .ZN(n8919) );
  AOI211_X1 U10118 ( .C1(n8921), .C2(n8742), .A(n10350), .B(n8733), .ZN(n8920)
         );
  NAND2_X1 U10119 ( .A1(n8920), .A2(n8854), .ZN(n8736) );
  AOI22_X1 U10120 ( .A1(n8858), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8734), .B2(
        n8856), .ZN(n8735) );
  OAI211_X1 U10121 ( .C1(n4748), .C2(n8861), .A(n8736), .B(n8735), .ZN(n8737)
         );
  AOI21_X1 U10122 ( .B1(n8919), .B2(n8896), .A(n8737), .ZN(n8738) );
  OAI21_X1 U10123 ( .B1(n8923), .B2(n8865), .A(n8738), .ZN(P2_U3271) );
  AOI21_X1 U10124 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8928) );
  INV_X1 U10125 ( .A(n8742), .ZN(n8743) );
  AOI21_X1 U10126 ( .B1(n8924), .B2(n4752), .A(n8743), .ZN(n8925) );
  AOI22_X1 U10127 ( .A1(n8858), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8744), .B2(
        n8856), .ZN(n8745) );
  OAI21_X1 U10128 ( .B1(n8746), .B2(n8861), .A(n8745), .ZN(n8754) );
  AOI211_X1 U10129 ( .C1(n8748), .C2(n8747), .A(n8847), .B(n4517), .ZN(n8752)
         );
  OAI22_X1 U10130 ( .A1(n8750), .A2(n8852), .B1(n8749), .B2(n8850), .ZN(n8751)
         );
  NOR2_X1 U10131 ( .A1(n8752), .A2(n8751), .ZN(n8927) );
  NOR2_X1 U10132 ( .A1(n8927), .A2(n8858), .ZN(n8753) );
  AOI211_X1 U10133 ( .C1(n8925), .C2(n8891), .A(n8754), .B(n8753), .ZN(n8755)
         );
  OAI21_X1 U10134 ( .B1(n8865), .B2(n8928), .A(n8755), .ZN(P2_U3272) );
  XNOR2_X1 U10135 ( .A(n8756), .B(n8758), .ZN(n8757) );
  AOI222_X1 U10136 ( .A1(n8878), .A2(n8757), .B1(n8795), .B2(n8871), .C1(n7993), .C2(n8873), .ZN(n8933) );
  OR2_X1 U10137 ( .A1(n4600), .A2(n8758), .ZN(n8929) );
  NAND3_X1 U10138 ( .A1(n8929), .A2(n8759), .A3(n8760), .ZN(n8767) );
  AOI21_X1 U10139 ( .B1(n8930), .B2(n8769), .A(n8761), .ZN(n8931) );
  AOI22_X1 U10140 ( .A1(n8858), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8762), .B2(
        n8856), .ZN(n8763) );
  OAI21_X1 U10141 ( .B1(n8764), .B2(n8861), .A(n8763), .ZN(n8765) );
  AOI21_X1 U10142 ( .B1(n8931), .B2(n8891), .A(n8765), .ZN(n8766) );
  OAI211_X1 U10143 ( .C1(n8858), .C2(n8933), .A(n8767), .B(n8766), .ZN(
        P2_U3273) );
  XNOR2_X1 U10144 ( .A(n8768), .B(n8777), .ZN(n8938) );
  INV_X1 U10145 ( .A(n8787), .ZN(n8771) );
  INV_X1 U10146 ( .A(n8769), .ZN(n8770) );
  AOI21_X1 U10147 ( .B1(n6200), .B2(n8771), .A(n8770), .ZN(n8935) );
  INV_X1 U10148 ( .A(n8772), .ZN(n8773) );
  AOI22_X1 U10149 ( .A1(n8858), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8773), .B2(
        n8856), .ZN(n8774) );
  OAI21_X1 U10150 ( .B1(n8775), .B2(n8861), .A(n8774), .ZN(n8784) );
  OAI211_X1 U10151 ( .C1(n8778), .C2(n8777), .A(n8776), .B(n8878), .ZN(n8782)
         );
  AOI22_X1 U10152 ( .A1(n8780), .A2(n8873), .B1(n8871), .B2(n8779), .ZN(n8781)
         );
  AND2_X1 U10153 ( .A1(n8782), .A2(n8781), .ZN(n8937) );
  NOR2_X1 U10154 ( .A1(n8937), .A2(n8858), .ZN(n8783) );
  AOI211_X1 U10155 ( .C1(n8935), .C2(n8891), .A(n8784), .B(n8783), .ZN(n8785)
         );
  OAI21_X1 U10156 ( .B1(n8865), .B2(n8938), .A(n8785), .ZN(P2_U3274) );
  XNOR2_X1 U10157 ( .A(n8786), .B(n8792), .ZN(n8943) );
  AOI21_X1 U10158 ( .B1(n8939), .B2(n8801), .A(n8787), .ZN(n8940) );
  INV_X1 U10159 ( .A(n8788), .ZN(n8789) );
  AOI22_X1 U10160 ( .A1(n8858), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8789), .B2(
        n8856), .ZN(n8790) );
  OAI21_X1 U10161 ( .B1(n8791), .B2(n8861), .A(n8790), .ZN(n8798) );
  XNOR2_X1 U10162 ( .A(n8793), .B(n8792), .ZN(n8796) );
  AOI222_X1 U10163 ( .A1(n8878), .A2(n8796), .B1(n8795), .B2(n8873), .C1(n8794), .C2(n8871), .ZN(n8942) );
  NOR2_X1 U10164 ( .A1(n8942), .A2(n8858), .ZN(n8797) );
  AOI211_X1 U10165 ( .C1(n8940), .C2(n8891), .A(n8798), .B(n8797), .ZN(n8799)
         );
  OAI21_X1 U10166 ( .B1(n8865), .B2(n8943), .A(n8799), .ZN(P2_U3275) );
  XNOR2_X1 U10167 ( .A(n8800), .B(n8808), .ZN(n8948) );
  INV_X1 U10168 ( .A(n8822), .ZN(n8803) );
  INV_X1 U10169 ( .A(n8801), .ZN(n8802) );
  AOI21_X1 U10170 ( .B1(n8944), .B2(n8803), .A(n8802), .ZN(n8945) );
  INV_X1 U10171 ( .A(n8804), .ZN(n8805) );
  AOI22_X1 U10172 ( .A1(n8858), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8805), .B2(
        n8856), .ZN(n8806) );
  OAI21_X1 U10173 ( .B1(n8807), .B2(n8861), .A(n8806), .ZN(n8815) );
  AOI211_X1 U10174 ( .C1(n8809), .C2(n8808), .A(n8847), .B(n4539), .ZN(n8813)
         );
  OAI22_X1 U10175 ( .A1(n8811), .A2(n8852), .B1(n8810), .B2(n8850), .ZN(n8812)
         );
  NOR2_X1 U10176 ( .A1(n8813), .A2(n8812), .ZN(n8947) );
  NOR2_X1 U10177 ( .A1(n8947), .A2(n8858), .ZN(n8814) );
  AOI211_X1 U10178 ( .C1(n8945), .C2(n8891), .A(n8815), .B(n8814), .ZN(n8816)
         );
  OAI21_X1 U10179 ( .B1(n8865), .B2(n8948), .A(n8816), .ZN(P2_U3276) );
  XNOR2_X1 U10180 ( .A(n8817), .B(n8818), .ZN(n8953) );
  AOI22_X1 U10181 ( .A1(n8951), .A2(n8886), .B1(n8858), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8827) );
  XOR2_X1 U10182 ( .A(n8819), .B(n8818), .Z(n8820) );
  OAI222_X1 U10183 ( .A1(n8852), .A2(n8821), .B1(n8850), .B2(n8851), .C1(n8847), .C2(n8820), .ZN(n8949) );
  AOI211_X1 U10184 ( .C1(n8951), .C2(n8829), .A(n10350), .B(n8822), .ZN(n8950)
         );
  INV_X1 U10185 ( .A(n8950), .ZN(n8824) );
  OAI22_X1 U10186 ( .A1(n8824), .A2(n4460), .B1(n8882), .B2(n8823), .ZN(n8825)
         );
  OAI21_X1 U10187 ( .B1(n8949), .B2(n8825), .A(n8896), .ZN(n8826) );
  OAI211_X1 U10188 ( .C1(n8953), .C2(n8865), .A(n8827), .B(n8826), .ZN(
        P2_U3277) );
  XOR2_X1 U10189 ( .A(n8834), .B(n8828), .Z(n8958) );
  INV_X1 U10190 ( .A(n8829), .ZN(n8830) );
  AOI21_X1 U10191 ( .B1(n8954), .B2(n4747), .A(n8830), .ZN(n8955) );
  AOI22_X1 U10192 ( .A1(n8858), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8831), .B2(
        n8856), .ZN(n8832) );
  OAI21_X1 U10193 ( .B1(n8833), .B2(n8861), .A(n8832), .ZN(n8839) );
  XOR2_X1 U10194 ( .A(n8835), .B(n8834), .Z(n8837) );
  AOI222_X1 U10195 ( .A1(n8878), .A2(n8837), .B1(n8836), .B2(n8873), .C1(n8874), .C2(n8871), .ZN(n8957) );
  NOR2_X1 U10196 ( .A1(n8957), .A2(n8858), .ZN(n8838) );
  AOI211_X1 U10197 ( .C1(n8955), .C2(n8891), .A(n8839), .B(n8838), .ZN(n8840)
         );
  OAI21_X1 U10198 ( .B1(n8865), .B2(n8958), .A(n8840), .ZN(P2_U3278) );
  OAI21_X1 U10199 ( .B1(n4538), .B2(n8845), .A(n8841), .ZN(n8842) );
  INV_X1 U10200 ( .A(n8842), .ZN(n8963) );
  NAND2_X1 U10201 ( .A1(n8843), .A2(n8844), .ZN(n8846) );
  XNOR2_X1 U10202 ( .A(n8846), .B(n8845), .ZN(n8848) );
  OAI222_X1 U10203 ( .A1(n8852), .A2(n8851), .B1(n8850), .B2(n8849), .C1(n8848), .C2(n8847), .ZN(n8959) );
  INV_X1 U10204 ( .A(n8961), .ZN(n8862) );
  AOI211_X1 U10205 ( .C1(n8961), .C2(n8890), .A(n10350), .B(n8853), .ZN(n8960)
         );
  NAND2_X1 U10206 ( .A1(n8960), .A2(n8854), .ZN(n8860) );
  INV_X1 U10207 ( .A(n8855), .ZN(n8857) );
  AOI22_X1 U10208 ( .A1(n8858), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8857), .B2(
        n8856), .ZN(n8859) );
  OAI211_X1 U10209 ( .C1(n8862), .C2(n8861), .A(n8860), .B(n8859), .ZN(n8863)
         );
  AOI21_X1 U10210 ( .B1(n8959), .B2(n8896), .A(n8863), .ZN(n8864) );
  OAI21_X1 U10211 ( .B1(n8963), .B2(n8865), .A(n8864), .ZN(P2_U3279) );
  AND2_X1 U10212 ( .A1(n8866), .A2(n8870), .ZN(n8868) );
  OR2_X1 U10213 ( .A1(n8868), .A2(n8867), .ZN(n8967) );
  OAI21_X1 U10214 ( .B1(n8870), .B2(n8869), .A(n8843), .ZN(n8879) );
  NAND2_X1 U10215 ( .A1(n8872), .A2(n8871), .ZN(n8876) );
  NAND2_X1 U10216 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  NAND2_X1 U10217 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  AOI21_X1 U10218 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8880) );
  OAI21_X1 U10219 ( .B1(n8967), .B2(n8881), .A(n8880), .ZN(n8969) );
  OAI22_X1 U10220 ( .A1(n8896), .A2(n8884), .B1(n8883), .B2(n8882), .ZN(n8885)
         );
  AOI21_X1 U10221 ( .B1(n8964), .B2(n8886), .A(n8885), .ZN(n8893) );
  OR2_X1 U10222 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  AND2_X1 U10223 ( .A1(n8890), .A2(n8889), .ZN(n8965) );
  NAND2_X1 U10224 ( .A1(n8965), .A2(n8891), .ZN(n8892) );
  OAI211_X1 U10225 ( .C1(n8967), .C2(n8894), .A(n8893), .B(n8892), .ZN(n8895)
         );
  AOI21_X1 U10226 ( .B1(n8969), .B2(n8896), .A(n8895), .ZN(n8897) );
  INV_X1 U10227 ( .A(n8897), .ZN(P2_U3280) );
  AOI21_X1 U10228 ( .B1(n8683), .B2(n9980), .A(n9979), .ZN(n8898) );
  OAI21_X1 U10229 ( .B1(n8899), .B2(n10350), .A(n8898), .ZN(n8990) );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8990), .S(n10370), .Z(
        P2_U3551) );
  AOI22_X1 U10231 ( .A1(n8905), .A2(n8985), .B1(n9980), .B2(n8904), .ZN(n8906)
         );
  OAI211_X1 U10232 ( .C1(n8981), .C2(n8908), .A(n8907), .B(n8906), .ZN(n8992)
         );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8992), .S(n10370), .Z(
        P2_U3548) );
  AOI22_X1 U10234 ( .A1(n8910), .A2(n8985), .B1(n9980), .B2(n8909), .ZN(n8911)
         );
  OAI211_X1 U10235 ( .C1(n8913), .C2(n8981), .A(n8912), .B(n8911), .ZN(n8993)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8993), .S(n10370), .Z(
        P2_U3547) );
  AOI211_X1 U10237 ( .C1(n9980), .C2(n8916), .A(n8915), .B(n8914), .ZN(n8917)
         );
  OAI21_X1 U10238 ( .B1(n8918), .B2(n8981), .A(n8917), .ZN(n8994) );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8994), .S(n10370), .Z(
        P2_U3546) );
  AOI211_X1 U10240 ( .C1(n9980), .C2(n8921), .A(n8920), .B(n8919), .ZN(n8922)
         );
  OAI21_X1 U10241 ( .B1(n8923), .B2(n8981), .A(n8922), .ZN(n8995) );
  MUX2_X1 U10242 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8995), .S(n10370), .Z(
        P2_U3545) );
  AOI22_X1 U10243 ( .A1(n8925), .A2(n8985), .B1(n9980), .B2(n8924), .ZN(n8926)
         );
  OAI211_X1 U10244 ( .C1(n8928), .C2(n8981), .A(n8927), .B(n8926), .ZN(n8996)
         );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8996), .S(n10370), .Z(
        P2_U3544) );
  NAND3_X1 U10246 ( .A1(n8929), .A2(n8759), .A3(n10354), .ZN(n8934) );
  AOI22_X1 U10247 ( .A1(n8931), .A2(n8985), .B1(n9980), .B2(n8930), .ZN(n8932)
         );
  NAND3_X1 U10248 ( .A1(n8934), .A2(n8933), .A3(n8932), .ZN(n8997) );
  MUX2_X1 U10249 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8997), .S(n10370), .Z(
        P2_U3543) );
  AOI22_X1 U10250 ( .A1(n8935), .A2(n8985), .B1(n9980), .B2(n6200), .ZN(n8936)
         );
  OAI211_X1 U10251 ( .C1(n8938), .C2(n8981), .A(n8937), .B(n8936), .ZN(n8998)
         );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8998), .S(n10370), .Z(
        P2_U3542) );
  AOI22_X1 U10253 ( .A1(n8940), .A2(n8985), .B1(n9980), .B2(n8939), .ZN(n8941)
         );
  OAI211_X1 U10254 ( .C1(n8943), .C2(n8981), .A(n8942), .B(n8941), .ZN(n8999)
         );
  MUX2_X1 U10255 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8999), .S(n10370), .Z(
        P2_U3541) );
  AOI22_X1 U10256 ( .A1(n8945), .A2(n8985), .B1(n9980), .B2(n8944), .ZN(n8946)
         );
  OAI211_X1 U10257 ( .C1(n8948), .C2(n8981), .A(n8947), .B(n8946), .ZN(n9000)
         );
  MUX2_X1 U10258 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9000), .S(n10370), .Z(
        P2_U3540) );
  AOI211_X1 U10259 ( .C1(n9980), .C2(n8951), .A(n8950), .B(n8949), .ZN(n8952)
         );
  OAI21_X1 U10260 ( .B1(n8981), .B2(n8953), .A(n8952), .ZN(n9001) );
  MUX2_X1 U10261 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9001), .S(n10370), .Z(
        P2_U3539) );
  AOI22_X1 U10262 ( .A1(n8955), .A2(n8985), .B1(n9980), .B2(n8954), .ZN(n8956)
         );
  OAI211_X1 U10263 ( .C1(n8958), .C2(n8981), .A(n8957), .B(n8956), .ZN(n9002)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9002), .S(n10370), .Z(
        P2_U3538) );
  AOI211_X1 U10265 ( .C1(n9980), .C2(n8961), .A(n8960), .B(n8959), .ZN(n8962)
         );
  OAI21_X1 U10266 ( .B1(n8963), .B2(n8981), .A(n8962), .ZN(n9003) );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9003), .S(n10370), .Z(
        P2_U3537) );
  AOI22_X1 U10268 ( .A1(n8965), .A2(n8985), .B1(n9980), .B2(n8964), .ZN(n8966)
         );
  OAI21_X1 U10269 ( .B1(n8967), .B2(n10335), .A(n8966), .ZN(n8968) );
  NOR2_X1 U10270 ( .A1(n8969), .A2(n8968), .ZN(n9004) );
  MUX2_X1 U10271 ( .A(n9810), .B(n9004), .S(n10370), .Z(n8970) );
  INV_X1 U10272 ( .A(n8970), .ZN(P2_U3536) );
  INV_X1 U10273 ( .A(n8971), .ZN(n8976) );
  AOI22_X1 U10274 ( .A1(n8973), .A2(n8985), .B1(n9980), .B2(n8972), .ZN(n8974)
         );
  OAI211_X1 U10275 ( .C1(n8976), .C2(n8981), .A(n8975), .B(n8974), .ZN(n9007)
         );
  MUX2_X1 U10276 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9007), .S(n10370), .Z(
        P2_U3535) );
  AOI22_X1 U10277 ( .A1(n8978), .A2(n8985), .B1(n9980), .B2(n8977), .ZN(n8979)
         );
  OAI211_X1 U10278 ( .C1(n8982), .C2(n8981), .A(n8980), .B(n8979), .ZN(n9008)
         );
  MUX2_X1 U10279 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9008), .S(n10370), .Z(
        P2_U3534) );
  INV_X1 U10280 ( .A(n8983), .ZN(n8989) );
  AOI22_X1 U10281 ( .A1(n8986), .A2(n8985), .B1(n9980), .B2(n8984), .ZN(n8987)
         );
  OAI211_X1 U10282 ( .C1(n10335), .C2(n8989), .A(n8988), .B(n8987), .ZN(n9009)
         );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9009), .S(n10370), .Z(
        P2_U3533) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8990), .S(n10358), .Z(
        P2_U3519) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8991), .S(n10358), .Z(
        P2_U3517) );
  MUX2_X1 U10286 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8992), .S(n10358), .Z(
        P2_U3516) );
  MUX2_X1 U10287 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8993), .S(n10358), .Z(
        P2_U3515) );
  MUX2_X1 U10288 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8994), .S(n10358), .Z(
        P2_U3514) );
  MUX2_X1 U10289 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8995), .S(n10358), .Z(
        P2_U3513) );
  MUX2_X1 U10290 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8996), .S(n10358), .Z(
        P2_U3512) );
  MUX2_X1 U10291 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8997), .S(n10358), .Z(
        P2_U3511) );
  MUX2_X1 U10292 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8998), .S(n10358), .Z(
        P2_U3510) );
  MUX2_X1 U10293 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8999), .S(n10358), .Z(
        P2_U3509) );
  MUX2_X1 U10294 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9000), .S(n10358), .Z(
        P2_U3508) );
  MUX2_X1 U10295 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9001), .S(n10358), .Z(
        P2_U3507) );
  MUX2_X1 U10296 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9002), .S(n10358), .Z(
        P2_U3505) );
  MUX2_X1 U10297 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9003), .S(n10358), .Z(
        P2_U3502) );
  INV_X1 U10298 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9005) );
  MUX2_X1 U10299 ( .A(n9005), .B(n9004), .S(n10358), .Z(n9006) );
  INV_X1 U10300 ( .A(n9006), .ZN(P2_U3499) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9007), .S(n10358), .Z(
        P2_U3496) );
  MUX2_X1 U10302 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9008), .S(n10358), .Z(
        P2_U3493) );
  MUX2_X1 U10303 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9009), .S(n10358), .Z(
        P2_U3490) );
  INV_X1 U10304 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9010) );
  MUX2_X1 U10305 ( .A(P2_REG0_REG_3__SCAN_IN), .B(n9011), .S(n10358), .Z(
        P2_U3460) );
  INV_X1 U10306 ( .A(n8160), .ZN(n9885) );
  NAND3_X1 U10307 ( .A1(n9012), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9014) );
  OAI22_X1 U10308 ( .A1(n4562), .A2(n9014), .B1(n9013), .B2(n9018), .ZN(n9015)
         );
  INV_X1 U10309 ( .A(n9015), .ZN(n9016) );
  OAI21_X1 U10310 ( .B1(n9885), .B2(n8454), .A(n9016), .ZN(P2_U3327) );
  INV_X1 U10311 ( .A(n9017), .ZN(n9886) );
  OAI222_X1 U10312 ( .A1(n8454), .A2(n9886), .B1(P2_U3152), .B2(n9020), .C1(
        n9019), .C2(n9018), .ZN(P2_U3329) );
  INV_X1 U10313 ( .A(n9021), .ZN(n9022) );
  MUX2_X1 U10314 ( .A(n9022), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10315 ( .A(n9023), .ZN(n9025) );
  NAND2_X1 U10316 ( .A1(n9025), .A2(n9024), .ZN(n9027) );
  XNOR2_X1 U10317 ( .A(n9027), .B(n9026), .ZN(n9033) );
  OAI22_X1 U10318 ( .A1(n9141), .A2(n9324), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9028), .ZN(n9029) );
  AOI21_X1 U10319 ( .B1(n9138), .B2(n9290), .A(n9029), .ZN(n9030) );
  OAI21_X1 U10320 ( .B1(n9153), .B2(n9326), .A(n9030), .ZN(n9031) );
  AOI21_X1 U10321 ( .B1(n9480), .B2(n9168), .A(n9031), .ZN(n9032) );
  OAI21_X1 U10322 ( .B1(n9033), .B2(n9172), .A(n9032), .ZN(P1_U3214) );
  NAND2_X1 U10323 ( .A1(n9034), .A2(n9135), .ZN(n9035) );
  INV_X1 U10324 ( .A(n9108), .ZN(n9038) );
  OAI21_X1 U10325 ( .B1(n9036), .B2(n9038), .A(n9035), .ZN(n9037) );
  OAI21_X1 U10326 ( .B1(n9109), .B2(n9038), .A(n9037), .ZN(n9039) );
  NAND2_X1 U10327 ( .A1(n9039), .A2(n9115), .ZN(n9044) );
  NAND2_X1 U10328 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U10329 ( .A1(n9162), .A2(n9395), .ZN(n9040) );
  OAI211_X1 U10330 ( .C1(n9164), .C2(n9041), .A(n9229), .B(n9040), .ZN(n9042)
         );
  AOI21_X1 U10331 ( .B1(n9391), .B2(n9166), .A(n9042), .ZN(n9043) );
  OAI211_X1 U10332 ( .C1(n4815), .C2(n9123), .A(n9044), .B(n9043), .ZN(
        P1_U3217) );
  INV_X1 U10333 ( .A(n9060), .ZN(n9053) );
  NAND2_X1 U10334 ( .A1(n9451), .A2(n5814), .ZN(n9047) );
  NAND2_X1 U10335 ( .A1(n9257), .A2(n9045), .ZN(n9046) );
  NAND2_X1 U10336 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  XNOR2_X1 U10337 ( .A(n9048), .B(n5374), .ZN(n9051) );
  AOI22_X1 U10338 ( .A1(n9451), .A2(n9045), .B1(n9049), .B2(n9257), .ZN(n9050)
         );
  XNOR2_X1 U10339 ( .A(n9051), .B(n9050), .ZN(n9062) );
  AND2_X1 U10340 ( .A1(n9062), .A2(n9115), .ZN(n9052) );
  NAND2_X1 U10341 ( .A1(n9053), .A2(n9052), .ZN(n9066) );
  AOI22_X1 U10342 ( .A1(n9246), .A2(n9138), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9055) );
  NAND2_X1 U10343 ( .A1(n9239), .A2(n9166), .ZN(n9054) );
  OAI211_X1 U10344 ( .C1(n9151), .C2(n9141), .A(n9055), .B(n9054), .ZN(n9056)
         );
  AOI21_X1 U10345 ( .B1(n9451), .B2(n9168), .A(n9056), .ZN(n9065) );
  INV_X1 U10346 ( .A(n9062), .ZN(n9059) );
  INV_X1 U10347 ( .A(n9061), .ZN(n9057) );
  AND2_X1 U10348 ( .A1(n9057), .A2(n9115), .ZN(n9058) );
  NAND2_X1 U10349 ( .A1(n9060), .A2(n5073), .ZN(n9064) );
  NAND3_X1 U10350 ( .A1(n9062), .A2(n9061), .A3(n9115), .ZN(n9063) );
  NAND4_X1 U10351 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(
        P1_U3218) );
  XOR2_X1 U10352 ( .A(n9067), .B(n9068), .Z(n9074) );
  OAI22_X1 U10353 ( .A1(n9164), .A2(n9324), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9069), .ZN(n9070) );
  AOI21_X1 U10354 ( .B1(n9162), .B2(n9396), .A(n9070), .ZN(n9071) );
  OAI21_X1 U10355 ( .B1(n9153), .B2(n9356), .A(n9071), .ZN(n9072) );
  AOI21_X1 U10356 ( .B1(n9489), .B2(n9168), .A(n9072), .ZN(n9073) );
  OAI21_X1 U10357 ( .B1(n9074), .B2(n9172), .A(n9073), .ZN(P1_U3221) );
  XOR2_X1 U10358 ( .A(n9076), .B(n9075), .Z(n9081) );
  NAND2_X1 U10359 ( .A1(n9291), .A2(n9138), .ZN(n9078) );
  AOI22_X1 U10360 ( .A1(n9290), .A2(n9162), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9077) );
  OAI211_X1 U10361 ( .C1(n9153), .C2(n9284), .A(n9078), .B(n9077), .ZN(n9079)
         );
  AOI21_X1 U10362 ( .B1(n9465), .B2(n9168), .A(n9079), .ZN(n9080) );
  OAI21_X1 U10363 ( .B1(n9081), .B2(n9172), .A(n9080), .ZN(P1_U3223) );
  INV_X1 U10364 ( .A(n9083), .ZN(n9084) );
  AOI21_X1 U10365 ( .B1(n9082), .B2(n9085), .A(n9084), .ZN(n9091) );
  NAND2_X1 U10366 ( .A1(n9166), .A2(n9994), .ZN(n9088) );
  NOR2_X1 U10367 ( .A1(n9086), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10156) );
  AOI21_X1 U10368 ( .B1(n9162), .B2(n9987), .A(n10156), .ZN(n9087) );
  OAI211_X1 U10369 ( .C1(n9142), .C2(n9164), .A(n9088), .B(n9087), .ZN(n9089)
         );
  AOI21_X1 U10370 ( .B1(n10009), .B2(n9168), .A(n9089), .ZN(n9090) );
  OAI21_X1 U10371 ( .B1(n9091), .B2(n9172), .A(n9090), .ZN(P1_U3224) );
  OAI21_X1 U10372 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9095) );
  NAND2_X1 U10373 ( .A1(n9095), .A2(n9115), .ZN(n9099) );
  NAND2_X1 U10374 ( .A1(n9162), .A2(n9175), .ZN(n9096) );
  NAND2_X1 U10375 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10164)
         );
  OAI211_X1 U10376 ( .C1(n9164), .C2(n9424), .A(n9096), .B(n10164), .ZN(n9097)
         );
  AOI21_X1 U10377 ( .B1(n9429), .B2(n9166), .A(n9097), .ZN(n9098) );
  OAI211_X1 U10378 ( .C1(n9433), .C2(n9123), .A(n9099), .B(n9098), .ZN(
        P1_U3226) );
  XOR2_X1 U10379 ( .A(n9101), .B(n9100), .Z(n9107) );
  AOI22_X1 U10380 ( .A1(n9305), .A2(n9162), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9103) );
  NAND2_X1 U10381 ( .A1(n9166), .A2(n9311), .ZN(n9102) );
  OAI211_X1 U10382 ( .C1(n9104), .C2(n9164), .A(n9103), .B(n9102), .ZN(n9105)
         );
  AOI21_X1 U10383 ( .B1(n9471), .B2(n9168), .A(n9105), .ZN(n9106) );
  OAI21_X1 U10384 ( .B1(n9107), .B2(n9172), .A(n9106), .ZN(P1_U3227) );
  INV_X1 U10385 ( .A(n9493), .ZN(n9378) );
  NAND2_X1 U10386 ( .A1(n9109), .A2(n9108), .ZN(n9113) );
  AND2_X1 U10387 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  OAI21_X1 U10388 ( .B1(n9114), .B2(n9113), .A(n9112), .ZN(n9116) );
  NAND2_X1 U10389 ( .A1(n9116), .A2(n9115), .ZN(n9122) );
  INV_X1 U10390 ( .A(n9117), .ZN(n9376) );
  AOI22_X1 U10391 ( .A1(n9138), .A2(n9381), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9118) );
  OAI21_X1 U10392 ( .B1(n9119), .B2(n9141), .A(n9118), .ZN(n9120) );
  AOI21_X1 U10393 ( .B1(n9376), .B2(n9166), .A(n9120), .ZN(n9121) );
  OAI211_X1 U10394 ( .C1(n9378), .C2(n9123), .A(n9122), .B(n9121), .ZN(
        P1_U3231) );
  INV_X1 U10395 ( .A(n9124), .ZN(n9128) );
  NAND2_X1 U10396 ( .A1(n4478), .A2(n4523), .ZN(n9126) );
  AOI22_X1 U10397 ( .A1(n9128), .A2(n9127), .B1(n9126), .B2(n9125), .ZN(n9133)
         );
  AOI22_X1 U10398 ( .A1(n9162), .A2(n9381), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9130) );
  NAND2_X1 U10399 ( .A1(n9305), .A2(n9138), .ZN(n9129) );
  OAI211_X1 U10400 ( .C1(n9153), .C2(n9341), .A(n9130), .B(n9129), .ZN(n9131)
         );
  AOI21_X1 U10401 ( .B1(n9485), .B2(n9168), .A(n9131), .ZN(n9132) );
  OAI21_X1 U10402 ( .B1(n9133), .B2(n9172), .A(n9132), .ZN(P1_U3233) );
  NAND2_X1 U10403 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  XOR2_X1 U10404 ( .A(n9137), .B(n9136), .Z(n9145) );
  NAND2_X1 U10405 ( .A1(n9166), .A2(n9405), .ZN(n9140) );
  NOR2_X1 U10406 ( .A1(n9824), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10183) );
  AOI21_X1 U10407 ( .B1(n9138), .B2(n9412), .A(n10183), .ZN(n9139) );
  OAI211_X1 U10408 ( .C1(n9142), .C2(n9141), .A(n9140), .B(n9139), .ZN(n9143)
         );
  AOI21_X1 U10409 ( .B1(n9503), .B2(n9168), .A(n9143), .ZN(n9144) );
  OAI21_X1 U10410 ( .B1(n9145), .B2(n9172), .A(n9144), .ZN(P1_U3236) );
  INV_X1 U10411 ( .A(n9146), .ZN(n9147) );
  NOR2_X1 U10412 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  XNOR2_X1 U10413 ( .A(n9150), .B(n9149), .ZN(n9157) );
  NOR2_X1 U10414 ( .A1(n9151), .A2(n9164), .ZN(n9155) );
  AOI22_X1 U10415 ( .A1(n9306), .A2(n9162), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9152) );
  OAI21_X1 U10416 ( .B1(n9153), .B2(n9267), .A(n9152), .ZN(n9154) );
  AOI211_X1 U10417 ( .C1(n9460), .C2(n9168), .A(n9155), .B(n9154), .ZN(n9156)
         );
  OAI21_X1 U10418 ( .B1(n9157), .B2(n9172), .A(n9156), .ZN(P1_U3238) );
  XNOR2_X1 U10419 ( .A(n9160), .B(n9159), .ZN(n9161) );
  XNOR2_X1 U10420 ( .A(n9158), .B(n9161), .ZN(n9173) );
  NAND2_X1 U10421 ( .A1(n9162), .A2(n9176), .ZN(n9163) );
  NAND2_X1 U10422 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10140)
         );
  OAI211_X1 U10423 ( .C1(n9164), .C2(n9422), .A(n9163), .B(n10140), .ZN(n9165)
         );
  AOI21_X1 U10424 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9171) );
  NAND2_X1 U10425 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  OAI211_X1 U10426 ( .C1(n9173), .C2(n9172), .A(n9171), .B(n9170), .ZN(
        P1_U3239) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9174), .S(n10079), .Z(
        P1_U3585) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9246), .S(n10079), .Z(
        P1_U3584) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9257), .S(n10079), .Z(
        P1_U3583) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9275), .S(n10079), .Z(
        P1_U3582) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9291), .S(n10079), .Z(
        P1_U3581) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9306), .S(n10079), .Z(
        P1_U3580) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9290), .S(n10079), .Z(
        P1_U3579) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9305), .S(n10079), .Z(
        P1_U3578) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9365), .S(n10079), .Z(
        P1_U3577) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9381), .S(n10079), .Z(
        P1_U3576) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9396), .S(n10079), .Z(
        P1_U3575) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9412), .S(n10079), .Z(
        P1_U3574) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9395), .S(n10079), .Z(
        P1_U3573) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9989), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9175), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9987), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9176), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9177), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9178), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9179), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9180), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9181), .S(n10079), .Z(
        P1_U3564) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9182), .S(n10079), .Z(
        P1_U3563) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9183), .S(n10079), .Z(
        P1_U3562) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9184), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9185), .S(n10079), .Z(
        P1_U3560) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9186), .S(n10079), .Z(
        P1_U3559) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9187), .S(n10079), .Z(
        P1_U3558) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9188), .S(n10079), .Z(
        P1_U3557) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6837), .S(n10079), .Z(
        P1_U3556) );
  NAND2_X1 U10457 ( .A1(n10120), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9191) );
  OAI21_X1 U10458 ( .B1(n10120), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9191), .ZN(
        n10116) );
  NOR2_X1 U10459 ( .A1(n9192), .A2(n9210), .ZN(n9193) );
  NOR2_X1 U10460 ( .A1(n7840), .A2(n10129), .ZN(n10128) );
  NOR2_X1 U10461 ( .A1(n9194), .A2(n9212), .ZN(n9195) );
  XNOR2_X1 U10462 ( .A(n9194), .B(n9212), .ZN(n10143) );
  NOR2_X1 U10463 ( .A1(n10142), .A2(n10143), .ZN(n10141) );
  NAND2_X1 U10464 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10157), .ZN(n9196) );
  OAI21_X1 U10465 ( .B1(n10157), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9196), .ZN(
        n10153) );
  NOR2_X1 U10466 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  AOI21_X1 U10467 ( .B1(n10157), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10152), 
        .ZN(n10167) );
  NAND2_X1 U10468 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10170), .ZN(n9197) );
  OAI21_X1 U10469 ( .B1(n10170), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9197), .ZN(
        n10166) );
  NOR2_X1 U10470 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  INV_X1 U10471 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U10472 ( .A1(n10185), .A2(n9199), .ZN(n9198) );
  AOI21_X1 U10473 ( .B1(n10185), .B2(n9199), .A(n9198), .ZN(n10180) );
  INV_X1 U10474 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9218) );
  XNOR2_X1 U10475 ( .A(n10185), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10188) );
  INV_X1 U10476 ( .A(n10170), .ZN(n9216) );
  INV_X1 U10477 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9215) );
  XOR2_X1 U10478 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10170), .Z(n10174) );
  INV_X1 U10479 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U10480 ( .A1(n10157), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9200) );
  AOI21_X1 U10481 ( .B1(n10157), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9200), .ZN(
        n10159) );
  INV_X1 U10482 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10030) );
  OR2_X1 U10483 ( .A1(n10120), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9208) );
  AOI21_X1 U10484 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n10122) );
  INV_X1 U10485 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9204) );
  OR2_X1 U10486 ( .A1(n10120), .A2(n9204), .ZN(n9206) );
  NAND2_X1 U10487 ( .A1(n10120), .A2(n9204), .ZN(n9205) );
  AND2_X1 U10488 ( .A1(n9206), .A2(n9205), .ZN(n10123) );
  NOR2_X1 U10489 ( .A1(n10122), .A2(n10123), .ZN(n10121) );
  INV_X1 U10490 ( .A(n10121), .ZN(n9207) );
  NOR2_X1 U10491 ( .A1(n9210), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9209) );
  AOI21_X1 U10492 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9210), .A(n9209), .ZN(
        n10135) );
  NOR2_X1 U10493 ( .A1(n10134), .A2(n10135), .ZN(n10133) );
  AOI21_X1 U10494 ( .B1(n9210), .B2(n10030), .A(n10133), .ZN(n9211) );
  NAND2_X1 U10495 ( .A1(n10146), .A2(n9211), .ZN(n9213) );
  XNOR2_X1 U10496 ( .A(n9212), .B(n9211), .ZN(n10148) );
  NAND2_X1 U10497 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10148), .ZN(n10147) );
  NAND2_X1 U10498 ( .A1(n9213), .A2(n10147), .ZN(n10160) );
  NAND2_X1 U10499 ( .A1(n10159), .A2(n10160), .ZN(n10158) );
  OAI21_X1 U10500 ( .B1(n9214), .B2(n10015), .A(n10158), .ZN(n10173) );
  NAND2_X1 U10501 ( .A1(n10174), .A2(n10173), .ZN(n10171) );
  OAI21_X1 U10502 ( .B1(n9216), .B2(n9215), .A(n10171), .ZN(n10187) );
  NOR2_X1 U10503 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  AOI21_X1 U10504 ( .B1(n9218), .B2(n9217), .A(n10186), .ZN(n9220) );
  INV_X1 U10505 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9219) );
  XOR2_X1 U10506 ( .A(n9220), .B(n9219), .Z(n9222) );
  OAI22_X1 U10507 ( .A1(n9226), .A2(n10178), .B1(n9222), .B2(n10190), .ZN(
        n9221) );
  INV_X1 U10508 ( .A(n9221), .ZN(n9228) );
  NAND2_X1 U10509 ( .A1(n9222), .A2(n10172), .ZN(n9223) );
  NAND2_X1 U10510 ( .A1(n9223), .A2(n10074), .ZN(n9224) );
  AOI21_X1 U10511 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9227) );
  MUX2_X1 U10512 ( .A(n9228), .B(n9227), .S(n9342), .Z(n9232) );
  INV_X1 U10513 ( .A(n9229), .ZN(n9230) );
  AOI21_X1 U10514 ( .B1(n10101), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9230), .ZN(
        n9231) );
  NAND2_X1 U10515 ( .A1(n9232), .A2(n9231), .ZN(P1_U3260) );
  AOI21_X1 U10516 ( .B1(n9244), .B2(n9234), .A(n9233), .ZN(n9235) );
  INV_X1 U10517 ( .A(n9235), .ZN(n9454) );
  INV_X1 U10518 ( .A(n9250), .ZN(n9238) );
  INV_X1 U10519 ( .A(n9236), .ZN(n9237) );
  AOI211_X1 U10520 ( .C1(n9451), .C2(n9238), .A(n10265), .B(n9237), .ZN(n9450)
         );
  AOI22_X1 U10521 ( .A1(n9239), .A2(n9993), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10216), .ZN(n9240) );
  OAI21_X1 U10522 ( .B1(n9241), .B2(n9432), .A(n9240), .ZN(n9248) );
  AND2_X1 U10523 ( .A1(n9254), .A2(n9242), .ZN(n9245) );
  OAI21_X1 U10524 ( .B1(n9245), .B2(n9244), .A(n9243), .ZN(n9247) );
  XOR2_X1 U10525 ( .A(n9255), .B(n9249), .Z(n9459) );
  AOI21_X1 U10526 ( .B1(n9455), .B2(n9264), .A(n9250), .ZN(n9456) );
  AOI22_X1 U10527 ( .A1(n9251), .A2(n9993), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10216), .ZN(n9252) );
  OAI21_X1 U10528 ( .B1(n9253), .B2(n9432), .A(n9252), .ZN(n9261) );
  OAI211_X1 U10529 ( .C1(n9256), .C2(n9255), .A(n9254), .B(n9985), .ZN(n9259)
         );
  AOI22_X1 U10530 ( .A1(n9257), .A2(n9990), .B1(n9988), .B2(n9291), .ZN(n9258)
         );
  AND2_X1 U10531 ( .A1(n9259), .A2(n9258), .ZN(n9458) );
  NOR2_X1 U10532 ( .A1(n9458), .A2(n10216), .ZN(n9260) );
  AOI211_X1 U10533 ( .C1(n10212), .C2(n9456), .A(n9261), .B(n9260), .ZN(n9262)
         );
  OAI21_X1 U10534 ( .B1(n9459), .B2(n10004), .A(n9262), .ZN(P1_U3264) );
  XNOR2_X1 U10535 ( .A(n9263), .B(n9274), .ZN(n9464) );
  INV_X1 U10536 ( .A(n9283), .ZN(n9266) );
  INV_X1 U10537 ( .A(n9264), .ZN(n9265) );
  AOI21_X1 U10538 ( .B1(n9460), .B2(n9266), .A(n9265), .ZN(n9461) );
  INV_X1 U10539 ( .A(n9267), .ZN(n9268) );
  AOI22_X1 U10540 ( .A1(n9268), .A2(n9993), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10216), .ZN(n9269) );
  OAI21_X1 U10541 ( .B1(n9270), .B2(n9432), .A(n9269), .ZN(n9278) );
  NAND2_X1 U10542 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  XOR2_X1 U10543 ( .A(n9274), .B(n9273), .Z(n9276) );
  AOI222_X1 U10544 ( .A1(n9985), .A2(n9276), .B1(n9275), .B2(n9990), .C1(n9306), .C2(n9988), .ZN(n9463) );
  NOR2_X1 U10545 ( .A1(n9463), .A2(n10216), .ZN(n9277) );
  AOI211_X1 U10546 ( .C1(n9461), .C2(n10212), .A(n9278), .B(n9277), .ZN(n9279)
         );
  OAI21_X1 U10547 ( .B1(n10004), .B2(n9464), .A(n9279), .ZN(P1_U3265) );
  OAI21_X1 U10548 ( .B1(n9280), .B2(n9288), .A(n9281), .ZN(n9282) );
  INV_X1 U10549 ( .A(n9282), .ZN(n9469) );
  AOI21_X1 U10550 ( .B1(n9465), .B2(n9309), .A(n9283), .ZN(n9466) );
  INV_X1 U10551 ( .A(n9465), .ZN(n9287) );
  INV_X1 U10552 ( .A(n9284), .ZN(n9285) );
  AOI22_X1 U10553 ( .A1(n9285), .A2(n9993), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n10216), .ZN(n9286) );
  OAI21_X1 U10554 ( .B1(n9287), .B2(n9432), .A(n9286), .ZN(n9294) );
  XNOR2_X1 U10555 ( .A(n9289), .B(n9288), .ZN(n9292) );
  AOI222_X1 U10556 ( .A1(n9985), .A2(n9292), .B1(n9291), .B2(n9990), .C1(n9290), .C2(n9988), .ZN(n9468) );
  NOR2_X1 U10557 ( .A1(n9468), .A2(n10216), .ZN(n9293) );
  AOI211_X1 U10558 ( .C1(n9466), .C2(n10212), .A(n9294), .B(n9293), .ZN(n9295)
         );
  OAI21_X1 U10559 ( .B1(n9469), .B2(n10004), .A(n9295), .ZN(P1_U3266) );
  AND2_X1 U10560 ( .A1(n9296), .A2(n9302), .ZN(n9297) );
  NOR2_X1 U10561 ( .A1(n9298), .A2(n9297), .ZN(n9470) );
  INV_X1 U10562 ( .A(n9470), .ZN(n9316) );
  AOI22_X1 U10563 ( .A1(n9471), .A2(n10213), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10216), .ZN(n9315) );
  INV_X1 U10564 ( .A(n9300), .ZN(n9301) );
  OR2_X1 U10565 ( .A1(n9299), .A2(n9301), .ZN(n9303) );
  XNOR2_X1 U10566 ( .A(n9303), .B(n9302), .ZN(n9304) );
  NAND2_X1 U10567 ( .A1(n9304), .A2(n9985), .ZN(n9308) );
  AOI22_X1 U10568 ( .A1(n9306), .A2(n9990), .B1(n9988), .B2(n9305), .ZN(n9307)
         );
  NAND2_X1 U10569 ( .A1(n9308), .A2(n9307), .ZN(n9475) );
  OAI211_X1 U10570 ( .C1(n9310), .C2(n4525), .A(n9999), .B(n9309), .ZN(n9473)
         );
  INV_X1 U10571 ( .A(n9311), .ZN(n9312) );
  OAI22_X1 U10572 ( .A1(n9473), .A2(n9342), .B1(n10221), .B2(n9312), .ZN(n9313) );
  OAI21_X1 U10573 ( .B1(n9475), .B2(n9313), .A(n10207), .ZN(n9314) );
  OAI211_X1 U10574 ( .C1(n9316), .C2(n10004), .A(n9315), .B(n9314), .ZN(
        P1_U3267) );
  XNOR2_X1 U10575 ( .A(n9317), .B(n9318), .ZN(n9482) );
  NOR2_X1 U10576 ( .A1(n9320), .A2(n9319), .ZN(n9322) );
  AOI21_X1 U10577 ( .B1(n9322), .B2(n9321), .A(n9299), .ZN(n9323) );
  OAI222_X1 U10578 ( .A1(n9425), .A2(n9325), .B1(n9423), .B2(n9324), .C1(n9421), .C2(n9323), .ZN(n9478) );
  INV_X1 U10579 ( .A(n9480), .ZN(n9330) );
  AOI211_X1 U10580 ( .C1(n9480), .C2(n9339), .A(n10265), .B(n4525), .ZN(n9479)
         );
  NAND2_X1 U10581 ( .A1(n9479), .A2(n9428), .ZN(n9329) );
  INV_X1 U10582 ( .A(n9326), .ZN(n9327) );
  AOI22_X1 U10583 ( .A1(n9327), .A2(n9993), .B1(n10216), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9328) );
  OAI211_X1 U10584 ( .C1(n9330), .C2(n9432), .A(n9329), .B(n9328), .ZN(n9331)
         );
  AOI21_X1 U10585 ( .B1(n9478), .B2(n10207), .A(n9331), .ZN(n9332) );
  OAI21_X1 U10586 ( .B1(n9482), .B2(n10004), .A(n9332), .ZN(P1_U3268) );
  XNOR2_X1 U10587 ( .A(n9333), .B(n9334), .ZN(n9487) );
  AOI22_X1 U10588 ( .A1(n9485), .A2(n10213), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10216), .ZN(n9346) );
  XNOR2_X1 U10589 ( .A(n9335), .B(n9334), .ZN(n9336) );
  OAI222_X1 U10590 ( .A1(n9425), .A2(n9338), .B1(n9423), .B2(n9337), .C1(n9336), .C2(n9421), .ZN(n9483) );
  INV_X1 U10591 ( .A(n9339), .ZN(n9340) );
  AOI211_X1 U10592 ( .C1(n9485), .C2(n9353), .A(n10265), .B(n9340), .ZN(n9484)
         );
  INV_X1 U10593 ( .A(n9484), .ZN(n9343) );
  OAI22_X1 U10594 ( .A1(n9343), .A2(n9342), .B1(n10221), .B2(n9341), .ZN(n9344) );
  OAI21_X1 U10595 ( .B1(n9483), .B2(n9344), .A(n10207), .ZN(n9345) );
  OAI211_X1 U10596 ( .C1(n9487), .C2(n10004), .A(n9346), .B(n9345), .ZN(
        P1_U3269) );
  NAND2_X1 U10597 ( .A1(n9401), .A2(n9347), .ZN(n9349) );
  NAND2_X1 U10598 ( .A1(n9349), .A2(n9348), .ZN(n9352) );
  OAI21_X1 U10599 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9492) );
  INV_X1 U10600 ( .A(n9375), .ZN(n9355) );
  INV_X1 U10601 ( .A(n9353), .ZN(n9354) );
  AOI211_X1 U10602 ( .C1(n9489), .C2(n9355), .A(n10265), .B(n9354), .ZN(n9488)
         );
  INV_X1 U10603 ( .A(n9356), .ZN(n9357) );
  AOI22_X1 U10604 ( .A1(n10216), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9357), 
        .B2(n9993), .ZN(n9358) );
  OAI21_X1 U10605 ( .B1(n9359), .B2(n9432), .A(n9358), .ZN(n9368) );
  AND2_X1 U10606 ( .A1(n9361), .A2(n9360), .ZN(n9364) );
  OAI21_X1 U10607 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9366) );
  AOI222_X1 U10608 ( .A1(n9985), .A2(n9366), .B1(n9396), .B2(n9988), .C1(n9365), .C2(n9990), .ZN(n9491) );
  NOR2_X1 U10609 ( .A1(n9491), .A2(n10216), .ZN(n9367) );
  AOI211_X1 U10610 ( .C1(n9488), .C2(n9428), .A(n9368), .B(n9367), .ZN(n9369)
         );
  OAI21_X1 U10611 ( .B1(n10004), .B2(n9492), .A(n9369), .ZN(P1_U3270) );
  NAND2_X1 U10612 ( .A1(n9401), .A2(n9410), .ZN(n9387) );
  NAND2_X1 U10613 ( .A1(n9387), .A2(n9370), .ZN(n9372) );
  AND2_X1 U10614 ( .A1(n9372), .A2(n9371), .ZN(n9374) );
  XNOR2_X1 U10615 ( .A(n9374), .B(n9373), .ZN(n9497) );
  AOI21_X1 U10616 ( .B1(n9493), .B2(n9389), .A(n9375), .ZN(n9494) );
  AOI22_X1 U10617 ( .A1(n10216), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9376), 
        .B2(n9993), .ZN(n9377) );
  OAI21_X1 U10618 ( .B1(n9378), .B2(n9432), .A(n9377), .ZN(n9384) );
  XNOR2_X1 U10619 ( .A(n9380), .B(n9379), .ZN(n9382) );
  AOI222_X1 U10620 ( .A1(n9985), .A2(n9382), .B1(n9381), .B2(n9990), .C1(n9412), .C2(n9988), .ZN(n9496) );
  NOR2_X1 U10621 ( .A1(n9496), .A2(n10216), .ZN(n9383) );
  AOI211_X1 U10622 ( .C1(n9494), .C2(n10212), .A(n9384), .B(n9383), .ZN(n9385)
         );
  OAI21_X1 U10623 ( .B1(n10004), .B2(n9497), .A(n9385), .ZN(P1_U3271) );
  NAND2_X1 U10624 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  XOR2_X1 U10625 ( .A(n9394), .B(n9388), .Z(n9502) );
  INV_X1 U10626 ( .A(n9389), .ZN(n9390) );
  AOI21_X1 U10627 ( .B1(n9498), .B2(n9402), .A(n9390), .ZN(n9499) );
  AOI22_X1 U10628 ( .A1(n10216), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9391), 
        .B2(n9993), .ZN(n9392) );
  OAI21_X1 U10629 ( .B1(n4815), .B2(n9432), .A(n9392), .ZN(n9399) );
  XNOR2_X1 U10630 ( .A(n9393), .B(n9394), .ZN(n9397) );
  AOI222_X1 U10631 ( .A1(n9985), .A2(n9397), .B1(n9396), .B2(n9990), .C1(n9395), .C2(n9988), .ZN(n9501) );
  NOR2_X1 U10632 ( .A1(n9501), .A2(n10216), .ZN(n9398) );
  AOI211_X1 U10633 ( .C1(n9499), .C2(n10212), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OAI21_X1 U10634 ( .B1(n10004), .B2(n9502), .A(n9400), .ZN(P1_U3272) );
  XNOR2_X1 U10635 ( .A(n9401), .B(n9410), .ZN(n9507) );
  INV_X1 U10636 ( .A(n9426), .ZN(n9404) );
  INV_X1 U10637 ( .A(n9402), .ZN(n9403) );
  AOI21_X1 U10638 ( .B1(n9503), .B2(n9404), .A(n9403), .ZN(n9504) );
  AOI22_X1 U10639 ( .A1(n10216), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9405), 
        .B2(n9993), .ZN(n9406) );
  OAI21_X1 U10640 ( .B1(n9407), .B2(n9432), .A(n9406), .ZN(n9415) );
  NAND2_X1 U10641 ( .A1(n9409), .A2(n9408), .ZN(n9411) );
  XNOR2_X1 U10642 ( .A(n9411), .B(n9410), .ZN(n9413) );
  AOI222_X1 U10643 ( .A1(n9985), .A2(n9413), .B1(n9989), .B2(n9988), .C1(n9412), .C2(n9990), .ZN(n9506) );
  NOR2_X1 U10644 ( .A1(n9506), .A2(n10216), .ZN(n9414) );
  AOI211_X1 U10645 ( .C1(n9504), .C2(n10212), .A(n9415), .B(n9414), .ZN(n9416)
         );
  OAI21_X1 U10646 ( .B1(n10004), .B2(n9507), .A(n9416), .ZN(P1_U3273) );
  XOR2_X1 U10647 ( .A(n9417), .B(n9418), .Z(n9513) );
  XNOR2_X1 U10648 ( .A(n9419), .B(n9418), .ZN(n9420) );
  OAI222_X1 U10649 ( .A1(n9425), .A2(n9424), .B1(n9423), .B2(n9422), .C1(n9421), .C2(n9420), .ZN(n9508) );
  INV_X1 U10650 ( .A(n10002), .ZN(n9427) );
  AOI211_X1 U10651 ( .C1(n9510), .C2(n9427), .A(n10265), .B(n9426), .ZN(n9509)
         );
  NAND2_X1 U10652 ( .A1(n9509), .A2(n9428), .ZN(n9431) );
  AOI22_X1 U10653 ( .A1(n10216), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9429), 
        .B2(n9993), .ZN(n9430) );
  OAI211_X1 U10654 ( .C1(n9433), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9434)
         );
  AOI21_X1 U10655 ( .B1(n9508), .B2(n10207), .A(n9434), .ZN(n9435) );
  OAI21_X1 U10656 ( .B1(n9513), .B2(n10004), .A(n9435), .ZN(P1_U3274) );
  NAND2_X1 U10657 ( .A1(n9436), .A2(n9999), .ZN(n9437) );
  OAI211_X1 U10658 ( .C1(n9438), .C2(n10263), .A(n9437), .B(n9441), .ZN(n9514)
         );
  MUX2_X1 U10659 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9514), .S(n4456), .Z(
        P1_U3554) );
  NAND3_X1 U10660 ( .A1(n9440), .A2(n9999), .A3(n9439), .ZN(n9442) );
  OAI211_X1 U10661 ( .C1(n9443), .C2(n10263), .A(n9442), .B(n9441), .ZN(n9515)
         );
  MUX2_X1 U10662 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9515), .S(n4456), .Z(
        P1_U3553) );
  AOI22_X1 U10663 ( .A1(n9445), .A2(n9999), .B1(n9511), .B2(n9444), .ZN(n9446)
         );
  OAI21_X1 U10664 ( .B1(n9449), .B2(n10016), .A(n9448), .ZN(n9516) );
  MUX2_X1 U10665 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9516), .S(n4456), .Z(
        P1_U3552) );
  AOI21_X1 U10666 ( .B1(n9511), .B2(n9451), .A(n9450), .ZN(n9452) );
  OAI211_X1 U10667 ( .C1(n9454), .C2(n10016), .A(n9453), .B(n9452), .ZN(n9517)
         );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9517), .S(n4456), .Z(
        P1_U3551) );
  AOI22_X1 U10669 ( .A1(n9456), .A2(n9999), .B1(n9511), .B2(n9455), .ZN(n9457)
         );
  OAI211_X1 U10670 ( .C1(n9459), .C2(n10016), .A(n9458), .B(n9457), .ZN(n9518)
         );
  MUX2_X1 U10671 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9518), .S(n4456), .Z(
        P1_U3550) );
  AOI22_X1 U10672 ( .A1(n9461), .A2(n9999), .B1(n9511), .B2(n9460), .ZN(n9462)
         );
  OAI211_X1 U10673 ( .C1(n9464), .C2(n10016), .A(n9463), .B(n9462), .ZN(n9519)
         );
  MUX2_X1 U10674 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9519), .S(n4456), .Z(
        P1_U3549) );
  AOI22_X1 U10675 ( .A1(n9466), .A2(n9999), .B1(n9511), .B2(n9465), .ZN(n9467)
         );
  OAI211_X1 U10676 ( .C1(n9469), .C2(n10016), .A(n9468), .B(n9467), .ZN(n9520)
         );
  MUX2_X1 U10677 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9520), .S(n4456), .Z(
        P1_U3548) );
  NAND2_X1 U10678 ( .A1(n9470), .A2(n10252), .ZN(n9477) );
  NAND2_X1 U10679 ( .A1(n9471), .A2(n9511), .ZN(n9472) );
  NAND2_X1 U10680 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  NOR2_X1 U10681 ( .A1(n9475), .A2(n9474), .ZN(n9476) );
  NAND2_X1 U10682 ( .A1(n9477), .A2(n9476), .ZN(n9521) );
  MUX2_X1 U10683 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9521), .S(n4456), .Z(
        P1_U3547) );
  AOI211_X1 U10684 ( .C1(n9511), .C2(n9480), .A(n9479), .B(n9478), .ZN(n9481)
         );
  OAI21_X1 U10685 ( .B1(n10016), .B2(n9482), .A(n9481), .ZN(n9522) );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9522), .S(n4456), .Z(
        P1_U3546) );
  AOI211_X1 U10687 ( .C1(n9511), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9486)
         );
  OAI21_X1 U10688 ( .B1(n10016), .B2(n9487), .A(n9486), .ZN(n9523) );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9523), .S(n4456), .Z(
        P1_U3545) );
  AOI21_X1 U10690 ( .B1(n9511), .B2(n9489), .A(n9488), .ZN(n9490) );
  OAI211_X1 U10691 ( .C1(n9492), .C2(n10016), .A(n9491), .B(n9490), .ZN(n9524)
         );
  MUX2_X1 U10692 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9524), .S(n4456), .Z(
        P1_U3544) );
  AOI22_X1 U10693 ( .A1(n9494), .A2(n9999), .B1(n9511), .B2(n9493), .ZN(n9495)
         );
  OAI211_X1 U10694 ( .C1(n9497), .C2(n10016), .A(n9496), .B(n9495), .ZN(n9525)
         );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9525), .S(n4456), .Z(
        P1_U3543) );
  AOI22_X1 U10696 ( .A1(n9499), .A2(n9999), .B1(n9511), .B2(n9498), .ZN(n9500)
         );
  OAI211_X1 U10697 ( .C1(n9502), .C2(n10016), .A(n9501), .B(n9500), .ZN(n9526)
         );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9526), .S(n4456), .Z(
        P1_U3542) );
  AOI22_X1 U10699 ( .A1(n9504), .A2(n9999), .B1(n9511), .B2(n9503), .ZN(n9505)
         );
  OAI211_X1 U10700 ( .C1(n9507), .C2(n10016), .A(n9506), .B(n9505), .ZN(n9527)
         );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9527), .S(n4456), .Z(
        P1_U3541) );
  AOI211_X1 U10702 ( .C1(n9511), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9512)
         );
  OAI21_X1 U10703 ( .B1(n10016), .B2(n9513), .A(n9512), .ZN(n9528) );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9528), .S(n4456), .Z(
        P1_U3540) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9514), .S(n10273), .Z(
        P1_U3522) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9515), .S(n10273), .Z(
        P1_U3521) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9516), .S(n10273), .Z(
        P1_U3520) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9517), .S(n10273), .Z(
        P1_U3519) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9518), .S(n10273), .Z(
        P1_U3518) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9519), .S(n10273), .Z(
        P1_U3517) );
  MUX2_X1 U10711 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9520), .S(n10273), .Z(
        P1_U3516) );
  MUX2_X1 U10712 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9521), .S(n10273), .Z(
        P1_U3515) );
  MUX2_X1 U10713 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9522), .S(n10273), .Z(
        P1_U3514) );
  MUX2_X1 U10714 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9523), .S(n10273), .Z(
        P1_U3513) );
  MUX2_X1 U10715 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9524), .S(n10273), .Z(
        P1_U3512) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9525), .S(n10273), .Z(
        P1_U3511) );
  MUX2_X1 U10717 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9526), .S(n10273), .Z(
        P1_U3510) );
  MUX2_X1 U10718 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9527), .S(n10273), .Z(
        P1_U3508) );
  MUX2_X1 U10719 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9528), .S(n10273), .Z(
        n9880) );
  AOI22_X1 U10720 ( .A1(SI_23_), .A2(keyinput179), .B1(P1_IR_REG_10__SCAN_IN), 
        .B2(keyinput175), .ZN(n9529) );
  OAI221_X1 U10721 ( .B1(SI_23_), .B2(keyinput179), .C1(P1_IR_REG_10__SCAN_IN), 
        .C2(keyinput175), .A(n9529), .ZN(n9536) );
  AOI22_X1 U10722 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(keyinput213), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(keyinput181), .ZN(n9530) );
  OAI221_X1 U10723 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(keyinput213), .C1(
        P1_DATAO_REG_1__SCAN_IN), .C2(keyinput181), .A(n9530), .ZN(n9535) );
  AOI22_X1 U10724 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput200), .B1(
        P1_D_REG_16__SCAN_IN), .B2(keyinput171), .ZN(n9531) );
  OAI221_X1 U10725 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput200), .C1(
        P1_D_REG_16__SCAN_IN), .C2(keyinput171), .A(n9531), .ZN(n9534) );
  AOI22_X1 U10726 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(keyinput186), .B1(
        P1_REG2_REG_21__SCAN_IN), .B2(keyinput198), .ZN(n9532) );
  OAI221_X1 U10727 ( .B1(P2_REG2_REG_22__SCAN_IN), .B2(keyinput186), .C1(
        P1_REG2_REG_21__SCAN_IN), .C2(keyinput198), .A(n9532), .ZN(n9533) );
  NOR4_X1 U10728 ( .A1(n9536), .A2(n9535), .A3(n9534), .A4(n9533), .ZN(n9564)
         );
  AOI22_X1 U10729 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput143), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput202), .ZN(n9537) );
  OAI221_X1 U10730 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput143), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput202), .A(n9537), .ZN(n9544) );
  AOI22_X1 U10731 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput148), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(keyinput252), .ZN(n9538) );
  OAI221_X1 U10732 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput148), .C1(
        P1_DATAO_REG_24__SCAN_IN), .C2(keyinput252), .A(n9538), .ZN(n9543) );
  AOI22_X1 U10733 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput146), .B1(
        P1_REG1_REG_14__SCAN_IN), .B2(keyinput194), .ZN(n9539) );
  OAI221_X1 U10734 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput146), .C1(
        P1_REG1_REG_14__SCAN_IN), .C2(keyinput194), .A(n9539), .ZN(n9542) );
  AOI22_X1 U10735 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput253), .B1(
        P1_REG1_REG_13__SCAN_IN), .B2(keyinput210), .ZN(n9540) );
  OAI221_X1 U10736 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput253), .C1(
        P1_REG1_REG_13__SCAN_IN), .C2(keyinput210), .A(n9540), .ZN(n9541) );
  NOR4_X1 U10737 ( .A1(n9544), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n9563)
         );
  AOI22_X1 U10738 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput132), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput247), .ZN(n9545) );
  OAI221_X1 U10739 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput132), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput247), .A(n9545), .ZN(n9552) );
  AOI22_X1 U10740 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput196), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput250), .ZN(n9546) );
  OAI221_X1 U10741 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput196), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput250), .A(n9546), .ZN(n9551) );
  AOI22_X1 U10742 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput193), .B1(
        P1_REG1_REG_10__SCAN_IN), .B2(keyinput208), .ZN(n9547) );
  OAI221_X1 U10743 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput193), .C1(
        P1_REG1_REG_10__SCAN_IN), .C2(keyinput208), .A(n9547), .ZN(n9550) );
  AOI22_X1 U10744 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(keyinput137), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput185), .ZN(n9548) );
  OAI221_X1 U10745 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(keyinput137), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput185), .A(n9548), .ZN(n9549) );
  NOR4_X1 U10746 ( .A1(n9552), .A2(n9551), .A3(n9550), .A4(n9549), .ZN(n9562)
         );
  AOI22_X1 U10747 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput230), .B1(
        P1_REG1_REG_28__SCAN_IN), .B2(keyinput160), .ZN(n9553) );
  OAI221_X1 U10748 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput230), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput160), .A(n9553), .ZN(n9560) );
  AOI22_X1 U10749 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(keyinput205), .B1(
        P2_REG0_REG_23__SCAN_IN), .B2(keyinput246), .ZN(n9554) );
  OAI221_X1 U10750 ( .B1(P2_REG0_REG_29__SCAN_IN), .B2(keyinput205), .C1(
        P2_REG0_REG_23__SCAN_IN), .C2(keyinput246), .A(n9554), .ZN(n9559) );
  AOI22_X1 U10751 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(keyinput220), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput209), .ZN(n9555) );
  OAI221_X1 U10752 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(keyinput220), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput209), .A(n9555), .ZN(n9558) );
  AOI22_X1 U10753 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput222), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput140), .ZN(n9556) );
  OAI221_X1 U10754 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput222), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput140), .A(n9556), .ZN(n9557) );
  NOR4_X1 U10755 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n9561)
         );
  NAND4_X1 U10756 ( .A1(n9564), .A2(n9563), .A3(n9562), .A4(n9561), .ZN(n9624)
         );
  AOI22_X1 U10757 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput190), .B1(SI_21_), 
        .B2(keyinput177), .ZN(n9565) );
  OAI221_X1 U10758 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput190), .C1(SI_21_), 
        .C2(keyinput177), .A(n9565), .ZN(n9572) );
  AOI22_X1 U10759 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput214), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput197), .ZN(n9566) );
  OAI221_X1 U10760 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput214), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput197), .A(n9566), .ZN(n9571) );
  AOI22_X1 U10761 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput164), .B1(
        P1_REG2_REG_17__SCAN_IN), .B2(keyinput223), .ZN(n9567) );
  OAI221_X1 U10762 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput164), .C1(
        P1_REG2_REG_17__SCAN_IN), .C2(keyinput223), .A(n9567), .ZN(n9570) );
  AOI22_X1 U10763 ( .A1(P2_D_REG_18__SCAN_IN), .A2(keyinput128), .B1(
        P1_D_REG_24__SCAN_IN), .B2(keyinput229), .ZN(n9568) );
  OAI221_X1 U10764 ( .B1(P2_D_REG_18__SCAN_IN), .B2(keyinput128), .C1(
        P1_D_REG_24__SCAN_IN), .C2(keyinput229), .A(n9568), .ZN(n9569) );
  NOR4_X1 U10765 ( .A1(n9572), .A2(n9571), .A3(n9570), .A4(n9569), .ZN(n9600)
         );
  AOI22_X1 U10766 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput234), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput221), .ZN(n9573) );
  OAI221_X1 U10767 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput234), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput221), .A(n9573), .ZN(n9580) );
  AOI22_X1 U10768 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput167), .B1(
        P2_IR_REG_0__SCAN_IN), .B2(keyinput226), .ZN(n9574) );
  OAI221_X1 U10769 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput167), .C1(
        P2_IR_REG_0__SCAN_IN), .C2(keyinput226), .A(n9574), .ZN(n9579) );
  AOI22_X1 U10770 ( .A1(P1_REG0_REG_22__SCAN_IN), .A2(keyinput191), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput178), .ZN(n9575) );
  OAI221_X1 U10771 ( .B1(P1_REG0_REG_22__SCAN_IN), .B2(keyinput191), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput178), .A(n9575), .ZN(n9578) );
  AOI22_X1 U10772 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput224), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput215), .ZN(n9576) );
  OAI221_X1 U10773 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput224), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput215), .A(n9576), .ZN(n9577) );
  NOR4_X1 U10774 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n9599)
         );
  AOI22_X1 U10775 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput192), .B1(
        P2_IR_REG_3__SCAN_IN), .B2(keyinput243), .ZN(n9581) );
  OAI221_X1 U10776 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput192), .C1(
        P2_IR_REG_3__SCAN_IN), .C2(keyinput243), .A(n9581), .ZN(n9588) );
  AOI22_X1 U10777 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput130), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput187), .ZN(n9582) );
  OAI221_X1 U10778 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput130), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput187), .A(n9582), .ZN(n9587) );
  AOI22_X1 U10779 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(keyinput233), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput183), .ZN(n9583) );
  OAI221_X1 U10780 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(keyinput233), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput183), .A(n9583), .ZN(n9586) );
  AOI22_X1 U10781 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput170), .B1(
        P1_D_REG_27__SCAN_IN), .B2(keyinput225), .ZN(n9584) );
  OAI221_X1 U10782 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput170), .C1(
        P1_D_REG_27__SCAN_IN), .C2(keyinput225), .A(n9584), .ZN(n9585) );
  NOR4_X1 U10783 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(n9598)
         );
  AOI22_X1 U10784 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput141), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput227), .ZN(n9589) );
  OAI221_X1 U10785 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput141), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput227), .A(n9589), .ZN(n9596) );
  AOI22_X1 U10786 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(keyinput237), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput206), .ZN(n9590) );
  OAI221_X1 U10787 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(keyinput237), .C1(
        P1_D_REG_23__SCAN_IN), .C2(keyinput206), .A(n9590), .ZN(n9595) );
  AOI22_X1 U10788 ( .A1(P2_D_REG_7__SCAN_IN), .A2(keyinput242), .B1(
        P1_REG2_REG_28__SCAN_IN), .B2(keyinput212), .ZN(n9591) );
  OAI221_X1 U10789 ( .B1(P2_D_REG_7__SCAN_IN), .B2(keyinput242), .C1(
        P1_REG2_REG_28__SCAN_IN), .C2(keyinput212), .A(n9591), .ZN(n9594) );
  AOI22_X1 U10790 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput203), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput138), .ZN(n9592) );
  OAI221_X1 U10791 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput203), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput138), .A(n9592), .ZN(n9593) );
  NOR4_X1 U10792 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9597)
         );
  NAND4_X1 U10793 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9623)
         );
  AOI22_X1 U10794 ( .A1(n9748), .A2(keyinput139), .B1(n9602), .B2(keyinput161), 
        .ZN(n9601) );
  OAI221_X1 U10795 ( .B1(n9748), .B2(keyinput139), .C1(n9602), .C2(keyinput161), .A(n9601), .ZN(n9610) );
  AOI22_X1 U10796 ( .A1(n9741), .A2(keyinput235), .B1(n9813), .B2(keyinput152), 
        .ZN(n9603) );
  OAI221_X1 U10797 ( .B1(n9741), .B2(keyinput235), .C1(n9813), .C2(keyinput152), .A(n9603), .ZN(n9609) );
  INV_X1 U10798 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10298) );
  XNOR2_X1 U10799 ( .A(n10298), .B(keyinput231), .ZN(n9608) );
  XOR2_X1 U10800 ( .A(n9791), .B(keyinput154), .Z(n9606) );
  XNOR2_X1 U10801 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput180), .ZN(n9605) );
  XNOR2_X1 U10802 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput188), .ZN(n9604) );
  NAND3_X1 U10803 ( .A1(n9606), .A2(n9605), .A3(n9604), .ZN(n9607) );
  OR4_X1 U10804 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n9622)
         );
  AOI22_X1 U10805 ( .A1(n9811), .A2(keyinput195), .B1(n6309), .B2(keyinput168), 
        .ZN(n9611) );
  OAI221_X1 U10806 ( .B1(n9811), .B2(keyinput195), .C1(n6309), .C2(keyinput168), .A(n9611), .ZN(n9620) );
  INV_X1 U10807 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U10808 ( .A1(n10024), .A2(keyinput238), .B1(keyinput182), .B2(
        n10209), .ZN(n9612) );
  OAI221_X1 U10809 ( .B1(n10024), .B2(keyinput238), .C1(n10209), .C2(
        keyinput182), .A(n9612), .ZN(n9619) );
  INV_X1 U10810 ( .A(SI_24_), .ZN(n9614) );
  INV_X1 U10811 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U10812 ( .A1(n9614), .A2(keyinput249), .B1(keyinput232), .B2(n10220), .ZN(n9613) );
  OAI221_X1 U10813 ( .B1(n9614), .B2(keyinput249), .C1(n10220), .C2(
        keyinput232), .A(n9613), .ZN(n9618) );
  AOI22_X1 U10814 ( .A1(n9616), .A2(keyinput189), .B1(n5110), .B2(keyinput228), 
        .ZN(n9615) );
  OAI221_X1 U10815 ( .B1(n9616), .B2(keyinput189), .C1(n5110), .C2(keyinput228), .A(n9615), .ZN(n9617) );
  OR4_X1 U10816 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n9621)
         );
  NOR4_X1 U10817 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(n9647)
         );
  AOI22_X1 U10818 ( .A1(n7067), .A2(keyinput239), .B1(n9626), .B2(keyinput211), 
        .ZN(n9625) );
  OAI221_X1 U10819 ( .B1(n7067), .B2(keyinput239), .C1(n9626), .C2(keyinput211), .A(n9625), .ZN(n9634) );
  AOI22_X1 U10820 ( .A1(n9798), .A2(keyinput176), .B1(n9816), .B2(keyinput244), 
        .ZN(n9627) );
  OAI221_X1 U10821 ( .B1(n9798), .B2(keyinput176), .C1(n9816), .C2(keyinput244), .A(n9627), .ZN(n9633) );
  AOI22_X1 U10822 ( .A1(n9629), .A2(keyinput162), .B1(n10228), .B2(keyinput163), .ZN(n9628) );
  OAI221_X1 U10823 ( .B1(n9629), .B2(keyinput162), .C1(n10228), .C2(
        keyinput163), .A(n9628), .ZN(n9632) );
  AOI22_X1 U10824 ( .A1(n6018), .A2(keyinput204), .B1(n7969), .B2(keyinput201), 
        .ZN(n9630) );
  OAI221_X1 U10825 ( .B1(n6018), .B2(keyinput204), .C1(n7969), .C2(keyinput201), .A(n9630), .ZN(n9631) );
  NOR4_X1 U10826 ( .A1(n9634), .A2(n9633), .A3(n9632), .A4(n9631), .ZN(n9646)
         );
  AOI22_X1 U10827 ( .A1(n5957), .A2(keyinput169), .B1(keyinput217), .B2(n6901), 
        .ZN(n9635) );
  OAI221_X1 U10828 ( .B1(n5957), .B2(keyinput169), .C1(n6901), .C2(keyinput217), .A(n9635), .ZN(n9644) );
  AOI22_X1 U10829 ( .A1(n9815), .A2(keyinput172), .B1(n9637), .B2(keyinput251), 
        .ZN(n9636) );
  OAI221_X1 U10830 ( .B1(n9815), .B2(keyinput172), .C1(n9637), .C2(keyinput251), .A(n9636), .ZN(n9643) );
  INV_X1 U10831 ( .A(SI_29_), .ZN(n9818) );
  AOI22_X1 U10832 ( .A1(n9818), .A2(keyinput145), .B1(n9639), .B2(keyinput156), 
        .ZN(n9638) );
  OAI221_X1 U10833 ( .B1(n9818), .B2(keyinput145), .C1(n9639), .C2(keyinput156), .A(n9638), .ZN(n9642) );
  INV_X1 U10834 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9730) );
  AOI22_X1 U10835 ( .A1(n9728), .A2(keyinput174), .B1(keyinput165), .B2(n9730), 
        .ZN(n9640) );
  OAI221_X1 U10836 ( .B1(n9728), .B2(keyinput174), .C1(n9730), .C2(keyinput165), .A(n9640), .ZN(n9641) );
  NOR4_X1 U10837 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n9645)
         );
  NAND3_X1 U10838 ( .A1(n9647), .A2(n9646), .A3(n9645), .ZN(n9878) );
  AOI22_X1 U10839 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput218), .B1(
        P2_IR_REG_10__SCAN_IN), .B2(keyinput151), .ZN(n9648) );
  OAI221_X1 U10840 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput218), .C1(
        P2_IR_REG_10__SCAN_IN), .C2(keyinput151), .A(n9648), .ZN(n9656) );
  AOI22_X1 U10841 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput135), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput248), .ZN(n9649) );
  OAI221_X1 U10842 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput135), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput248), .A(n9649), .ZN(n9655) );
  AOI22_X1 U10843 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput142), .B1(n9651), 
        .B2(keyinput245), .ZN(n9650) );
  OAI221_X1 U10844 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput142), .C1(n9651), .C2(keyinput245), .A(n9650), .ZN(n9654) );
  AOI22_X1 U10845 ( .A1(n5951), .A2(keyinput147), .B1(n6232), .B2(keyinput254), 
        .ZN(n9652) );
  OAI221_X1 U10846 ( .B1(n5951), .B2(keyinput147), .C1(n6232), .C2(keyinput254), .A(n9652), .ZN(n9653) );
  NOR4_X1 U10847 ( .A1(n9656), .A2(n9655), .A3(n9654), .A4(n9653), .ZN(n9690)
         );
  INV_X1 U10848 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U10849 ( .A1(n10296), .A2(keyinput136), .B1(n9658), .B2(keyinput134), .ZN(n9657) );
  OAI221_X1 U10850 ( .B1(n10296), .B2(keyinput136), .C1(n9658), .C2(
        keyinput134), .A(n9657), .ZN(n9668) );
  INV_X1 U10851 ( .A(SI_1_), .ZN(n9660) );
  INV_X1 U10852 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U10853 ( .A1(n9660), .A2(keyinput144), .B1(keyinput133), .B2(n9944), 
        .ZN(n9659) );
  OAI221_X1 U10854 ( .B1(n9660), .B2(keyinput144), .C1(n9944), .C2(keyinput133), .A(n9659), .ZN(n9667) );
  AOI22_X1 U10855 ( .A1(n5845), .A2(keyinput199), .B1(n9662), .B2(keyinput207), 
        .ZN(n9661) );
  OAI221_X1 U10856 ( .B1(n5845), .B2(keyinput199), .C1(n9662), .C2(keyinput207), .A(n9661), .ZN(n9666) );
  INV_X1 U10857 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9664) );
  AOI22_X1 U10858 ( .A1(n9785), .A2(keyinput159), .B1(n9664), .B2(keyinput153), 
        .ZN(n9663) );
  OAI221_X1 U10859 ( .B1(n9785), .B2(keyinput159), .C1(n9664), .C2(keyinput153), .A(n9663), .ZN(n9665) );
  NOR4_X1 U10860 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n9689)
         );
  INV_X1 U10861 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10295) );
  INV_X1 U10862 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U10863 ( .A1(n10295), .A2(keyinput173), .B1(n10223), .B2(
        keyinput184), .ZN(n9669) );
  OAI221_X1 U10864 ( .B1(n10295), .B2(keyinput173), .C1(n10223), .C2(
        keyinput184), .A(n9669), .ZN(n9677) );
  INV_X1 U10865 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9732) );
  INV_X1 U10866 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U10867 ( .A1(n9732), .A2(keyinput157), .B1(n10253), .B2(keyinput131), .ZN(n9670) );
  OAI221_X1 U10868 ( .B1(n9732), .B2(keyinput157), .C1(n10253), .C2(
        keyinput131), .A(n9670), .ZN(n9676) );
  AOI22_X1 U10869 ( .A1(n9787), .A2(keyinput155), .B1(n6166), .B2(keyinput216), 
        .ZN(n9671) );
  OAI221_X1 U10870 ( .B1(n9787), .B2(keyinput155), .C1(n6166), .C2(keyinput216), .A(n9671), .ZN(n9675) );
  INV_X1 U10871 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U10872 ( .A1(n9673), .A2(keyinput158), .B1(n9735), .B2(keyinput166), 
        .ZN(n9672) );
  OAI221_X1 U10873 ( .B1(n9673), .B2(keyinput158), .C1(n9735), .C2(keyinput166), .A(n9672), .ZN(n9674) );
  NOR4_X1 U10874 ( .A1(n9677), .A2(n9676), .A3(n9675), .A4(n9674), .ZN(n9688)
         );
  INV_X1 U10875 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U10876 ( .A1(n10294), .A2(keyinput129), .B1(keyinput255), .B2(n9889), .ZN(n9678) );
  OAI221_X1 U10877 ( .B1(n10294), .B2(keyinput129), .C1(n9889), .C2(
        keyinput255), .A(n9678), .ZN(n9686) );
  AOI22_X1 U10878 ( .A1(n10229), .A2(keyinput236), .B1(keyinput149), .B2(n9680), .ZN(n9679) );
  OAI221_X1 U10879 ( .B1(n10229), .B2(keyinput236), .C1(n9680), .C2(
        keyinput149), .A(n9679), .ZN(n9685) );
  AOI22_X1 U10880 ( .A1(n5922), .A2(keyinput150), .B1(keyinput241), .B2(n9828), 
        .ZN(n9681) );
  OAI221_X1 U10881 ( .B1(n5922), .B2(keyinput150), .C1(n9828), .C2(keyinput241), .A(n9681), .ZN(n9684) );
  AOI22_X1 U10882 ( .A1(n9013), .A2(keyinput240), .B1(n10304), .B2(keyinput219), .ZN(n9682) );
  OAI221_X1 U10883 ( .B1(n9013), .B2(keyinput240), .C1(n10304), .C2(
        keyinput219), .A(n9682), .ZN(n9683) );
  NOR4_X1 U10884 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n9687)
         );
  NAND4_X1 U10885 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n9877)
         );
  OAI22_X1 U10886 ( .A1(P1_D_REG_15__SCAN_IN), .A2(keyinput35), .B1(keyinput41), .B2(P2_IR_REG_2__SCAN_IN), .ZN(n9691) );
  AOI221_X1 U10887 ( .B1(P1_D_REG_15__SCAN_IN), .B2(keyinput35), .C1(
        P2_IR_REG_2__SCAN_IN), .C2(keyinput41), .A(n9691), .ZN(n9698) );
  OAI22_X1 U10888 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput14), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput34), .ZN(n9692) );
  AOI221_X1 U10889 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput14), .C1(
        keyinput34), .C2(P2_REG3_REG_24__SCAN_IN), .A(n9692), .ZN(n9697) );
  OAI22_X1 U10890 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput6), .B1(
        P2_IR_REG_26__SCAN_IN), .B2(keyinput22), .ZN(n9693) );
  AOI221_X1 U10891 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput6), .C1(
        keyinput22), .C2(P2_IR_REG_26__SCAN_IN), .A(n9693), .ZN(n9696) );
  OAI22_X1 U10892 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput25), .B1(
        P2_IR_REG_5__SCAN_IN), .B2(keyinput76), .ZN(n9694) );
  AOI221_X1 U10893 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput25), .C1(
        keyinput76), .C2(P2_IR_REG_5__SCAN_IN), .A(n9694), .ZN(n9695) );
  NAND4_X1 U10894 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9726)
         );
  OAI22_X1 U10895 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(keyinput70), .B1(
        keyinput28), .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9699) );
  AOI221_X1 U10896 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(keyinput70), .C1(
        P1_DATAO_REG_30__SCAN_IN), .C2(keyinput28), .A(n9699), .ZN(n9706) );
  OAI22_X1 U10897 ( .A1(SI_25_), .A2(keyinput79), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(keyinput73), .ZN(n9700) );
  AOI221_X1 U10898 ( .B1(SI_25_), .B2(keyinput79), .C1(keyinput73), .C2(
        P1_REG3_REG_2__SCAN_IN), .A(n9700), .ZN(n9705) );
  OAI22_X1 U10899 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(keyinput23), .B1(
        keyinput125), .B2(P2_REG1_REG_4__SCAN_IN), .ZN(n9701) );
  AOI221_X1 U10900 ( .B1(P2_IR_REG_10__SCAN_IN), .B2(keyinput23), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput125), .A(n9701), .ZN(n9704) );
  OAI22_X1 U10901 ( .A1(P2_D_REG_18__SCAN_IN), .A2(keyinput0), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput112), .ZN(n9702) );
  AOI221_X1 U10902 ( .B1(P2_D_REG_18__SCAN_IN), .B2(keyinput0), .C1(
        keyinput112), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n9702), .ZN(n9703) );
  NAND4_X1 U10903 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n9725)
         );
  OAI22_X1 U10904 ( .A1(SI_21_), .A2(keyinput49), .B1(P2_D_REG_1__SCAN_IN), 
        .B2(keyinput91), .ZN(n9707) );
  AOI221_X1 U10905 ( .B1(SI_21_), .B2(keyinput49), .C1(keyinput91), .C2(
        P2_D_REG_1__SCAN_IN), .A(n9707), .ZN(n9714) );
  OAI22_X1 U10906 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput68), .B1(
        P2_IR_REG_22__SCAN_IN), .B2(keyinput18), .ZN(n9708) );
  AOI221_X1 U10907 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput68), .C1(
        keyinput18), .C2(P2_IR_REG_22__SCAN_IN), .A(n9708), .ZN(n9713) );
  OAI22_X1 U10908 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput50), .B1(
        P2_REG2_REG_22__SCAN_IN), .B2(keyinput58), .ZN(n9709) );
  AOI221_X1 U10909 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput50), .C1(
        keyinput58), .C2(P2_REG2_REG_22__SCAN_IN), .A(n9709), .ZN(n9712) );
  OAI22_X1 U10910 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput47), .B1(
        keyinput93), .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n9710) );
  AOI221_X1 U10911 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput47), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput93), .A(n9710), .ZN(n9711) );
  NAND4_X1 U10912 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n9724)
         );
  OAI22_X1 U10913 ( .A1(P1_D_REG_27__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG1_REG_2__SCAN_IN), .B2(keyinput9), .ZN(n9715) );
  AOI221_X1 U10914 ( .B1(P1_D_REG_27__SCAN_IN), .B2(keyinput97), .C1(keyinput9), .C2(P1_REG1_REG_2__SCAN_IN), .A(n9715), .ZN(n9722) );
  OAI22_X1 U10915 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(keyinput124), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput12), .ZN(n9716) );
  AOI221_X1 U10916 ( .B1(P1_DATAO_REG_24__SCAN_IN), .B2(keyinput124), .C1(
        keyinput12), .C2(P2_REG3_REG_7__SCAN_IN), .A(n9716), .ZN(n9721) );
  OAI22_X1 U10917 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput72), .B1(keyinput90), .B2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9717) );
  AOI221_X1 U10918 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput72), .C1(
        P2_ADDR_REG_17__SCAN_IN), .C2(keyinput90), .A(n9717), .ZN(n9720) );
  OAI22_X1 U10919 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput108), .B1(
        P2_D_REG_12__SCAN_IN), .B2(keyinput64), .ZN(n9718) );
  AOI221_X1 U10920 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput108), .C1(
        keyinput64), .C2(P2_D_REG_12__SCAN_IN), .A(n9718), .ZN(n9719) );
  NAND4_X1 U10921 ( .A1(n9722), .A2(n9721), .A3(n9720), .A4(n9719), .ZN(n9723)
         );
  NOR4_X1 U10922 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n9838)
         );
  AOI22_X1 U10923 ( .A1(n9204), .A2(keyinput82), .B1(n9728), .B2(keyinput46), 
        .ZN(n9727) );
  OAI221_X1 U10924 ( .B1(n9204), .B2(keyinput82), .C1(n9728), .C2(keyinput46), 
        .A(n9727), .ZN(n9739) );
  INV_X1 U10925 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U10926 ( .A1(n10297), .A2(keyinput114), .B1(keyinput37), .B2(n9730), 
        .ZN(n9729) );
  OAI221_X1 U10927 ( .B1(n10297), .B2(keyinput114), .C1(n9730), .C2(keyinput37), .A(n9729), .ZN(n9738) );
  AOI22_X1 U10928 ( .A1(n9732), .A2(keyinput29), .B1(n10253), .B2(keyinput3), 
        .ZN(n9731) );
  OAI221_X1 U10929 ( .B1(n9732), .B2(keyinput29), .C1(n10253), .C2(keyinput3), 
        .A(n9731), .ZN(n9737) );
  AOI22_X1 U10930 ( .A1(n9735), .A2(keyinput38), .B1(keyinput94), .B2(n9734), 
        .ZN(n9733) );
  OAI221_X1 U10931 ( .B1(n9735), .B2(keyinput38), .C1(n9734), .C2(keyinput94), 
        .A(n9733), .ZN(n9736) );
  NOR4_X1 U10932 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9837)
         );
  AOI22_X1 U10933 ( .A1(n9944), .A2(keyinput5), .B1(n9741), .B2(keyinput107), 
        .ZN(n9740) );
  OAI221_X1 U10934 ( .B1(n9944), .B2(keyinput5), .C1(n9741), .C2(keyinput107), 
        .A(n9740), .ZN(n9746) );
  INV_X1 U10935 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U10936 ( .A1(n10375), .A2(keyinput102), .B1(n9743), .B2(keyinput118), .ZN(n9742) );
  OAI221_X1 U10937 ( .B1(n10375), .B2(keyinput102), .C1(n9743), .C2(
        keyinput118), .A(n9742), .ZN(n9745) );
  XNOR2_X1 U10938 ( .A(n10223), .B(keyinput56), .ZN(n9744) );
  NOR3_X1 U10939 ( .A1(n9746), .A2(n9745), .A3(n9744), .ZN(n9777) );
  AOI22_X1 U10940 ( .A1(n9748), .A2(keyinput11), .B1(keyinput54), .B2(n10209), 
        .ZN(n9747) );
  OAI221_X1 U10941 ( .B1(n9748), .B2(keyinput11), .C1(n10209), .C2(keyinput54), 
        .A(n9747), .ZN(n9751) );
  AOI22_X1 U10942 ( .A1(n10024), .A2(keyinput110), .B1(keyinput1), .B2(n10294), 
        .ZN(n9749) );
  OAI221_X1 U10943 ( .B1(n10024), .B2(keyinput110), .C1(n10294), .C2(keyinput1), .A(n9749), .ZN(n9750) );
  NOR2_X1 U10944 ( .A1(n9751), .A2(n9750), .ZN(n9776) );
  INV_X1 U10945 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U10946 ( .A1(n9754), .A2(keyinput10), .B1(keyinput122), .B2(n9753), 
        .ZN(n9752) );
  OAI221_X1 U10947 ( .B1(n9754), .B2(keyinput10), .C1(n9753), .C2(keyinput122), 
        .A(n9752), .ZN(n9755) );
  INV_X1 U10948 ( .A(n9755), .ZN(n9771) );
  XNOR2_X1 U10949 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput55), .ZN(n9758) );
  XNOR2_X1 U10950 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput83), .ZN(n9757) );
  XNOR2_X1 U10951 ( .A(keyinput13), .B(P2_REG0_REG_3__SCAN_IN), .ZN(n9756) );
  AND3_X1 U10952 ( .A1(n9758), .A2(n9757), .A3(n9756), .ZN(n9770) );
  XNOR2_X1 U10953 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput60), .ZN(n9762) );
  XNOR2_X1 U10954 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput87), .ZN(n9761) );
  XNOR2_X1 U10955 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput57), .ZN(n9760) );
  XNOR2_X1 U10956 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput62), .ZN(n9759) );
  NAND4_X1 U10957 ( .A1(n9762), .A2(n9761), .A3(n9760), .A4(n9759), .ZN(n9768)
         );
  XNOR2_X1 U10958 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput127), .ZN(n9766)
         );
  XNOR2_X1 U10959 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput7), .ZN(n9765) );
  XNOR2_X1 U10960 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput53), .ZN(n9764) );
  XNOR2_X1 U10961 ( .A(keyinput81), .B(P2_REG2_REG_21__SCAN_IN), .ZN(n9763) );
  NAND4_X1 U10962 ( .A1(n9766), .A2(n9765), .A3(n9764), .A4(n9763), .ZN(n9767)
         );
  NOR2_X1 U10963 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  AND3_X1 U10964 ( .A1(n9771), .A2(n9770), .A3(n9769), .ZN(n9775) );
  XNOR2_X1 U10965 ( .A(n10295), .B(keyinput45), .ZN(n9773) );
  XNOR2_X1 U10966 ( .A(n10296), .B(keyinput8), .ZN(n9772) );
  NOR2_X1 U10967 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  NAND4_X1 U10968 ( .A1(n9777), .A2(n9776), .A3(n9775), .A4(n9774), .ZN(n9808)
         );
  AOI22_X1 U10969 ( .A1(n6039), .A2(keyinput39), .B1(keyinput2), .B2(n9779), 
        .ZN(n9778) );
  OAI221_X1 U10970 ( .B1(n6039), .B2(keyinput39), .C1(n9779), .C2(keyinput2), 
        .A(n9778), .ZN(n9783) );
  AOI22_X1 U10971 ( .A1(n9781), .A2(keyinput59), .B1(keyinput103), .B2(n10298), 
        .ZN(n9780) );
  OAI221_X1 U10972 ( .B1(n9781), .B2(keyinput59), .C1(n10298), .C2(keyinput103), .A(n9780), .ZN(n9782) );
  NOR2_X1 U10973 ( .A1(n9783), .A2(n9782), .ZN(n9806) );
  AOI22_X1 U10974 ( .A1(n9785), .A2(keyinput31), .B1(n10030), .B2(keyinput66), 
        .ZN(n9784) );
  OAI221_X1 U10975 ( .B1(n9785), .B2(keyinput31), .C1(n10030), .C2(keyinput66), 
        .A(n9784), .ZN(n9789) );
  AOI22_X1 U10976 ( .A1(n9787), .A2(keyinput27), .B1(n10233), .B2(keyinput69), 
        .ZN(n9786) );
  OAI221_X1 U10977 ( .B1(n9787), .B2(keyinput27), .C1(n10233), .C2(keyinput69), 
        .A(n9786), .ZN(n9788) );
  NOR2_X1 U10978 ( .A1(n9789), .A2(n9788), .ZN(n9805) );
  AOI22_X1 U10979 ( .A1(n9791), .A2(keyinput26), .B1(n5845), .B2(keyinput71), 
        .ZN(n9790) );
  OAI221_X1 U10980 ( .B1(n9791), .B2(keyinput26), .C1(n5845), .C2(keyinput71), 
        .A(n9790), .ZN(n9795) );
  AOI22_X1 U10981 ( .A1(n9793), .A2(keyinput32), .B1(keyinput105), .B2(n6179), 
        .ZN(n9792) );
  OAI221_X1 U10982 ( .B1(n9793), .B2(keyinput32), .C1(n6179), .C2(keyinput105), 
        .A(n9792), .ZN(n9794) );
  NOR2_X1 U10983 ( .A1(n9795), .A2(n9794), .ZN(n9804) );
  INV_X1 U10984 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10985 ( .A1(n9798), .A2(keyinput48), .B1(keyinput115), .B2(n9797), 
        .ZN(n9796) );
  OAI221_X1 U10986 ( .B1(n9798), .B2(keyinput48), .C1(n9797), .C2(keyinput115), 
        .A(n9796), .ZN(n9802) );
  AOI22_X1 U10987 ( .A1(n10410), .A2(keyinput75), .B1(n9800), .B2(keyinput63), 
        .ZN(n9799) );
  OAI221_X1 U10988 ( .B1(n10410), .B2(keyinput75), .C1(n9800), .C2(keyinput63), 
        .A(n9799), .ZN(n9801) );
  NOR2_X1 U10989 ( .A1(n9802), .A2(n9801), .ZN(n9803) );
  NAND4_X1 U10990 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n9807)
         );
  NOR2_X1 U10991 ( .A1(n9808), .A2(n9807), .ZN(n9836) );
  AOI22_X1 U10992 ( .A1(n9811), .A2(keyinput67), .B1(keyinput85), .B2(n9810), 
        .ZN(n9809) );
  OAI221_X1 U10993 ( .B1(n9811), .B2(keyinput67), .C1(n9810), .C2(keyinput85), 
        .A(n9809), .ZN(n9822) );
  AOI22_X1 U10994 ( .A1(n5110), .A2(keyinput100), .B1(keyinput24), .B2(n9813), 
        .ZN(n9812) );
  OAI221_X1 U10995 ( .B1(n5110), .B2(keyinput100), .C1(n9813), .C2(keyinput24), 
        .A(n9812), .ZN(n9821) );
  AOI22_X1 U10996 ( .A1(n9816), .A2(keyinput116), .B1(keyinput44), .B2(n9815), 
        .ZN(n9814) );
  OAI221_X1 U10997 ( .B1(n9816), .B2(keyinput116), .C1(n9815), .C2(keyinput44), 
        .A(n9814), .ZN(n9820) );
  AOI22_X1 U10998 ( .A1(n9818), .A2(keyinput17), .B1(n6901), .B2(keyinput89), 
        .ZN(n9817) );
  OAI221_X1 U10999 ( .B1(n9818), .B2(keyinput17), .C1(n6901), .C2(keyinput89), 
        .A(n9817), .ZN(n9819) );
  NOR4_X1 U11000 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(n9834)
         );
  INV_X1 U11001 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U11002 ( .A1(n10226), .A2(keyinput101), .B1(keyinput109), .B2(n9824), .ZN(n9823) );
  OAI221_X1 U11003 ( .B1(n10226), .B2(keyinput101), .C1(n9824), .C2(
        keyinput109), .A(n9823), .ZN(n9832) );
  INV_X1 U11004 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10227) );
  INV_X1 U11005 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U11006 ( .A1(n10227), .A2(keyinput43), .B1(keyinput36), .B2(n10318), 
        .ZN(n9825) );
  OAI221_X1 U11007 ( .B1(n10227), .B2(keyinput43), .C1(n10318), .C2(keyinput36), .A(n9825), .ZN(n9831) );
  AOI22_X1 U11008 ( .A1(n7067), .A2(keyinput111), .B1(n7795), .B2(keyinput65), 
        .ZN(n9826) );
  OAI221_X1 U11009 ( .B1(n7067), .B2(keyinput111), .C1(n7795), .C2(keyinput65), 
        .A(n9826), .ZN(n9830) );
  AOI22_X1 U11010 ( .A1(n9828), .A2(keyinput113), .B1(n6309), .B2(keyinput40), 
        .ZN(n9827) );
  OAI221_X1 U11011 ( .B1(n9828), .B2(keyinput113), .C1(n6309), .C2(keyinput40), 
        .A(n9827), .ZN(n9829) );
  NOR4_X1 U11012 ( .A1(n9832), .A2(n9831), .A3(n9830), .A4(n9829), .ZN(n9833)
         );
  AND2_X1 U11013 ( .A1(n9834), .A2(n9833), .ZN(n9835) );
  AND4_X1 U11014 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n9876)
         );
  OAI22_X1 U11015 ( .A1(SI_1_), .A2(keyinput16), .B1(keyinput77), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n9839) );
  AOI221_X1 U11016 ( .B1(SI_1_), .B2(keyinput16), .C1(P2_REG0_REG_29__SCAN_IN), 
        .C2(keyinput77), .A(n9839), .ZN(n9846) );
  OAI22_X1 U11017 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(keyinput88), .B1(
        keyinput42), .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9840) );
  AOI221_X1 U11018 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(keyinput88), .C1(
        P2_DATAO_REG_30__SCAN_IN), .C2(keyinput42), .A(n9840), .ZN(n9845) );
  OAI22_X1 U11019 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput20), .B1(
        keyinput84), .B2(P1_REG2_REG_28__SCAN_IN), .ZN(n9841) );
  AOI221_X1 U11020 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput20), .C1(
        P1_REG2_REG_28__SCAN_IN), .C2(keyinput84), .A(n9841), .ZN(n9844) );
  OAI22_X1 U11021 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput106), .B1(
        keyinput117), .B2(P2_REG1_REG_15__SCAN_IN), .ZN(n9842) );
  AOI221_X1 U11022 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput106), .C1(
        P2_REG1_REG_15__SCAN_IN), .C2(keyinput117), .A(n9842), .ZN(n9843) );
  NAND4_X1 U11023 ( .A1(n9846), .A2(n9845), .A3(n9844), .A4(n9843), .ZN(n9874)
         );
  OAI22_X1 U11024 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(keyinput80), .B1(
        keyinput30), .B2(P1_REG2_REG_31__SCAN_IN), .ZN(n9847) );
  AOI221_X1 U11025 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(keyinput80), .C1(
        P1_REG2_REG_31__SCAN_IN), .C2(keyinput30), .A(n9847), .ZN(n9854) );
  OAI22_X1 U11026 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput95), .B1(
        P2_D_REG_19__SCAN_IN), .B2(keyinput4), .ZN(n9848) );
  AOI221_X1 U11027 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput95), .C1(
        keyinput4), .C2(P2_D_REG_19__SCAN_IN), .A(n9848), .ZN(n9853) );
  OAI22_X1 U11028 ( .A1(SI_23_), .A2(keyinput51), .B1(keyinput104), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9849) );
  AOI221_X1 U11029 ( .B1(SI_23_), .B2(keyinput51), .C1(P1_REG3_REG_0__SCAN_IN), 
        .C2(keyinput104), .A(n9849), .ZN(n9852) );
  OAI22_X1 U11030 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(keyinput98), .B1(keyinput92), .B2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9850) );
  AOI221_X1 U11031 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(keyinput98), .C1(
        P2_ADDR_REG_6__SCAN_IN), .C2(keyinput92), .A(n9850), .ZN(n9851) );
  NAND4_X1 U11032 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n9851), .ZN(n9873)
         );
  OAI22_X1 U11033 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput123), .B1(
        keyinput19), .B2(P2_REG0_REG_2__SCAN_IN), .ZN(n9855) );
  AOI221_X1 U11034 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput123), .C1(
        P2_REG0_REG_2__SCAN_IN), .C2(keyinput19), .A(n9855), .ZN(n9862) );
  OAI22_X1 U11035 ( .A1(P1_D_REG_12__SCAN_IN), .A2(keyinput119), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput78), .ZN(n9856) );
  AOI221_X1 U11036 ( .B1(P1_D_REG_12__SCAN_IN), .B2(keyinput119), .C1(
        keyinput78), .C2(P1_D_REG_23__SCAN_IN), .A(n9856), .ZN(n9861) );
  OAI22_X1 U11037 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput74), .B1(
        keyinput15), .B2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9857) );
  AOI221_X1 U11038 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput74), .C1(
        P1_ADDR_REG_13__SCAN_IN), .C2(keyinput15), .A(n9857), .ZN(n9860) );
  OAI22_X1 U11039 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput99), .B1(
        keyinput61), .B2(P2_REG1_REG_13__SCAN_IN), .ZN(n9858) );
  AOI221_X1 U11040 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput99), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput61), .A(n9858), .ZN(n9859) );
  NAND4_X1 U11041 ( .A1(n9862), .A2(n9861), .A3(n9860), .A4(n9859), .ZN(n9872)
         );
  OAI22_X1 U11042 ( .A1(SI_24_), .A2(keyinput121), .B1(keyinput21), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n9863) );
  AOI221_X1 U11043 ( .B1(SI_24_), .B2(keyinput121), .C1(
        P2_REG1_REG_14__SCAN_IN), .C2(keyinput21), .A(n9863), .ZN(n9870) );
  OAI22_X1 U11044 ( .A1(P1_D_REG_28__SCAN_IN), .A2(keyinput120), .B1(
        P2_REG0_REG_8__SCAN_IN), .B2(keyinput96), .ZN(n9864) );
  AOI221_X1 U11045 ( .B1(P1_D_REG_28__SCAN_IN), .B2(keyinput120), .C1(
        keyinput96), .C2(P2_REG0_REG_8__SCAN_IN), .A(n9864), .ZN(n9869) );
  OAI22_X1 U11046 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput52), .B1(keyinput33), .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9865) );
  AOI221_X1 U11047 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput52), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput33), .A(n9865), .ZN(n9868) );
  OAI22_X1 U11048 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput126), .B1(
        P2_ADDR_REG_11__SCAN_IN), .B2(keyinput86), .ZN(n9866) );
  AOI221_X1 U11049 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput126), .C1(
        keyinput86), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n9866), .ZN(n9867) );
  NAND4_X1 U11050 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n9871)
         );
  NOR4_X1 U11051 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n9875)
         );
  OAI211_X1 U11052 ( .C1(n9878), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9879)
         );
  XNOR2_X1 U11053 ( .A(n9880), .B(n9879), .ZN(P1_U3505) );
  MUX2_X1 U11054 ( .A(P1_D_REG_0__SCAN_IN), .B(n9881), .S(n10234), .Z(P1_U3440) );
  NOR4_X1 U11055 ( .A1(n9882), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5390), .A4(
        P1_U3084), .ZN(n9883) );
  AOI21_X1 U11056 ( .B1(n9892), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9883), .ZN(
        n9884) );
  OAI21_X1 U11057 ( .B1(n9885), .B2(n4459), .A(n9884), .ZN(P1_U3322) );
  OAI222_X1 U11058 ( .A1(n9890), .A2(n9889), .B1(P1_U3084), .B2(n9887), .C1(
        n4459), .C2(n9886), .ZN(P1_U3324) );
  AOI21_X1 U11059 ( .B1(n9892), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9891), .ZN(
        n9893) );
  OAI21_X1 U11060 ( .B1(n9894), .B2(n4459), .A(n9893), .ZN(P1_U3325) );
  AOI22_X1 U11061 ( .A1(n10101), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(n10184), 
        .B2(n9895), .ZN(n9906) );
  AOI21_X1 U11062 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9899) );
  NAND2_X1 U11063 ( .A1(n10106), .A2(n9899), .ZN(n9904) );
  OAI211_X1 U11064 ( .C1(n9902), .C2(n9901), .A(n10172), .B(n9900), .ZN(n9903)
         );
  NAND4_X1 U11065 ( .A1(n9906), .A2(n9905), .A3(n9904), .A4(n9903), .ZN(
        P1_U3244) );
  INV_X1 U11066 ( .A(n9907), .ZN(n9911) );
  NAND2_X1 U11067 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9908) );
  NAND2_X1 U11068 ( .A1(n9909), .A2(n9908), .ZN(n9910) );
  NAND3_X1 U11069 ( .A1(n10282), .A2(n9911), .A3(n9910), .ZN(n9916) );
  INV_X1 U11070 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9951) );
  OAI22_X1 U11071 ( .A1(n9913), .A2(n9951), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9912), .ZN(n9914) );
  INV_X1 U11072 ( .A(n9914), .ZN(n9915) );
  OAI211_X1 U11073 ( .C1(n10283), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9918)
         );
  INV_X1 U11074 ( .A(n9918), .ZN(n9923) );
  NOR2_X1 U11075 ( .A1(n10290), .A2(n10359), .ZN(n9921) );
  OAI211_X1 U11076 ( .C1(n9921), .C2(n9920), .A(n10281), .B(n9919), .ZN(n9922)
         );
  NAND2_X1 U11077 ( .A1(n9923), .A2(n9922), .ZN(P2_U3246) );
  AOI22_X1 U11078 ( .A1(n10287), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9936) );
  AOI211_X1 U11079 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9928)
         );
  AOI21_X1 U11080 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n9935) );
  OAI211_X1 U11081 ( .C1(n9933), .C2(n9932), .A(n10281), .B(n9931), .ZN(n9934)
         );
  NAND3_X1 U11082 ( .A1(n9936), .A2(n9935), .A3(n9934), .ZN(P2_U3247) );
  INV_X1 U11083 ( .A(n9937), .ZN(n10270) );
  OAI21_X1 U11084 ( .B1(n9939), .B2(n10263), .A(n9938), .ZN(n9940) );
  AOI21_X1 U11085 ( .B1(n9941), .B2(n10270), .A(n9940), .ZN(n9942) );
  AND2_X1 U11086 ( .A1(n9943), .A2(n9942), .ZN(n9945) );
  AOI22_X1 U11087 ( .A1(n10273), .A2(n9945), .B1(n9944), .B2(n10271), .ZN(
        P1_U3484) );
  AOI22_X1 U11088 ( .A1(n4456), .A2(n9945), .B1(n6658), .B2(n10279), .ZN(
        P1_U3533) );
  INV_X1 U11089 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U11090 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9946) );
  AOI21_X1 U11091 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9946), .ZN(n10378) );
  NOR2_X1 U11092 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9947) );
  AOI21_X1 U11093 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9947), .ZN(n10381) );
  NOR2_X1 U11094 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9948) );
  AOI21_X1 U11095 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9948), .ZN(n10384) );
  NOR2_X1 U11096 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9949) );
  AOI21_X1 U11097 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9949), .ZN(n10387) );
  NOR2_X1 U11098 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n9950) );
  AOI21_X1 U11099 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9950), .ZN(n10390) );
  NOR2_X1 U11100 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9957) );
  XNOR2_X1 U11101 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10418) );
  NAND2_X1 U11102 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9955) );
  XOR2_X1 U11103 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10416) );
  NAND2_X1 U11104 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9953) );
  XOR2_X1 U11105 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10414) );
  AOI21_X1 U11106 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10371) );
  NAND3_X1 U11107 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10373) );
  OAI21_X1 U11108 ( .B1(n10371), .B2(n9951), .A(n10373), .ZN(n10413) );
  NAND2_X1 U11109 ( .A1(n10414), .A2(n10413), .ZN(n9952) );
  NAND2_X1 U11110 ( .A1(n9953), .A2(n9952), .ZN(n10415) );
  NAND2_X1 U11111 ( .A1(n10416), .A2(n10415), .ZN(n9954) );
  NAND2_X1 U11112 ( .A1(n9955), .A2(n9954), .ZN(n10417) );
  NOR2_X1 U11113 ( .A1(n10418), .A2(n10417), .ZN(n9956) );
  NOR2_X1 U11114 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  NOR2_X1 U11115 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9958), .ZN(n10402) );
  AND2_X1 U11116 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9958), .ZN(n10401) );
  NOR2_X1 U11117 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10401), .ZN(n9959) );
  NOR2_X1 U11118 ( .A1(n10402), .A2(n9959), .ZN(n9960) );
  NAND2_X1 U11119 ( .A1(n9960), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9962) );
  XOR2_X1 U11120 ( .A(n9960), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10400) );
  NAND2_X1 U11121 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10400), .ZN(n9961) );
  NAND2_X1 U11122 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  NAND2_X1 U11123 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9963), .ZN(n9965) );
  XOR2_X1 U11124 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9963), .Z(n10412) );
  NAND2_X1 U11125 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10412), .ZN(n9964) );
  NAND2_X1 U11126 ( .A1(n9965), .A2(n9964), .ZN(n9966) );
  NAND2_X1 U11127 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9966), .ZN(n9968) );
  XOR2_X1 U11128 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9966), .Z(n10411) );
  NAND2_X1 U11129 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10411), .ZN(n9967) );
  NAND2_X1 U11130 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  AND2_X1 U11131 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9969), .ZN(n9970) );
  XNOR2_X1 U11132 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9969), .ZN(n10409) );
  NOR2_X1 U11133 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  NAND2_X1 U11134 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9971) );
  OAI21_X1 U11135 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9971), .ZN(n10398) );
  NAND2_X1 U11136 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9972) );
  OAI21_X1 U11137 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9972), .ZN(n10395) );
  NOR2_X1 U11138 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9973) );
  AOI21_X1 U11139 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9973), .ZN(n10392) );
  NAND2_X1 U11140 ( .A1(n10393), .A2(n10392), .ZN(n10391) );
  NAND2_X1 U11141 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  NAND2_X1 U11142 ( .A1(n10387), .A2(n10386), .ZN(n10385) );
  OAI21_X1 U11143 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10385), .ZN(n10383) );
  NAND2_X1 U11144 ( .A1(n10384), .A2(n10383), .ZN(n10382) );
  OAI21_X1 U11145 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10382), .ZN(n10380) );
  NAND2_X1 U11146 ( .A1(n10381), .A2(n10380), .ZN(n10379) );
  OAI21_X1 U11147 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10379), .ZN(n10377) );
  NAND2_X1 U11148 ( .A1(n10378), .A2(n10377), .ZN(n10376) );
  NOR2_X1 U11149 ( .A1(n10406), .A2(n10405), .ZN(n9974) );
  NAND2_X1 U11150 ( .A1(n10406), .A2(n10405), .ZN(n10404) );
  OAI21_X1 U11151 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9974), .A(n10404), .ZN(
        n9976) );
  XOR2_X1 U11152 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9975) );
  XNOR2_X1 U11153 ( .A(n9976), .B(n9975), .ZN(ADD_1071_U4) );
  NOR2_X1 U11154 ( .A1(n9977), .A2(n10350), .ZN(n9978) );
  AOI22_X1 U11155 ( .A1(n10370), .A2(n9982), .B1(n6281), .B2(n10368), .ZN(
        P2_U3550) );
  INV_X1 U11156 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11157 ( .A1(n10358), .A2(n9982), .B1(n9981), .B2(n10356), .ZN(
        P2_U3518) );
  XNOR2_X1 U11158 ( .A(n9984), .B(n9983), .ZN(n9986) );
  NAND2_X1 U11159 ( .A1(n9986), .A2(n9985), .ZN(n9992) );
  AOI22_X1 U11160 ( .A1(n9990), .A2(n9989), .B1(n9988), .B2(n9987), .ZN(n9991)
         );
  AOI222_X1 U11161 ( .A1(n10009), .A2(n10213), .B1(n9994), .B2(n9993), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(n10216), .ZN(n10007) );
  OAI21_X1 U11162 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n10008) );
  NAND2_X1 U11163 ( .A1(n9998), .A2(n10009), .ZN(n10000) );
  NAND2_X1 U11164 ( .A1(n10000), .A2(n9999), .ZN(n10001) );
  OR2_X1 U11165 ( .A1(n10002), .A2(n10001), .ZN(n10010) );
  OAI22_X1 U11166 ( .A1(n10008), .A2(n10004), .B1(n10010), .B2(n10003), .ZN(
        n10005) );
  INV_X1 U11167 ( .A(n10005), .ZN(n10006) );
  OAI211_X1 U11168 ( .C1(n10216), .C2(n10011), .A(n10007), .B(n10006), .ZN(
        P1_U3275) );
  INV_X1 U11169 ( .A(n10008), .ZN(n10014) );
  INV_X1 U11170 ( .A(n10009), .ZN(n10012) );
  OAI211_X1 U11171 ( .C1(n10012), .C2(n10263), .A(n10011), .B(n10010), .ZN(
        n10013) );
  AOI21_X1 U11172 ( .B1(n10014), .B2(n10252), .A(n10013), .ZN(n10044) );
  AOI22_X1 U11173 ( .A1(n4456), .A2(n10044), .B1(n10015), .B2(n10279), .ZN(
        P1_U3539) );
  NOR2_X1 U11174 ( .A1(n10017), .A2(n10016), .ZN(n10023) );
  OAI211_X1 U11175 ( .C1(n10020), .C2(n10263), .A(n10019), .B(n10018), .ZN(
        n10021) );
  AOI21_X1 U11176 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10046) );
  AOI22_X1 U11177 ( .A1(n4456), .A2(n10046), .B1(n10024), .B2(n10279), .ZN(
        P1_U3538) );
  OAI211_X1 U11178 ( .C1(n10027), .C2(n10263), .A(n10026), .B(n10025), .ZN(
        n10028) );
  AOI21_X1 U11179 ( .B1(n10252), .B2(n10029), .A(n10028), .ZN(n10048) );
  AOI22_X1 U11180 ( .A1(n4456), .A2(n10048), .B1(n10030), .B2(n10279), .ZN(
        P1_U3537) );
  OAI22_X1 U11181 ( .A1(n10032), .A2(n10265), .B1(n10031), .B2(n10263), .ZN(
        n10033) );
  AOI21_X1 U11182 ( .B1(n10034), .B2(n10270), .A(n10033), .ZN(n10035) );
  AND2_X1 U11183 ( .A1(n10036), .A2(n10035), .ZN(n10050) );
  AOI22_X1 U11184 ( .A1(n4456), .A2(n10050), .B1(n9204), .B2(n10279), .ZN(
        P1_U3536) );
  OAI22_X1 U11185 ( .A1(n10038), .A2(n10265), .B1(n10037), .B2(n10263), .ZN(
        n10040) );
  AOI211_X1 U11186 ( .C1(n10041), .C2(n10252), .A(n10040), .B(n10039), .ZN(
        n10052) );
  AOI22_X1 U11187 ( .A1(n4456), .A2(n10052), .B1(n10042), .B2(n10279), .ZN(
        P1_U3534) );
  INV_X1 U11188 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U11189 ( .A1(n10273), .A2(n10044), .B1(n10043), .B2(n10271), .ZN(
        P1_U3502) );
  INV_X1 U11190 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10045) );
  AOI22_X1 U11191 ( .A1(n10273), .A2(n10046), .B1(n10045), .B2(n10271), .ZN(
        P1_U3499) );
  INV_X1 U11192 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11193 ( .A1(n10273), .A2(n10048), .B1(n10047), .B2(n10271), .ZN(
        P1_U3496) );
  INV_X1 U11194 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U11195 ( .A1(n10273), .A2(n10050), .B1(n10049), .B2(n10271), .ZN(
        P1_U3493) );
  INV_X1 U11196 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11197 ( .A1(n10273), .A2(n10052), .B1(n10051), .B2(n10271), .ZN(
        P1_U3487) );
  XNOR2_X1 U11198 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11199 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U11200 ( .C1(n10076), .C2(n10054), .A(n10053), .B(n10178), .ZN(
        n10055) );
  AOI21_X1 U11201 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n10055), 
        .ZN(n10064) );
  AOI22_X1 U11202 ( .A1(n10101), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n10184), 
        .B2(n10056), .ZN(n10063) );
  NOR2_X1 U11203 ( .A1(n10058), .A2(n10057), .ZN(n10061) );
  OAI211_X1 U11204 ( .C1(n10061), .C2(n10060), .A(n10172), .B(n10059), .ZN(
        n10062) );
  NAND3_X1 U11205 ( .A1(n10064), .A2(n10063), .A3(n10062), .ZN(P1_U3242) );
  INV_X1 U11206 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10085) );
  AOI21_X1 U11207 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10083) );
  NAND2_X1 U11208 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10072) );
  OAI211_X1 U11209 ( .C1(n10070), .C2(n10069), .A(n10172), .B(n10068), .ZN(
        n10071) );
  OAI211_X1 U11210 ( .C1(n10074), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10082) );
  MUX2_X1 U11211 ( .A(n10077), .B(n10076), .S(n10075), .Z(n10080) );
  OAI211_X1 U11212 ( .C1(n10080), .C2(n5886), .A(n10079), .B(n10078), .ZN(
        n10097) );
  INV_X1 U11213 ( .A(n10097), .ZN(n10081) );
  AOI211_X1 U11214 ( .C1(n10106), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10084) );
  OAI21_X1 U11215 ( .B1(n10193), .B2(n10085), .A(n10084), .ZN(P1_U3243) );
  INV_X1 U11216 ( .A(n10086), .ZN(n10090) );
  XNOR2_X1 U11217 ( .A(n10088), .B(n10087), .ZN(n10089) );
  AOI22_X1 U11218 ( .A1(n10090), .A2(n10184), .B1(n10106), .B2(n10089), .ZN(
        n10099) );
  AOI21_X1 U11219 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10094) );
  NOR2_X1 U11220 ( .A1(n10190), .A2(n10094), .ZN(n10095) );
  AOI211_X1 U11221 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n10101), .A(n10096), .B(
        n10095), .ZN(n10098) );
  NAND3_X1 U11222 ( .A1(n10099), .A2(n10098), .A3(n10097), .ZN(P1_U3245) );
  AOI22_X1 U11223 ( .A1(n10101), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n10184), 
        .B2(n10100), .ZN(n10114) );
  INV_X1 U11224 ( .A(n10102), .ZN(n10113) );
  OAI21_X1 U11225 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10107) );
  NAND2_X1 U11226 ( .A1(n10107), .A2(n10106), .ZN(n10112) );
  OAI211_X1 U11227 ( .C1(n10110), .C2(n10109), .A(n10172), .B(n10108), .ZN(
        n10111) );
  NAND4_X1 U11228 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        P1_U3249) );
  INV_X1 U11229 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10127) );
  AOI211_X1 U11230 ( .C1(n10117), .C2(n10116), .A(n10115), .B(n10178), .ZN(
        n10118) );
  AOI211_X1 U11231 ( .C1(n10184), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10126) );
  AOI21_X1 U11232 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10124) );
  OR2_X1 U11233 ( .A1(n10190), .A2(n10124), .ZN(n10125) );
  OAI211_X1 U11234 ( .C1(n10193), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        P1_U3254) );
  INV_X1 U11235 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10139) );
  AOI211_X1 U11236 ( .C1(n10129), .C2(n7840), .A(n10128), .B(n10178), .ZN(
        n10130) );
  AOI211_X1 U11237 ( .C1(n10184), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10138) );
  AOI21_X1 U11238 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10136) );
  OR2_X1 U11239 ( .A1(n10190), .A2(n10136), .ZN(n10137) );
  OAI211_X1 U11240 ( .C1(n10139), .C2(n10193), .A(n10138), .B(n10137), .ZN(
        P1_U3255) );
  INV_X1 U11241 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10151) );
  INV_X1 U11242 ( .A(n10140), .ZN(n10145) );
  AOI211_X1 U11243 ( .C1(n10143), .C2(n10142), .A(n10141), .B(n10178), .ZN(
        n10144) );
  AOI211_X1 U11244 ( .C1(n10184), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10150) );
  OAI211_X1 U11245 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10148), .A(n10172), 
        .B(n10147), .ZN(n10149) );
  OAI211_X1 U11246 ( .C1(n10151), .C2(n10193), .A(n10150), .B(n10149), .ZN(
        P1_U3256) );
  INV_X1 U11247 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10163) );
  AOI211_X1 U11248 ( .C1(n10154), .C2(n10153), .A(n10152), .B(n10178), .ZN(
        n10155) );
  AOI211_X1 U11249 ( .C1(n10184), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10162) );
  OAI211_X1 U11250 ( .C1(n10160), .C2(n10159), .A(n10172), .B(n10158), .ZN(
        n10161) );
  OAI211_X1 U11251 ( .C1(n10163), .C2(n10193), .A(n10162), .B(n10161), .ZN(
        P1_U3257) );
  INV_X1 U11252 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10177) );
  INV_X1 U11253 ( .A(n10164), .ZN(n10169) );
  AOI211_X1 U11254 ( .C1(n10167), .C2(n10166), .A(n10165), .B(n10178), .ZN(
        n10168) );
  AOI211_X1 U11255 ( .C1(n10184), .C2(n10170), .A(n10169), .B(n10168), .ZN(
        n10176) );
  OAI211_X1 U11256 ( .C1(n10174), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10175) );
  OAI211_X1 U11257 ( .C1(n10177), .C2(n10193), .A(n10176), .B(n10175), .ZN(
        P1_U3258) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10194) );
  AOI211_X1 U11259 ( .C1(n10181), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10182) );
  AOI211_X1 U11260 ( .C1(n10185), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        n10192) );
  AOI21_X1 U11261 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(n10189) );
  OR2_X1 U11262 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  OAI211_X1 U11263 ( .C1(n10194), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        P1_U3259) );
  INV_X1 U11264 ( .A(n10195), .ZN(n10205) );
  OAI22_X1 U11265 ( .A1(n10221), .A2(n10198), .B1(n10197), .B2(n10196), .ZN(
        n10199) );
  AOI21_X1 U11266 ( .B1(n10201), .B2(n10200), .A(n10199), .ZN(n10202) );
  OAI211_X1 U11267 ( .C1(n10205), .C2(n10204), .A(n10203), .B(n10202), .ZN(
        n10206) );
  INV_X1 U11268 ( .A(n10206), .ZN(n10208) );
  AOI22_X1 U11269 ( .A1(n10216), .A2(n10209), .B1(n10208), .B2(n10207), .ZN(
        P1_U3286) );
  INV_X1 U11270 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10210) );
  OR2_X1 U11271 ( .A1(n10207), .A2(n10210), .ZN(n10215) );
  OAI21_X1 U11272 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n10214) );
  OAI211_X1 U11273 ( .C1(n10217), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n10218) );
  INV_X1 U11274 ( .A(n10218), .ZN(n10219) );
  OAI21_X1 U11275 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(P1_U3291) );
  AND2_X1 U11276 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10231), .ZN(P1_U3292) );
  AND2_X1 U11277 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10231), .ZN(P1_U3293) );
  NOR2_X1 U11278 ( .A1(n10230), .A2(n10223), .ZN(P1_U3294) );
  NOR2_X1 U11279 ( .A1(n10230), .A2(n10224), .ZN(P1_U3295) );
  NOR2_X1 U11280 ( .A1(n10230), .A2(n10225), .ZN(P1_U3296) );
  AND2_X1 U11281 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10231), .ZN(P1_U3297) );
  AND2_X1 U11282 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10231), .ZN(P1_U3298) );
  NOR2_X1 U11283 ( .A1(n10230), .A2(n10226), .ZN(P1_U3299) );
  AND2_X1 U11284 ( .A1(n10231), .A2(P1_D_REG_23__SCAN_IN), .ZN(P1_U3300) );
  AND2_X1 U11285 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10231), .ZN(P1_U3301) );
  AND2_X1 U11286 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10231), .ZN(P1_U3302) );
  AND2_X1 U11287 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10231), .ZN(P1_U3303) );
  AND2_X1 U11288 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10231), .ZN(P1_U3304) );
  AND2_X1 U11289 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10231), .ZN(P1_U3305) );
  AND2_X1 U11290 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10231), .ZN(P1_U3306) );
  NOR2_X1 U11291 ( .A1(n10230), .A2(n10227), .ZN(P1_U3307) );
  NOR2_X1 U11292 ( .A1(n10230), .A2(n10228), .ZN(P1_U3308) );
  AND2_X1 U11293 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10231), .ZN(P1_U3309) );
  AND2_X1 U11294 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10231), .ZN(P1_U3310) );
  AND2_X1 U11295 ( .A1(n10231), .A2(P1_D_REG_12__SCAN_IN), .ZN(P1_U3311) );
  AND2_X1 U11296 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10231), .ZN(P1_U3312) );
  NOR2_X1 U11297 ( .A1(n10230), .A2(n10229), .ZN(P1_U3313) );
  AND2_X1 U11298 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10231), .ZN(P1_U3314) );
  AND2_X1 U11299 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10231), .ZN(P1_U3315) );
  AND2_X1 U11300 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10231), .ZN(P1_U3316) );
  AND2_X1 U11301 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10231), .ZN(P1_U3317) );
  AND2_X1 U11302 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10231), .ZN(P1_U3318) );
  AND2_X1 U11303 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10231), .ZN(P1_U3319) );
  AND2_X1 U11304 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10231), .ZN(P1_U3320) );
  AND2_X1 U11305 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10231), .ZN(P1_U3321) );
  OAI21_X1 U11306 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(P1_U3441) );
  OAI22_X1 U11307 ( .A1(n10236), .A2(n10265), .B1(n10235), .B2(n10263), .ZN(
        n10238) );
  AOI211_X1 U11308 ( .C1(n10270), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10275) );
  INV_X1 U11309 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11310 ( .A1(n10273), .A2(n10275), .B1(n10240), .B2(n10271), .ZN(
        P1_U3460) );
  OAI22_X1 U11311 ( .A1(n10242), .A2(n10265), .B1(n10241), .B2(n10263), .ZN(
        n10244) );
  AOI211_X1 U11312 ( .C1(n10270), .C2(n10245), .A(n10244), .B(n10243), .ZN(
        n10276) );
  INV_X1 U11313 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U11314 ( .A1(n10273), .A2(n10276), .B1(n10246), .B2(n10271), .ZN(
        P1_U3466) );
  OAI22_X1 U11315 ( .A1(n10248), .A2(n10265), .B1(n10247), .B2(n10263), .ZN(
        n10250) );
  AOI211_X1 U11316 ( .C1(n10252), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        n10277) );
  AOI22_X1 U11317 ( .A1(n10273), .A2(n10277), .B1(n10253), .B2(n10271), .ZN(
        P1_U3472) );
  INV_X1 U11318 ( .A(n10254), .ZN(n10259) );
  OAI21_X1 U11319 ( .B1(n10256), .B2(n10263), .A(n10255), .ZN(n10258) );
  AOI211_X1 U11320 ( .C1(n10270), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        n10278) );
  INV_X1 U11321 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U11322 ( .A1(n10273), .A2(n10278), .B1(n10260), .B2(n10271), .ZN(
        P1_U3478) );
  INV_X1 U11323 ( .A(n10261), .ZN(n10269) );
  INV_X1 U11324 ( .A(n10262), .ZN(n10264) );
  OAI22_X1 U11325 ( .A1(n10266), .A2(n10265), .B1(n10264), .B2(n10263), .ZN(
        n10268) );
  AOI211_X1 U11326 ( .C1(n10270), .C2(n10269), .A(n10268), .B(n10267), .ZN(
        n10280) );
  INV_X1 U11327 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U11328 ( .A1(n10273), .A2(n10280), .B1(n10272), .B2(n10271), .ZN(
        P1_U3481) );
  AOI22_X1 U11329 ( .A1(n4456), .A2(n10275), .B1(n10274), .B2(n10279), .ZN(
        P1_U3525) );
  AOI22_X1 U11330 ( .A1(n4456), .A2(n10276), .B1(n6535), .B2(n10279), .ZN(
        P1_U3527) );
  AOI22_X1 U11331 ( .A1(n4456), .A2(n10277), .B1(n6537), .B2(n10279), .ZN(
        P1_U3529) );
  AOI22_X1 U11332 ( .A1(n4456), .A2(n10278), .B1(n6528), .B2(n10279), .ZN(
        P1_U3531) );
  AOI22_X1 U11333 ( .A1(n4456), .A2(n10280), .B1(n6541), .B2(n10279), .ZN(
        P1_U3532) );
  AOI22_X1 U11334 ( .A1(n10282), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10281), .ZN(n10291) );
  NAND2_X1 U11335 ( .A1(n10282), .A2(n5939), .ZN(n10284) );
  OAI211_X1 U11336 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10285), .A(n10284), .B(
        n10283), .ZN(n10286) );
  INV_X1 U11337 ( .A(n10286), .ZN(n10289) );
  AOI22_X1 U11338 ( .A1(n10287), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10288) );
  OAI221_X1 U11339 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10291), .C1(n10290), .C2(
        n10289), .A(n10288), .ZN(P2_U3245) );
  AND2_X1 U11340 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10303), .ZN(P2_U3297) );
  AND2_X1 U11341 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10303), .ZN(P2_U3298) );
  AND2_X1 U11342 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10303), .ZN(P2_U3299) );
  NOR2_X1 U11343 ( .A1(n10299), .A2(n10294), .ZN(P2_U3300) );
  AND2_X1 U11344 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10303), .ZN(P2_U3301) );
  AND2_X1 U11345 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10303), .ZN(P2_U3302) );
  AND2_X1 U11346 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10303), .ZN(P2_U3303) );
  AND2_X1 U11347 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10303), .ZN(P2_U3304) );
  AND2_X1 U11348 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10303), .ZN(P2_U3305) );
  AND2_X1 U11349 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10303), .ZN(P2_U3306) );
  AND2_X1 U11350 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10303), .ZN(P2_U3307) );
  AND2_X1 U11351 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10303), .ZN(P2_U3308) );
  AND2_X1 U11352 ( .A1(n10303), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3309) );
  AND2_X1 U11353 ( .A1(n10303), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3310) );
  NOR2_X1 U11354 ( .A1(n10299), .A2(n10295), .ZN(P2_U3311) );
  AND2_X1 U11355 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10303), .ZN(P2_U3312) );
  AND2_X1 U11356 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10303), .ZN(P2_U3313) );
  AND2_X1 U11357 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10303), .ZN(P2_U3314) );
  AND2_X1 U11358 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10303), .ZN(P2_U3315) );
  AND2_X1 U11359 ( .A1(n10303), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3316) );
  AND2_X1 U11360 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10303), .ZN(P2_U3317) );
  AND2_X1 U11361 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10303), .ZN(P2_U3318) );
  NOR2_X1 U11362 ( .A1(n10299), .A2(n10296), .ZN(P2_U3319) );
  AND2_X1 U11363 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10303), .ZN(P2_U3320) );
  NOR2_X1 U11364 ( .A1(n10299), .A2(n10297), .ZN(P2_U3321) );
  NOR2_X1 U11365 ( .A1(n10299), .A2(n10298), .ZN(P2_U3322) );
  AND2_X1 U11366 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10303), .ZN(P2_U3323) );
  AND2_X1 U11367 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10303), .ZN(P2_U3324) );
  AND2_X1 U11368 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10303), .ZN(P2_U3325) );
  AND2_X1 U11369 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10303), .ZN(P2_U3326) );
  AOI22_X1 U11370 ( .A1(n10306), .A2(n10301), .B1(n10300), .B2(n10303), .ZN(
        P2_U3437) );
  INV_X1 U11371 ( .A(n10302), .ZN(n10305) );
  AOI22_X1 U11372 ( .A1(n10306), .A2(n10305), .B1(n10304), .B2(n10303), .ZN(
        P2_U3438) );
  AOI22_X1 U11373 ( .A1(n10309), .A2(n10354), .B1(n10308), .B2(n10307), .ZN(
        n10310) );
  AND2_X1 U11374 ( .A1(n10311), .A2(n10310), .ZN(n10360) );
  INV_X1 U11375 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U11376 ( .A1(n10358), .A2(n10360), .B1(n10312), .B2(n10356), .ZN(
        P2_U3451) );
  OAI22_X1 U11377 ( .A1(n10313), .A2(n10350), .B1(n6741), .B2(n10348), .ZN(
        n10316) );
  INV_X1 U11378 ( .A(n10314), .ZN(n10315) );
  AOI211_X1 U11379 ( .C1(n10354), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        n10361) );
  AOI22_X1 U11380 ( .A1(n10358), .A2(n10361), .B1(n10318), .B2(n10356), .ZN(
        P2_U3454) );
  OAI22_X1 U11381 ( .A1(n10319), .A2(n10350), .B1(n4457), .B2(n10348), .ZN(
        n10321) );
  AOI211_X1 U11382 ( .C1(n10354), .C2(n10322), .A(n10321), .B(n10320), .ZN(
        n10363) );
  AOI22_X1 U11383 ( .A1(n10358), .A2(n10363), .B1(n5951), .B2(n10356), .ZN(
        P2_U3457) );
  OAI22_X1 U11384 ( .A1(n10324), .A2(n10350), .B1(n10323), .B2(n10348), .ZN(
        n10326) );
  AOI211_X1 U11385 ( .C1(n10354), .C2(n10327), .A(n10326), .B(n10325), .ZN(
        n10364) );
  INV_X1 U11386 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U11387 ( .A1(n10358), .A2(n10364), .B1(n10328), .B2(n10356), .ZN(
        P2_U3463) );
  OAI22_X1 U11388 ( .A1(n10330), .A2(n10350), .B1(n10329), .B2(n10348), .ZN(
        n10332) );
  AOI211_X1 U11389 ( .C1(n10354), .C2(n10333), .A(n10332), .B(n10331), .ZN(
        n10365) );
  INV_X1 U11390 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U11391 ( .A1(n10358), .A2(n10365), .B1(n10334), .B2(n10356), .ZN(
        P2_U3469) );
  NOR2_X1 U11392 ( .A1(n10336), .A2(n10335), .ZN(n10340) );
  OAI22_X1 U11393 ( .A1(n10338), .A2(n10350), .B1(n10337), .B2(n10348), .ZN(
        n10339) );
  NOR3_X1 U11394 ( .A1(n10341), .A2(n10340), .A3(n10339), .ZN(n10366) );
  AOI22_X1 U11395 ( .A1(n10358), .A2(n10366), .B1(n6027), .B2(n10356), .ZN(
        P2_U3475) );
  OAI22_X1 U11396 ( .A1(n10343), .A2(n10350), .B1(n10342), .B2(n10348), .ZN(
        n10344) );
  AOI211_X1 U11397 ( .C1(n10346), .C2(n10354), .A(n10345), .B(n10344), .ZN(
        n10367) );
  INV_X1 U11398 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U11399 ( .A1(n10358), .A2(n10367), .B1(n10347), .B2(n10356), .ZN(
        P2_U3481) );
  OAI22_X1 U11400 ( .A1(n10351), .A2(n10350), .B1(n10349), .B2(n10348), .ZN(
        n10353) );
  AOI211_X1 U11401 ( .C1(n10355), .C2(n10354), .A(n10353), .B(n10352), .ZN(
        n10369) );
  INV_X1 U11402 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U11403 ( .A1(n10358), .A2(n10369), .B1(n10357), .B2(n10356), .ZN(
        P2_U3487) );
  AOI22_X1 U11404 ( .A1(n10370), .A2(n10360), .B1(n10359), .B2(n10368), .ZN(
        P2_U3520) );
  AOI22_X1 U11405 ( .A1(n10370), .A2(n10361), .B1(n6898), .B2(n10368), .ZN(
        P2_U3521) );
  AOI22_X1 U11406 ( .A1(n10370), .A2(n10363), .B1(n10362), .B2(n10368), .ZN(
        P2_U3522) );
  AOI22_X1 U11407 ( .A1(n10370), .A2(n10364), .B1(n6900), .B2(n10368), .ZN(
        P2_U3524) );
  AOI22_X1 U11408 ( .A1(n10370), .A2(n10365), .B1(n7078), .B2(n10368), .ZN(
        P2_U3526) );
  AOI22_X1 U11409 ( .A1(n10370), .A2(n10366), .B1(n7113), .B2(n10368), .ZN(
        P2_U3528) );
  AOI22_X1 U11410 ( .A1(n10370), .A2(n10367), .B1(n7115), .B2(n10368), .ZN(
        P2_U3530) );
  AOI22_X1 U11411 ( .A1(n10370), .A2(n10369), .B1(n6076), .B2(n10368), .ZN(
        P2_U3532) );
  INV_X1 U11412 ( .A(n10371), .ZN(n10372) );
  NAND2_X1 U11413 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  XNOR2_X1 U11414 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10374), .ZN(ADD_1071_U5)
         );
  AOI22_X1 U11415 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n6648), .B2(n10375), .ZN(ADD_1071_U46) );
  OAI21_X1 U11416 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(ADD_1071_U56) );
  OAI21_X1 U11417 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(ADD_1071_U57) );
  OAI21_X1 U11418 ( .B1(n10384), .B2(n10383), .A(n10382), .ZN(ADD_1071_U58) );
  OAI21_X1 U11419 ( .B1(n10387), .B2(n10386), .A(n10385), .ZN(ADD_1071_U59) );
  OAI21_X1 U11420 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(ADD_1071_U60) );
  OAI21_X1 U11421 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(ADD_1071_U61) );
  AOI21_X1 U11422 ( .B1(n10396), .B2(n10395), .A(n10394), .ZN(ADD_1071_U62) );
  AOI21_X1 U11423 ( .B1(n10399), .B2(n10398), .A(n10397), .ZN(ADD_1071_U63) );
  XOR2_X1 U11424 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10400), .Z(ADD_1071_U50) );
  NOR2_X1 U11425 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  XOR2_X1 U11426 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10403), .Z(ADD_1071_U51) );
  OAI21_X1 U11427 ( .B1(n10406), .B2(n10405), .A(n10404), .ZN(n10407) );
  XNOR2_X1 U11428 ( .A(n10407), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11429 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(ADD_1071_U47) );
  XOR2_X1 U11430 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10411), .Z(ADD_1071_U48) );
  XOR2_X1 U11431 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10412), .Z(ADD_1071_U49) );
  XOR2_X1 U11432 ( .A(n10414), .B(n10413), .Z(ADD_1071_U54) );
  XOR2_X1 U11433 ( .A(n10416), .B(n10415), .Z(ADD_1071_U53) );
  XNOR2_X1 U11434 ( .A(n10418), .B(n10417), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4984 ( .A(n5948), .Z(n4466) );
  CLKBUF_X1 U5162 ( .A(n5128), .Z(n6555) );
endmodule

